VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2433.460 2924.800 2434.660 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2903.340 2924.800 2904.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3410.620 2.400 3411.820 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 2.400 3124.860 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2836.020 2.400 2837.220 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 2.400 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 2.400 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1974.460 2.400 1975.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 2.400 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 2.400 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 2.400 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 2.400 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 2.400 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 2.400 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 2.400 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 2.400 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1964.260 2924.800 1965.460 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2198.860 2924.800 2200.060 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 2.400 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 2.400 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 2.400 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 2.400 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 2.400 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 2.400 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 2.400 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 2.400 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 2.400 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 2.400 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 2.400 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 2.400 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.220 2.400 3340.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 2.400 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 2.400 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2476.980 2.400 2478.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 2.400 2190.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 2.400 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 2.400 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 2.400 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 2.400 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 2.400 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 2.400 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 2.400 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 2.400 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 656.565 24.565 659.495 24.735 ;
        RECT 650.585 24.055 650.755 24.395 ;
        RECT 650.585 23.885 652.595 24.055 ;
        RECT 656.565 23.885 656.735 24.565 ;
      LAYER mcon ;
        RECT 659.325 24.565 659.495 24.735 ;
        RECT 650.585 24.225 650.755 24.395 ;
        RECT 652.425 23.885 652.595 24.055 ;
      LAYER met1 ;
        RECT 659.265 24.720 659.555 24.765 ;
        RECT 1331.770 24.720 1332.090 24.780 ;
        RECT 659.265 24.580 1332.090 24.720 ;
        RECT 659.265 24.535 659.555 24.580 ;
        RECT 1331.770 24.520 1332.090 24.580 ;
        RECT 633.030 24.380 633.350 24.440 ;
        RECT 650.525 24.380 650.815 24.425 ;
        RECT 633.030 24.240 650.815 24.380 ;
        RECT 633.030 24.180 633.350 24.240 ;
        RECT 650.525 24.195 650.815 24.240 ;
        RECT 652.365 24.040 652.655 24.085 ;
        RECT 656.505 24.040 656.795 24.085 ;
        RECT 652.365 23.900 656.795 24.040 ;
        RECT 652.365 23.855 652.655 23.900 ;
        RECT 656.505 23.855 656.795 23.900 ;
      LAYER via ;
        RECT 1331.800 24.520 1332.060 24.780 ;
        RECT 633.060 24.180 633.320 24.440 ;
      LAYER met2 ;
        RECT 1336.010 1600.450 1336.290 1604.000 ;
        RECT 1331.860 1600.310 1336.290 1600.450 ;
        RECT 1331.860 24.810 1332.000 1600.310 ;
        RECT 1336.010 1600.000 1336.290 1600.310 ;
        RECT 1331.800 24.490 1332.060 24.810 ;
        RECT 633.060 24.150 633.320 24.470 ;
        RECT 633.120 2.400 633.260 24.150 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 24.380 651.290 24.440 ;
        RECT 1359.370 24.380 1359.690 24.440 ;
        RECT 650.970 24.240 1359.690 24.380 ;
        RECT 650.970 24.180 651.290 24.240 ;
        RECT 1359.370 24.180 1359.690 24.240 ;
      LAYER via ;
        RECT 651.000 24.180 651.260 24.440 ;
        RECT 1359.400 24.180 1359.660 24.440 ;
      LAYER met2 ;
        RECT 1365.450 1600.450 1365.730 1604.000 ;
        RECT 1359.460 1600.310 1365.730 1600.450 ;
        RECT 1359.460 24.470 1359.600 1600.310 ;
        RECT 1365.450 1600.000 1365.730 1600.310 ;
        RECT 651.000 24.150 651.260 24.470 ;
        RECT 1359.400 24.150 1359.660 24.470 ;
        RECT 651.060 2.400 651.200 24.150 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1346.130 1600.450 1346.410 1604.000 ;
        RECT 1345.660 1600.310 1346.410 1600.450 ;
        RECT 1345.660 25.685 1345.800 1600.310 ;
        RECT 1346.130 1600.000 1346.410 1600.310 ;
        RECT 639.030 25.315 639.310 25.685 ;
        RECT 1345.590 25.315 1345.870 25.685 ;
        RECT 639.100 2.400 639.240 25.315 ;
        RECT 638.890 -4.800 639.450 2.400 ;
      LAYER via2 ;
        RECT 639.030 25.360 639.310 25.640 ;
        RECT 1345.590 25.360 1345.870 25.640 ;
      LAYER met3 ;
        RECT 639.005 25.650 639.335 25.665 ;
        RECT 1345.565 25.650 1345.895 25.665 ;
        RECT 639.005 25.350 1345.895 25.650 ;
        RECT 639.005 25.335 639.335 25.350 ;
        RECT 1345.565 25.335 1345.895 25.350 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 24.040 657.270 24.100 ;
        RECT 1373.170 24.040 1373.490 24.100 ;
        RECT 656.950 23.900 1373.490 24.040 ;
        RECT 656.950 23.840 657.270 23.900 ;
        RECT 1373.170 23.840 1373.490 23.900 ;
      LAYER via ;
        RECT 656.980 23.840 657.240 24.100 ;
        RECT 1373.200 23.840 1373.460 24.100 ;
      LAYER met2 ;
        RECT 1375.110 1600.450 1375.390 1604.000 ;
        RECT 1373.260 1600.310 1375.390 1600.450 ;
        RECT 1373.260 24.130 1373.400 1600.310 ;
        RECT 1375.110 1600.000 1375.390 1600.310 ;
        RECT 656.980 23.810 657.240 24.130 ;
        RECT 1373.200 23.810 1373.460 24.130 ;
        RECT 657.040 2.400 657.180 23.810 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1394.430 1600.450 1394.710 1604.000 ;
        RECT 1393.960 1600.310 1394.710 1600.450 ;
        RECT 1393.960 24.325 1394.100 1600.310 ;
        RECT 1394.430 1600.000 1394.710 1600.310 ;
        RECT 674.450 23.955 674.730 24.325 ;
        RECT 1393.890 23.955 1394.170 24.325 ;
        RECT 674.520 2.400 674.660 23.955 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 674.450 24.000 674.730 24.280 ;
        RECT 1393.890 24.000 1394.170 24.280 ;
      LAYER met3 ;
        RECT 674.425 24.290 674.755 24.305 ;
        RECT 1393.865 24.290 1394.195 24.305 ;
        RECT 674.425 23.990 1394.195 24.290 ;
        RECT 674.425 23.975 674.755 23.990 ;
        RECT 1393.865 23.975 1394.195 23.990 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1355.790 1600.450 1356.070 1604.000 ;
        RECT 1352.560 1600.310 1356.070 1600.450 ;
        RECT 1352.560 26.365 1352.700 1600.310 ;
        RECT 1355.790 1600.000 1356.070 1600.310 ;
        RECT 645.010 25.995 645.290 26.365 ;
        RECT 1352.490 25.995 1352.770 26.365 ;
        RECT 645.080 2.400 645.220 25.995 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 645.010 26.040 645.290 26.320 ;
        RECT 1352.490 26.040 1352.770 26.320 ;
      LAYER met3 ;
        RECT 644.985 26.330 645.315 26.345 ;
        RECT 1352.465 26.330 1352.795 26.345 ;
        RECT 644.985 26.030 1352.795 26.330 ;
        RECT 644.985 26.015 645.315 26.030 ;
        RECT 1352.465 26.015 1352.795 26.030 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1384.770 1600.450 1385.050 1604.000 ;
        RECT 1380.160 1600.310 1385.050 1600.450 ;
        RECT 1380.160 25.005 1380.300 1600.310 ;
        RECT 1384.770 1600.000 1385.050 1600.310 ;
        RECT 662.950 24.635 663.230 25.005 ;
        RECT 1380.090 24.635 1380.370 25.005 ;
        RECT 663.020 2.400 663.160 24.635 ;
        RECT 662.810 -4.800 663.370 2.400 ;
      LAYER via2 ;
        RECT 662.950 24.680 663.230 24.960 ;
        RECT 1380.090 24.680 1380.370 24.960 ;
      LAYER met3 ;
        RECT 662.925 24.970 663.255 24.985 ;
        RECT 1380.065 24.970 1380.395 24.985 ;
        RECT 662.925 24.670 1380.395 24.970 ;
        RECT 662.925 24.655 663.255 24.670 ;
        RECT 1380.065 24.655 1380.395 24.670 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1569.130 2794.700 1569.450 2794.760 ;
        RECT 2069.610 2794.700 2069.930 2794.760 ;
        RECT 1566.460 2794.560 2069.930 2794.700 ;
        RECT 972.050 2794.360 972.370 2794.420 ;
        RECT 1566.460 2794.360 1566.600 2794.560 ;
        RECT 1569.130 2794.500 1569.450 2794.560 ;
        RECT 2069.610 2794.500 2069.930 2794.560 ;
        RECT 972.050 2794.220 1566.600 2794.360 ;
        RECT 972.050 2794.160 972.370 2794.220 ;
        RECT 2069.610 2792.320 2069.930 2792.380 ;
        RECT 2215.430 2792.320 2215.750 2792.380 ;
        RECT 2069.610 2792.180 2215.750 2792.320 ;
        RECT 2069.610 2792.120 2069.930 2792.180 ;
        RECT 2215.430 2792.120 2215.750 2792.180 ;
        RECT 2069.610 2068.120 2069.930 2068.180 ;
        RECT 2100.890 2068.120 2101.210 2068.180 ;
        RECT 2069.610 2067.980 2101.210 2068.120 ;
        RECT 2069.610 2067.920 2069.930 2067.980 ;
        RECT 2100.890 2067.920 2101.210 2067.980 ;
        RECT 1718.170 1593.820 1718.490 1593.880 ;
        RECT 2100.890 1593.820 2101.210 1593.880 ;
        RECT 2265.570 1593.820 2265.890 1593.880 ;
        RECT 1718.170 1593.680 2265.890 1593.820 ;
        RECT 1718.170 1593.620 1718.490 1593.680 ;
        RECT 2100.890 1593.620 2101.210 1593.680 ;
        RECT 2265.570 1593.620 2265.890 1593.680 ;
        RECT 306.890 1590.420 307.210 1590.480 ;
        RECT 1718.170 1590.420 1718.490 1590.480 ;
        RECT 306.890 1590.280 1718.490 1590.420 ;
        RECT 306.890 1590.220 307.210 1590.280 ;
        RECT 1718.170 1590.220 1718.490 1590.280 ;
        RECT 2.830 14.860 3.150 14.920 ;
        RECT 306.890 14.860 307.210 14.920 ;
        RECT 2.830 14.720 307.210 14.860 ;
        RECT 2.830 14.660 3.150 14.720 ;
        RECT 306.890 14.660 307.210 14.720 ;
      LAYER via ;
        RECT 972.080 2794.160 972.340 2794.420 ;
        RECT 1569.160 2794.500 1569.420 2794.760 ;
        RECT 2069.640 2794.500 2069.900 2794.760 ;
        RECT 2069.640 2792.120 2069.900 2792.380 ;
        RECT 2215.460 2792.120 2215.720 2792.380 ;
        RECT 2069.640 2067.920 2069.900 2068.180 ;
        RECT 2100.920 2067.920 2101.180 2068.180 ;
        RECT 1718.200 1593.620 1718.460 1593.880 ;
        RECT 2100.920 1593.620 2101.180 1593.880 ;
        RECT 2265.600 1593.620 2265.860 1593.880 ;
        RECT 306.920 1590.220 307.180 1590.480 ;
        RECT 1718.200 1590.220 1718.460 1590.480 ;
        RECT 2.860 14.660 3.120 14.920 ;
        RECT 306.920 14.660 307.180 14.920 ;
      LAYER met2 ;
        RECT 1569.160 2794.645 1569.420 2794.790 ;
        RECT 972.080 2794.130 972.340 2794.450 ;
        RECT 1569.150 2794.275 1569.430 2794.645 ;
        RECT 2069.640 2794.470 2069.900 2794.790 ;
        RECT 972.140 2793.965 972.280 2794.130 ;
        RECT 972.070 2793.595 972.350 2793.965 ;
        RECT 2069.700 2792.410 2069.840 2794.470 ;
        RECT 2215.450 2794.275 2215.730 2794.645 ;
        RECT 2215.520 2792.410 2215.660 2794.275 ;
        RECT 2069.640 2792.090 2069.900 2792.410 ;
        RECT 2215.460 2792.090 2215.720 2792.410 ;
        RECT 2069.700 2069.765 2069.840 2792.090 ;
        RECT 2069.630 2069.395 2069.910 2069.765 ;
        RECT 2069.700 2068.210 2069.840 2069.395 ;
        RECT 2069.640 2067.890 2069.900 2068.210 ;
        RECT 2100.920 2067.890 2101.180 2068.210 ;
        RECT 2100.980 2064.325 2101.120 2067.890 ;
        RECT 2100.910 2063.955 2101.190 2064.325 ;
        RECT 304.690 1600.450 304.970 1604.000 ;
        RECT 304.690 1600.310 307.120 1600.450 ;
        RECT 304.690 1600.000 304.970 1600.310 ;
        RECT 306.980 1590.510 307.120 1600.310 ;
        RECT 2100.980 1593.910 2101.120 2063.955 ;
        RECT 1718.200 1593.765 1718.460 1593.910 ;
        RECT 1718.190 1593.395 1718.470 1593.765 ;
        RECT 2100.920 1593.590 2101.180 1593.910 ;
        RECT 2265.600 1593.765 2265.860 1593.910 ;
        RECT 2265.590 1593.395 2265.870 1593.765 ;
        RECT 1718.260 1590.510 1718.400 1593.395 ;
        RECT 306.920 1590.190 307.180 1590.510 ;
        RECT 1718.200 1590.190 1718.460 1590.510 ;
        RECT 306.980 14.950 307.120 1590.190 ;
        RECT 2.860 14.630 3.120 14.950 ;
        RECT 306.920 14.630 307.180 14.950 ;
        RECT 2.920 2.400 3.060 14.630 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 1569.150 2794.320 1569.430 2794.600 ;
        RECT 972.070 2793.640 972.350 2793.920 ;
        RECT 2215.450 2794.320 2215.730 2794.600 ;
        RECT 2069.630 2069.440 2069.910 2069.720 ;
        RECT 2100.910 2064.000 2101.190 2064.280 ;
        RECT 1718.190 1593.440 1718.470 1593.720 ;
        RECT 2265.590 1593.440 2265.870 1593.720 ;
      LAYER met3 ;
        RECT 1569.125 2794.620 1569.455 2794.625 ;
        RECT 1568.870 2794.610 1569.455 2794.620 ;
        RECT 1568.670 2794.310 1569.455 2794.610 ;
        RECT 1568.870 2794.300 1569.455 2794.310 ;
        RECT 1569.125 2794.295 1569.455 2794.300 ;
        RECT 2215.425 2794.620 2215.755 2794.625 ;
        RECT 2215.425 2794.610 2216.010 2794.620 ;
        RECT 2215.425 2794.310 2216.210 2794.610 ;
        RECT 2215.425 2794.300 2216.010 2794.310 ;
        RECT 2215.425 2794.295 2215.755 2794.300 ;
        RECT 972.045 2793.940 972.375 2793.945 ;
        RECT 321.350 2793.930 321.730 2793.940 ;
        RECT 971.790 2793.930 972.375 2793.940 ;
        RECT 321.350 2793.630 972.375 2793.930 ;
        RECT 321.350 2793.620 321.730 2793.630 ;
        RECT 971.790 2793.620 972.375 2793.630 ;
        RECT 972.045 2793.615 972.375 2793.620 ;
        RECT 2069.605 2069.740 2069.935 2069.745 ;
        RECT 2069.350 2069.730 2069.935 2069.740 ;
        RECT 2069.150 2069.430 2069.935 2069.730 ;
        RECT 2069.350 2069.420 2069.935 2069.430 ;
        RECT 2069.605 2069.415 2069.935 2069.420 ;
        RECT 2100.885 2064.290 2101.215 2064.305 ;
        RECT 2614.910 2064.290 2615.290 2064.300 ;
        RECT 2100.885 2063.990 2615.290 2064.290 ;
        RECT 2100.885 2063.975 2101.215 2063.990 ;
        RECT 2614.910 2063.980 2615.290 2063.990 ;
        RECT 1718.165 1593.730 1718.495 1593.745 ;
        RECT 1719.750 1593.730 1720.130 1593.740 ;
        RECT 1718.165 1593.430 1720.130 1593.730 ;
        RECT 1718.165 1593.415 1718.495 1593.430 ;
        RECT 1719.750 1593.420 1720.130 1593.430 ;
        RECT 2265.565 1593.730 2265.895 1593.745 ;
        RECT 2266.230 1593.730 2266.610 1593.740 ;
        RECT 2265.565 1593.430 2266.610 1593.730 ;
        RECT 2265.565 1593.415 2265.895 1593.430 ;
        RECT 2266.230 1593.420 2266.610 1593.430 ;
      LAYER via3 ;
        RECT 1568.900 2794.300 1569.220 2794.620 ;
        RECT 2215.660 2794.300 2215.980 2794.620 ;
        RECT 321.380 2793.620 321.700 2793.940 ;
        RECT 971.820 2793.620 972.140 2793.940 ;
        RECT 2069.380 2069.420 2069.700 2069.740 ;
        RECT 2614.940 2063.980 2615.260 2064.300 ;
        RECT 1719.780 1593.420 1720.100 1593.740 ;
        RECT 2266.260 1593.420 2266.580 1593.740 ;
      LAYER met4 ;
        RECT 319.015 2801.750 319.315 2804.600 ;
        RECT 969.015 2801.750 969.315 2804.600 ;
        RECT 1569.015 2801.750 1569.315 2804.600 ;
        RECT 2219.015 2801.750 2219.315 2804.600 ;
        RECT 319.015 2801.450 321.690 2801.750 ;
        RECT 319.015 2800.000 319.315 2801.450 ;
        RECT 321.390 2793.945 321.690 2801.450 ;
        RECT 969.015 2801.450 972.130 2801.750 ;
        RECT 969.015 2800.000 969.315 2801.450 ;
        RECT 971.830 2793.945 972.130 2801.450 ;
        RECT 1568.910 2800.000 1569.315 2801.750 ;
        RECT 2215.670 2801.450 2219.315 2801.750 ;
        RECT 1568.910 2794.625 1569.210 2800.000 ;
        RECT 2215.670 2794.625 2215.970 2801.450 ;
        RECT 2219.015 2800.000 2219.315 2801.450 ;
        RECT 1568.895 2794.295 1569.225 2794.625 ;
        RECT 2215.655 2794.295 2215.985 2794.625 ;
        RECT 321.375 2793.615 321.705 2793.945 ;
        RECT 971.815 2793.615 972.145 2793.945 ;
        RECT 2069.375 2069.415 2069.705 2069.745 ;
        RECT 2067.165 2055.450 2067.465 2056.235 ;
        RECT 2069.390 2055.450 2069.690 2069.415 ;
        RECT 2614.935 2063.975 2615.265 2064.305 ;
        RECT 2067.165 2055.150 2069.690 2055.450 ;
        RECT 2614.950 2055.450 2615.250 2063.975 ;
        RECT 2617.865 2055.450 2618.165 2056.235 ;
        RECT 2614.950 2055.150 2618.165 2055.450 ;
        RECT 2067.165 2051.635 2067.465 2055.150 ;
        RECT 2617.865 2051.635 2618.165 2055.150 ;
        RECT 1718.315 1603.250 1718.615 1604.600 ;
        RECT 1718.315 1602.950 1720.090 1603.250 ;
        RECT 1718.315 1600.000 1718.615 1602.950 ;
        RECT 1719.790 1593.745 1720.090 1602.950 ;
        RECT 2269.015 1601.550 2269.315 1604.600 ;
        RECT 2266.270 1601.250 2269.315 1601.550 ;
        RECT 2266.270 1593.745 2266.570 1601.250 ;
        RECT 2269.015 1600.000 2269.315 1601.250 ;
        RECT 1719.775 1593.415 1720.105 1593.745 ;
        RECT 2266.255 1593.415 2266.585 1593.745 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 34.185 14.365 34.355 15.895 ;
      LAYER mcon ;
        RECT 34.185 15.725 34.355 15.895 ;
      LAYER met1 ;
        RECT 8.350 15.880 8.670 15.940 ;
        RECT 34.125 15.880 34.415 15.925 ;
        RECT 8.350 15.740 34.415 15.880 ;
        RECT 8.350 15.680 8.670 15.740 ;
        RECT 34.125 15.695 34.415 15.740 ;
        RECT 34.125 14.520 34.415 14.565 ;
        RECT 34.125 14.380 294.700 14.520 ;
        RECT 34.125 14.335 34.415 14.380 ;
        RECT 294.560 14.180 294.700 14.380 ;
        RECT 311.030 14.180 311.350 14.240 ;
        RECT 294.560 14.040 311.350 14.180 ;
        RECT 311.030 13.980 311.350 14.040 ;
      LAYER via ;
        RECT 8.380 15.680 8.640 15.940 ;
        RECT 311.060 13.980 311.320 14.240 ;
      LAYER met2 ;
        RECT 314.350 1600.450 314.630 1604.000 ;
        RECT 311.120 1600.310 314.630 1600.450 ;
        RECT 8.380 15.650 8.640 15.970 ;
        RECT 8.440 2.400 8.580 15.650 ;
        RECT 311.120 14.270 311.260 1600.310 ;
        RECT 314.350 1600.000 314.630 1600.310 ;
        RECT 311.060 13.950 311.320 14.270 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 292.705 14.025 292.875 16.915 ;
      LAYER mcon ;
        RECT 292.705 16.745 292.875 16.915 ;
      LAYER met1 ;
        RECT 292.645 16.900 292.935 16.945 ;
        RECT 318.390 16.900 318.710 16.960 ;
        RECT 292.645 16.760 318.710 16.900 ;
        RECT 292.645 16.715 292.935 16.760 ;
        RECT 318.390 16.700 318.710 16.760 ;
        RECT 14.330 14.180 14.650 14.240 ;
        RECT 292.645 14.180 292.935 14.225 ;
        RECT 14.330 14.040 292.935 14.180 ;
        RECT 14.330 13.980 14.650 14.040 ;
        RECT 292.645 13.995 292.935 14.040 ;
      LAYER via ;
        RECT 318.420 16.700 318.680 16.960 ;
        RECT 14.360 13.980 14.620 14.240 ;
      LAYER met2 ;
        RECT 324.010 1600.450 324.290 1604.000 ;
        RECT 318.480 1600.310 324.290 1600.450 ;
        RECT 318.480 16.990 318.620 1600.310 ;
        RECT 324.010 1600.000 324.290 1600.310 ;
        RECT 318.420 16.670 318.680 16.990 ;
        RECT 14.360 13.950 14.620 14.270 ;
        RECT 14.420 2.400 14.560 13.950 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 15.880 38.570 15.940 ;
        RECT 38.250 15.740 342.080 15.880 ;
        RECT 38.250 15.680 38.570 15.740 ;
        RECT 341.940 15.200 342.080 15.740 ;
        RECT 359.790 15.540 360.110 15.600 ;
        RECT 352.520 15.400 360.110 15.540 ;
        RECT 352.520 15.200 352.660 15.400 ;
        RECT 359.790 15.340 360.110 15.400 ;
        RECT 341.940 15.060 352.660 15.200 ;
      LAYER via ;
        RECT 38.280 15.680 38.540 15.940 ;
        RECT 359.820 15.340 360.080 15.600 ;
      LAYER met2 ;
        RECT 362.650 1600.450 362.930 1604.000 ;
        RECT 359.880 1600.310 362.930 1600.450 ;
        RECT 38.280 15.650 38.540 15.970 ;
        RECT 38.340 2.400 38.480 15.650 ;
        RECT 359.880 15.630 360.020 1600.310 ;
        RECT 362.650 1600.000 362.930 1600.310 ;
        RECT 359.820 15.310 360.080 15.630 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 241.110 20.980 241.430 21.040 ;
        RECT 690.070 20.980 690.390 21.040 ;
        RECT 241.110 20.840 690.390 20.980 ;
        RECT 241.110 20.780 241.430 20.840 ;
        RECT 690.070 20.780 690.390 20.840 ;
      LAYER via ;
        RECT 241.140 20.780 241.400 21.040 ;
        RECT 690.100 20.780 690.360 21.040 ;
      LAYER met2 ;
        RECT 693.850 1600.450 694.130 1604.000 ;
        RECT 690.160 1600.310 694.130 1600.450 ;
        RECT 690.160 21.070 690.300 1600.310 ;
        RECT 693.850 1600.000 694.130 1600.310 ;
        RECT 241.140 20.750 241.400 21.070 ;
        RECT 690.100 20.750 690.360 21.070 ;
        RECT 241.200 10.610 241.340 20.750 ;
        RECT 240.740 10.470 241.340 10.610 ;
        RECT 240.740 2.400 240.880 10.470 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 21.320 258.450 21.380 ;
        RECT 717.670 21.320 717.990 21.380 ;
        RECT 258.130 21.180 717.990 21.320 ;
        RECT 258.130 21.120 258.450 21.180 ;
        RECT 717.670 21.120 717.990 21.180 ;
      LAYER via ;
        RECT 258.160 21.120 258.420 21.380 ;
        RECT 717.700 21.120 717.960 21.380 ;
      LAYER met2 ;
        RECT 722.830 1600.450 723.110 1604.000 ;
        RECT 717.760 1600.310 723.110 1600.450 ;
        RECT 717.760 21.410 717.900 1600.310 ;
        RECT 722.830 1600.000 723.110 1600.310 ;
        RECT 258.160 21.090 258.420 21.410 ;
        RECT 717.700 21.090 717.960 21.410 ;
        RECT 258.220 2.400 258.360 21.090 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 21.660 276.390 21.720 ;
        RECT 752.170 21.660 752.490 21.720 ;
        RECT 276.070 21.520 752.490 21.660 ;
        RECT 276.070 21.460 276.390 21.520 ;
        RECT 752.170 21.460 752.490 21.520 ;
      LAYER via ;
        RECT 276.100 21.460 276.360 21.720 ;
        RECT 752.200 21.460 752.460 21.720 ;
      LAYER met2 ;
        RECT 752.270 1600.380 752.550 1604.000 ;
        RECT 752.260 1600.000 752.550 1600.380 ;
        RECT 752.260 21.750 752.400 1600.000 ;
        RECT 276.100 21.430 276.360 21.750 ;
        RECT 752.200 21.430 752.460 21.750 ;
        RECT 276.160 2.400 276.300 21.430 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 22.000 294.330 22.060 ;
        RECT 779.770 22.000 780.090 22.060 ;
        RECT 294.010 21.860 780.090 22.000 ;
        RECT 294.010 21.800 294.330 21.860 ;
        RECT 779.770 21.800 780.090 21.860 ;
      LAYER via ;
        RECT 294.040 21.800 294.300 22.060 ;
        RECT 779.800 21.800 780.060 22.060 ;
      LAYER met2 ;
        RECT 781.250 1600.450 781.530 1604.000 ;
        RECT 779.860 1600.310 781.530 1600.450 ;
        RECT 779.860 22.090 780.000 1600.310 ;
        RECT 781.250 1600.000 781.530 1600.310 ;
        RECT 294.040 21.770 294.300 22.090 ;
        RECT 779.800 21.770 780.060 22.090 ;
        RECT 294.100 2.400 294.240 21.770 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 22.340 312.270 22.400 ;
        RECT 807.370 22.340 807.690 22.400 ;
        RECT 311.950 22.200 807.690 22.340 ;
        RECT 311.950 22.140 312.270 22.200 ;
        RECT 807.370 22.140 807.690 22.200 ;
      LAYER via ;
        RECT 311.980 22.140 312.240 22.400 ;
        RECT 807.400 22.140 807.660 22.400 ;
      LAYER met2 ;
        RECT 810.690 1600.450 810.970 1604.000 ;
        RECT 807.460 1600.310 810.970 1600.450 ;
        RECT 807.460 22.430 807.600 1600.310 ;
        RECT 810.690 1600.000 810.970 1600.310 ;
        RECT 311.980 22.110 312.240 22.430 ;
        RECT 807.400 22.110 807.660 22.430 ;
        RECT 312.040 2.400 312.180 22.110 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 22.680 330.210 22.740 ;
        RECT 834.970 22.680 835.290 22.740 ;
        RECT 329.890 22.540 835.290 22.680 ;
        RECT 329.890 22.480 330.210 22.540 ;
        RECT 834.970 22.480 835.290 22.540 ;
      LAYER via ;
        RECT 329.920 22.480 330.180 22.740 ;
        RECT 835.000 22.480 835.260 22.740 ;
      LAYER met2 ;
        RECT 839.670 1600.450 839.950 1604.000 ;
        RECT 835.060 1600.310 839.950 1600.450 ;
        RECT 835.060 22.770 835.200 1600.310 ;
        RECT 839.670 1600.000 839.950 1600.310 ;
        RECT 329.920 22.450 330.180 22.770 ;
        RECT 835.000 22.450 835.260 22.770 ;
        RECT 329.980 2.400 330.120 22.450 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 23.020 347.690 23.080 ;
        RECT 862.570 23.020 862.890 23.080 ;
        RECT 347.370 22.880 862.890 23.020 ;
        RECT 347.370 22.820 347.690 22.880 ;
        RECT 862.570 22.820 862.890 22.880 ;
      LAYER via ;
        RECT 347.400 22.820 347.660 23.080 ;
        RECT 862.600 22.820 862.860 23.080 ;
      LAYER met2 ;
        RECT 869.110 1600.450 869.390 1604.000 ;
        RECT 862.660 1600.310 869.390 1600.450 ;
        RECT 862.660 23.110 862.800 1600.310 ;
        RECT 869.110 1600.000 869.390 1600.310 ;
        RECT 347.400 22.790 347.660 23.110 ;
        RECT 862.600 22.790 862.860 23.110 ;
        RECT 347.460 2.400 347.600 22.790 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 23.360 365.630 23.420 ;
        RECT 897.070 23.360 897.390 23.420 ;
        RECT 365.310 23.220 897.390 23.360 ;
        RECT 365.310 23.160 365.630 23.220 ;
        RECT 897.070 23.160 897.390 23.220 ;
      LAYER via ;
        RECT 365.340 23.160 365.600 23.420 ;
        RECT 897.100 23.160 897.360 23.420 ;
      LAYER met2 ;
        RECT 898.090 1600.450 898.370 1604.000 ;
        RECT 897.160 1600.310 898.370 1600.450 ;
        RECT 897.160 23.450 897.300 1600.310 ;
        RECT 898.090 1600.000 898.370 1600.310 ;
        RECT 365.340 23.130 365.600 23.450 ;
        RECT 897.100 23.130 897.360 23.450 ;
        RECT 365.400 2.400 365.540 23.130 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 23.700 383.570 23.760 ;
        RECT 924.670 23.700 924.990 23.760 ;
        RECT 383.250 23.560 924.990 23.700 ;
        RECT 383.250 23.500 383.570 23.560 ;
        RECT 924.670 23.500 924.990 23.560 ;
      LAYER via ;
        RECT 383.280 23.500 383.540 23.760 ;
        RECT 924.700 23.500 924.960 23.760 ;
      LAYER met2 ;
        RECT 927.530 1600.450 927.810 1604.000 ;
        RECT 924.760 1600.310 927.810 1600.450 ;
        RECT 924.760 23.790 924.900 1600.310 ;
        RECT 927.530 1600.000 927.810 1600.310 ;
        RECT 383.280 23.470 383.540 23.790 ;
        RECT 924.700 23.470 924.960 23.790 ;
        RECT 383.340 2.400 383.480 23.470 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 27.440 401.510 27.500 ;
        RECT 952.270 27.440 952.590 27.500 ;
        RECT 401.190 27.300 952.590 27.440 ;
        RECT 401.190 27.240 401.510 27.300 ;
        RECT 952.270 27.240 952.590 27.300 ;
      LAYER via ;
        RECT 401.220 27.240 401.480 27.500 ;
        RECT 952.300 27.240 952.560 27.500 ;
      LAYER met2 ;
        RECT 956.510 1600.450 956.790 1604.000 ;
        RECT 952.360 1600.310 956.790 1600.450 ;
        RECT 952.360 27.530 952.500 1600.310 ;
        RECT 956.510 1600.000 956.790 1600.310 ;
        RECT 401.220 27.210 401.480 27.530 ;
        RECT 952.300 27.210 952.560 27.530 ;
        RECT 401.280 2.400 401.420 27.210 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 276.145 13.345 276.315 16.915 ;
        RECT 317.545 14.705 319.095 14.875 ;
        RECT 323.985 14.705 324.155 16.915 ;
        RECT 317.545 14.025 317.715 14.705 ;
      LAYER mcon ;
        RECT 276.145 16.745 276.315 16.915 ;
        RECT 323.985 16.745 324.155 16.915 ;
        RECT 318.925 14.705 319.095 14.875 ;
      LAYER met1 ;
        RECT 62.170 16.900 62.490 16.960 ;
        RECT 276.085 16.900 276.375 16.945 ;
        RECT 62.170 16.760 276.375 16.900 ;
        RECT 62.170 16.700 62.490 16.760 ;
        RECT 276.085 16.715 276.375 16.760 ;
        RECT 323.925 16.900 324.215 16.945 ;
        RECT 323.925 16.760 384.860 16.900 ;
        RECT 323.925 16.715 324.215 16.760 ;
        RECT 384.720 16.560 384.860 16.760 ;
        RECT 400.730 16.560 401.050 16.620 ;
        RECT 384.720 16.420 401.050 16.560 ;
        RECT 400.730 16.360 401.050 16.420 ;
        RECT 318.865 14.860 319.155 14.905 ;
        RECT 323.925 14.860 324.215 14.905 ;
        RECT 318.865 14.720 324.215 14.860 ;
        RECT 318.865 14.675 319.155 14.720 ;
        RECT 323.925 14.675 324.215 14.720 ;
        RECT 317.485 14.180 317.775 14.225 ;
        RECT 311.580 14.040 317.775 14.180 ;
        RECT 276.085 13.500 276.375 13.545 ;
        RECT 311.580 13.500 311.720 14.040 ;
        RECT 317.485 13.995 317.775 14.040 ;
        RECT 276.085 13.360 311.720 13.500 ;
        RECT 276.085 13.315 276.375 13.360 ;
      LAYER via ;
        RECT 62.200 16.700 62.460 16.960 ;
        RECT 400.760 16.360 401.020 16.620 ;
      LAYER met2 ;
        RECT 401.750 1600.450 402.030 1604.000 ;
        RECT 400.820 1600.310 402.030 1600.450 ;
        RECT 62.200 16.670 62.460 16.990 ;
        RECT 62.260 2.400 62.400 16.670 ;
        RECT 400.820 16.650 400.960 1600.310 ;
        RECT 401.750 1600.000 402.030 1600.310 ;
        RECT 400.760 16.330 401.020 16.650 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 27.100 419.450 27.160 ;
        RECT 979.870 27.100 980.190 27.160 ;
        RECT 419.130 26.960 980.190 27.100 ;
        RECT 419.130 26.900 419.450 26.960 ;
        RECT 979.870 26.900 980.190 26.960 ;
      LAYER via ;
        RECT 419.160 26.900 419.420 27.160 ;
        RECT 979.900 26.900 980.160 27.160 ;
      LAYER met2 ;
        RECT 985.950 1600.450 986.230 1604.000 ;
        RECT 979.960 1600.310 986.230 1600.450 ;
        RECT 979.960 27.190 980.100 1600.310 ;
        RECT 985.950 1600.000 986.230 1600.310 ;
        RECT 419.160 26.870 419.420 27.190 ;
        RECT 979.900 26.870 980.160 27.190 ;
        RECT 419.220 2.400 419.360 26.870 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 26.760 436.930 26.820 ;
        RECT 1014.370 26.760 1014.690 26.820 ;
        RECT 436.610 26.620 1014.690 26.760 ;
        RECT 436.610 26.560 436.930 26.620 ;
        RECT 1014.370 26.560 1014.690 26.620 ;
      LAYER via ;
        RECT 436.640 26.560 436.900 26.820 ;
        RECT 1014.400 26.560 1014.660 26.820 ;
      LAYER met2 ;
        RECT 1014.930 1600.450 1015.210 1604.000 ;
        RECT 1014.460 1600.310 1015.210 1600.450 ;
        RECT 1014.460 26.850 1014.600 1600.310 ;
        RECT 1014.930 1600.000 1015.210 1600.310 ;
        RECT 436.640 26.530 436.900 26.850 ;
        RECT 1014.400 26.530 1014.660 26.850 ;
        RECT 436.700 2.400 436.840 26.530 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 455.010 26.420 455.330 26.480 ;
        RECT 1041.970 26.420 1042.290 26.480 ;
        RECT 455.010 26.280 1042.290 26.420 ;
        RECT 455.010 26.220 455.330 26.280 ;
        RECT 1041.970 26.220 1042.290 26.280 ;
      LAYER via ;
        RECT 455.040 26.220 455.300 26.480 ;
        RECT 1042.000 26.220 1042.260 26.480 ;
      LAYER met2 ;
        RECT 1044.370 1600.450 1044.650 1604.000 ;
        RECT 1042.060 1600.310 1044.650 1600.450 ;
        RECT 1042.060 26.510 1042.200 1600.310 ;
        RECT 1044.370 1600.000 1044.650 1600.310 ;
        RECT 455.040 26.190 455.300 26.510 ;
        RECT 1042.000 26.190 1042.260 26.510 ;
        RECT 455.100 13.330 455.240 26.190 ;
        RECT 454.640 13.190 455.240 13.330 ;
        RECT 454.640 2.400 454.780 13.190 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 26.080 472.810 26.140 ;
        RECT 1069.570 26.080 1069.890 26.140 ;
        RECT 472.490 25.940 1069.890 26.080 ;
        RECT 472.490 25.880 472.810 25.940 ;
        RECT 1069.570 25.880 1069.890 25.940 ;
      LAYER via ;
        RECT 472.520 25.880 472.780 26.140 ;
        RECT 1069.600 25.880 1069.860 26.140 ;
      LAYER met2 ;
        RECT 1073.350 1600.450 1073.630 1604.000 ;
        RECT 1069.660 1600.310 1073.630 1600.450 ;
        RECT 1069.660 26.170 1069.800 1600.310 ;
        RECT 1073.350 1600.000 1073.630 1600.310 ;
        RECT 472.520 25.850 472.780 26.170 ;
        RECT 1069.600 25.850 1069.860 26.170 ;
        RECT 472.580 2.400 472.720 25.850 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 490.430 25.740 490.750 25.800 ;
        RECT 1097.170 25.740 1097.490 25.800 ;
        RECT 490.430 25.600 1097.490 25.740 ;
        RECT 490.430 25.540 490.750 25.600 ;
        RECT 1097.170 25.540 1097.490 25.600 ;
      LAYER via ;
        RECT 490.460 25.540 490.720 25.800 ;
        RECT 1097.200 25.540 1097.460 25.800 ;
      LAYER met2 ;
        RECT 1102.790 1600.450 1103.070 1604.000 ;
        RECT 1097.260 1600.310 1103.070 1600.450 ;
        RECT 1097.260 25.830 1097.400 1600.310 ;
        RECT 1102.790 1600.000 1103.070 1600.310 ;
        RECT 490.460 25.510 490.720 25.830 ;
        RECT 1097.200 25.510 1097.460 25.830 ;
        RECT 490.520 2.400 490.660 25.510 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 25.400 508.230 25.460 ;
        RECT 1131.670 25.400 1131.990 25.460 ;
        RECT 507.910 25.260 1131.990 25.400 ;
        RECT 507.910 25.200 508.230 25.260 ;
        RECT 1131.670 25.200 1131.990 25.260 ;
      LAYER via ;
        RECT 507.940 25.200 508.200 25.460 ;
        RECT 1131.700 25.200 1131.960 25.460 ;
      LAYER met2 ;
        RECT 1131.770 1600.380 1132.050 1604.000 ;
        RECT 1131.760 1600.000 1132.050 1600.380 ;
        RECT 1131.760 25.490 1131.900 1600.000 ;
        RECT 507.940 25.170 508.200 25.490 ;
        RECT 1131.700 25.170 1131.960 25.490 ;
        RECT 508.000 2.400 508.140 25.170 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 25.060 526.170 25.120 ;
        RECT 1159.270 25.060 1159.590 25.120 ;
        RECT 525.850 24.920 1159.590 25.060 ;
        RECT 525.850 24.860 526.170 24.920 ;
        RECT 1159.270 24.860 1159.590 24.920 ;
      LAYER via ;
        RECT 525.880 24.860 526.140 25.120 ;
        RECT 1159.300 24.860 1159.560 25.120 ;
      LAYER met2 ;
        RECT 1161.210 1600.450 1161.490 1604.000 ;
        RECT 1159.360 1600.310 1161.490 1600.450 ;
        RECT 1159.360 25.150 1159.500 1600.310 ;
        RECT 1161.210 1600.000 1161.490 1600.310 ;
        RECT 525.880 24.830 526.140 25.150 ;
        RECT 1159.300 24.830 1159.560 25.150 ;
        RECT 525.940 2.400 526.080 24.830 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1190.190 1600.450 1190.470 1604.000 ;
        RECT 1186.960 1600.310 1190.470 1600.450 ;
        RECT 1186.960 27.725 1187.100 1600.310 ;
        RECT 1190.190 1600.000 1190.470 1600.310 ;
        RECT 543.810 27.355 544.090 27.725 ;
        RECT 1186.890 27.355 1187.170 27.725 ;
        RECT 543.880 2.400 544.020 27.355 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 543.810 27.400 544.090 27.680 ;
        RECT 1186.890 27.400 1187.170 27.680 ;
      LAYER met3 ;
        RECT 543.785 27.690 544.115 27.705 ;
        RECT 1186.865 27.690 1187.195 27.705 ;
        RECT 543.785 27.390 1187.195 27.690 ;
        RECT 543.785 27.375 544.115 27.390 ;
        RECT 1186.865 27.375 1187.195 27.390 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1219.170 1600.450 1219.450 1604.000 ;
        RECT 1214.560 1600.310 1219.450 1600.450 ;
        RECT 1214.560 27.045 1214.700 1600.310 ;
        RECT 1219.170 1600.000 1219.450 1600.310 ;
        RECT 561.750 26.675 562.030 27.045 ;
        RECT 1214.490 26.675 1214.770 27.045 ;
        RECT 561.820 2.400 561.960 26.675 ;
        RECT 561.610 -4.800 562.170 2.400 ;
      LAYER via2 ;
        RECT 561.750 26.720 562.030 27.000 ;
        RECT 1214.490 26.720 1214.770 27.000 ;
      LAYER met3 ;
        RECT 561.725 27.010 562.055 27.025 ;
        RECT 1214.465 27.010 1214.795 27.025 ;
        RECT 561.725 26.710 1214.795 27.010 ;
        RECT 561.725 26.695 562.055 26.710 ;
        RECT 1214.465 26.695 1214.795 26.710 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 665.690 1593.820 666.010 1593.880 ;
        RECT 1248.510 1593.820 1248.830 1593.880 ;
        RECT 665.690 1593.680 1248.830 1593.820 ;
        RECT 665.690 1593.620 666.010 1593.680 ;
        RECT 1248.510 1593.620 1248.830 1593.680 ;
      LAYER via ;
        RECT 665.720 1593.620 665.980 1593.880 ;
        RECT 1248.540 1593.620 1248.800 1593.880 ;
      LAYER met2 ;
        RECT 1248.610 1600.380 1248.890 1604.000 ;
        RECT 1248.600 1600.000 1248.890 1600.380 ;
        RECT 1248.600 1593.910 1248.740 1600.000 ;
        RECT 665.720 1593.590 665.980 1593.910 ;
        RECT 1248.540 1593.590 1248.800 1593.910 ;
        RECT 665.780 24.325 665.920 1593.590 ;
        RECT 579.690 23.955 579.970 24.325 ;
        RECT 665.710 23.955 665.990 24.325 ;
        RECT 579.760 2.400 579.900 23.955 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 579.690 24.000 579.970 24.280 ;
        RECT 665.710 24.000 665.990 24.280 ;
      LAYER met3 ;
        RECT 579.665 24.290 579.995 24.305 ;
        RECT 665.685 24.290 666.015 24.305 ;
        RECT 579.665 23.990 666.015 24.290 ;
        RECT 579.665 23.975 579.995 23.990 ;
        RECT 665.685 23.975 666.015 23.990 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 19.960 86.410 20.020 ;
        RECT 434.770 19.960 435.090 20.020 ;
        RECT 86.090 19.820 435.090 19.960 ;
        RECT 86.090 19.760 86.410 19.820 ;
        RECT 434.770 19.760 435.090 19.820 ;
      LAYER via ;
        RECT 86.120 19.760 86.380 20.020 ;
        RECT 434.800 19.760 435.060 20.020 ;
      LAYER met2 ;
        RECT 440.850 1600.450 441.130 1604.000 ;
        RECT 434.860 1600.310 441.130 1600.450 ;
        RECT 434.860 20.050 435.000 1600.310 ;
        RECT 440.850 1600.000 441.130 1600.310 ;
        RECT 86.120 19.730 86.380 20.050 ;
        RECT 434.800 19.730 435.060 20.050 ;
        RECT 86.180 2.400 86.320 19.730 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 17.920 597.470 17.980 ;
        RECT 1276.570 17.920 1276.890 17.980 ;
        RECT 597.150 17.780 1276.890 17.920 ;
        RECT 597.150 17.720 597.470 17.780 ;
        RECT 1276.570 17.720 1276.890 17.780 ;
      LAYER via ;
        RECT 597.180 17.720 597.440 17.980 ;
        RECT 1276.600 17.720 1276.860 17.980 ;
      LAYER met2 ;
        RECT 1277.590 1600.450 1277.870 1604.000 ;
        RECT 1276.660 1600.310 1277.870 1600.450 ;
        RECT 1276.660 18.010 1276.800 1600.310 ;
        RECT 1277.590 1600.000 1277.870 1600.310 ;
        RECT 597.180 17.690 597.440 18.010 ;
        RECT 1276.600 17.690 1276.860 18.010 ;
        RECT 597.240 2.400 597.380 17.690 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 651.890 1591.440 652.210 1591.500 ;
        RECT 1306.930 1591.440 1307.250 1591.500 ;
        RECT 651.890 1591.300 1307.250 1591.440 ;
        RECT 651.890 1591.240 652.210 1591.300 ;
        RECT 1306.930 1591.240 1307.250 1591.300 ;
        RECT 615.090 24.040 615.410 24.100 ;
        RECT 651.890 24.040 652.210 24.100 ;
        RECT 615.090 23.900 652.210 24.040 ;
        RECT 615.090 23.840 615.410 23.900 ;
        RECT 651.890 23.840 652.210 23.900 ;
      LAYER via ;
        RECT 651.920 1591.240 652.180 1591.500 ;
        RECT 1306.960 1591.240 1307.220 1591.500 ;
        RECT 615.120 23.840 615.380 24.100 ;
        RECT 651.920 23.840 652.180 24.100 ;
      LAYER met2 ;
        RECT 1307.030 1600.380 1307.310 1604.000 ;
        RECT 1307.020 1600.000 1307.310 1600.380 ;
        RECT 1307.020 1591.530 1307.160 1600.000 ;
        RECT 651.920 1591.210 652.180 1591.530 ;
        RECT 1306.960 1591.210 1307.220 1591.530 ;
        RECT 651.980 24.130 652.120 1591.210 ;
        RECT 615.120 23.810 615.380 24.130 ;
        RECT 651.920 23.810 652.180 24.130 ;
        RECT 615.180 2.400 615.320 23.810 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 476.170 19.280 476.490 19.340 ;
        RECT 110.560 19.140 476.490 19.280 ;
        RECT 109.550 18.940 109.870 19.000 ;
        RECT 110.560 18.940 110.700 19.140 ;
        RECT 476.170 19.080 476.490 19.140 ;
        RECT 109.550 18.800 110.700 18.940 ;
        RECT 109.550 18.740 109.870 18.800 ;
      LAYER via ;
        RECT 109.580 18.740 109.840 19.000 ;
        RECT 476.200 19.080 476.460 19.340 ;
      LAYER met2 ;
        RECT 479.490 1600.450 479.770 1604.000 ;
        RECT 476.260 1600.310 479.770 1600.450 ;
        RECT 476.260 19.370 476.400 1600.310 ;
        RECT 479.490 1600.000 479.770 1600.310 ;
        RECT 476.200 19.050 476.460 19.370 ;
        RECT 109.580 18.710 109.840 19.030 ;
        RECT 109.640 2.400 109.780 18.710 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 18.260 133.790 18.320 ;
        RECT 517.570 18.260 517.890 18.320 ;
        RECT 133.470 18.120 517.890 18.260 ;
        RECT 133.470 18.060 133.790 18.120 ;
        RECT 517.570 18.060 517.890 18.120 ;
      LAYER via ;
        RECT 133.500 18.060 133.760 18.320 ;
        RECT 517.600 18.060 517.860 18.320 ;
      LAYER met2 ;
        RECT 518.590 1600.450 518.870 1604.000 ;
        RECT 517.660 1600.310 518.870 1600.450 ;
        RECT 517.660 18.350 517.800 1600.310 ;
        RECT 518.590 1600.000 518.870 1600.310 ;
        RECT 133.500 18.030 133.760 18.350 ;
        RECT 517.600 18.030 517.860 18.350 ;
        RECT 133.560 2.400 133.700 18.030 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 179.545 17.085 179.715 17.935 ;
      LAYER mcon ;
        RECT 179.545 17.765 179.715 17.935 ;
      LAYER met1 ;
        RECT 545.170 18.260 545.490 18.320 ;
        RECT 519.500 18.120 545.490 18.260 ;
        RECT 179.485 17.920 179.775 17.965 ;
        RECT 519.500 17.920 519.640 18.120 ;
        RECT 545.170 18.060 545.490 18.120 ;
        RECT 179.485 17.780 519.640 17.920 ;
        RECT 179.485 17.735 179.775 17.780 ;
        RECT 150.950 17.240 151.270 17.300 ;
        RECT 179.485 17.240 179.775 17.285 ;
        RECT 150.950 17.100 179.775 17.240 ;
        RECT 150.950 17.040 151.270 17.100 ;
        RECT 179.485 17.055 179.775 17.100 ;
      LAYER via ;
        RECT 545.200 18.060 545.460 18.320 ;
        RECT 150.980 17.040 151.240 17.300 ;
      LAYER met2 ;
        RECT 547.570 1600.450 547.850 1604.000 ;
        RECT 545.260 1600.310 547.850 1600.450 ;
        RECT 545.260 18.350 545.400 1600.310 ;
        RECT 547.570 1600.000 547.850 1600.310 ;
        RECT 545.200 18.030 545.460 18.350 ;
        RECT 150.980 17.010 151.240 17.330 ;
        RECT 151.040 8.570 151.180 17.010 ;
        RECT 151.040 8.430 151.640 8.570 ;
        RECT 151.500 2.400 151.640 8.430 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 17.580 169.670 17.640 ;
        RECT 572.770 17.580 573.090 17.640 ;
        RECT 169.350 17.440 573.090 17.580 ;
        RECT 169.350 17.380 169.670 17.440 ;
        RECT 572.770 17.380 573.090 17.440 ;
      LAYER via ;
        RECT 169.380 17.380 169.640 17.640 ;
        RECT 572.800 17.380 573.060 17.640 ;
      LAYER met2 ;
        RECT 577.010 1600.450 577.290 1604.000 ;
        RECT 572.860 1600.310 577.290 1600.450 ;
        RECT 572.860 17.670 573.000 1600.310 ;
        RECT 577.010 1600.000 577.290 1600.310 ;
        RECT 169.380 17.350 169.640 17.670 ;
        RECT 572.800 17.350 573.060 17.670 ;
        RECT 169.440 2.400 169.580 17.350 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 24.040 187.150 24.100 ;
        RECT 600.370 24.040 600.690 24.100 ;
        RECT 186.830 23.900 600.690 24.040 ;
        RECT 186.830 23.840 187.150 23.900 ;
        RECT 600.370 23.840 600.690 23.900 ;
      LAYER via ;
        RECT 186.860 23.840 187.120 24.100 ;
        RECT 600.400 23.840 600.660 24.100 ;
      LAYER met2 ;
        RECT 605.990 1600.450 606.270 1604.000 ;
        RECT 600.460 1600.310 606.270 1600.450 ;
        RECT 600.460 24.130 600.600 1600.310 ;
        RECT 605.990 1600.000 606.270 1600.310 ;
        RECT 186.860 23.810 187.120 24.130 ;
        RECT 600.400 23.810 600.660 24.130 ;
        RECT 186.920 2.400 187.060 23.810 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 635.430 1600.450 635.710 1604.000 ;
        RECT 634.960 1600.310 635.710 1600.450 ;
        RECT 634.960 19.565 635.100 1600.310 ;
        RECT 635.430 1600.000 635.710 1600.310 ;
        RECT 204.790 19.195 205.070 19.565 ;
        RECT 634.890 19.195 635.170 19.565 ;
        RECT 204.860 2.400 205.000 19.195 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 204.790 19.240 205.070 19.520 ;
        RECT 634.890 19.240 635.170 19.520 ;
      LAYER met3 ;
        RECT 204.765 19.530 205.095 19.545 ;
        RECT 634.865 19.530 635.195 19.545 ;
        RECT 204.765 19.230 635.195 19.530 ;
        RECT 204.765 19.215 205.095 19.230 ;
        RECT 634.865 19.215 635.195 19.230 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 655.185 1587.545 655.355 1593.835 ;
      LAYER mcon ;
        RECT 655.185 1593.665 655.355 1593.835 ;
      LAYER met1 ;
        RECT 655.125 1593.820 655.415 1593.865 ;
        RECT 664.310 1593.820 664.630 1593.880 ;
        RECT 655.125 1593.680 664.630 1593.820 ;
        RECT 655.125 1593.635 655.415 1593.680 ;
        RECT 664.310 1593.620 664.630 1593.680 ;
        RECT 617.390 1587.700 617.710 1587.760 ;
        RECT 655.125 1587.700 655.415 1587.745 ;
        RECT 617.390 1587.560 655.415 1587.700 ;
        RECT 617.390 1587.500 617.710 1587.560 ;
        RECT 655.125 1587.515 655.415 1587.560 ;
      LAYER via ;
        RECT 664.340 1593.620 664.600 1593.880 ;
        RECT 617.420 1587.500 617.680 1587.760 ;
      LAYER met2 ;
        RECT 664.410 1600.380 664.690 1604.000 ;
        RECT 664.400 1600.000 664.690 1600.380 ;
        RECT 664.400 1593.910 664.540 1600.000 ;
        RECT 664.340 1593.590 664.600 1593.910 ;
        RECT 617.420 1587.470 617.680 1587.790 ;
        RECT 617.480 20.245 617.620 1587.470 ;
        RECT 222.730 19.875 223.010 20.245 ;
        RECT 617.410 19.875 617.690 20.245 ;
        RECT 222.800 2.400 222.940 19.875 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 222.730 19.920 223.010 20.200 ;
        RECT 617.410 19.920 617.690 20.200 ;
      LAYER met3 ;
        RECT 222.705 20.210 223.035 20.225 ;
        RECT 617.385 20.210 617.715 20.225 ;
        RECT 222.705 19.910 617.715 20.210 ;
        RECT 222.705 19.895 223.035 19.910 ;
        RECT 617.385 19.895 617.715 19.910 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 15.200 20.630 15.260 ;
        RECT 331.730 15.200 332.050 15.260 ;
        RECT 20.310 15.060 332.050 15.200 ;
        RECT 20.310 15.000 20.630 15.060 ;
        RECT 331.730 15.000 332.050 15.060 ;
      LAYER via ;
        RECT 20.340 15.000 20.600 15.260 ;
        RECT 331.760 15.000 332.020 15.260 ;
      LAYER met2 ;
        RECT 333.670 1600.450 333.950 1604.000 ;
        RECT 331.820 1600.310 333.950 1600.450 ;
        RECT 331.820 15.290 331.960 1600.310 ;
        RECT 333.670 1600.000 333.950 1600.310 ;
        RECT 20.340 14.970 20.600 15.290 ;
        RECT 331.760 14.970 332.020 15.290 ;
        RECT 20.400 2.400 20.540 14.970 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.670 16.560 372.990 16.620 ;
        RECT 365.400 16.420 372.990 16.560 ;
        RECT 44.230 16.220 44.550 16.280 ;
        RECT 365.400 16.220 365.540 16.420 ;
        RECT 372.670 16.360 372.990 16.420 ;
        RECT 44.230 16.080 365.540 16.220 ;
        RECT 44.230 16.020 44.550 16.080 ;
      LAYER via ;
        RECT 44.260 16.020 44.520 16.280 ;
        RECT 372.700 16.360 372.960 16.620 ;
      LAYER met2 ;
        RECT 372.770 1600.380 373.050 1604.000 ;
        RECT 372.760 1600.000 373.050 1600.380 ;
        RECT 372.760 16.650 372.900 1600.000 ;
        RECT 372.700 16.330 372.960 16.650 ;
        RECT 44.260 15.990 44.520 16.310 ;
        RECT 44.320 2.400 44.460 15.990 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 246.630 30.840 246.950 30.900 ;
        RECT 696.970 30.840 697.290 30.900 ;
        RECT 246.630 30.700 697.290 30.840 ;
        RECT 246.630 30.640 246.950 30.700 ;
        RECT 696.970 30.640 697.290 30.700 ;
      LAYER via ;
        RECT 246.660 30.640 246.920 30.900 ;
        RECT 697.000 30.640 697.260 30.900 ;
      LAYER met2 ;
        RECT 703.510 1600.450 703.790 1604.000 ;
        RECT 697.060 1600.310 703.790 1600.450 ;
        RECT 697.060 30.930 697.200 1600.310 ;
        RECT 703.510 1600.000 703.790 1600.310 ;
        RECT 246.660 30.610 246.920 30.930 ;
        RECT 697.000 30.610 697.260 30.930 ;
        RECT 246.720 2.400 246.860 30.610 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 268.710 1588.720 269.030 1588.780 ;
        RECT 732.850 1588.720 733.170 1588.780 ;
        RECT 268.710 1588.580 733.170 1588.720 ;
        RECT 268.710 1588.520 269.030 1588.580 ;
        RECT 732.850 1588.520 733.170 1588.580 ;
      LAYER via ;
        RECT 268.740 1588.520 269.000 1588.780 ;
        RECT 732.880 1588.520 733.140 1588.780 ;
      LAYER met2 ;
        RECT 732.950 1600.380 733.230 1604.000 ;
        RECT 732.940 1600.000 733.230 1600.380 ;
        RECT 732.940 1588.810 733.080 1600.000 ;
        RECT 268.740 1588.490 269.000 1588.810 ;
        RECT 732.880 1588.490 733.140 1588.810 ;
        RECT 268.800 17.410 268.940 1588.490 ;
        RECT 264.200 17.270 268.940 17.410 ;
        RECT 264.200 2.400 264.340 17.270 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 761.930 1600.450 762.210 1604.000 ;
        RECT 759.160 1600.310 762.210 1600.450 ;
        RECT 759.160 17.525 759.300 1600.310 ;
        RECT 761.930 1600.000 762.210 1600.310 ;
        RECT 282.070 17.155 282.350 17.525 ;
        RECT 759.090 17.155 759.370 17.525 ;
        RECT 282.140 2.400 282.280 17.155 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 282.070 17.200 282.350 17.480 ;
        RECT 759.090 17.200 759.370 17.480 ;
      LAYER met3 ;
        RECT 282.045 17.490 282.375 17.505 ;
        RECT 759.065 17.490 759.395 17.505 ;
        RECT 282.045 17.190 759.395 17.490 ;
        RECT 282.045 17.175 282.375 17.190 ;
        RECT 759.065 17.175 759.395 17.190 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 624.290 1587.360 624.610 1587.420 ;
        RECT 790.810 1587.360 791.130 1587.420 ;
        RECT 624.290 1587.220 791.130 1587.360 ;
        RECT 624.290 1587.160 624.610 1587.220 ;
        RECT 790.810 1587.160 791.130 1587.220 ;
        RECT 299.990 24.380 300.310 24.440 ;
        RECT 624.290 24.380 624.610 24.440 ;
        RECT 299.990 24.240 624.610 24.380 ;
        RECT 299.990 24.180 300.310 24.240 ;
        RECT 624.290 24.180 624.610 24.240 ;
      LAYER via ;
        RECT 624.320 1587.160 624.580 1587.420 ;
        RECT 790.840 1587.160 791.100 1587.420 ;
        RECT 300.020 24.180 300.280 24.440 ;
        RECT 624.320 24.180 624.580 24.440 ;
      LAYER met2 ;
        RECT 790.910 1600.380 791.190 1604.000 ;
        RECT 790.900 1600.000 791.190 1600.380 ;
        RECT 790.900 1587.450 791.040 1600.000 ;
        RECT 624.320 1587.130 624.580 1587.450 ;
        RECT 790.840 1587.130 791.100 1587.450 ;
        RECT 624.380 24.470 624.520 1587.130 ;
        RECT 300.020 24.150 300.280 24.470 ;
        RECT 624.320 24.150 624.580 24.470 ;
        RECT 300.080 2.400 300.220 24.150 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 14.180 318.250 14.240 ;
        RECT 814.270 14.180 814.590 14.240 ;
        RECT 317.930 14.040 814.590 14.180 ;
        RECT 317.930 13.980 318.250 14.040 ;
        RECT 814.270 13.980 814.590 14.040 ;
      LAYER via ;
        RECT 317.960 13.980 318.220 14.240 ;
        RECT 814.300 13.980 814.560 14.240 ;
      LAYER met2 ;
        RECT 820.350 1600.450 820.630 1604.000 ;
        RECT 814.360 1600.310 820.630 1600.450 ;
        RECT 814.360 14.270 814.500 1600.310 ;
        RECT 820.350 1600.000 820.630 1600.310 ;
        RECT 317.960 13.950 318.220 14.270 ;
        RECT 814.300 13.950 814.560 14.270 ;
        RECT 318.020 2.400 318.160 13.950 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 658.790 1587.700 659.110 1587.760 ;
        RECT 849.230 1587.700 849.550 1587.760 ;
        RECT 658.790 1587.560 849.550 1587.700 ;
        RECT 658.790 1587.500 659.110 1587.560 ;
        RECT 849.230 1587.500 849.550 1587.560 ;
        RECT 335.870 24.720 336.190 24.780 ;
        RECT 658.790 24.720 659.110 24.780 ;
        RECT 335.870 24.580 659.110 24.720 ;
        RECT 335.870 24.520 336.190 24.580 ;
        RECT 658.790 24.520 659.110 24.580 ;
      LAYER via ;
        RECT 658.820 1587.500 659.080 1587.760 ;
        RECT 849.260 1587.500 849.520 1587.760 ;
        RECT 335.900 24.520 336.160 24.780 ;
        RECT 658.820 24.520 659.080 24.780 ;
      LAYER met2 ;
        RECT 849.330 1600.380 849.610 1604.000 ;
        RECT 849.320 1600.000 849.610 1600.380 ;
        RECT 849.320 1587.790 849.460 1600.000 ;
        RECT 658.820 1587.470 659.080 1587.790 ;
        RECT 849.260 1587.470 849.520 1587.790 ;
        RECT 658.880 24.810 659.020 1587.470 ;
        RECT 335.900 24.490 336.160 24.810 ;
        RECT 658.820 24.490 659.080 24.810 ;
        RECT 335.960 2.400 336.100 24.490 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 353.350 15.200 353.670 15.260 ;
        RECT 876.370 15.200 876.690 15.260 ;
        RECT 353.350 15.060 876.690 15.200 ;
        RECT 353.350 15.000 353.670 15.060 ;
        RECT 876.370 15.000 876.690 15.060 ;
      LAYER via ;
        RECT 353.380 15.000 353.640 15.260 ;
        RECT 876.400 15.000 876.660 15.260 ;
      LAYER met2 ;
        RECT 878.770 1600.450 879.050 1604.000 ;
        RECT 876.460 1600.310 879.050 1600.450 ;
        RECT 876.460 15.290 876.600 1600.310 ;
        RECT 878.770 1600.000 879.050 1600.310 ;
        RECT 353.380 14.970 353.640 15.290 ;
        RECT 876.400 14.970 876.660 15.290 ;
        RECT 353.440 2.400 353.580 14.970 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 371.290 2.960 371.610 3.020 ;
        RECT 372.210 2.960 372.530 3.020 ;
        RECT 371.290 2.820 372.530 2.960 ;
        RECT 371.290 2.760 371.610 2.820 ;
        RECT 372.210 2.760 372.530 2.820 ;
      LAYER via ;
        RECT 371.320 2.760 371.580 3.020 ;
        RECT 372.240 2.760 372.500 3.020 ;
      LAYER met2 ;
        RECT 907.750 1600.380 908.030 1604.000 ;
        RECT 907.740 1600.000 908.030 1600.380 ;
        RECT 907.740 1592.405 907.880 1600.000 ;
        RECT 372.230 1592.035 372.510 1592.405 ;
        RECT 907.670 1592.035 907.950 1592.405 ;
        RECT 372.300 3.050 372.440 1592.035 ;
        RECT 371.320 2.730 371.580 3.050 ;
        RECT 372.240 2.730 372.500 3.050 ;
        RECT 371.380 2.400 371.520 2.730 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 372.230 1592.080 372.510 1592.360 ;
        RECT 907.670 1592.080 907.950 1592.360 ;
      LAYER met3 ;
        RECT 372.205 1592.370 372.535 1592.385 ;
        RECT 907.645 1592.370 907.975 1592.385 ;
        RECT 372.205 1592.070 907.975 1592.370 ;
        RECT 372.205 1592.055 372.535 1592.070 ;
        RECT 907.645 1592.055 907.975 1592.070 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 389.230 15.880 389.550 15.940 ;
        RECT 931.570 15.880 931.890 15.940 ;
        RECT 389.230 15.740 931.890 15.880 ;
        RECT 389.230 15.680 389.550 15.740 ;
        RECT 931.570 15.680 931.890 15.740 ;
      LAYER via ;
        RECT 389.260 15.680 389.520 15.940 ;
        RECT 931.600 15.680 931.860 15.940 ;
      LAYER met2 ;
        RECT 937.190 1600.450 937.470 1604.000 ;
        RECT 931.660 1600.310 937.470 1600.450 ;
        RECT 931.660 15.970 931.800 1600.310 ;
        RECT 937.190 1600.000 937.470 1600.310 ;
        RECT 389.260 15.650 389.520 15.970 ;
        RECT 931.600 15.650 931.860 15.970 ;
        RECT 389.320 2.400 389.460 15.650 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 407.170 20.300 407.490 20.360 ;
        RECT 413.150 20.300 413.470 20.360 ;
        RECT 407.170 20.160 413.470 20.300 ;
        RECT 407.170 20.100 407.490 20.160 ;
        RECT 413.150 20.100 413.470 20.160 ;
      LAYER via ;
        RECT 407.200 20.100 407.460 20.360 ;
        RECT 413.180 20.100 413.440 20.360 ;
      LAYER met2 ;
        RECT 966.170 1600.380 966.450 1604.000 ;
        RECT 966.160 1600.000 966.450 1600.380 ;
        RECT 966.160 1591.725 966.300 1600.000 ;
        RECT 413.170 1591.355 413.450 1591.725 ;
        RECT 966.090 1591.355 966.370 1591.725 ;
        RECT 413.240 20.390 413.380 1591.355 ;
        RECT 407.200 20.070 407.460 20.390 ;
        RECT 413.180 20.070 413.440 20.390 ;
        RECT 407.260 2.400 407.400 20.070 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 413.170 1591.400 413.450 1591.680 ;
        RECT 966.090 1591.400 966.370 1591.680 ;
      LAYER met3 ;
        RECT 413.145 1591.690 413.475 1591.705 ;
        RECT 966.065 1591.690 966.395 1591.705 ;
        RECT 413.145 1591.390 966.395 1591.690 ;
        RECT 413.145 1591.375 413.475 1591.390 ;
        RECT 966.065 1591.375 966.395 1591.390 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 82.945 19.805 83.115 20.655 ;
        RECT 276.145 20.485 276.315 22.695 ;
        RECT 323.985 20.485 324.155 22.695 ;
      LAYER mcon ;
        RECT 276.145 22.525 276.315 22.695 ;
        RECT 82.945 20.485 83.115 20.655 ;
        RECT 323.985 22.525 324.155 22.695 ;
      LAYER met1 ;
        RECT 276.085 22.680 276.375 22.725 ;
        RECT 323.925 22.680 324.215 22.725 ;
        RECT 276.085 22.540 324.215 22.680 ;
        RECT 276.085 22.495 276.375 22.540 ;
        RECT 323.925 22.495 324.215 22.540 ;
        RECT 82.885 20.640 83.175 20.685 ;
        RECT 276.085 20.640 276.375 20.685 ;
        RECT 82.885 20.500 276.375 20.640 ;
        RECT 82.885 20.455 83.175 20.500 ;
        RECT 276.085 20.455 276.375 20.500 ;
        RECT 323.925 20.640 324.215 20.685 ;
        RECT 406.710 20.640 407.030 20.700 ;
        RECT 323.925 20.500 407.030 20.640 ;
        RECT 323.925 20.455 324.215 20.500 ;
        RECT 406.710 20.440 407.030 20.500 ;
        RECT 68.150 19.960 68.470 20.020 ;
        RECT 82.885 19.960 83.175 20.005 ;
        RECT 68.150 19.820 83.175 19.960 ;
        RECT 68.150 19.760 68.470 19.820 ;
        RECT 82.885 19.775 83.175 19.820 ;
      LAYER via ;
        RECT 406.740 20.440 407.000 20.700 ;
        RECT 68.180 19.760 68.440 20.020 ;
      LAYER met2 ;
        RECT 411.410 1600.450 411.690 1604.000 ;
        RECT 407.260 1600.310 411.690 1600.450 ;
        RECT 407.260 20.810 407.400 1600.310 ;
        RECT 411.410 1600.000 411.690 1600.310 ;
        RECT 406.800 20.730 407.400 20.810 ;
        RECT 406.740 20.670 407.400 20.730 ;
        RECT 406.740 20.410 407.000 20.670 ;
        RECT 68.180 19.730 68.440 20.050 ;
        RECT 68.240 2.400 68.380 19.730 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 456.465 16.065 456.635 19.635 ;
      LAYER mcon ;
        RECT 456.465 19.465 456.635 19.635 ;
      LAYER met1 ;
        RECT 424.650 19.620 424.970 19.680 ;
        RECT 456.405 19.620 456.695 19.665 ;
        RECT 424.650 19.480 456.695 19.620 ;
        RECT 424.650 19.420 424.970 19.480 ;
        RECT 456.405 19.435 456.695 19.480 ;
        RECT 456.405 16.220 456.695 16.265 ;
        RECT 993.670 16.220 993.990 16.280 ;
        RECT 456.405 16.080 993.990 16.220 ;
        RECT 456.405 16.035 456.695 16.080 ;
        RECT 993.670 16.020 993.990 16.080 ;
      LAYER via ;
        RECT 424.680 19.420 424.940 19.680 ;
        RECT 993.700 16.020 993.960 16.280 ;
      LAYER met2 ;
        RECT 995.610 1600.450 995.890 1604.000 ;
        RECT 993.760 1600.310 995.890 1600.450 ;
        RECT 424.680 19.390 424.940 19.710 ;
        RECT 424.740 2.400 424.880 19.390 ;
        RECT 993.760 16.310 993.900 1600.310 ;
        RECT 995.610 1600.000 995.890 1600.310 ;
        RECT 993.700 15.990 993.960 16.310 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1021.270 16.900 1021.590 16.960 ;
        RECT 455.560 16.760 1021.590 16.900 ;
        RECT 442.590 16.560 442.910 16.620 ;
        RECT 455.560 16.560 455.700 16.760 ;
        RECT 1021.270 16.700 1021.590 16.760 ;
        RECT 442.590 16.420 455.700 16.560 ;
        RECT 442.590 16.360 442.910 16.420 ;
      LAYER via ;
        RECT 442.620 16.360 442.880 16.620 ;
        RECT 1021.300 16.700 1021.560 16.960 ;
      LAYER met2 ;
        RECT 1024.590 1600.450 1024.870 1604.000 ;
        RECT 1021.360 1600.310 1024.870 1600.450 ;
        RECT 1021.360 16.990 1021.500 1600.310 ;
        RECT 1024.590 1600.000 1024.870 1600.310 ;
        RECT 1021.300 16.670 1021.560 16.990 ;
        RECT 442.620 16.330 442.880 16.650 ;
        RECT 442.680 2.400 442.820 16.330 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 1593.480 462.230 1593.540 ;
        RECT 1053.930 1593.480 1054.250 1593.540 ;
        RECT 461.910 1593.340 1054.250 1593.480 ;
        RECT 461.910 1593.280 462.230 1593.340 ;
        RECT 1053.930 1593.280 1054.250 1593.340 ;
      LAYER via ;
        RECT 461.940 1593.280 462.200 1593.540 ;
        RECT 1053.960 1593.280 1054.220 1593.540 ;
      LAYER met2 ;
        RECT 1054.030 1600.380 1054.310 1604.000 ;
        RECT 1054.020 1600.000 1054.310 1600.380 ;
        RECT 1054.020 1593.570 1054.160 1600.000 ;
        RECT 461.940 1593.250 462.200 1593.570 ;
        RECT 1053.960 1593.250 1054.220 1593.570 ;
        RECT 462.000 16.730 462.140 1593.250 ;
        RECT 460.620 16.590 462.140 16.730 ;
        RECT 460.620 2.400 460.760 16.590 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 488.665 1592.985 490.675 1593.155 ;
      LAYER mcon ;
        RECT 490.505 1592.985 490.675 1593.155 ;
      LAYER met1 ;
        RECT 482.610 1593.140 482.930 1593.200 ;
        RECT 488.605 1593.140 488.895 1593.185 ;
        RECT 482.610 1593.000 488.895 1593.140 ;
        RECT 482.610 1592.940 482.930 1593.000 ;
        RECT 488.605 1592.955 488.895 1593.000 ;
        RECT 490.445 1593.140 490.735 1593.185 ;
        RECT 1082.910 1593.140 1083.230 1593.200 ;
        RECT 490.445 1593.000 1083.230 1593.140 ;
        RECT 490.445 1592.955 490.735 1593.000 ;
        RECT 1082.910 1592.940 1083.230 1593.000 ;
        RECT 478.470 18.600 478.790 18.660 ;
        RECT 482.610 18.600 482.930 18.660 ;
        RECT 478.470 18.460 482.930 18.600 ;
        RECT 478.470 18.400 478.790 18.460 ;
        RECT 482.610 18.400 482.930 18.460 ;
      LAYER via ;
        RECT 482.640 1592.940 482.900 1593.200 ;
        RECT 1082.940 1592.940 1083.200 1593.200 ;
        RECT 478.500 18.400 478.760 18.660 ;
        RECT 482.640 18.400 482.900 18.660 ;
      LAYER met2 ;
        RECT 1083.010 1600.380 1083.290 1604.000 ;
        RECT 1083.000 1600.000 1083.290 1600.380 ;
        RECT 1083.000 1593.230 1083.140 1600.000 ;
        RECT 482.640 1592.910 482.900 1593.230 ;
        RECT 1082.940 1592.910 1083.200 1593.230 ;
        RECT 482.700 18.690 482.840 1592.910 ;
        RECT 478.500 18.370 478.760 18.690 ;
        RECT 482.640 18.370 482.900 18.690 ;
        RECT 478.560 2.400 478.700 18.370 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.410 19.960 496.730 20.020 ;
        RECT 1110.970 19.960 1111.290 20.020 ;
        RECT 496.410 19.820 1111.290 19.960 ;
        RECT 496.410 19.760 496.730 19.820 ;
        RECT 1110.970 19.760 1111.290 19.820 ;
      LAYER via ;
        RECT 496.440 19.760 496.700 20.020 ;
        RECT 1111.000 19.760 1111.260 20.020 ;
      LAYER met2 ;
        RECT 1112.450 1600.450 1112.730 1604.000 ;
        RECT 1111.060 1600.310 1112.730 1600.450 ;
        RECT 1111.060 20.050 1111.200 1600.310 ;
        RECT 1112.450 1600.000 1112.730 1600.310 ;
        RECT 496.440 19.730 496.700 20.050 ;
        RECT 1111.000 19.730 1111.260 20.050 ;
        RECT 496.500 2.400 496.640 19.730 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 513.890 19.620 514.210 19.680 ;
        RECT 1138.570 19.620 1138.890 19.680 ;
        RECT 513.890 19.480 1138.890 19.620 ;
        RECT 513.890 19.420 514.210 19.480 ;
        RECT 1138.570 19.420 1138.890 19.480 ;
      LAYER via ;
        RECT 513.920 19.420 514.180 19.680 ;
        RECT 1138.600 19.420 1138.860 19.680 ;
      LAYER met2 ;
        RECT 1141.430 1600.450 1141.710 1604.000 ;
        RECT 1138.660 1600.310 1141.710 1600.450 ;
        RECT 1138.660 19.710 1138.800 1600.310 ;
        RECT 1141.430 1600.000 1141.710 1600.310 ;
        RECT 513.920 19.390 514.180 19.710 ;
        RECT 1138.600 19.390 1138.860 19.710 ;
        RECT 513.980 2.400 514.120 19.390 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 538.270 1592.460 538.590 1592.520 ;
        RECT 1170.770 1592.460 1171.090 1592.520 ;
        RECT 538.270 1592.320 1171.090 1592.460 ;
        RECT 538.270 1592.260 538.590 1592.320 ;
        RECT 1170.770 1592.260 1171.090 1592.320 ;
        RECT 531.830 17.920 532.150 17.980 ;
        RECT 537.810 17.920 538.130 17.980 ;
        RECT 531.830 17.780 538.130 17.920 ;
        RECT 531.830 17.720 532.150 17.780 ;
        RECT 537.810 17.720 538.130 17.780 ;
      LAYER via ;
        RECT 538.300 1592.260 538.560 1592.520 ;
        RECT 1170.800 1592.260 1171.060 1592.520 ;
        RECT 531.860 17.720 532.120 17.980 ;
        RECT 537.840 17.720 538.100 17.980 ;
      LAYER met2 ;
        RECT 1170.870 1600.380 1171.150 1604.000 ;
        RECT 1170.860 1600.000 1171.150 1600.380 ;
        RECT 1170.860 1592.550 1171.000 1600.000 ;
        RECT 538.300 1592.230 538.560 1592.550 ;
        RECT 1170.800 1592.230 1171.060 1592.550 ;
        RECT 538.360 1591.610 538.500 1592.230 ;
        RECT 537.900 1591.470 538.500 1591.610 ;
        RECT 537.900 18.010 538.040 1591.470 ;
        RECT 531.860 17.690 532.120 18.010 ;
        RECT 537.840 17.690 538.100 18.010 ;
        RECT 531.920 2.400 532.060 17.690 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 1592.120 551.930 1592.180 ;
        RECT 1199.750 1592.120 1200.070 1592.180 ;
        RECT 551.610 1591.980 1200.070 1592.120 ;
        RECT 551.610 1591.920 551.930 1591.980 ;
        RECT 1199.750 1591.920 1200.070 1591.980 ;
      LAYER via ;
        RECT 551.640 1591.920 551.900 1592.180 ;
        RECT 1199.780 1591.920 1200.040 1592.180 ;
      LAYER met2 ;
        RECT 1199.850 1600.380 1200.130 1604.000 ;
        RECT 1199.840 1600.000 1200.130 1600.380 ;
        RECT 1199.840 1592.210 1199.980 1600.000 ;
        RECT 551.640 1591.890 551.900 1592.210 ;
        RECT 1199.780 1591.890 1200.040 1592.210 ;
        RECT 551.700 16.730 551.840 1591.890 ;
        RECT 549.860 16.590 551.840 16.730 ;
        RECT 549.860 2.400 550.000 16.590 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 567.710 18.600 568.030 18.660 ;
        RECT 1228.270 18.600 1228.590 18.660 ;
        RECT 567.710 18.460 1228.590 18.600 ;
        RECT 567.710 18.400 568.030 18.460 ;
        RECT 1228.270 18.400 1228.590 18.460 ;
      LAYER via ;
        RECT 567.740 18.400 568.000 18.660 ;
        RECT 1228.300 18.400 1228.560 18.660 ;
      LAYER met2 ;
        RECT 1229.290 1600.450 1229.570 1604.000 ;
        RECT 1228.360 1600.310 1229.570 1600.450 ;
        RECT 1228.360 18.690 1228.500 1600.310 ;
        RECT 1229.290 1600.000 1229.570 1600.310 ;
        RECT 567.740 18.370 568.000 18.690 ;
        RECT 1228.300 18.370 1228.560 18.690 ;
        RECT 567.800 2.400 567.940 18.370 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 585.650 18.260 585.970 18.320 ;
        RECT 1255.870 18.260 1256.190 18.320 ;
        RECT 585.650 18.120 1256.190 18.260 ;
        RECT 585.650 18.060 585.970 18.120 ;
        RECT 1255.870 18.060 1256.190 18.120 ;
      LAYER via ;
        RECT 585.680 18.060 585.940 18.320 ;
        RECT 1255.900 18.060 1256.160 18.320 ;
      LAYER met2 ;
        RECT 1258.270 1600.450 1258.550 1604.000 ;
        RECT 1255.960 1600.310 1258.550 1600.450 ;
        RECT 1255.960 18.350 1256.100 1600.310 ;
        RECT 1258.270 1600.000 1258.550 1600.310 ;
        RECT 585.680 18.030 585.940 18.350 ;
        RECT 1255.900 18.030 1256.160 18.350 ;
        RECT 585.740 2.400 585.880 18.030 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 424.265 19.465 424.435 20.655 ;
      LAYER mcon ;
        RECT 424.265 20.485 424.435 20.655 ;
      LAYER met1 ;
        RECT 424.205 20.640 424.495 20.685 ;
        RECT 448.570 20.640 448.890 20.700 ;
        RECT 424.205 20.500 448.890 20.640 ;
        RECT 424.205 20.455 424.495 20.500 ;
        RECT 448.570 20.440 448.890 20.500 ;
        RECT 91.610 19.620 91.930 19.680 ;
        RECT 424.205 19.620 424.495 19.665 ;
        RECT 91.610 19.480 424.495 19.620 ;
        RECT 91.610 19.420 91.930 19.480 ;
        RECT 424.205 19.435 424.495 19.480 ;
      LAYER via ;
        RECT 448.600 20.440 448.860 20.700 ;
        RECT 91.640 19.420 91.900 19.680 ;
      LAYER met2 ;
        RECT 450.510 1600.450 450.790 1604.000 ;
        RECT 448.660 1600.310 450.790 1600.450 ;
        RECT 448.660 20.730 448.800 1600.310 ;
        RECT 450.510 1600.000 450.790 1600.310 ;
        RECT 448.600 20.410 448.860 20.730 ;
        RECT 91.640 19.390 91.900 19.710 ;
        RECT 91.700 2.400 91.840 19.390 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 603.130 17.580 603.450 17.640 ;
        RECT 1283.470 17.580 1283.790 17.640 ;
        RECT 603.130 17.440 1283.790 17.580 ;
        RECT 603.130 17.380 603.450 17.440 ;
        RECT 1283.470 17.380 1283.790 17.440 ;
      LAYER via ;
        RECT 603.160 17.380 603.420 17.640 ;
        RECT 1283.500 17.380 1283.760 17.640 ;
      LAYER met2 ;
        RECT 1287.710 1600.450 1287.990 1604.000 ;
        RECT 1283.560 1600.310 1287.990 1600.450 ;
        RECT 1283.560 17.670 1283.700 1600.310 ;
        RECT 1287.710 1600.000 1287.990 1600.310 ;
        RECT 603.160 17.350 603.420 17.670 ;
        RECT 1283.500 17.350 1283.760 17.670 ;
        RECT 603.220 2.400 603.360 17.350 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 621.070 17.240 621.390 17.300 ;
        RECT 1311.070 17.240 1311.390 17.300 ;
        RECT 621.070 17.100 1311.390 17.240 ;
        RECT 621.070 17.040 621.390 17.100 ;
        RECT 1311.070 17.040 1311.390 17.100 ;
      LAYER via ;
        RECT 621.100 17.040 621.360 17.300 ;
        RECT 1311.100 17.040 1311.360 17.300 ;
      LAYER met2 ;
        RECT 1316.690 1600.450 1316.970 1604.000 ;
        RECT 1311.160 1600.310 1316.970 1600.450 ;
        RECT 1311.160 17.330 1311.300 1600.310 ;
        RECT 1316.690 1600.000 1316.970 1600.310 ;
        RECT 621.100 17.010 621.360 17.330 ;
        RECT 1311.100 17.010 1311.360 17.330 ;
        RECT 621.160 2.400 621.300 17.010 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 116.910 1592.800 117.230 1592.860 ;
        RECT 489.510 1592.800 489.830 1592.860 ;
        RECT 116.910 1592.660 489.830 1592.800 ;
        RECT 116.910 1592.600 117.230 1592.660 ;
        RECT 489.510 1592.600 489.830 1592.660 ;
      LAYER via ;
        RECT 116.940 1592.600 117.200 1592.860 ;
        RECT 489.540 1592.600 489.800 1592.860 ;
      LAYER met2 ;
        RECT 489.610 1600.380 489.890 1604.000 ;
        RECT 489.600 1600.000 489.890 1600.380 ;
        RECT 489.600 1592.890 489.740 1600.000 ;
        RECT 116.940 1592.570 117.200 1592.890 ;
        RECT 489.540 1592.570 489.800 1592.890 ;
        RECT 117.000 24.210 117.140 1592.570 ;
        RECT 115.620 24.070 117.140 24.210 ;
        RECT 115.620 2.400 115.760 24.070 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 144.510 1592.120 144.830 1592.180 ;
        RECT 528.150 1592.120 528.470 1592.180 ;
        RECT 144.510 1591.980 528.470 1592.120 ;
        RECT 144.510 1591.920 144.830 1591.980 ;
        RECT 528.150 1591.920 528.470 1591.980 ;
        RECT 139.450 17.580 139.770 17.640 ;
        RECT 144.510 17.580 144.830 17.640 ;
        RECT 139.450 17.440 144.830 17.580 ;
        RECT 139.450 17.380 139.770 17.440 ;
        RECT 144.510 17.380 144.830 17.440 ;
      LAYER via ;
        RECT 144.540 1591.920 144.800 1592.180 ;
        RECT 528.180 1591.920 528.440 1592.180 ;
        RECT 139.480 17.380 139.740 17.640 ;
        RECT 144.540 17.380 144.800 17.640 ;
      LAYER met2 ;
        RECT 528.250 1600.380 528.530 1604.000 ;
        RECT 528.240 1600.000 528.530 1600.380 ;
        RECT 528.240 1592.210 528.380 1600.000 ;
        RECT 144.540 1591.890 144.800 1592.210 ;
        RECT 528.180 1591.890 528.440 1592.210 ;
        RECT 144.600 17.670 144.740 1591.890 ;
        RECT 139.480 17.350 139.740 17.670 ;
        RECT 144.540 17.350 144.800 17.670 ;
        RECT 139.540 2.400 139.680 17.350 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 1591.780 158.630 1591.840 ;
        RECT 557.590 1591.780 557.910 1591.840 ;
        RECT 158.310 1591.640 557.910 1591.780 ;
        RECT 158.310 1591.580 158.630 1591.640 ;
        RECT 557.590 1591.580 557.910 1591.640 ;
      LAYER via ;
        RECT 158.340 1591.580 158.600 1591.840 ;
        RECT 557.620 1591.580 557.880 1591.840 ;
      LAYER met2 ;
        RECT 557.690 1600.380 557.970 1604.000 ;
        RECT 557.680 1600.000 557.970 1600.380 ;
        RECT 557.680 1591.870 557.820 1600.000 ;
        RECT 158.340 1591.550 158.600 1591.870 ;
        RECT 557.620 1591.550 557.880 1591.870 ;
        RECT 158.400 17.410 158.540 1591.550 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 179.010 1591.100 179.330 1591.160 ;
        RECT 586.570 1591.100 586.890 1591.160 ;
        RECT 179.010 1590.960 586.890 1591.100 ;
        RECT 179.010 1590.900 179.330 1590.960 ;
        RECT 586.570 1590.900 586.890 1590.960 ;
        RECT 174.870 17.920 175.190 17.980 ;
        RECT 179.010 17.920 179.330 17.980 ;
        RECT 174.870 17.780 179.330 17.920 ;
        RECT 174.870 17.720 175.190 17.780 ;
        RECT 179.010 17.720 179.330 17.780 ;
      LAYER via ;
        RECT 179.040 1590.900 179.300 1591.160 ;
        RECT 586.600 1590.900 586.860 1591.160 ;
        RECT 174.900 17.720 175.160 17.980 ;
        RECT 179.040 17.720 179.300 17.980 ;
      LAYER met2 ;
        RECT 586.670 1600.380 586.950 1604.000 ;
        RECT 586.660 1600.000 586.950 1600.380 ;
        RECT 586.660 1591.190 586.800 1600.000 ;
        RECT 179.040 1590.870 179.300 1591.190 ;
        RECT 586.600 1590.870 586.860 1591.190 ;
        RECT 179.100 18.010 179.240 1590.870 ;
        RECT 174.900 17.690 175.160 18.010 ;
        RECT 179.040 17.690 179.300 18.010 ;
        RECT 174.960 2.400 175.100 17.690 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.350 1587.700 192.670 1587.760 ;
        RECT 616.010 1587.700 616.330 1587.760 ;
        RECT 192.350 1587.560 616.330 1587.700 ;
        RECT 192.350 1587.500 192.670 1587.560 ;
        RECT 616.010 1587.500 616.330 1587.560 ;
      LAYER via ;
        RECT 192.380 1587.500 192.640 1587.760 ;
        RECT 616.040 1587.500 616.300 1587.760 ;
      LAYER met2 ;
        RECT 616.110 1600.380 616.390 1604.000 ;
        RECT 616.100 1600.000 616.390 1600.380 ;
        RECT 616.100 1587.790 616.240 1600.000 ;
        RECT 192.380 1587.470 192.640 1587.790 ;
        RECT 616.040 1587.470 616.300 1587.790 ;
        RECT 192.440 24.210 192.580 1587.470 ;
        RECT 192.440 24.070 193.040 24.210 ;
        RECT 192.900 2.400 193.040 24.070 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 213.510 1591.440 213.830 1591.500 ;
        RECT 644.990 1591.440 645.310 1591.500 ;
        RECT 213.510 1591.300 645.310 1591.440 ;
        RECT 213.510 1591.240 213.830 1591.300 ;
        RECT 644.990 1591.240 645.310 1591.300 ;
      LAYER via ;
        RECT 213.540 1591.240 213.800 1591.500 ;
        RECT 645.020 1591.240 645.280 1591.500 ;
      LAYER met2 ;
        RECT 645.090 1600.380 645.370 1604.000 ;
        RECT 645.080 1600.000 645.370 1600.380 ;
        RECT 645.080 1591.530 645.220 1600.000 ;
        RECT 213.540 1591.210 213.800 1591.530 ;
        RECT 645.020 1591.210 645.280 1591.530 ;
        RECT 213.600 24.210 213.740 1591.210 ;
        RECT 210.840 24.070 213.740 24.210 ;
        RECT 210.840 2.400 210.980 24.070 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 674.530 1600.450 674.810 1604.000 ;
        RECT 669.460 1600.310 674.810 1600.450 ;
        RECT 669.460 18.885 669.600 1600.310 ;
        RECT 674.530 1600.000 674.810 1600.310 ;
        RECT 228.710 18.515 228.990 18.885 ;
        RECT 669.390 18.515 669.670 18.885 ;
        RECT 228.780 2.400 228.920 18.515 ;
        RECT 228.570 -4.800 229.130 2.400 ;
      LAYER via2 ;
        RECT 228.710 18.560 228.990 18.840 ;
        RECT 669.390 18.560 669.670 18.840 ;
      LAYER met3 ;
        RECT 228.685 18.850 229.015 18.865 ;
        RECT 669.365 18.850 669.695 18.865 ;
        RECT 228.685 18.550 669.695 18.850 ;
        RECT 228.685 18.535 229.015 18.550 ;
        RECT 669.365 18.535 669.695 18.550 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 348.365 15.725 348.535 16.575 ;
      LAYER mcon ;
        RECT 348.365 16.405 348.535 16.575 ;
      LAYER met1 ;
        RECT 50.210 16.560 50.530 16.620 ;
        RECT 348.305 16.560 348.595 16.605 ;
        RECT 50.210 16.420 348.595 16.560 ;
        RECT 50.210 16.360 50.530 16.420 ;
        RECT 348.305 16.375 348.595 16.420 ;
        RECT 348.305 15.880 348.595 15.925 ;
        RECT 380.030 15.880 380.350 15.940 ;
        RECT 348.305 15.740 380.350 15.880 ;
        RECT 348.305 15.695 348.595 15.740 ;
        RECT 380.030 15.680 380.350 15.740 ;
      LAYER via ;
        RECT 50.240 16.360 50.500 16.620 ;
        RECT 380.060 15.680 380.320 15.940 ;
      LAYER met2 ;
        RECT 382.430 1600.450 382.710 1604.000 ;
        RECT 380.120 1600.310 382.710 1600.450 ;
        RECT 50.240 16.330 50.500 16.650 ;
        RECT 50.300 2.400 50.440 16.330 ;
        RECT 380.120 15.970 380.260 1600.310 ;
        RECT 382.430 1600.000 382.710 1600.310 ;
        RECT 380.060 15.650 380.320 15.970 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 1588.380 255.230 1588.440 ;
        RECT 713.070 1588.380 713.390 1588.440 ;
        RECT 254.910 1588.240 713.390 1588.380 ;
        RECT 254.910 1588.180 255.230 1588.240 ;
        RECT 713.070 1588.180 713.390 1588.240 ;
      LAYER via ;
        RECT 254.940 1588.180 255.200 1588.440 ;
        RECT 713.100 1588.180 713.360 1588.440 ;
      LAYER met2 ;
        RECT 713.170 1600.380 713.450 1604.000 ;
        RECT 713.160 1600.000 713.450 1600.380 ;
        RECT 713.160 1588.470 713.300 1600.000 ;
        RECT 254.940 1588.150 255.200 1588.470 ;
        RECT 713.100 1588.150 713.360 1588.470 ;
        RECT 255.000 17.410 255.140 1588.150 ;
        RECT 252.700 17.270 255.140 17.410 ;
        RECT 252.700 2.400 252.840 17.270 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 742.610 1600.450 742.890 1604.000 ;
        RECT 738.460 1600.310 742.890 1600.450 ;
        RECT 738.460 18.205 738.600 1600.310 ;
        RECT 742.610 1600.000 742.890 1600.310 ;
        RECT 270.110 17.835 270.390 18.205 ;
        RECT 738.390 17.835 738.670 18.205 ;
        RECT 270.180 2.400 270.320 17.835 ;
        RECT 269.970 -4.800 270.530 2.400 ;
      LAYER via2 ;
        RECT 270.110 17.880 270.390 18.160 ;
        RECT 738.390 17.880 738.670 18.160 ;
      LAYER met3 ;
        RECT 270.085 18.170 270.415 18.185 ;
        RECT 738.365 18.170 738.695 18.185 ;
        RECT 270.085 17.870 738.695 18.170 ;
        RECT 270.085 17.855 270.415 17.870 ;
        RECT 738.365 17.855 738.695 17.870 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 1589.060 289.730 1589.120 ;
        RECT 771.490 1589.060 771.810 1589.120 ;
        RECT 289.410 1588.920 771.810 1589.060 ;
        RECT 289.410 1588.860 289.730 1588.920 ;
        RECT 771.490 1588.860 771.810 1588.920 ;
      LAYER via ;
        RECT 289.440 1588.860 289.700 1589.120 ;
        RECT 771.520 1588.860 771.780 1589.120 ;
      LAYER met2 ;
        RECT 771.590 1600.380 771.870 1604.000 ;
        RECT 771.580 1600.000 771.870 1600.380 ;
        RECT 771.580 1589.150 771.720 1600.000 ;
        RECT 289.440 1588.830 289.700 1589.150 ;
        RECT 771.520 1588.830 771.780 1589.150 ;
        RECT 289.500 3.130 289.640 1588.830 ;
        RECT 288.120 2.990 289.640 3.130 ;
        RECT 288.120 2.400 288.260 2.990 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 14.520 306.290 14.580 ;
        RECT 800.470 14.520 800.790 14.580 ;
        RECT 305.970 14.380 800.790 14.520 ;
        RECT 305.970 14.320 306.290 14.380 ;
        RECT 800.470 14.320 800.790 14.380 ;
      LAYER via ;
        RECT 306.000 14.320 306.260 14.580 ;
        RECT 800.500 14.320 800.760 14.580 ;
      LAYER met2 ;
        RECT 801.030 1600.450 801.310 1604.000 ;
        RECT 800.560 1600.310 801.310 1600.450 ;
        RECT 800.560 14.610 800.700 1600.310 ;
        RECT 801.030 1600.000 801.310 1600.310 ;
        RECT 306.000 14.290 306.260 14.610 ;
        RECT 800.500 14.290 800.760 14.610 ;
        RECT 306.060 2.400 306.200 14.290 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 830.010 1600.380 830.290 1604.000 ;
        RECT 830.000 1600.000 830.290 1600.380 ;
        RECT 830.000 1593.085 830.140 1600.000 ;
        RECT 323.930 1592.715 324.210 1593.085 ;
        RECT 829.930 1592.715 830.210 1593.085 ;
        RECT 324.000 2.400 324.140 1592.715 ;
        RECT 323.790 -4.800 324.350 2.400 ;
      LAYER via2 ;
        RECT 323.930 1592.760 324.210 1593.040 ;
        RECT 829.930 1592.760 830.210 1593.040 ;
      LAYER met3 ;
        RECT 323.905 1593.050 324.235 1593.065 ;
        RECT 829.905 1593.050 830.235 1593.065 ;
        RECT 323.905 1592.750 830.235 1593.050 ;
        RECT 323.905 1592.735 324.235 1592.750 ;
        RECT 829.905 1592.735 830.235 1592.750 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 14.860 341.710 14.920 ;
        RECT 855.670 14.860 855.990 14.920 ;
        RECT 341.390 14.720 855.990 14.860 ;
        RECT 341.390 14.660 341.710 14.720 ;
        RECT 855.670 14.660 855.990 14.720 ;
      LAYER via ;
        RECT 341.420 14.660 341.680 14.920 ;
        RECT 855.700 14.660 855.960 14.920 ;
      LAYER met2 ;
        RECT 859.450 1600.450 859.730 1604.000 ;
        RECT 855.760 1600.310 859.730 1600.450 ;
        RECT 855.760 14.950 855.900 1600.310 ;
        RECT 859.450 1600.000 859.730 1600.310 ;
        RECT 341.420 14.630 341.680 14.950 ;
        RECT 855.700 14.630 855.960 14.950 ;
        RECT 341.480 2.400 341.620 14.630 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 1589.400 365.170 1589.460 ;
        RECT 888.330 1589.400 888.650 1589.460 ;
        RECT 364.850 1589.260 888.650 1589.400 ;
        RECT 364.850 1589.200 365.170 1589.260 ;
        RECT 888.330 1589.200 888.650 1589.260 ;
        RECT 359.330 16.560 359.650 16.620 ;
        RECT 364.850 16.560 365.170 16.620 ;
        RECT 359.330 16.420 365.170 16.560 ;
        RECT 359.330 16.360 359.650 16.420 ;
        RECT 364.850 16.360 365.170 16.420 ;
      LAYER via ;
        RECT 364.880 1589.200 365.140 1589.460 ;
        RECT 888.360 1589.200 888.620 1589.460 ;
        RECT 359.360 16.360 359.620 16.620 ;
        RECT 364.880 16.360 365.140 16.620 ;
      LAYER met2 ;
        RECT 888.430 1600.380 888.710 1604.000 ;
        RECT 888.420 1600.000 888.710 1600.380 ;
        RECT 888.420 1589.490 888.560 1600.000 ;
        RECT 364.880 1589.170 365.140 1589.490 ;
        RECT 888.360 1589.170 888.620 1589.490 ;
        RECT 364.940 16.650 365.080 1589.170 ;
        RECT 359.360 16.330 359.620 16.650 ;
        RECT 364.880 16.330 365.140 16.650 ;
        RECT 359.420 2.400 359.560 16.330 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 377.270 15.540 377.590 15.600 ;
        RECT 917.770 15.540 918.090 15.600 ;
        RECT 377.270 15.400 918.090 15.540 ;
        RECT 377.270 15.340 377.590 15.400 ;
        RECT 917.770 15.340 918.090 15.400 ;
      LAYER via ;
        RECT 377.300 15.340 377.560 15.600 ;
        RECT 917.800 15.340 918.060 15.600 ;
      LAYER met2 ;
        RECT 917.870 1600.380 918.150 1604.000 ;
        RECT 917.860 1600.000 918.150 1600.380 ;
        RECT 917.860 15.630 918.000 1600.000 ;
        RECT 377.300 15.310 377.560 15.630 ;
        RECT 917.800 15.310 918.060 15.630 ;
        RECT 377.360 2.400 377.500 15.310 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 399.810 1589.740 400.130 1589.800 ;
        RECT 946.750 1589.740 947.070 1589.800 ;
        RECT 399.810 1589.600 947.070 1589.740 ;
        RECT 399.810 1589.540 400.130 1589.600 ;
        RECT 946.750 1589.540 947.070 1589.600 ;
        RECT 395.210 16.900 395.530 16.960 ;
        RECT 399.810 16.900 400.130 16.960 ;
        RECT 395.210 16.760 400.130 16.900 ;
        RECT 395.210 16.700 395.530 16.760 ;
        RECT 399.810 16.700 400.130 16.760 ;
      LAYER via ;
        RECT 399.840 1589.540 400.100 1589.800 ;
        RECT 946.780 1589.540 947.040 1589.800 ;
        RECT 395.240 16.700 395.500 16.960 ;
        RECT 399.840 16.700 400.100 16.960 ;
      LAYER met2 ;
        RECT 946.850 1600.380 947.130 1604.000 ;
        RECT 946.840 1600.000 947.130 1600.380 ;
        RECT 946.840 1589.830 946.980 1600.000 ;
        RECT 399.840 1589.510 400.100 1589.830 ;
        RECT 946.780 1589.510 947.040 1589.830 ;
        RECT 399.900 16.990 400.040 1589.510 ;
        RECT 395.240 16.670 395.500 16.990 ;
        RECT 399.840 16.670 400.100 16.990 ;
        RECT 395.300 2.400 395.440 16.670 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 975.830 1600.380 976.110 1604.000 ;
        RECT 975.820 1600.000 976.110 1600.380 ;
        RECT 975.820 1591.045 975.960 1600.000 ;
        RECT 413.630 1590.675 413.910 1591.045 ;
        RECT 975.750 1590.675 976.030 1591.045 ;
        RECT 413.700 17.410 413.840 1590.675 ;
        RECT 413.240 17.270 413.840 17.410 ;
        RECT 413.240 2.400 413.380 17.270 ;
        RECT 413.030 -4.800 413.590 2.400 ;
      LAYER via2 ;
        RECT 413.630 1590.720 413.910 1591.000 ;
        RECT 975.750 1590.720 976.030 1591.000 ;
      LAYER met3 ;
        RECT 413.605 1591.010 413.935 1591.025 ;
        RECT 975.725 1591.010 976.055 1591.025 ;
        RECT 413.605 1590.710 976.055 1591.010 ;
        RECT 413.605 1590.695 413.935 1590.710 ;
        RECT 975.725 1590.695 976.055 1590.710 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 400.345 16.745 400.515 20.315 ;
      LAYER mcon ;
        RECT 400.345 20.145 400.515 20.315 ;
      LAYER met1 ;
        RECT 74.130 20.300 74.450 20.360 ;
        RECT 276.530 20.300 276.850 20.360 ;
        RECT 74.130 20.160 276.850 20.300 ;
        RECT 74.130 20.100 74.450 20.160 ;
        RECT 276.530 20.100 276.850 20.160 ;
        RECT 323.450 20.300 323.770 20.360 ;
        RECT 400.285 20.300 400.575 20.345 ;
        RECT 323.450 20.160 400.575 20.300 ;
        RECT 323.450 20.100 323.770 20.160 ;
        RECT 400.285 20.115 400.575 20.160 ;
        RECT 400.285 16.900 400.575 16.945 ;
        RECT 420.970 16.900 421.290 16.960 ;
        RECT 400.285 16.760 421.290 16.900 ;
        RECT 400.285 16.715 400.575 16.760 ;
        RECT 420.970 16.700 421.290 16.760 ;
      LAYER via ;
        RECT 74.160 20.100 74.420 20.360 ;
        RECT 276.560 20.100 276.820 20.360 ;
        RECT 323.480 20.100 323.740 20.360 ;
        RECT 421.000 16.700 421.260 16.960 ;
      LAYER met2 ;
        RECT 421.070 1600.380 421.350 1604.000 ;
        RECT 421.060 1600.000 421.350 1600.380 ;
        RECT 276.550 20.555 276.830 20.925 ;
        RECT 323.470 20.555 323.750 20.925 ;
        RECT 276.620 20.390 276.760 20.555 ;
        RECT 323.540 20.390 323.680 20.555 ;
        RECT 74.160 20.070 74.420 20.390 ;
        RECT 276.560 20.070 276.820 20.390 ;
        RECT 323.480 20.070 323.740 20.390 ;
        RECT 74.220 2.400 74.360 20.070 ;
        RECT 421.060 16.990 421.200 1600.000 ;
        RECT 421.000 16.670 421.260 16.990 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 276.550 20.600 276.830 20.880 ;
        RECT 323.470 20.600 323.750 20.880 ;
      LAYER met3 ;
        RECT 276.525 20.890 276.855 20.905 ;
        RECT 323.445 20.890 323.775 20.905 ;
        RECT 276.525 20.590 323.775 20.890 ;
        RECT 276.525 20.575 276.855 20.590 ;
        RECT 323.445 20.575 323.775 20.590 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1000.570 16.560 1000.890 16.620 ;
        RECT 456.020 16.420 1000.890 16.560 ;
        RECT 430.630 16.220 430.950 16.280 ;
        RECT 456.020 16.220 456.160 16.420 ;
        RECT 1000.570 16.360 1000.890 16.420 ;
        RECT 430.630 16.080 456.160 16.220 ;
        RECT 430.630 16.020 430.950 16.080 ;
      LAYER via ;
        RECT 430.660 16.020 430.920 16.280 ;
        RECT 1000.600 16.360 1000.860 16.620 ;
      LAYER met2 ;
        RECT 1005.270 1600.450 1005.550 1604.000 ;
        RECT 1000.660 1600.310 1005.550 1600.450 ;
        RECT 1000.660 16.650 1000.800 1600.310 ;
        RECT 1005.270 1600.000 1005.550 1600.310 ;
        RECT 1000.600 16.330 1000.860 16.650 ;
        RECT 430.660 15.990 430.920 16.310 ;
        RECT 430.720 2.400 430.860 15.990 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 454.550 1590.080 454.870 1590.140 ;
        RECT 1034.150 1590.080 1034.470 1590.140 ;
        RECT 454.550 1589.940 1034.470 1590.080 ;
        RECT 454.550 1589.880 454.870 1589.940 ;
        RECT 1034.150 1589.880 1034.470 1589.940 ;
        RECT 448.570 16.900 448.890 16.960 ;
        RECT 454.550 16.900 454.870 16.960 ;
        RECT 448.570 16.760 454.870 16.900 ;
        RECT 448.570 16.700 448.890 16.760 ;
        RECT 454.550 16.700 454.870 16.760 ;
      LAYER via ;
        RECT 454.580 1589.880 454.840 1590.140 ;
        RECT 1034.180 1589.880 1034.440 1590.140 ;
        RECT 448.600 16.700 448.860 16.960 ;
        RECT 454.580 16.700 454.840 16.960 ;
      LAYER met2 ;
        RECT 1034.250 1600.380 1034.530 1604.000 ;
        RECT 1034.240 1600.000 1034.530 1600.380 ;
        RECT 1034.240 1590.170 1034.380 1600.000 ;
        RECT 454.580 1589.850 454.840 1590.170 ;
        RECT 1034.180 1589.850 1034.440 1590.170 ;
        RECT 454.640 16.990 454.780 1589.850 ;
        RECT 448.600 16.670 448.860 16.990 ;
        RECT 454.580 16.670 454.840 16.990 ;
        RECT 448.660 2.400 448.800 16.670 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 466.510 20.640 466.830 20.700 ;
        RECT 1062.670 20.640 1062.990 20.700 ;
        RECT 466.510 20.500 1062.990 20.640 ;
        RECT 466.510 20.440 466.830 20.500 ;
        RECT 1062.670 20.440 1062.990 20.500 ;
      LAYER via ;
        RECT 466.540 20.440 466.800 20.700 ;
        RECT 1062.700 20.440 1062.960 20.700 ;
      LAYER met2 ;
        RECT 1063.690 1600.450 1063.970 1604.000 ;
        RECT 1062.760 1600.310 1063.970 1600.450 ;
        RECT 1062.760 20.730 1062.900 1600.310 ;
        RECT 1063.690 1600.000 1063.970 1600.310 ;
        RECT 466.540 20.410 466.800 20.730 ;
        RECT 1062.700 20.410 1062.960 20.730 ;
        RECT 466.600 2.400 466.740 20.410 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 489.970 1592.800 490.290 1592.860 ;
        RECT 1092.570 1592.800 1092.890 1592.860 ;
        RECT 489.970 1592.660 1092.890 1592.800 ;
        RECT 489.970 1592.600 490.290 1592.660 ;
        RECT 1092.570 1592.600 1092.890 1592.660 ;
        RECT 484.450 18.600 484.770 18.660 ;
        RECT 489.510 18.600 489.830 18.660 ;
        RECT 484.450 18.460 489.830 18.600 ;
        RECT 484.450 18.400 484.770 18.460 ;
        RECT 489.510 18.400 489.830 18.460 ;
      LAYER via ;
        RECT 490.000 1592.600 490.260 1592.860 ;
        RECT 1092.600 1592.600 1092.860 1592.860 ;
        RECT 484.480 18.400 484.740 18.660 ;
        RECT 489.540 18.400 489.800 18.660 ;
      LAYER met2 ;
        RECT 1092.670 1600.380 1092.950 1604.000 ;
        RECT 1092.660 1600.000 1092.950 1600.380 ;
        RECT 1092.660 1592.890 1092.800 1600.000 ;
        RECT 490.000 1592.570 490.260 1592.890 ;
        RECT 1092.600 1592.570 1092.860 1592.890 ;
        RECT 490.060 1592.290 490.200 1592.570 ;
        RECT 489.600 1592.150 490.200 1592.290 ;
        RECT 489.600 18.690 489.740 1592.150 ;
        RECT 484.480 18.370 484.740 18.690 ;
        RECT 489.540 18.370 489.800 18.690 ;
        RECT 484.540 2.400 484.680 18.370 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 541.565 19.125 541.735 20.315 ;
      LAYER mcon ;
        RECT 541.565 20.145 541.735 20.315 ;
      LAYER met1 ;
        RECT 541.505 20.300 541.795 20.345 ;
        RECT 1117.870 20.300 1118.190 20.360 ;
        RECT 541.505 20.160 1118.190 20.300 ;
        RECT 541.505 20.115 541.795 20.160 ;
        RECT 1117.870 20.100 1118.190 20.160 ;
        RECT 502.390 19.280 502.710 19.340 ;
        RECT 541.505 19.280 541.795 19.325 ;
        RECT 502.390 19.140 541.795 19.280 ;
        RECT 502.390 19.080 502.710 19.140 ;
        RECT 541.505 19.095 541.795 19.140 ;
      LAYER via ;
        RECT 1117.900 20.100 1118.160 20.360 ;
        RECT 502.420 19.080 502.680 19.340 ;
      LAYER met2 ;
        RECT 1122.110 1600.450 1122.390 1604.000 ;
        RECT 1117.960 1600.310 1122.390 1600.450 ;
        RECT 1117.960 20.390 1118.100 1600.310 ;
        RECT 1122.110 1600.000 1122.390 1600.310 ;
        RECT 1117.900 20.070 1118.160 20.390 ;
        RECT 502.420 19.050 502.680 19.370 ;
        RECT 502.480 2.400 502.620 19.050 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 17.920 520.190 17.980 ;
        RECT 524.010 17.920 524.330 17.980 ;
        RECT 519.870 17.780 524.330 17.920 ;
        RECT 519.870 17.720 520.190 17.780 ;
        RECT 524.010 17.720 524.330 17.780 ;
      LAYER via ;
        RECT 519.900 17.720 520.160 17.980 ;
        RECT 524.040 17.720 524.300 17.980 ;
      LAYER met2 ;
        RECT 1151.090 1600.380 1151.370 1604.000 ;
        RECT 1151.080 1600.000 1151.370 1600.380 ;
        RECT 1151.080 1590.365 1151.220 1600.000 ;
        RECT 524.030 1589.995 524.310 1590.365 ;
        RECT 1151.010 1589.995 1151.290 1590.365 ;
        RECT 524.100 18.010 524.240 1589.995 ;
        RECT 519.900 17.690 520.160 18.010 ;
        RECT 524.040 17.690 524.300 18.010 ;
        RECT 519.960 2.400 520.100 17.690 ;
        RECT 519.750 -4.800 520.310 2.400 ;
      LAYER via2 ;
        RECT 524.030 1590.040 524.310 1590.320 ;
        RECT 1151.010 1590.040 1151.290 1590.320 ;
      LAYER met3 ;
        RECT 524.005 1590.330 524.335 1590.345 ;
        RECT 1150.985 1590.330 1151.315 1590.345 ;
        RECT 524.005 1590.030 1151.315 1590.330 ;
        RECT 524.005 1590.015 524.335 1590.030 ;
        RECT 1150.985 1590.015 1151.315 1590.030 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1179.970 19.280 1180.290 19.340 ;
        RECT 549.400 19.140 1180.290 19.280 ;
        RECT 537.350 18.940 537.670 19.000 ;
        RECT 549.400 18.940 549.540 19.140 ;
        RECT 1179.970 19.080 1180.290 19.140 ;
        RECT 537.350 18.800 549.540 18.940 ;
        RECT 537.350 18.740 537.670 18.800 ;
      LAYER via ;
        RECT 537.380 18.740 537.640 19.000 ;
        RECT 1180.000 19.080 1180.260 19.340 ;
      LAYER met2 ;
        RECT 1180.530 1600.450 1180.810 1604.000 ;
        RECT 1180.060 1600.310 1180.810 1600.450 ;
        RECT 1180.060 19.370 1180.200 1600.310 ;
        RECT 1180.530 1600.000 1180.810 1600.310 ;
        RECT 1180.000 19.050 1180.260 19.370 ;
        RECT 537.380 18.710 537.640 19.030 ;
        RECT 537.440 9.930 537.580 18.710 ;
        RECT 537.440 9.790 538.040 9.930 ;
        RECT 537.900 2.400 538.040 9.790 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 558.510 1591.780 558.830 1591.840 ;
        RECT 1209.410 1591.780 1209.730 1591.840 ;
        RECT 558.510 1591.640 1209.730 1591.780 ;
        RECT 558.510 1591.580 558.830 1591.640 ;
        RECT 1209.410 1591.580 1209.730 1591.640 ;
        RECT 555.750 17.920 556.070 17.980 ;
        RECT 558.510 17.920 558.830 17.980 ;
        RECT 555.750 17.780 558.830 17.920 ;
        RECT 555.750 17.720 556.070 17.780 ;
        RECT 558.510 17.720 558.830 17.780 ;
      LAYER via ;
        RECT 558.540 1591.580 558.800 1591.840 ;
        RECT 1209.440 1591.580 1209.700 1591.840 ;
        RECT 555.780 17.720 556.040 17.980 ;
        RECT 558.540 17.720 558.800 17.980 ;
      LAYER met2 ;
        RECT 1209.510 1600.380 1209.790 1604.000 ;
        RECT 1209.500 1600.000 1209.790 1600.380 ;
        RECT 1209.500 1591.870 1209.640 1600.000 ;
        RECT 558.540 1591.550 558.800 1591.870 ;
        RECT 1209.440 1591.550 1209.700 1591.870 ;
        RECT 558.600 18.010 558.740 1591.550 ;
        RECT 555.780 17.690 556.040 18.010 ;
        RECT 558.540 17.690 558.800 18.010 ;
        RECT 555.840 2.400 555.980 17.690 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 573.690 18.940 574.010 19.000 ;
        RECT 1235.170 18.940 1235.490 19.000 ;
        RECT 573.690 18.800 1235.490 18.940 ;
        RECT 573.690 18.740 574.010 18.800 ;
        RECT 1235.170 18.740 1235.490 18.800 ;
      LAYER via ;
        RECT 573.720 18.740 573.980 19.000 ;
        RECT 1235.200 18.740 1235.460 19.000 ;
      LAYER met2 ;
        RECT 1238.950 1600.450 1239.230 1604.000 ;
        RECT 1235.260 1600.310 1239.230 1600.450 ;
        RECT 1235.260 19.030 1235.400 1600.310 ;
        RECT 1238.950 1600.000 1239.230 1600.310 ;
        RECT 573.720 18.710 573.980 19.030 ;
        RECT 1235.200 18.710 1235.460 19.030 ;
        RECT 573.780 2.400 573.920 18.710 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 593.010 1591.100 593.330 1591.160 ;
        RECT 1267.830 1591.100 1268.150 1591.160 ;
        RECT 593.010 1590.960 1268.150 1591.100 ;
        RECT 593.010 1590.900 593.330 1590.960 ;
        RECT 1267.830 1590.900 1268.150 1590.960 ;
      LAYER via ;
        RECT 593.040 1590.900 593.300 1591.160 ;
        RECT 1267.860 1590.900 1268.120 1591.160 ;
      LAYER met2 ;
        RECT 1267.930 1600.380 1268.210 1604.000 ;
        RECT 1267.920 1600.000 1268.210 1600.380 ;
        RECT 1267.920 1591.190 1268.060 1600.000 ;
        RECT 593.040 1590.870 593.300 1591.190 ;
        RECT 1267.860 1590.870 1268.120 1591.190 ;
        RECT 593.100 16.730 593.240 1590.870 ;
        RECT 591.260 16.590 593.240 16.730 ;
        RECT 591.260 2.400 591.400 16.590 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 103.110 1593.480 103.430 1593.540 ;
        RECT 460.070 1593.480 460.390 1593.540 ;
        RECT 103.110 1593.340 460.390 1593.480 ;
        RECT 103.110 1593.280 103.430 1593.340 ;
        RECT 460.070 1593.280 460.390 1593.340 ;
        RECT 97.590 19.280 97.910 19.340 ;
        RECT 103.110 19.280 103.430 19.340 ;
        RECT 97.590 19.140 103.430 19.280 ;
        RECT 97.590 19.080 97.910 19.140 ;
        RECT 103.110 19.080 103.430 19.140 ;
      LAYER via ;
        RECT 103.140 1593.280 103.400 1593.540 ;
        RECT 460.100 1593.280 460.360 1593.540 ;
        RECT 97.620 19.080 97.880 19.340 ;
        RECT 103.140 19.080 103.400 19.340 ;
      LAYER met2 ;
        RECT 460.170 1600.380 460.450 1604.000 ;
        RECT 460.160 1600.000 460.450 1600.380 ;
        RECT 460.160 1593.570 460.300 1600.000 ;
        RECT 103.140 1593.250 103.400 1593.570 ;
        RECT 460.100 1593.250 460.360 1593.570 ;
        RECT 103.200 19.370 103.340 1593.250 ;
        RECT 97.620 19.050 97.880 19.370 ;
        RECT 103.140 19.050 103.400 19.370 ;
        RECT 97.680 2.400 97.820 19.050 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1297.370 1600.380 1297.650 1604.000 ;
        RECT 1297.360 1600.000 1297.650 1600.380 ;
        RECT 1297.360 16.845 1297.500 1600.000 ;
        RECT 609.130 16.475 609.410 16.845 ;
        RECT 1297.290 16.475 1297.570 16.845 ;
        RECT 609.200 2.400 609.340 16.475 ;
        RECT 608.990 -4.800 609.550 2.400 ;
      LAYER via2 ;
        RECT 609.130 16.520 609.410 16.800 ;
        RECT 1297.290 16.520 1297.570 16.800 ;
      LAYER met3 ;
        RECT 609.105 16.810 609.435 16.825 ;
        RECT 1297.265 16.810 1297.595 16.825 ;
        RECT 609.105 16.510 1297.595 16.810 ;
        RECT 609.105 16.495 609.435 16.510 ;
        RECT 1297.265 16.495 1297.595 16.510 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.510 1590.760 627.830 1590.820 ;
        RECT 1326.250 1590.760 1326.570 1590.820 ;
        RECT 627.510 1590.620 1326.570 1590.760 ;
        RECT 627.510 1590.560 627.830 1590.620 ;
        RECT 1326.250 1590.560 1326.570 1590.620 ;
      LAYER via ;
        RECT 627.540 1590.560 627.800 1590.820 ;
        RECT 1326.280 1590.560 1326.540 1590.820 ;
      LAYER met2 ;
        RECT 1326.350 1600.380 1326.630 1604.000 ;
        RECT 1326.340 1600.000 1326.630 1600.380 ;
        RECT 1326.340 1590.850 1326.480 1600.000 ;
        RECT 627.540 1590.530 627.800 1590.850 ;
        RECT 1326.280 1590.530 1326.540 1590.850 ;
        RECT 627.600 17.410 627.740 1590.530 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 478.085 18.445 478.255 19.295 ;
      LAYER mcon ;
        RECT 478.085 19.125 478.255 19.295 ;
      LAYER met1 ;
        RECT 478.025 19.280 478.315 19.325 ;
        RECT 496.870 19.280 497.190 19.340 ;
        RECT 478.025 19.140 497.190 19.280 ;
        RECT 478.025 19.095 478.315 19.140 ;
        RECT 496.870 19.080 497.190 19.140 ;
        RECT 121.510 18.600 121.830 18.660 ;
        RECT 478.025 18.600 478.315 18.645 ;
        RECT 121.510 18.460 478.315 18.600 ;
        RECT 121.510 18.400 121.830 18.460 ;
        RECT 478.025 18.415 478.315 18.460 ;
      LAYER via ;
        RECT 496.900 19.080 497.160 19.340 ;
        RECT 121.540 18.400 121.800 18.660 ;
      LAYER met2 ;
        RECT 499.270 1600.450 499.550 1604.000 ;
        RECT 496.960 1600.310 499.550 1600.450 ;
        RECT 496.960 19.370 497.100 1600.310 ;
        RECT 499.270 1600.000 499.550 1600.310 ;
        RECT 496.900 19.050 497.160 19.370 ;
        RECT 121.540 18.370 121.800 18.690 ;
        RECT 121.600 2.400 121.740 18.370 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 151.410 1592.460 151.730 1592.520 ;
        RECT 537.810 1592.460 538.130 1592.520 ;
        RECT 151.410 1592.320 538.130 1592.460 ;
        RECT 151.410 1592.260 151.730 1592.320 ;
        RECT 537.810 1592.260 538.130 1592.320 ;
        RECT 145.430 17.580 145.750 17.640 ;
        RECT 151.410 17.580 151.730 17.640 ;
        RECT 145.430 17.440 151.730 17.580 ;
        RECT 145.430 17.380 145.750 17.440 ;
        RECT 151.410 17.380 151.730 17.440 ;
      LAYER via ;
        RECT 151.440 1592.260 151.700 1592.520 ;
        RECT 537.840 1592.260 538.100 1592.520 ;
        RECT 145.460 17.380 145.720 17.640 ;
        RECT 151.440 17.380 151.700 17.640 ;
      LAYER met2 ;
        RECT 537.910 1600.380 538.190 1604.000 ;
        RECT 537.900 1600.000 538.190 1600.380 ;
        RECT 537.900 1592.550 538.040 1600.000 ;
        RECT 151.440 1592.230 151.700 1592.550 ;
        RECT 537.840 1592.230 538.100 1592.550 ;
        RECT 151.500 17.670 151.640 1592.230 ;
        RECT 145.460 17.350 145.720 17.670 ;
        RECT 151.440 17.350 151.700 17.670 ;
        RECT 145.520 2.400 145.660 17.350 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 165.210 1587.360 165.530 1587.420 ;
        RECT 567.250 1587.360 567.570 1587.420 ;
        RECT 165.210 1587.220 567.570 1587.360 ;
        RECT 165.210 1587.160 165.530 1587.220 ;
        RECT 567.250 1587.160 567.570 1587.220 ;
      LAYER via ;
        RECT 165.240 1587.160 165.500 1587.420 ;
        RECT 567.280 1587.160 567.540 1587.420 ;
      LAYER met2 ;
        RECT 567.350 1600.380 567.630 1604.000 ;
        RECT 567.340 1600.000 567.630 1600.380 ;
        RECT 567.340 1587.450 567.480 1600.000 ;
        RECT 165.240 1587.130 165.500 1587.450 ;
        RECT 567.280 1587.130 567.540 1587.450 ;
        RECT 165.300 17.410 165.440 1587.130 ;
        RECT 163.460 17.270 165.440 17.410 ;
        RECT 163.460 2.400 163.600 17.270 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 17.240 181.170 17.300 ;
        RECT 593.470 17.240 593.790 17.300 ;
        RECT 180.850 17.100 593.790 17.240 ;
        RECT 180.850 17.040 181.170 17.100 ;
        RECT 593.470 17.040 593.790 17.100 ;
      LAYER via ;
        RECT 180.880 17.040 181.140 17.300 ;
        RECT 593.500 17.040 593.760 17.300 ;
      LAYER met2 ;
        RECT 596.330 1600.450 596.610 1604.000 ;
        RECT 593.560 1600.310 596.610 1600.450 ;
        RECT 593.560 17.330 593.700 1600.310 ;
        RECT 596.330 1600.000 596.610 1600.310 ;
        RECT 180.880 17.010 181.140 17.330 ;
        RECT 593.500 17.010 593.760 17.330 ;
        RECT 180.940 2.400 181.080 17.010 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 199.710 1590.760 200.030 1590.820 ;
        RECT 625.670 1590.760 625.990 1590.820 ;
        RECT 199.710 1590.620 625.990 1590.760 ;
        RECT 199.710 1590.560 200.030 1590.620 ;
        RECT 625.670 1590.560 625.990 1590.620 ;
      LAYER via ;
        RECT 199.740 1590.560 200.000 1590.820 ;
        RECT 625.700 1590.560 625.960 1590.820 ;
      LAYER met2 ;
        RECT 625.770 1600.380 626.050 1604.000 ;
        RECT 625.760 1600.000 626.050 1600.380 ;
        RECT 625.760 1590.850 625.900 1600.000 ;
        RECT 199.740 1590.530 200.000 1590.850 ;
        RECT 625.700 1590.530 625.960 1590.850 ;
        RECT 199.800 24.210 199.940 1590.530 ;
        RECT 198.880 24.070 199.940 24.210 ;
        RECT 198.880 2.400 199.020 24.070 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 220.410 1593.820 220.730 1593.880 ;
        RECT 654.650 1593.820 654.970 1593.880 ;
        RECT 220.410 1593.680 654.970 1593.820 ;
        RECT 220.410 1593.620 220.730 1593.680 ;
        RECT 654.650 1593.620 654.970 1593.680 ;
      LAYER via ;
        RECT 220.440 1593.620 220.700 1593.880 ;
        RECT 654.680 1593.620 654.940 1593.880 ;
      LAYER met2 ;
        RECT 654.750 1600.380 655.030 1604.000 ;
        RECT 654.740 1600.000 655.030 1600.380 ;
        RECT 654.740 1593.910 654.880 1600.000 ;
        RECT 220.440 1593.590 220.700 1593.910 ;
        RECT 654.680 1593.590 654.940 1593.910 ;
        RECT 220.500 24.210 220.640 1593.590 ;
        RECT 216.820 24.070 220.640 24.210 ;
        RECT 216.820 2.400 216.960 24.070 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 240.650 1588.040 240.970 1588.100 ;
        RECT 684.090 1588.040 684.410 1588.100 ;
        RECT 240.650 1587.900 684.410 1588.040 ;
        RECT 240.650 1587.840 240.970 1587.900 ;
        RECT 684.090 1587.840 684.410 1587.900 ;
        RECT 234.670 20.980 234.990 21.040 ;
        RECT 240.650 20.980 240.970 21.040 ;
        RECT 234.670 20.840 240.970 20.980 ;
        RECT 234.670 20.780 234.990 20.840 ;
        RECT 240.650 20.780 240.970 20.840 ;
      LAYER via ;
        RECT 240.680 1587.840 240.940 1588.100 ;
        RECT 684.120 1587.840 684.380 1588.100 ;
        RECT 234.700 20.780 234.960 21.040 ;
        RECT 240.680 20.780 240.940 21.040 ;
      LAYER met2 ;
        RECT 684.190 1600.380 684.470 1604.000 ;
        RECT 684.180 1600.000 684.470 1600.380 ;
        RECT 684.180 1588.130 684.320 1600.000 ;
        RECT 240.680 1587.810 240.940 1588.130 ;
        RECT 684.120 1587.810 684.380 1588.130 ;
        RECT 240.740 21.070 240.880 1587.810 ;
        RECT 234.700 20.750 234.960 21.070 ;
        RECT 240.680 20.750 240.940 21.070 ;
        RECT 234.760 2.400 234.900 20.750 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 61.710 1589.740 62.030 1589.800 ;
        RECT 391.990 1589.740 392.310 1589.800 ;
        RECT 61.710 1589.600 392.310 1589.740 ;
        RECT 61.710 1589.540 62.030 1589.600 ;
        RECT 391.990 1589.540 392.310 1589.600 ;
        RECT 56.190 17.580 56.510 17.640 ;
        RECT 61.710 17.580 62.030 17.640 ;
        RECT 56.190 17.440 62.030 17.580 ;
        RECT 56.190 17.380 56.510 17.440 ;
        RECT 61.710 17.380 62.030 17.440 ;
      LAYER via ;
        RECT 61.740 1589.540 62.000 1589.800 ;
        RECT 392.020 1589.540 392.280 1589.800 ;
        RECT 56.220 17.380 56.480 17.640 ;
        RECT 61.740 17.380 62.000 17.640 ;
      LAYER met2 ;
        RECT 392.090 1600.380 392.370 1604.000 ;
        RECT 392.080 1600.000 392.370 1600.380 ;
        RECT 392.080 1589.830 392.220 1600.000 ;
        RECT 61.740 1589.510 62.000 1589.830 ;
        RECT 392.020 1589.510 392.280 1589.830 ;
        RECT 61.800 17.670 61.940 1589.510 ;
        RECT 56.220 17.350 56.480 17.670 ;
        RECT 61.740 17.350 62.000 17.670 ;
        RECT 56.280 2.400 56.420 17.350 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 82.410 1590.080 82.730 1590.140 ;
        RECT 431.090 1590.080 431.410 1590.140 ;
        RECT 82.410 1589.940 431.410 1590.080 ;
        RECT 82.410 1589.880 82.730 1589.940 ;
        RECT 431.090 1589.880 431.410 1589.940 ;
        RECT 80.110 17.580 80.430 17.640 ;
        RECT 82.410 17.580 82.730 17.640 ;
        RECT 80.110 17.440 82.730 17.580 ;
        RECT 80.110 17.380 80.430 17.440 ;
        RECT 82.410 17.380 82.730 17.440 ;
      LAYER via ;
        RECT 82.440 1589.880 82.700 1590.140 ;
        RECT 431.120 1589.880 431.380 1590.140 ;
        RECT 80.140 17.380 80.400 17.640 ;
        RECT 82.440 17.380 82.700 17.640 ;
      LAYER met2 ;
        RECT 431.190 1600.380 431.470 1604.000 ;
        RECT 431.180 1600.000 431.470 1600.380 ;
        RECT 431.180 1590.170 431.320 1600.000 ;
        RECT 82.440 1589.850 82.700 1590.170 ;
        RECT 431.120 1589.850 431.380 1590.170 ;
        RECT 82.500 17.670 82.640 1589.850 ;
        RECT 80.140 17.350 80.400 17.670 ;
        RECT 82.440 17.350 82.700 17.670 ;
        RECT 80.200 2.400 80.340 17.350 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 1593.140 110.330 1593.200 ;
        RECT 469.730 1593.140 470.050 1593.200 ;
        RECT 110.010 1593.000 470.050 1593.140 ;
        RECT 110.010 1592.940 110.330 1593.000 ;
        RECT 469.730 1592.940 470.050 1593.000 ;
        RECT 103.570 19.280 103.890 19.340 ;
        RECT 110.010 19.280 110.330 19.340 ;
        RECT 103.570 19.140 110.330 19.280 ;
        RECT 103.570 19.080 103.890 19.140 ;
        RECT 110.010 19.080 110.330 19.140 ;
      LAYER via ;
        RECT 110.040 1592.940 110.300 1593.200 ;
        RECT 469.760 1592.940 470.020 1593.200 ;
        RECT 103.600 19.080 103.860 19.340 ;
        RECT 110.040 19.080 110.300 19.340 ;
      LAYER met2 ;
        RECT 469.830 1600.380 470.110 1604.000 ;
        RECT 469.820 1600.000 470.110 1600.380 ;
        RECT 469.820 1593.230 469.960 1600.000 ;
        RECT 110.040 1592.910 110.300 1593.230 ;
        RECT 469.760 1592.910 470.020 1593.230 ;
        RECT 110.100 19.370 110.240 1592.910 ;
        RECT 103.600 19.050 103.860 19.370 ;
        RECT 110.040 19.050 110.300 19.370 ;
        RECT 103.660 2.400 103.800 19.050 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 127.490 18.940 127.810 19.000 ;
        RECT 503.770 18.940 504.090 19.000 ;
        RECT 127.490 18.800 504.090 18.940 ;
        RECT 127.490 18.740 127.810 18.800 ;
        RECT 503.770 18.740 504.090 18.800 ;
      LAYER via ;
        RECT 127.520 18.740 127.780 19.000 ;
        RECT 503.800 18.740 504.060 19.000 ;
      LAYER met2 ;
        RECT 508.930 1600.450 509.210 1604.000 ;
        RECT 503.860 1600.310 509.210 1600.450 ;
        RECT 503.860 19.030 504.000 1600.310 ;
        RECT 508.930 1600.000 509.210 1600.310 ;
        RECT 127.520 18.710 127.780 19.030 ;
        RECT 503.800 18.710 504.060 19.030 ;
        RECT 127.580 2.400 127.720 18.710 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 27.210 1589.400 27.530 1589.460 ;
        RECT 343.230 1589.400 343.550 1589.460 ;
        RECT 27.210 1589.260 343.550 1589.400 ;
        RECT 27.210 1589.200 27.530 1589.260 ;
        RECT 343.230 1589.200 343.550 1589.260 ;
        RECT 26.290 2.960 26.610 3.020 ;
        RECT 27.210 2.960 27.530 3.020 ;
        RECT 26.290 2.820 27.530 2.960 ;
        RECT 26.290 2.760 26.610 2.820 ;
        RECT 27.210 2.760 27.530 2.820 ;
      LAYER via ;
        RECT 27.240 1589.200 27.500 1589.460 ;
        RECT 343.260 1589.200 343.520 1589.460 ;
        RECT 26.320 2.760 26.580 3.020 ;
        RECT 27.240 2.760 27.500 3.020 ;
      LAYER met2 ;
        RECT 343.330 1600.380 343.610 1604.000 ;
        RECT 343.320 1600.000 343.610 1600.380 ;
        RECT 343.320 1589.490 343.460 1600.000 ;
        RECT 27.240 1589.170 27.500 1589.490 ;
        RECT 343.260 1589.170 343.520 1589.490 ;
        RECT 27.300 3.050 27.440 1589.170 ;
        RECT 26.320 2.730 26.580 3.050 ;
        RECT 27.240 2.730 27.500 3.050 ;
        RECT 26.380 2.400 26.520 2.730 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 341.465 15.385 342.555 15.555 ;
      LAYER mcon ;
        RECT 342.385 15.385 342.555 15.555 ;
      LAYER met1 ;
        RECT 32.270 15.540 32.590 15.600 ;
        RECT 341.405 15.540 341.695 15.585 ;
        RECT 32.270 15.400 341.695 15.540 ;
        RECT 32.270 15.340 32.590 15.400 ;
        RECT 341.405 15.355 341.695 15.400 ;
        RECT 342.325 15.540 342.615 15.585 ;
        RECT 351.970 15.540 352.290 15.600 ;
        RECT 342.325 15.400 352.290 15.540 ;
        RECT 342.325 15.355 342.615 15.400 ;
        RECT 351.970 15.340 352.290 15.400 ;
      LAYER via ;
        RECT 32.300 15.340 32.560 15.600 ;
        RECT 352.000 15.340 352.260 15.600 ;
      LAYER met2 ;
        RECT 352.990 1600.450 353.270 1604.000 ;
        RECT 352.060 1600.310 353.270 1600.450 ;
        RECT 352.060 15.630 352.200 1600.310 ;
        RECT 352.990 1600.000 353.270 1600.310 ;
        RECT 32.300 15.310 32.560 15.630 ;
        RECT 352.000 15.310 352.260 15.630 ;
        RECT 32.360 2.400 32.500 15.310 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.480 3243.600 684.050 3244.660 ;
        RECT 1331.480 3243.600 1334.050 3244.660 ;
        RECT 1931.480 3243.600 1934.050 3244.660 ;
        RECT 2581.480 3243.600 2584.050 3244.660 ;
        RECT 2631.480 2043.600 2634.050 2044.660 ;
        RECT 1702.430 1611.575 1705.000 1612.635 ;
      LAYER via3 ;
        RECT 682.500 3243.620 684.020 3244.630 ;
        RECT 1332.500 3243.620 1334.020 3244.630 ;
        RECT 1932.500 3243.620 1934.020 3244.630 ;
        RECT 2582.500 3243.620 2584.020 3244.630 ;
        RECT 2632.500 2043.620 2634.020 2044.630 ;
        RECT 1702.460 1611.605 1703.980 1612.615 ;
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 364.020 3271.235 367.020 3529.000 ;
        RECT 382.020 3271.235 385.020 3538.400 ;
        RECT 400.020 3271.235 403.020 3547.800 ;
        RECT 418.020 3271.235 421.020 3557.200 ;
        RECT 544.020 3271.235 547.020 3529.000 ;
        RECT 562.020 3271.235 565.020 3538.400 ;
        RECT 580.020 3271.235 583.020 3547.800 ;
        RECT 598.020 3271.235 601.020 3557.200 ;
        RECT 682.470 2803.670 684.070 3244.680 ;
        RECT 382.020 2715.000 385.020 2785.000 ;
        RECT 400.020 2715.000 403.020 2785.000 ;
        RECT 418.020 2715.000 421.020 2785.000 ;
        RECT 562.020 2715.000 565.020 2785.000 ;
        RECT 580.020 2715.000 583.020 2785.000 ;
        RECT 598.020 2715.000 601.020 2785.000 ;
        RECT 724.020 2715.000 727.020 3529.000 ;
        RECT 742.020 2715.000 745.020 3538.400 ;
        RECT 760.020 2715.000 763.020 3547.800 ;
        RECT 778.020 2715.000 781.020 3557.200 ;
        RECT 904.020 2715.000 907.020 3529.000 ;
        RECT 922.020 2715.000 925.020 3538.400 ;
        RECT 940.020 3271.235 943.020 3547.800 ;
        RECT 958.020 3271.235 961.020 3557.200 ;
        RECT 1084.020 3271.235 1087.020 3529.000 ;
        RECT 1102.020 3271.235 1105.020 3538.400 ;
        RECT 1120.020 3271.235 1123.020 3547.800 ;
        RECT 1138.020 3271.235 1141.020 3557.200 ;
        RECT 1264.020 3271.235 1267.020 3529.000 ;
        RECT 1282.020 3271.235 1285.020 3538.400 ;
        RECT 1300.020 3271.235 1303.020 3547.800 ;
        RECT 1318.020 3271.235 1321.020 3557.200 ;
        RECT 1332.470 2803.670 1334.070 3244.680 ;
        RECT 940.020 2715.000 943.020 2785.000 ;
        RECT 958.020 2715.000 961.020 2785.000 ;
        RECT 1102.020 2715.000 1105.020 2785.000 ;
        RECT 1120.020 2715.000 1123.020 2785.000 ;
        RECT 1138.020 2715.000 1141.020 2785.000 ;
        RECT 1282.020 2715.000 1285.020 2785.000 ;
        RECT 1300.020 2715.000 1303.020 2785.000 ;
        RECT 1318.020 2715.000 1321.020 2785.000 ;
        RECT 321.040 1610.640 322.640 2688.240 ;
        RECT 364.020 -9.320 367.020 1585.000 ;
        RECT 382.020 -18.720 385.020 1585.000 ;
        RECT 400.020 -28.120 403.020 1585.000 ;
        RECT 418.020 -37.520 421.020 1585.000 ;
        RECT 544.020 -9.320 547.020 1585.000 ;
        RECT 562.020 -18.720 565.020 1585.000 ;
        RECT 580.020 -28.120 583.020 1585.000 ;
        RECT 598.020 -37.520 601.020 1585.000 ;
        RECT 724.020 -9.320 727.020 1585.000 ;
        RECT 742.020 -18.720 745.020 1585.000 ;
        RECT 760.020 -28.120 763.020 1585.000 ;
        RECT 778.020 -37.520 781.020 1585.000 ;
        RECT 904.020 -9.320 907.020 1585.000 ;
        RECT 922.020 -18.720 925.020 1585.000 ;
        RECT 940.020 -28.120 943.020 1585.000 ;
        RECT 958.020 -37.520 961.020 1585.000 ;
        RECT 1084.020 -9.320 1087.020 1585.000 ;
        RECT 1102.020 -18.720 1105.020 1585.000 ;
        RECT 1120.020 -28.120 1123.020 1585.000 ;
        RECT 1138.020 -37.520 1141.020 1585.000 ;
        RECT 1264.020 -9.320 1267.020 1585.000 ;
        RECT 1282.020 -18.720 1285.020 1585.000 ;
        RECT 1300.020 -28.120 1303.020 1585.000 ;
        RECT 1318.020 -37.520 1321.020 1585.000 ;
        RECT 1444.020 -9.320 1447.020 3529.000 ;
        RECT 1462.020 -18.720 1465.020 3538.400 ;
        RECT 1480.020 -28.120 1483.020 3547.800 ;
        RECT 1498.020 -37.520 1501.020 3557.200 ;
        RECT 1624.020 3271.235 1627.020 3529.000 ;
        RECT 1642.020 3271.235 1645.020 3538.400 ;
        RECT 1660.020 3271.235 1663.020 3547.800 ;
        RECT 1678.020 3271.235 1681.020 3557.200 ;
        RECT 1804.020 3271.235 1807.020 3529.000 ;
        RECT 1822.020 3271.235 1825.020 3538.400 ;
        RECT 1840.020 3271.235 1843.020 3547.800 ;
        RECT 1858.020 3271.235 1861.020 3557.200 ;
        RECT 1932.470 2803.670 1934.070 3244.680 ;
        RECT 1624.020 1515.000 1627.020 2785.000 ;
        RECT 1642.020 1515.000 1645.020 2785.000 ;
        RECT 1660.020 1515.000 1663.020 2785.000 ;
        RECT 1678.020 1515.000 1681.020 2785.000 ;
        RECT 1804.020 2071.235 1807.020 2785.000 ;
        RECT 1822.020 2071.235 1825.020 2785.000 ;
        RECT 1840.020 2071.235 1843.020 2785.000 ;
        RECT 1858.020 2071.235 1861.020 2785.000 ;
        RECT 1984.020 2071.235 1987.020 3529.000 ;
        RECT 2002.020 2071.235 2005.020 3538.400 ;
        RECT 2020.020 2071.235 2023.020 3547.800 ;
        RECT 2038.020 2071.235 2041.020 3557.200 ;
        RECT 1702.410 1611.555 1704.010 2052.565 ;
        RECT 2164.020 1515.000 2167.020 3529.000 ;
        RECT 2182.020 3271.235 2185.020 3538.400 ;
        RECT 2200.020 3271.235 2203.020 3547.800 ;
        RECT 2218.020 3271.235 2221.020 3557.200 ;
        RECT 2344.020 3271.235 2347.020 3529.000 ;
        RECT 2362.020 3271.235 2365.020 3538.400 ;
        RECT 2380.020 3271.235 2383.020 3547.800 ;
        RECT 2398.020 3271.235 2401.020 3557.200 ;
        RECT 2524.020 3271.235 2527.020 3529.000 ;
        RECT 2542.020 3271.235 2545.020 3538.400 ;
        RECT 2560.020 3271.235 2563.020 3547.800 ;
        RECT 2578.020 3271.235 2581.020 3557.200 ;
        RECT 2582.470 2803.670 2584.070 3244.680 ;
        RECT 2182.020 1515.000 2185.020 2785.000 ;
        RECT 2200.020 1515.000 2203.020 2785.000 ;
        RECT 2218.020 1515.000 2221.020 2785.000 ;
        RECT 2344.020 2071.235 2347.020 2785.000 ;
        RECT 2362.020 2071.235 2365.020 2785.000 ;
        RECT 2380.020 2071.235 2383.020 2785.000 ;
        RECT 2398.020 2071.235 2401.020 2785.000 ;
        RECT 2524.020 2071.235 2527.020 2785.000 ;
        RECT 2542.020 2071.235 2545.020 2785.000 ;
        RECT 2560.020 2071.235 2563.020 2785.000 ;
        RECT 2578.020 2071.235 2581.020 2785.000 ;
        RECT 2632.470 1603.670 2634.070 2044.680 ;
        RECT 1571.040 410.640 1572.640 1488.240 ;
        RECT 1624.020 -9.320 1627.020 385.000 ;
        RECT 1642.020 -18.720 1645.020 385.000 ;
        RECT 1660.020 -28.120 1663.020 385.000 ;
        RECT 1678.020 -37.520 1681.020 385.000 ;
        RECT 1804.020 -9.320 1807.020 385.000 ;
        RECT 1822.020 -18.720 1825.020 385.000 ;
        RECT 1840.020 -28.120 1843.020 385.000 ;
        RECT 1858.020 -37.520 1861.020 385.000 ;
        RECT 1984.020 -9.320 1987.020 385.000 ;
        RECT 2002.020 -18.720 2005.020 385.000 ;
        RECT 2020.020 -28.120 2023.020 385.000 ;
        RECT 2038.020 -37.520 2041.020 385.000 ;
        RECT 2164.020 -9.320 2167.020 385.000 ;
        RECT 2182.020 -18.720 2185.020 385.000 ;
        RECT 2200.020 -28.120 2203.020 385.000 ;
        RECT 2218.020 -37.520 2221.020 385.000 ;
        RECT 2344.020 -9.320 2347.020 385.000 ;
        RECT 2362.020 -18.720 2365.020 385.000 ;
        RECT 2380.020 -28.120 2383.020 385.000 ;
        RECT 2398.020 -37.520 2401.020 385.000 ;
        RECT 2524.020 -9.320 2527.020 385.000 ;
        RECT 2542.020 -18.720 2545.020 385.000 ;
        RECT 2560.020 -28.120 2563.020 385.000 ;
        RECT 2578.020 -37.520 2581.020 385.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 682.680 3125.090 683.860 3126.270 ;
        RECT 682.680 3123.490 683.860 3124.670 ;
        RECT 682.680 3107.090 683.860 3108.270 ;
        RECT 682.680 3105.490 683.860 3106.670 ;
        RECT 682.680 3089.090 683.860 3090.270 ;
        RECT 682.680 3087.490 683.860 3088.670 ;
        RECT 682.680 3071.090 683.860 3072.270 ;
        RECT 682.680 3069.490 683.860 3070.670 ;
        RECT 682.680 2945.090 683.860 2946.270 ;
        RECT 682.680 2943.490 683.860 2944.670 ;
        RECT 682.680 2927.090 683.860 2928.270 ;
        RECT 682.680 2925.490 683.860 2926.670 ;
        RECT 682.680 2909.090 683.860 2910.270 ;
        RECT 682.680 2907.490 683.860 2908.670 ;
        RECT 682.680 2891.090 683.860 2892.270 ;
        RECT 682.680 2889.490 683.860 2890.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 1332.680 3125.090 1333.860 3126.270 ;
        RECT 1332.680 3123.490 1333.860 3124.670 ;
        RECT 1332.680 3107.090 1333.860 3108.270 ;
        RECT 1332.680 3105.490 1333.860 3106.670 ;
        RECT 1332.680 3089.090 1333.860 3090.270 ;
        RECT 1332.680 3087.490 1333.860 3088.670 ;
        RECT 1332.680 3071.090 1333.860 3072.270 ;
        RECT 1332.680 3069.490 1333.860 3070.670 ;
        RECT 1332.680 2945.090 1333.860 2946.270 ;
        RECT 1332.680 2943.490 1333.860 2944.670 ;
        RECT 1332.680 2927.090 1333.860 2928.270 ;
        RECT 1332.680 2925.490 1333.860 2926.670 ;
        RECT 1332.680 2909.090 1333.860 2910.270 ;
        RECT 1332.680 2907.490 1333.860 2908.670 ;
        RECT 1332.680 2891.090 1333.860 2892.270 ;
        RECT 1332.680 2889.490 1333.860 2890.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 321.250 2585.090 322.430 2586.270 ;
        RECT 321.250 2583.490 322.430 2584.670 ;
        RECT 321.250 2567.090 322.430 2568.270 ;
        RECT 321.250 2565.490 322.430 2566.670 ;
        RECT 321.250 2549.090 322.430 2550.270 ;
        RECT 321.250 2547.490 322.430 2548.670 ;
        RECT 321.250 2531.090 322.430 2532.270 ;
        RECT 321.250 2529.490 322.430 2530.670 ;
        RECT 321.250 2405.090 322.430 2406.270 ;
        RECT 321.250 2403.490 322.430 2404.670 ;
        RECT 321.250 2387.090 322.430 2388.270 ;
        RECT 321.250 2385.490 322.430 2386.670 ;
        RECT 321.250 2369.090 322.430 2370.270 ;
        RECT 321.250 2367.490 322.430 2368.670 ;
        RECT 321.250 2351.090 322.430 2352.270 ;
        RECT 321.250 2349.490 322.430 2350.670 ;
        RECT 321.250 2225.090 322.430 2226.270 ;
        RECT 321.250 2223.490 322.430 2224.670 ;
        RECT 321.250 2207.090 322.430 2208.270 ;
        RECT 321.250 2205.490 322.430 2206.670 ;
        RECT 321.250 2189.090 322.430 2190.270 ;
        RECT 321.250 2187.490 322.430 2188.670 ;
        RECT 321.250 2171.090 322.430 2172.270 ;
        RECT 321.250 2169.490 322.430 2170.670 ;
        RECT 321.250 2045.090 322.430 2046.270 ;
        RECT 321.250 2043.490 322.430 2044.670 ;
        RECT 321.250 2027.090 322.430 2028.270 ;
        RECT 321.250 2025.490 322.430 2026.670 ;
        RECT 321.250 2009.090 322.430 2010.270 ;
        RECT 321.250 2007.490 322.430 2008.670 ;
        RECT 321.250 1991.090 322.430 1992.270 ;
        RECT 321.250 1989.490 322.430 1990.670 ;
        RECT 321.250 1865.090 322.430 1866.270 ;
        RECT 321.250 1863.490 322.430 1864.670 ;
        RECT 321.250 1847.090 322.430 1848.270 ;
        RECT 321.250 1845.490 322.430 1846.670 ;
        RECT 321.250 1829.090 322.430 1830.270 ;
        RECT 321.250 1827.490 322.430 1828.670 ;
        RECT 321.250 1811.090 322.430 1812.270 ;
        RECT 321.250 1809.490 322.430 1810.670 ;
        RECT 321.250 1685.090 322.430 1686.270 ;
        RECT 321.250 1683.490 322.430 1684.670 ;
        RECT 321.250 1667.090 322.430 1668.270 ;
        RECT 321.250 1665.490 322.430 1666.670 ;
        RECT 321.250 1649.090 322.430 1650.270 ;
        RECT 321.250 1647.490 322.430 1648.670 ;
        RECT 321.250 1631.090 322.430 1632.270 ;
        RECT 321.250 1629.490 322.430 1630.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1932.680 3125.090 1933.860 3126.270 ;
        RECT 1932.680 3123.490 1933.860 3124.670 ;
        RECT 1932.680 3107.090 1933.860 3108.270 ;
        RECT 1932.680 3105.490 1933.860 3106.670 ;
        RECT 1932.680 3089.090 1933.860 3090.270 ;
        RECT 1932.680 3087.490 1933.860 3088.670 ;
        RECT 1932.680 3071.090 1933.860 3072.270 ;
        RECT 1932.680 3069.490 1933.860 3070.670 ;
        RECT 1932.680 2945.090 1933.860 2946.270 ;
        RECT 1932.680 2943.490 1933.860 2944.670 ;
        RECT 1932.680 2927.090 1933.860 2928.270 ;
        RECT 1932.680 2925.490 1933.860 2926.670 ;
        RECT 1932.680 2909.090 1933.860 2910.270 ;
        RECT 1932.680 2907.490 1933.860 2908.670 ;
        RECT 1932.680 2891.090 1933.860 2892.270 ;
        RECT 1932.680 2889.490 1933.860 2890.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2582.680 3125.090 2583.860 3126.270 ;
        RECT 2582.680 3123.490 2583.860 3124.670 ;
        RECT 2582.680 3107.090 2583.860 3108.270 ;
        RECT 2582.680 3105.490 2583.860 3106.670 ;
        RECT 2582.680 3089.090 2583.860 3090.270 ;
        RECT 2582.680 3087.490 2583.860 3088.670 ;
        RECT 2582.680 3071.090 2583.860 3072.270 ;
        RECT 2582.680 3069.490 2583.860 3070.670 ;
        RECT 2582.680 2945.090 2583.860 2946.270 ;
        RECT 2582.680 2943.490 2583.860 2944.670 ;
        RECT 2582.680 2927.090 2583.860 2928.270 ;
        RECT 2582.680 2925.490 2583.860 2926.670 ;
        RECT 2582.680 2909.090 2583.860 2910.270 ;
        RECT 2582.680 2907.490 2583.860 2908.670 ;
        RECT 2582.680 2891.090 2583.860 2892.270 ;
        RECT 2582.680 2889.490 2583.860 2890.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1702.620 2045.090 1703.800 2046.270 ;
        RECT 1702.620 2043.490 1703.800 2044.670 ;
        RECT 1702.620 2027.090 1703.800 2028.270 ;
        RECT 1702.620 2025.490 1703.800 2026.670 ;
        RECT 1702.620 2009.090 1703.800 2010.270 ;
        RECT 1702.620 2007.490 1703.800 2008.670 ;
        RECT 1702.620 1991.090 1703.800 1992.270 ;
        RECT 1702.620 1989.490 1703.800 1990.670 ;
        RECT 1702.620 1865.090 1703.800 1866.270 ;
        RECT 1702.620 1863.490 1703.800 1864.670 ;
        RECT 1702.620 1847.090 1703.800 1848.270 ;
        RECT 1702.620 1845.490 1703.800 1846.670 ;
        RECT 1702.620 1829.090 1703.800 1830.270 ;
        RECT 1702.620 1827.490 1703.800 1828.670 ;
        RECT 1702.620 1811.090 1703.800 1812.270 ;
        RECT 1702.620 1809.490 1703.800 1810.670 ;
        RECT 1702.620 1685.090 1703.800 1686.270 ;
        RECT 1702.620 1683.490 1703.800 1684.670 ;
        RECT 1702.620 1667.090 1703.800 1668.270 ;
        RECT 1702.620 1665.490 1703.800 1666.670 ;
        RECT 1702.620 1649.090 1703.800 1650.270 ;
        RECT 1702.620 1647.490 1703.800 1648.670 ;
        RECT 1702.620 1631.090 1703.800 1632.270 ;
        RECT 1702.620 1629.490 1703.800 1630.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2632.680 2027.090 2633.860 2028.270 ;
        RECT 2632.680 2025.490 2633.860 2026.670 ;
        RECT 2632.680 2009.090 2633.860 2010.270 ;
        RECT 2632.680 2007.490 2633.860 2008.670 ;
        RECT 2632.680 1991.090 2633.860 1992.270 ;
        RECT 2632.680 1989.490 2633.860 1990.670 ;
        RECT 2632.680 1865.090 2633.860 1866.270 ;
        RECT 2632.680 1863.490 2633.860 1864.670 ;
        RECT 2632.680 1847.090 2633.860 1848.270 ;
        RECT 2632.680 1845.490 2633.860 1846.670 ;
        RECT 2632.680 1829.090 2633.860 1830.270 ;
        RECT 2632.680 1827.490 2633.860 1828.670 ;
        RECT 2632.680 1811.090 2633.860 1812.270 ;
        RECT 2632.680 1809.490 2633.860 1810.670 ;
        RECT 2632.680 1685.090 2633.860 1686.270 ;
        RECT 2632.680 1683.490 2633.860 1684.670 ;
        RECT 2632.680 1667.090 2633.860 1668.270 ;
        RECT 2632.680 1665.490 2633.860 1666.670 ;
        RECT 2632.680 1649.090 2633.860 1650.270 ;
        RECT 2632.680 1647.490 2633.860 1648.670 ;
        RECT 2632.680 1631.090 2633.860 1632.270 ;
        RECT 2632.680 1629.490 2633.860 1630.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1571.250 1469.090 1572.430 1470.270 ;
        RECT 1571.250 1467.490 1572.430 1468.670 ;
        RECT 1571.250 1451.090 1572.430 1452.270 ;
        RECT 1571.250 1449.490 1572.430 1450.670 ;
        RECT 1571.250 1325.090 1572.430 1326.270 ;
        RECT 1571.250 1323.490 1572.430 1324.670 ;
        RECT 1571.250 1307.090 1572.430 1308.270 ;
        RECT 1571.250 1305.490 1572.430 1306.670 ;
        RECT 1571.250 1289.090 1572.430 1290.270 ;
        RECT 1571.250 1287.490 1572.430 1288.670 ;
        RECT 1571.250 1271.090 1572.430 1272.270 ;
        RECT 1571.250 1269.490 1572.430 1270.670 ;
        RECT 1571.250 1145.090 1572.430 1146.270 ;
        RECT 1571.250 1143.490 1572.430 1144.670 ;
        RECT 1571.250 1127.090 1572.430 1128.270 ;
        RECT 1571.250 1125.490 1572.430 1126.670 ;
        RECT 1571.250 1109.090 1572.430 1110.270 ;
        RECT 1571.250 1107.490 1572.430 1108.670 ;
        RECT 1571.250 1091.090 1572.430 1092.270 ;
        RECT 1571.250 1089.490 1572.430 1090.670 ;
        RECT 1571.250 965.090 1572.430 966.270 ;
        RECT 1571.250 963.490 1572.430 964.670 ;
        RECT 1571.250 947.090 1572.430 948.270 ;
        RECT 1571.250 945.490 1572.430 946.670 ;
        RECT 1571.250 929.090 1572.430 930.270 ;
        RECT 1571.250 927.490 1572.430 928.670 ;
        RECT 1571.250 911.090 1572.430 912.270 ;
        RECT 1571.250 909.490 1572.430 910.670 ;
        RECT 1571.250 785.090 1572.430 786.270 ;
        RECT 1571.250 783.490 1572.430 784.670 ;
        RECT 1571.250 767.090 1572.430 768.270 ;
        RECT 1571.250 765.490 1572.430 766.670 ;
        RECT 1571.250 749.090 1572.430 750.270 ;
        RECT 1571.250 747.490 1572.430 748.670 ;
        RECT 1571.250 731.090 1572.430 732.270 ;
        RECT 1571.250 729.490 1572.430 730.670 ;
        RECT 1571.250 605.090 1572.430 606.270 ;
        RECT 1571.250 603.490 1572.430 604.670 ;
        RECT 1571.250 587.090 1572.430 588.270 ;
        RECT 1571.250 585.490 1572.430 586.670 ;
        RECT 1571.250 569.090 1572.430 570.270 ;
        RECT 1571.250 567.490 1572.430 568.670 ;
        RECT 1571.250 551.090 1572.430 552.270 ;
        RECT 1571.250 549.490 1572.430 550.670 ;
        RECT 1571.250 425.090 1572.430 426.270 ;
        RECT 1571.250 423.490 1572.430 424.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 682.470 3126.380 684.070 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 1332.470 3126.380 1334.070 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1932.470 3126.380 1934.070 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2582.470 3126.380 2584.070 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 682.470 3123.370 684.070 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 1332.470 3123.370 1334.070 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1932.470 3123.370 1934.070 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2582.470 3123.370 2584.070 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 682.470 3108.380 684.070 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 1332.470 3108.380 1334.070 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1932.470 3108.380 1934.070 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2582.470 3108.380 2584.070 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 682.470 3105.370 684.070 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 1332.470 3105.370 1334.070 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1932.470 3105.370 1934.070 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2582.470 3105.370 2584.070 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 682.470 3090.380 684.070 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1332.470 3090.380 1334.070 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1932.470 3090.380 1934.070 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2582.470 3090.380 2584.070 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 682.470 3087.370 684.070 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1332.470 3087.370 1334.070 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1932.470 3087.370 1934.070 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2582.470 3087.370 2584.070 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 682.470 3072.380 684.070 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1332.470 3072.380 1334.070 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1932.470 3072.380 1934.070 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2582.470 3072.380 2584.070 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 682.470 3069.370 684.070 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1332.470 3069.370 1334.070 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1932.470 3069.370 1934.070 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2582.470 3069.370 2584.070 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 682.470 2946.380 684.070 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 1332.470 2946.380 1334.070 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1932.470 2946.380 1934.070 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2582.470 2946.380 2584.070 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 682.470 2943.370 684.070 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 1332.470 2943.370 1334.070 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1932.470 2943.370 1934.070 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2582.470 2943.370 2584.070 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 682.470 2928.380 684.070 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 1332.470 2928.380 1334.070 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1932.470 2928.380 1934.070 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2582.470 2928.380 2584.070 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 682.470 2925.370 684.070 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 1332.470 2925.370 1334.070 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1932.470 2925.370 1934.070 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2582.470 2925.370 2584.070 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 682.470 2910.380 684.070 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1332.470 2910.380 1334.070 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1932.470 2910.380 1934.070 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2582.470 2910.380 2584.070 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 682.470 2907.370 684.070 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1332.470 2907.370 1334.070 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1932.470 2907.370 1934.070 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2582.470 2907.370 2584.070 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 682.470 2892.380 684.070 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1332.470 2892.380 1334.070 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1932.470 2892.380 1934.070 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2582.470 2892.380 2584.070 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 682.470 2889.370 684.070 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1332.470 2889.370 1334.070 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1932.470 2889.370 1934.070 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2582.470 2889.370 2584.070 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 321.040 2586.380 322.640 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 321.040 2583.370 322.640 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 321.040 2568.380 322.640 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 321.040 2565.370 322.640 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 321.040 2550.380 322.640 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 321.040 2547.370 322.640 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 321.040 2532.380 322.640 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 321.040 2529.370 322.640 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 321.040 2406.380 322.640 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 321.040 2403.370 322.640 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 321.040 2388.380 322.640 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 321.040 2385.370 322.640 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 321.040 2370.380 322.640 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 321.040 2367.370 322.640 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 321.040 2352.380 322.640 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 321.040 2349.370 322.640 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 321.040 2226.380 322.640 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 321.040 2223.370 322.640 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 321.040 2208.380 322.640 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 321.040 2205.370 322.640 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 321.040 2190.380 322.640 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 321.040 2187.370 322.640 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 321.040 2172.380 322.640 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 321.040 2169.370 322.640 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 321.040 2046.380 322.640 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1702.410 2046.380 1704.010 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 321.040 2043.370 322.640 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1702.410 2043.370 1704.010 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 321.040 2028.380 322.640 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1702.410 2028.380 1704.010 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2632.470 2028.380 2634.070 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 321.040 2025.370 322.640 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1702.410 2025.370 1704.010 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2632.470 2025.370 2634.070 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 321.040 2010.380 322.640 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1702.410 2010.380 1704.010 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2632.470 2010.380 2634.070 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 321.040 2007.370 322.640 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1702.410 2007.370 1704.010 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2632.470 2007.370 2634.070 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 321.040 1992.380 322.640 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1702.410 1992.380 1704.010 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2632.470 1992.380 2634.070 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 321.040 1989.370 322.640 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1702.410 1989.370 1704.010 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2632.470 1989.370 2634.070 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 321.040 1866.380 322.640 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1702.410 1866.380 1704.010 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2632.470 1866.380 2634.070 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 321.040 1863.370 322.640 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1702.410 1863.370 1704.010 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2632.470 1863.370 2634.070 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 321.040 1848.380 322.640 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1702.410 1848.380 1704.010 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2632.470 1848.380 2634.070 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 321.040 1845.370 322.640 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1702.410 1845.370 1704.010 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2632.470 1845.370 2634.070 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 321.040 1830.380 322.640 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1702.410 1830.380 1704.010 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2632.470 1830.380 2634.070 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 321.040 1827.370 322.640 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1702.410 1827.370 1704.010 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2632.470 1827.370 2634.070 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 321.040 1812.380 322.640 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1702.410 1812.380 1704.010 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2632.470 1812.380 2634.070 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 321.040 1809.370 322.640 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1702.410 1809.370 1704.010 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2632.470 1809.370 2634.070 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 321.040 1686.380 322.640 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1702.410 1686.380 1704.010 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2632.470 1686.380 2634.070 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 321.040 1683.370 322.640 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1702.410 1683.370 1704.010 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2632.470 1683.370 2634.070 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 321.040 1668.380 322.640 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1702.410 1668.380 1704.010 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2632.470 1668.380 2634.070 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 321.040 1665.370 322.640 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1702.410 1665.370 1704.010 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2632.470 1665.370 2634.070 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 321.040 1650.380 322.640 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1702.410 1650.380 1704.010 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2632.470 1650.380 2634.070 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 321.040 1647.370 322.640 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1702.410 1647.370 1704.010 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2632.470 1647.370 2634.070 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 321.040 1632.380 322.640 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1702.410 1632.380 1704.010 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2632.470 1632.380 2634.070 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 321.040 1629.370 322.640 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1702.410 1629.370 1704.010 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2632.470 1629.370 2634.070 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1571.040 1470.380 1572.640 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1571.040 1467.370 1572.640 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1571.040 1452.380 1572.640 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1571.040 1449.370 1572.640 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1571.040 1326.380 1572.640 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1571.040 1323.370 1572.640 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1571.040 1308.380 1572.640 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1571.040 1305.370 1572.640 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1571.040 1290.380 1572.640 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1571.040 1287.370 1572.640 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1571.040 1272.380 1572.640 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1571.040 1269.370 1572.640 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1571.040 1146.380 1572.640 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1571.040 1143.370 1572.640 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1571.040 1128.380 1572.640 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1571.040 1125.370 1572.640 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1571.040 1110.380 1572.640 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1571.040 1107.370 1572.640 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1571.040 1092.380 1572.640 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1571.040 1089.370 1572.640 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1571.040 966.380 1572.640 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1571.040 963.370 1572.640 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1571.040 948.380 1572.640 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1571.040 945.370 1572.640 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1571.040 930.380 1572.640 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1571.040 927.370 1572.640 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1571.040 912.380 1572.640 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1571.040 909.370 1572.640 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1571.040 786.380 1572.640 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1571.040 783.370 1572.640 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1571.040 768.380 1572.640 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1571.040 765.370 1572.640 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1571.040 750.380 1572.640 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1571.040 747.370 1572.640 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1571.040 732.380 1572.640 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1571.040 729.370 1572.640 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1571.040 606.380 1572.640 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1571.040 603.370 1572.640 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1571.040 588.380 1572.640 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1571.040 585.370 1572.640 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1571.040 570.380 1572.640 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1571.040 567.370 1572.640 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1571.040 552.380 1572.640 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1571.040 549.370 1572.640 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1571.040 426.380 1572.640 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1571.040 423.370 1572.640 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.040 3251.235 686.300 3252.140 ;
        RECT 1331.040 3251.235 1336.300 3252.140 ;
        RECT 1931.040 3251.235 1936.300 3252.140 ;
        RECT 2581.040 3251.235 2586.300 3252.140 ;
        RECT 681.480 3250.400 686.300 3251.235 ;
        RECT 1331.480 3250.400 1336.300 3251.235 ;
        RECT 1931.480 3250.400 1936.300 3251.235 ;
        RECT 2581.480 3250.400 2586.300 3251.235 ;
        RECT 2631.040 2051.235 2636.300 2052.140 ;
        RECT 2631.480 2050.400 2636.300 2051.235 ;
        RECT 1700.180 1605.000 1705.000 1605.835 ;
        RECT 1700.180 1604.095 1705.440 1605.000 ;
      LAYER via3 ;
        RECT 684.720 3250.440 686.240 3252.050 ;
        RECT 1334.720 3250.440 1336.240 3252.050 ;
        RECT 1934.720 3250.440 1936.240 3252.050 ;
        RECT 2584.720 3250.440 2586.240 3252.050 ;
        RECT 2634.720 2050.440 2636.240 2052.050 ;
        RECT 1700.240 1604.185 1701.760 1605.795 ;
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 292.020 3271.235 295.020 3538.400 ;
        RECT 310.020 3271.235 313.020 3547.800 ;
        RECT 328.020 3271.235 331.020 3557.200 ;
        RECT 454.020 3271.235 457.020 3529.000 ;
        RECT 472.020 3271.235 475.020 3538.400 ;
        RECT 490.020 3271.235 493.020 3547.800 ;
        RECT 508.020 3271.235 511.020 3557.200 ;
        RECT 634.020 3271.235 637.020 3529.000 ;
        RECT 652.020 3271.235 655.020 3538.400 ;
        RECT 670.020 3271.235 673.020 3547.800 ;
        RECT 688.020 3271.235 691.020 3557.200 ;
        RECT 684.690 2804.060 686.310 3252.140 ;
        RECT 814.020 2715.000 817.020 3529.000 ;
        RECT 832.020 2715.000 835.020 3538.400 ;
        RECT 850.020 2715.000 853.020 3547.800 ;
        RECT 868.020 2715.000 871.020 3557.200 ;
        RECT 994.020 3271.235 997.020 3529.000 ;
        RECT 1012.020 3271.235 1015.020 3538.400 ;
        RECT 1030.020 3271.235 1033.020 3547.800 ;
        RECT 1048.020 3271.235 1051.020 3557.200 ;
        RECT 1174.020 3271.235 1177.020 3529.000 ;
        RECT 1192.020 3271.235 1195.020 3538.400 ;
        RECT 1210.020 3271.235 1213.020 3547.800 ;
        RECT 1228.020 3271.235 1231.020 3557.200 ;
        RECT 1334.690 2804.060 1336.310 3252.140 ;
        RECT 1354.020 2715.000 1357.020 3529.000 ;
        RECT 1372.020 2715.000 1375.020 3538.400 ;
        RECT 1390.020 2715.000 1393.020 3547.800 ;
        RECT 1408.020 2715.000 1411.020 3557.200 ;
        RECT 1534.020 3271.235 1537.020 3529.000 ;
        RECT 1552.020 3271.235 1555.020 3538.400 ;
        RECT 1570.020 3271.235 1573.020 3547.800 ;
        RECT 1588.020 3271.235 1591.020 3557.200 ;
        RECT 1714.020 3271.235 1717.020 3529.000 ;
        RECT 1732.020 3271.235 1735.020 3538.400 ;
        RECT 1750.020 3271.235 1753.020 3547.800 ;
        RECT 1768.020 3271.235 1771.020 3557.200 ;
        RECT 1894.020 3271.235 1897.020 3529.000 ;
        RECT 1912.020 3271.235 1915.020 3538.400 ;
        RECT 1930.020 3271.235 1933.020 3547.800 ;
        RECT 1948.020 3271.235 1951.020 3557.200 ;
        RECT 1934.690 2804.060 1936.310 3252.140 ;
        RECT 397.840 1610.640 399.440 2688.240 ;
        RECT 292.020 -18.720 295.020 1585.000 ;
        RECT 310.020 -28.120 313.020 1585.000 ;
        RECT 328.020 -37.520 331.020 1585.000 ;
        RECT 454.020 -9.320 457.020 1585.000 ;
        RECT 472.020 -18.720 475.020 1585.000 ;
        RECT 490.020 -28.120 493.020 1585.000 ;
        RECT 508.020 -37.520 511.020 1585.000 ;
        RECT 634.020 -9.320 637.020 1585.000 ;
        RECT 652.020 -18.720 655.020 1585.000 ;
        RECT 670.020 -28.120 673.020 1585.000 ;
        RECT 688.020 -37.520 691.020 1585.000 ;
        RECT 814.020 -9.320 817.020 1585.000 ;
        RECT 832.020 -18.720 835.020 1585.000 ;
        RECT 850.020 -28.120 853.020 1585.000 ;
        RECT 868.020 -37.520 871.020 1585.000 ;
        RECT 994.020 -9.320 997.020 1585.000 ;
        RECT 1012.020 -18.720 1015.020 1585.000 ;
        RECT 1030.020 -28.120 1033.020 1585.000 ;
        RECT 1048.020 -37.520 1051.020 1585.000 ;
        RECT 1174.020 -9.320 1177.020 1585.000 ;
        RECT 1192.020 -18.720 1195.020 1585.000 ;
        RECT 1210.020 -28.120 1213.020 1585.000 ;
        RECT 1228.020 -37.520 1231.020 1585.000 ;
        RECT 1354.020 -9.320 1357.020 1585.000 ;
        RECT 1372.020 -18.720 1375.020 1585.000 ;
        RECT 1390.020 -28.120 1393.020 1585.000 ;
        RECT 1408.020 -37.520 1411.020 1585.000 ;
        RECT 1534.020 1515.000 1537.020 2785.000 ;
        RECT 1552.020 1515.000 1555.020 2785.000 ;
        RECT 1570.020 1515.000 1573.020 2785.000 ;
        RECT 1588.020 1515.000 1591.020 2785.000 ;
        RECT 1714.020 2071.235 1717.020 2785.000 ;
        RECT 1732.020 2071.235 1735.020 2785.000 ;
        RECT 1750.020 2071.235 1753.020 2785.000 ;
        RECT 1768.020 2071.235 1771.020 2785.000 ;
        RECT 1894.020 2071.235 1897.020 2785.000 ;
        RECT 1912.020 2071.235 1915.020 2785.000 ;
        RECT 1930.020 2071.235 1933.020 2785.000 ;
        RECT 1948.020 2071.235 1951.020 2785.000 ;
        RECT 2074.020 2071.235 2077.020 3529.000 ;
        RECT 2092.020 2071.235 2095.020 3538.400 ;
        RECT 1700.170 1604.095 1701.790 2052.175 ;
        RECT 1714.020 1515.000 1717.020 1585.000 ;
        RECT 1732.020 1515.000 1735.020 1585.000 ;
        RECT 1750.020 1515.000 1753.020 1585.000 ;
        RECT 1894.020 1515.000 1897.020 1585.000 ;
        RECT 1912.020 1515.000 1915.020 1585.000 ;
        RECT 1930.020 1515.000 1933.020 1585.000 ;
        RECT 2074.020 1515.000 2077.020 1585.000 ;
        RECT 2092.020 1515.000 2095.020 1585.000 ;
        RECT 2110.020 1515.000 2113.020 3547.800 ;
        RECT 2128.020 1515.000 2131.020 3557.200 ;
        RECT 2254.020 3271.235 2257.020 3529.000 ;
        RECT 2272.020 3271.235 2275.020 3538.400 ;
        RECT 2290.020 3271.235 2293.020 3547.800 ;
        RECT 2308.020 3271.235 2311.020 3557.200 ;
        RECT 2434.020 3271.235 2437.020 3529.000 ;
        RECT 2452.020 3271.235 2455.020 3538.400 ;
        RECT 2470.020 3271.235 2473.020 3547.800 ;
        RECT 2488.020 3271.235 2491.020 3557.200 ;
        RECT 2584.690 2804.060 2586.310 3252.140 ;
        RECT 2254.020 2071.235 2257.020 2785.000 ;
        RECT 2272.020 2071.235 2275.020 2785.000 ;
        RECT 2290.020 2071.235 2293.020 2785.000 ;
        RECT 2308.020 2071.235 2311.020 2785.000 ;
        RECT 2434.020 2071.235 2437.020 2785.000 ;
        RECT 2452.020 2071.235 2455.020 2785.000 ;
        RECT 2470.020 2071.235 2473.020 2785.000 ;
        RECT 2488.020 2071.235 2491.020 2785.000 ;
        RECT 2614.020 2071.235 2617.020 3529.000 ;
        RECT 2632.020 2071.235 2635.020 3538.400 ;
        RECT 2650.020 2071.235 2653.020 3547.800 ;
        RECT 2634.690 1604.060 2636.310 2052.140 ;
        RECT 2254.020 1515.000 2257.020 1585.000 ;
        RECT 2272.020 1515.000 2275.020 1585.000 ;
        RECT 2290.020 1515.000 2293.020 1585.000 ;
        RECT 2434.020 1515.000 2437.020 1585.000 ;
        RECT 2452.020 1515.000 2455.020 1585.000 ;
        RECT 2470.020 1515.000 2473.020 1585.000 ;
        RECT 2614.020 1515.000 2617.020 1585.000 ;
        RECT 2632.020 1515.000 2635.020 1585.000 ;
        RECT 2650.020 1515.000 2653.020 1585.000 ;
        RECT 1647.840 410.640 1649.440 1488.240 ;
        RECT 1534.020 -9.320 1537.020 385.000 ;
        RECT 1552.020 -18.720 1555.020 385.000 ;
        RECT 1570.020 -28.120 1573.020 385.000 ;
        RECT 1588.020 -37.520 1591.020 385.000 ;
        RECT 1714.020 -9.320 1717.020 385.000 ;
        RECT 1732.020 -18.720 1735.020 385.000 ;
        RECT 1750.020 -28.120 1753.020 385.000 ;
        RECT 1768.020 -37.520 1771.020 385.000 ;
        RECT 1894.020 -9.320 1897.020 385.000 ;
        RECT 1912.020 -18.720 1915.020 385.000 ;
        RECT 1930.020 -28.120 1933.020 385.000 ;
        RECT 1948.020 -37.520 1951.020 385.000 ;
        RECT 2074.020 -9.320 2077.020 385.000 ;
        RECT 2092.020 -18.720 2095.020 385.000 ;
        RECT 2110.020 -28.120 2113.020 385.000 ;
        RECT 2128.020 -37.520 2131.020 385.000 ;
        RECT 2254.020 -9.320 2257.020 385.000 ;
        RECT 2272.020 -18.720 2275.020 385.000 ;
        RECT 2290.020 -28.120 2293.020 385.000 ;
        RECT 2308.020 -37.520 2311.020 385.000 ;
        RECT 2434.020 -9.320 2437.020 385.000 ;
        RECT 2452.020 -18.720 2455.020 385.000 ;
        RECT 2470.020 -28.120 2473.020 385.000 ;
        RECT 2488.020 -37.520 2491.020 385.000 ;
        RECT 2614.020 -9.320 2617.020 385.000 ;
        RECT 2632.020 -18.720 2635.020 385.000 ;
        RECT 2650.020 -28.120 2653.020 385.000 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 684.910 3215.090 686.090 3216.270 ;
        RECT 684.910 3213.490 686.090 3214.670 ;
        RECT 684.910 3197.090 686.090 3198.270 ;
        RECT 684.910 3195.490 686.090 3196.670 ;
        RECT 684.910 3179.090 686.090 3180.270 ;
        RECT 684.910 3177.490 686.090 3178.670 ;
        RECT 684.910 3161.090 686.090 3162.270 ;
        RECT 684.910 3159.490 686.090 3160.670 ;
        RECT 684.910 3035.090 686.090 3036.270 ;
        RECT 684.910 3033.490 686.090 3034.670 ;
        RECT 684.910 3017.090 686.090 3018.270 ;
        RECT 684.910 3015.490 686.090 3016.670 ;
        RECT 684.910 2999.090 686.090 3000.270 ;
        RECT 684.910 2997.490 686.090 2998.670 ;
        RECT 684.910 2981.090 686.090 2982.270 ;
        RECT 684.910 2979.490 686.090 2980.670 ;
        RECT 684.910 2855.090 686.090 2856.270 ;
        RECT 684.910 2853.490 686.090 2854.670 ;
        RECT 684.910 2837.090 686.090 2838.270 ;
        RECT 684.910 2835.490 686.090 2836.670 ;
        RECT 684.910 2819.090 686.090 2820.270 ;
        RECT 684.910 2817.490 686.090 2818.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 1334.910 3215.090 1336.090 3216.270 ;
        RECT 1334.910 3213.490 1336.090 3214.670 ;
        RECT 1334.910 3197.090 1336.090 3198.270 ;
        RECT 1334.910 3195.490 1336.090 3196.670 ;
        RECT 1334.910 3179.090 1336.090 3180.270 ;
        RECT 1334.910 3177.490 1336.090 3178.670 ;
        RECT 1334.910 3161.090 1336.090 3162.270 ;
        RECT 1334.910 3159.490 1336.090 3160.670 ;
        RECT 1334.910 3035.090 1336.090 3036.270 ;
        RECT 1334.910 3033.490 1336.090 3034.670 ;
        RECT 1334.910 3017.090 1336.090 3018.270 ;
        RECT 1334.910 3015.490 1336.090 3016.670 ;
        RECT 1334.910 2999.090 1336.090 3000.270 ;
        RECT 1334.910 2997.490 1336.090 2998.670 ;
        RECT 1334.910 2981.090 1336.090 2982.270 ;
        RECT 1334.910 2979.490 1336.090 2980.670 ;
        RECT 1334.910 2855.090 1336.090 2856.270 ;
        RECT 1334.910 2853.490 1336.090 2854.670 ;
        RECT 1334.910 2837.090 1336.090 2838.270 ;
        RECT 1334.910 2835.490 1336.090 2836.670 ;
        RECT 1334.910 2819.090 1336.090 2820.270 ;
        RECT 1334.910 2817.490 1336.090 2818.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1934.910 3215.090 1936.090 3216.270 ;
        RECT 1934.910 3213.490 1936.090 3214.670 ;
        RECT 1934.910 3197.090 1936.090 3198.270 ;
        RECT 1934.910 3195.490 1936.090 3196.670 ;
        RECT 1934.910 3179.090 1936.090 3180.270 ;
        RECT 1934.910 3177.490 1936.090 3178.670 ;
        RECT 1934.910 3161.090 1936.090 3162.270 ;
        RECT 1934.910 3159.490 1936.090 3160.670 ;
        RECT 1934.910 3035.090 1936.090 3036.270 ;
        RECT 1934.910 3033.490 1936.090 3034.670 ;
        RECT 1934.910 3017.090 1936.090 3018.270 ;
        RECT 1934.910 3015.490 1936.090 3016.670 ;
        RECT 1934.910 2999.090 1936.090 3000.270 ;
        RECT 1934.910 2997.490 1936.090 2998.670 ;
        RECT 1934.910 2981.090 1936.090 2982.270 ;
        RECT 1934.910 2979.490 1936.090 2980.670 ;
        RECT 1934.910 2855.090 1936.090 2856.270 ;
        RECT 1934.910 2853.490 1936.090 2854.670 ;
        RECT 1934.910 2837.090 1936.090 2838.270 ;
        RECT 1934.910 2835.490 1936.090 2836.670 ;
        RECT 1934.910 2819.090 1936.090 2820.270 ;
        RECT 1934.910 2817.490 1936.090 2818.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 398.050 2675.090 399.230 2676.270 ;
        RECT 398.050 2673.490 399.230 2674.670 ;
        RECT 398.050 2657.090 399.230 2658.270 ;
        RECT 398.050 2655.490 399.230 2656.670 ;
        RECT 398.050 2639.090 399.230 2640.270 ;
        RECT 398.050 2637.490 399.230 2638.670 ;
        RECT 398.050 2621.090 399.230 2622.270 ;
        RECT 398.050 2619.490 399.230 2620.670 ;
        RECT 398.050 2495.090 399.230 2496.270 ;
        RECT 398.050 2493.490 399.230 2494.670 ;
        RECT 398.050 2477.090 399.230 2478.270 ;
        RECT 398.050 2475.490 399.230 2476.670 ;
        RECT 398.050 2459.090 399.230 2460.270 ;
        RECT 398.050 2457.490 399.230 2458.670 ;
        RECT 398.050 2441.090 399.230 2442.270 ;
        RECT 398.050 2439.490 399.230 2440.670 ;
        RECT 398.050 2315.090 399.230 2316.270 ;
        RECT 398.050 2313.490 399.230 2314.670 ;
        RECT 398.050 2297.090 399.230 2298.270 ;
        RECT 398.050 2295.490 399.230 2296.670 ;
        RECT 398.050 2279.090 399.230 2280.270 ;
        RECT 398.050 2277.490 399.230 2278.670 ;
        RECT 398.050 2261.090 399.230 2262.270 ;
        RECT 398.050 2259.490 399.230 2260.670 ;
        RECT 398.050 2135.090 399.230 2136.270 ;
        RECT 398.050 2133.490 399.230 2134.670 ;
        RECT 398.050 2117.090 399.230 2118.270 ;
        RECT 398.050 2115.490 399.230 2116.670 ;
        RECT 398.050 2099.090 399.230 2100.270 ;
        RECT 398.050 2097.490 399.230 2098.670 ;
        RECT 398.050 2081.090 399.230 2082.270 ;
        RECT 398.050 2079.490 399.230 2080.670 ;
        RECT 398.050 1955.090 399.230 1956.270 ;
        RECT 398.050 1953.490 399.230 1954.670 ;
        RECT 398.050 1937.090 399.230 1938.270 ;
        RECT 398.050 1935.490 399.230 1936.670 ;
        RECT 398.050 1919.090 399.230 1920.270 ;
        RECT 398.050 1917.490 399.230 1918.670 ;
        RECT 398.050 1901.090 399.230 1902.270 ;
        RECT 398.050 1899.490 399.230 1900.670 ;
        RECT 398.050 1775.090 399.230 1776.270 ;
        RECT 398.050 1773.490 399.230 1774.670 ;
        RECT 398.050 1757.090 399.230 1758.270 ;
        RECT 398.050 1755.490 399.230 1756.670 ;
        RECT 398.050 1739.090 399.230 1740.270 ;
        RECT 398.050 1737.490 399.230 1738.670 ;
        RECT 398.050 1721.090 399.230 1722.270 ;
        RECT 398.050 1719.490 399.230 1720.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1700.390 1955.090 1701.570 1956.270 ;
        RECT 1700.390 1953.490 1701.570 1954.670 ;
        RECT 1700.390 1937.090 1701.570 1938.270 ;
        RECT 1700.390 1935.490 1701.570 1936.670 ;
        RECT 1700.390 1919.090 1701.570 1920.270 ;
        RECT 1700.390 1917.490 1701.570 1918.670 ;
        RECT 1700.390 1901.090 1701.570 1902.270 ;
        RECT 1700.390 1899.490 1701.570 1900.670 ;
        RECT 1700.390 1775.090 1701.570 1776.270 ;
        RECT 1700.390 1773.490 1701.570 1774.670 ;
        RECT 1700.390 1757.090 1701.570 1758.270 ;
        RECT 1700.390 1755.490 1701.570 1756.670 ;
        RECT 1700.390 1739.090 1701.570 1740.270 ;
        RECT 1700.390 1737.490 1701.570 1738.670 ;
        RECT 1700.390 1721.090 1701.570 1722.270 ;
        RECT 1700.390 1719.490 1701.570 1720.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2584.910 3215.090 2586.090 3216.270 ;
        RECT 2584.910 3213.490 2586.090 3214.670 ;
        RECT 2584.910 3197.090 2586.090 3198.270 ;
        RECT 2584.910 3195.490 2586.090 3196.670 ;
        RECT 2584.910 3179.090 2586.090 3180.270 ;
        RECT 2584.910 3177.490 2586.090 3178.670 ;
        RECT 2584.910 3161.090 2586.090 3162.270 ;
        RECT 2584.910 3159.490 2586.090 3160.670 ;
        RECT 2584.910 3035.090 2586.090 3036.270 ;
        RECT 2584.910 3033.490 2586.090 3034.670 ;
        RECT 2584.910 3017.090 2586.090 3018.270 ;
        RECT 2584.910 3015.490 2586.090 3016.670 ;
        RECT 2584.910 2999.090 2586.090 3000.270 ;
        RECT 2584.910 2997.490 2586.090 2998.670 ;
        RECT 2584.910 2981.090 2586.090 2982.270 ;
        RECT 2584.910 2979.490 2586.090 2980.670 ;
        RECT 2584.910 2855.090 2586.090 2856.270 ;
        RECT 2584.910 2853.490 2586.090 2854.670 ;
        RECT 2584.910 2837.090 2586.090 2838.270 ;
        RECT 2584.910 2835.490 2586.090 2836.670 ;
        RECT 2584.910 2819.090 2586.090 2820.270 ;
        RECT 2584.910 2817.490 2586.090 2818.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2634.910 1955.090 2636.090 1956.270 ;
        RECT 2634.910 1953.490 2636.090 1954.670 ;
        RECT 2634.910 1937.090 2636.090 1938.270 ;
        RECT 2634.910 1935.490 2636.090 1936.670 ;
        RECT 2634.910 1919.090 2636.090 1920.270 ;
        RECT 2634.910 1917.490 2636.090 1918.670 ;
        RECT 2634.910 1901.090 2636.090 1902.270 ;
        RECT 2634.910 1899.490 2636.090 1900.670 ;
        RECT 2634.910 1775.090 2636.090 1776.270 ;
        RECT 2634.910 1773.490 2636.090 1774.670 ;
        RECT 2634.910 1757.090 2636.090 1758.270 ;
        RECT 2634.910 1755.490 2636.090 1756.670 ;
        RECT 2634.910 1739.090 2636.090 1740.270 ;
        RECT 2634.910 1737.490 2636.090 1738.670 ;
        RECT 2634.910 1721.090 2636.090 1722.270 ;
        RECT 2634.910 1719.490 2636.090 1720.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1648.050 1415.090 1649.230 1416.270 ;
        RECT 1648.050 1413.490 1649.230 1414.670 ;
        RECT 1648.050 1397.090 1649.230 1398.270 ;
        RECT 1648.050 1395.490 1649.230 1396.670 ;
        RECT 1648.050 1379.090 1649.230 1380.270 ;
        RECT 1648.050 1377.490 1649.230 1378.670 ;
        RECT 1648.050 1361.090 1649.230 1362.270 ;
        RECT 1648.050 1359.490 1649.230 1360.670 ;
        RECT 1648.050 1235.090 1649.230 1236.270 ;
        RECT 1648.050 1233.490 1649.230 1234.670 ;
        RECT 1648.050 1217.090 1649.230 1218.270 ;
        RECT 1648.050 1215.490 1649.230 1216.670 ;
        RECT 1648.050 1199.090 1649.230 1200.270 ;
        RECT 1648.050 1197.490 1649.230 1198.670 ;
        RECT 1648.050 1181.090 1649.230 1182.270 ;
        RECT 1648.050 1179.490 1649.230 1180.670 ;
        RECT 1648.050 1055.090 1649.230 1056.270 ;
        RECT 1648.050 1053.490 1649.230 1054.670 ;
        RECT 1648.050 1037.090 1649.230 1038.270 ;
        RECT 1648.050 1035.490 1649.230 1036.670 ;
        RECT 1648.050 1019.090 1649.230 1020.270 ;
        RECT 1648.050 1017.490 1649.230 1018.670 ;
        RECT 1648.050 1001.090 1649.230 1002.270 ;
        RECT 1648.050 999.490 1649.230 1000.670 ;
        RECT 1648.050 875.090 1649.230 876.270 ;
        RECT 1648.050 873.490 1649.230 874.670 ;
        RECT 1648.050 857.090 1649.230 858.270 ;
        RECT 1648.050 855.490 1649.230 856.670 ;
        RECT 1648.050 839.090 1649.230 840.270 ;
        RECT 1648.050 837.490 1649.230 838.670 ;
        RECT 1648.050 821.090 1649.230 822.270 ;
        RECT 1648.050 819.490 1649.230 820.670 ;
        RECT 1648.050 695.090 1649.230 696.270 ;
        RECT 1648.050 693.490 1649.230 694.670 ;
        RECT 1648.050 677.090 1649.230 678.270 ;
        RECT 1648.050 675.490 1649.230 676.670 ;
        RECT 1648.050 659.090 1649.230 660.270 ;
        RECT 1648.050 657.490 1649.230 658.670 ;
        RECT 1648.050 641.090 1649.230 642.270 ;
        RECT 1648.050 639.490 1649.230 640.670 ;
        RECT 1648.050 515.090 1649.230 516.270 ;
        RECT 1648.050 513.490 1649.230 514.670 ;
        RECT 1648.050 497.090 1649.230 498.270 ;
        RECT 1648.050 495.490 1649.230 496.670 ;
        RECT 1648.050 479.090 1649.230 480.270 ;
        RECT 1648.050 477.490 1649.230 478.670 ;
        RECT 1648.050 461.090 1649.230 462.270 ;
        RECT 1648.050 459.490 1649.230 460.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 684.690 3216.380 686.310 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1334.690 3216.380 1336.310 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1934.690 3216.380 1936.310 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2584.690 3216.380 2586.310 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 684.690 3213.370 686.310 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1334.690 3213.370 1336.310 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1934.690 3213.370 1936.310 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2584.690 3213.370 2586.310 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 684.690 3198.380 686.310 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1334.690 3198.380 1336.310 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1934.690 3198.380 1936.310 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2584.690 3198.380 2586.310 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 684.690 3195.370 686.310 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1334.690 3195.370 1336.310 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1934.690 3195.370 1936.310 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2584.690 3195.370 2586.310 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 684.690 3180.380 686.310 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1334.690 3180.380 1336.310 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1934.690 3180.380 1936.310 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2584.690 3180.380 2586.310 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 684.690 3177.370 686.310 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1334.690 3177.370 1336.310 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1934.690 3177.370 1936.310 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2584.690 3177.370 2586.310 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 684.690 3162.380 686.310 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 1334.690 3162.380 1336.310 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1934.690 3162.380 1936.310 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2584.690 3162.380 2586.310 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 684.690 3159.370 686.310 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 1334.690 3159.370 1336.310 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1934.690 3159.370 1936.310 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2584.690 3159.370 2586.310 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 684.690 3036.380 686.310 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1334.690 3036.380 1336.310 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1934.690 3036.380 1936.310 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2584.690 3036.380 2586.310 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 684.690 3033.370 686.310 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1334.690 3033.370 1336.310 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1934.690 3033.370 1936.310 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2584.690 3033.370 2586.310 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 684.690 3018.380 686.310 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1334.690 3018.380 1336.310 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1934.690 3018.380 1936.310 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2584.690 3018.380 2586.310 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 684.690 3015.370 686.310 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1334.690 3015.370 1336.310 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1934.690 3015.370 1936.310 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2584.690 3015.370 2586.310 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 684.690 3000.380 686.310 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1334.690 3000.380 1336.310 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1934.690 3000.380 1936.310 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2584.690 3000.380 2586.310 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 684.690 2997.370 686.310 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1334.690 2997.370 1336.310 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1934.690 2997.370 1936.310 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2584.690 2997.370 2586.310 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 684.690 2982.380 686.310 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 1334.690 2982.380 1336.310 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1934.690 2982.380 1936.310 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2584.690 2982.380 2586.310 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 684.690 2979.370 686.310 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 1334.690 2979.370 1336.310 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1934.690 2979.370 1936.310 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2584.690 2979.370 2586.310 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 684.690 2856.380 686.310 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1334.690 2856.380 1336.310 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1934.690 2856.380 1936.310 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2584.690 2856.380 2586.310 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 684.690 2853.370 686.310 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1334.690 2853.370 1336.310 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1934.690 2853.370 1936.310 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2584.690 2853.370 2586.310 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 684.690 2838.380 686.310 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1334.690 2838.380 1336.310 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1934.690 2838.380 1936.310 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2584.690 2838.380 2586.310 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 684.690 2835.370 686.310 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1334.690 2835.370 1336.310 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1934.690 2835.370 1936.310 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2584.690 2835.370 2586.310 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 684.690 2820.380 686.310 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1334.690 2820.380 1336.310 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1934.690 2820.380 1936.310 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2584.690 2820.380 2586.310 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 684.690 2817.370 686.310 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1334.690 2817.370 1336.310 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1934.690 2817.370 1936.310 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2584.690 2817.370 2586.310 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 397.840 2676.380 399.440 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 397.840 2673.370 399.440 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 397.840 2658.380 399.440 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 397.840 2655.370 399.440 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 397.840 2640.380 399.440 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 397.840 2637.370 399.440 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 397.840 2622.380 399.440 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 397.840 2619.370 399.440 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 397.840 2496.380 399.440 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 397.840 2493.370 399.440 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 397.840 2478.380 399.440 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 397.840 2475.370 399.440 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 397.840 2460.380 399.440 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 397.840 2457.370 399.440 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 397.840 2442.380 399.440 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 397.840 2439.370 399.440 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 397.840 2316.380 399.440 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 397.840 2313.370 399.440 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 397.840 2298.380 399.440 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 397.840 2295.370 399.440 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 397.840 2280.380 399.440 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 397.840 2277.370 399.440 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 397.840 2262.380 399.440 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 397.840 2259.370 399.440 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 397.840 2136.380 399.440 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 397.840 2133.370 399.440 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 397.840 2118.380 399.440 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 397.840 2115.370 399.440 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 397.840 2100.380 399.440 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 397.840 2097.370 399.440 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 397.840 2082.380 399.440 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 397.840 2079.370 399.440 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 397.840 1956.380 399.440 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1700.170 1956.380 1701.790 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2634.690 1956.380 2636.310 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 397.840 1953.370 399.440 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1700.170 1953.370 1701.790 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2634.690 1953.370 2636.310 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 397.840 1938.380 399.440 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1700.170 1938.380 1701.790 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2634.690 1938.380 2636.310 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 397.840 1935.370 399.440 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1700.170 1935.370 1701.790 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2634.690 1935.370 2636.310 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 397.840 1920.380 399.440 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1700.170 1920.380 1701.790 1920.390 ;
        RECT 2634.690 1920.380 2636.310 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 397.840 1917.370 399.440 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1700.170 1917.370 1701.790 1917.380 ;
        RECT 2634.690 1917.370 2636.310 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 397.840 1902.380 399.440 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1700.170 1902.380 1701.790 1902.390 ;
        RECT 2634.690 1902.380 2636.310 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 397.840 1899.370 399.440 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1700.170 1899.370 1701.790 1899.380 ;
        RECT 2634.690 1899.370 2636.310 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 397.840 1776.380 399.440 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1700.170 1776.380 1701.790 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2634.690 1776.380 2636.310 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 397.840 1773.370 399.440 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1700.170 1773.370 1701.790 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2634.690 1773.370 2636.310 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 397.840 1758.380 399.440 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1700.170 1758.380 1701.790 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2634.690 1758.380 2636.310 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 397.840 1755.370 399.440 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1700.170 1755.370 1701.790 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2634.690 1755.370 2636.310 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 397.840 1740.380 399.440 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1700.170 1740.380 1701.790 1740.390 ;
        RECT 2634.690 1740.380 2636.310 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 397.840 1737.370 399.440 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1700.170 1737.370 1701.790 1737.380 ;
        RECT 2634.690 1737.370 2636.310 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 397.840 1722.380 399.440 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1700.170 1722.380 1701.790 1722.390 ;
        RECT 2634.690 1722.380 2636.310 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 397.840 1719.370 399.440 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1700.170 1719.370 1701.790 1719.380 ;
        RECT 2634.690 1719.370 2636.310 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1647.840 1416.380 1649.440 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1647.840 1413.370 1649.440 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1647.840 1398.380 1649.440 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1647.840 1395.370 1649.440 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1647.840 1380.380 1649.440 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1647.840 1377.370 1649.440 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1647.840 1362.380 1649.440 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1647.840 1359.370 1649.440 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1647.840 1236.380 1649.440 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1647.840 1233.370 1649.440 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1647.840 1218.380 1649.440 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1647.840 1215.370 1649.440 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1647.840 1200.380 1649.440 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1647.840 1197.370 1649.440 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1647.840 1182.380 1649.440 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1647.840 1179.370 1649.440 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1647.840 1056.380 1649.440 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1647.840 1053.370 1649.440 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1647.840 1038.380 1649.440 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1647.840 1035.370 1649.440 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1647.840 1020.380 1649.440 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1647.840 1017.370 1649.440 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1647.840 1002.380 1649.440 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1647.840 999.370 1649.440 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1647.840 876.380 1649.440 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1647.840 873.370 1649.440 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1647.840 858.380 1649.440 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1647.840 855.370 1649.440 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1647.840 840.380 1649.440 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1647.840 837.370 1649.440 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1647.840 822.380 1649.440 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1647.840 819.370 1649.440 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1647.840 696.380 1649.440 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1647.840 693.370 1649.440 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1647.840 678.380 1649.440 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1647.840 675.370 1649.440 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1647.840 660.380 1649.440 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1647.840 657.370 1649.440 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1647.840 642.380 1649.440 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1647.840 639.370 1649.440 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1647.840 516.380 1649.440 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1647.840 513.370 1649.440 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1647.840 498.380 1649.440 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1647.840 495.370 1649.440 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1647.840 480.380 1649.440 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1647.840 477.370 1649.440 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1647.840 462.380 1649.440 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1647.840 459.370 1649.440 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 1304.245 3263.745 1304.415 3266.975 ;
        RECT 966.145 3251.505 966.315 3252.695 ;
        RECT 1013.985 3251.845 1014.155 3252.695 ;
        RECT 1062.745 3251.505 1062.915 3252.695 ;
        RECT 1110.585 3251.845 1110.755 3252.695 ;
        RECT 1159.345 3251.505 1159.515 3252.695 ;
        RECT 1207.185 3251.845 1207.355 3252.695 ;
        RECT 1255.945 3251.505 1256.115 3252.695 ;
        RECT 1303.785 3251.845 1303.955 3252.695 ;
        RECT 1400.845 3252.525 1401.015 3253.375 ;
        RECT 1365.885 3252.185 1366.515 3252.355 ;
        RECT 1448.685 3252.185 1448.855 3253.375 ;
        RECT 1594.045 3253.205 1594.215 3254.055 ;
        RECT 1559.085 3252.865 1559.715 3253.035 ;
        RECT 1641.885 3252.865 1642.055 3254.055 ;
        RECT 1690.645 3253.205 1690.815 3254.055 ;
        RECT 1655.685 3252.865 1656.315 3253.035 ;
        RECT 1738.485 3252.865 1738.655 3254.055 ;
        RECT 1787.245 3253.205 1787.415 3254.055 ;
        RECT 1752.285 3252.865 1752.915 3253.035 ;
        RECT 1835.085 3252.865 1835.255 3254.055 ;
        RECT 1849.345 3252.865 1849.975 3253.035 ;
        RECT 1462.485 3252.185 1463.115 3252.355 ;
      LAYER li1 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER li1 ;
        RECT 2028.745 3250.825 2028.915 3252.695 ;
        RECT 2125.345 3251.505 2125.515 3253.375 ;
        RECT 2173.645 3253.205 2173.815 3254.055 ;
        RECT 2221.485 3252.865 2221.655 3254.055 ;
        RECT 2270.245 3253.205 2270.415 3254.055 ;
        RECT 2235.285 3252.865 2235.915 3253.035 ;
        RECT 2318.085 3252.865 2318.255 3254.055 ;
        RECT 2366.845 3253.205 2367.015 3254.055 ;
        RECT 2331.885 3252.865 2332.515 3253.035 ;
        RECT 2414.685 3252.865 2414.855 3254.055 ;
        RECT 2463.445 3253.205 2463.615 3254.055 ;
        RECT 2428.485 3252.865 2429.115 3253.035 ;
        RECT 2511.285 3252.865 2511.455 3254.055 ;
        RECT 2525.545 3252.865 2526.175 3253.035 ;
      LAYER li1 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER li1 ;
        RECT 509.825 2793.525 514.595 2793.695 ;
        RECT 469.345 2789.445 469.515 2792.335 ;
        RECT 486.365 2789.615 486.535 2793.355 ;
        RECT 485.445 2789.445 486.535 2789.615 ;
        RECT 498.785 2789.445 498.955 2793.355 ;
        RECT 509.825 2793.185 509.995 2793.525 ;
        RECT 499.245 2789.445 499.415 2793.015 ;
        RECT 1042.965 2789.445 1043.135 2791.995 ;
        RECT 1111.045 2789.445 1111.215 2790.635 ;
        RECT 1158.885 2789.445 1159.055 2790.295 ;
        RECT 469.805 2789.105 474.575 2789.275 ;
        RECT 474.405 2788.425 474.575 2789.105 ;
        RECT 491.425 2788.425 491.595 2789.275 ;
        RECT 531.445 2787.405 531.615 2789.275 ;
        RECT 579.285 2787.405 579.455 2788.935 ;
        RECT 627.125 2787.405 627.295 2789.275 ;
        RECT 1628.545 2789.105 1628.715 2791.995 ;
        RECT 641.385 2787.745 642.015 2787.915 ;
        RECT 628.045 2784.345 628.215 2787.575 ;
        RECT 727.405 2712.265 727.575 2718.555 ;
        RECT 761.905 2711.925 762.075 2717.875 ;
        RECT 762.365 2712.605 762.535 2718.555 ;
        RECT 1083.905 2714.645 1084.075 2716.175 ;
      LAYER li1 ;
        RECT 305.520 1610.795 1395.115 2688.085 ;
      LAYER li1 ;
        RECT 1408.205 2069.325 1408.375 2106.895 ;
        RECT 1410.505 2088.025 1410.675 2157.895 ;
        RECT 1869.585 2063.545 1869.755 2065.075 ;
        RECT 1879.705 2064.565 1879.875 2067.455 ;
        RECT 1887.065 2064.905 1887.235 2066.095 ;
        RECT 1887.525 2063.715 1887.695 2066.095 ;
        RECT 1893.045 2065.585 1893.215 2067.115 ;
        RECT 1894.425 2066.095 1894.595 2067.115 ;
        RECT 1893.505 2065.925 1894.595 2066.095 ;
        RECT 1906.845 2064.905 1907.015 2068.135 ;
        RECT 1886.605 2063.545 1887.695 2063.715 ;
        RECT 1921.105 2062.865 1921.275 2064.735 ;
        RECT 1921.565 2063.545 1921.735 2066.775 ;
        RECT 1922.025 2063.545 1922.195 2067.115 ;
        RECT 1922.485 2065.585 1922.655 2069.155 ;
        RECT 1922.945 2068.985 1923.115 2070.175 ;
        RECT 1932.605 2067.965 1932.775 2069.155 ;
        RECT 1922.945 2065.245 1923.115 2067.115 ;
        RECT 1939.505 2063.205 1939.675 2065.075 ;
        RECT 1939.965 2063.205 1940.135 2068.135 ;
        RECT 1410.965 1931.965 1411.135 1980.075 ;
        RECT 1411.425 1835.745 1411.595 1849.515 ;
        RECT 1410.505 1787.125 1410.675 1834.555 ;
        RECT 1411.885 1642.285 1412.055 1690.395 ;
      LAYER li1 ;
        RECT 1705.000 1605.000 2081.480 2051.235 ;
        RECT 2255.000 1605.000 2631.480 2051.235 ;
        RECT 1555.520 410.795 2645.115 1488.085 ;
      LAYER mcon ;
        RECT 1304.245 3266.805 1304.415 3266.975 ;
        RECT 1594.045 3253.885 1594.215 3254.055 ;
        RECT 1400.845 3253.205 1401.015 3253.375 ;
        RECT 966.145 3252.525 966.315 3252.695 ;
        RECT 1013.985 3252.525 1014.155 3252.695 ;
        RECT 1062.745 3252.525 1062.915 3252.695 ;
        RECT 1110.585 3252.525 1110.755 3252.695 ;
        RECT 1159.345 3252.525 1159.515 3252.695 ;
        RECT 1207.185 3252.525 1207.355 3252.695 ;
        RECT 1255.945 3252.525 1256.115 3252.695 ;
        RECT 1303.785 3252.525 1303.955 3252.695 ;
        RECT 1448.685 3253.205 1448.855 3253.375 ;
        RECT 1641.885 3253.885 1642.055 3254.055 ;
        RECT 1690.645 3253.885 1690.815 3254.055 ;
        RECT 1738.485 3253.885 1738.655 3254.055 ;
        RECT 1787.245 3253.885 1787.415 3254.055 ;
        RECT 1835.085 3253.885 1835.255 3254.055 ;
        RECT 2173.645 3253.885 2173.815 3254.055 ;
        RECT 2125.345 3253.205 2125.515 3253.375 ;
        RECT 2221.485 3253.885 2221.655 3254.055 ;
        RECT 1559.545 3252.865 1559.715 3253.035 ;
        RECT 1656.145 3252.865 1656.315 3253.035 ;
        RECT 1752.745 3252.865 1752.915 3253.035 ;
        RECT 1849.805 3252.865 1849.975 3253.035 ;
        RECT 2028.745 3252.525 2028.915 3252.695 ;
        RECT 1366.345 3252.185 1366.515 3252.355 ;
        RECT 1462.945 3252.185 1463.115 3252.355 ;
        RECT 2270.245 3253.885 2270.415 3254.055 ;
        RECT 2318.085 3253.885 2318.255 3254.055 ;
        RECT 2366.845 3253.885 2367.015 3254.055 ;
        RECT 2414.685 3253.885 2414.855 3254.055 ;
        RECT 2463.445 3253.885 2463.615 3254.055 ;
        RECT 2511.285 3253.885 2511.455 3254.055 ;
        RECT 2235.745 3252.865 2235.915 3253.035 ;
        RECT 2332.345 3252.865 2332.515 3253.035 ;
        RECT 2428.945 3252.865 2429.115 3253.035 ;
        RECT 2526.005 3252.865 2526.175 3253.035 ;
        RECT 514.425 2793.525 514.595 2793.695 ;
        RECT 486.365 2793.185 486.535 2793.355 ;
        RECT 469.345 2792.165 469.515 2792.335 ;
        RECT 498.785 2793.185 498.955 2793.355 ;
        RECT 499.245 2792.845 499.415 2793.015 ;
        RECT 1042.965 2791.825 1043.135 2791.995 ;
        RECT 1628.545 2791.825 1628.715 2791.995 ;
        RECT 1111.045 2790.465 1111.215 2790.635 ;
        RECT 1158.885 2790.125 1159.055 2790.295 ;
        RECT 491.425 2789.105 491.595 2789.275 ;
        RECT 531.445 2789.105 531.615 2789.275 ;
        RECT 627.125 2789.105 627.295 2789.275 ;
        RECT 579.285 2788.765 579.455 2788.935 ;
        RECT 641.845 2787.745 642.015 2787.915 ;
        RECT 628.045 2787.405 628.215 2787.575 ;
        RECT 727.405 2718.385 727.575 2718.555 ;
        RECT 762.365 2718.385 762.535 2718.555 ;
        RECT 761.905 2717.705 762.075 2717.875 ;
        RECT 1083.905 2716.005 1084.075 2716.175 ;
        RECT 1410.505 2157.725 1410.675 2157.895 ;
        RECT 1408.205 2106.725 1408.375 2106.895 ;
        RECT 1922.945 2070.005 1923.115 2070.175 ;
        RECT 1922.485 2068.985 1922.655 2069.155 ;
        RECT 1932.605 2068.985 1932.775 2069.155 ;
        RECT 1906.845 2067.965 1907.015 2068.135 ;
        RECT 1879.705 2067.285 1879.875 2067.455 ;
        RECT 1869.585 2064.905 1869.755 2065.075 ;
        RECT 1893.045 2066.945 1893.215 2067.115 ;
        RECT 1887.065 2065.925 1887.235 2066.095 ;
        RECT 1887.525 2065.925 1887.695 2066.095 ;
        RECT 1894.425 2066.945 1894.595 2067.115 ;
        RECT 1922.025 2066.945 1922.195 2067.115 ;
        RECT 1921.565 2066.605 1921.735 2066.775 ;
        RECT 1921.105 2064.565 1921.275 2064.735 ;
        RECT 1939.965 2067.965 1940.135 2068.135 ;
        RECT 1922.945 2066.945 1923.115 2067.115 ;
        RECT 1939.505 2064.905 1939.675 2065.075 ;
        RECT 1410.965 1979.905 1411.135 1980.075 ;
        RECT 1411.425 1849.345 1411.595 1849.515 ;
        RECT 1410.505 1834.385 1410.675 1834.555 ;
        RECT 1411.885 1690.225 1412.055 1690.395 ;
      LAYER met1 ;
        RECT 1304.185 3266.960 1304.475 3267.005 ;
        RECT 1317.970 3266.960 1318.290 3267.020 ;
        RECT 1890.670 3266.960 1890.990 3267.020 ;
        RECT 1304.185 3266.820 1890.990 3266.960 ;
        RECT 1304.185 3266.775 1304.475 3266.820 ;
        RECT 1317.970 3266.760 1318.290 3266.820 ;
        RECT 1890.670 3266.760 1890.990 3266.820 ;
        RECT 1917.810 3266.960 1918.130 3267.020 ;
        RECT 2542.030 3266.960 2542.350 3267.020 ;
        RECT 1917.810 3266.820 2542.350 3266.960 ;
        RECT 1917.810 3266.760 1918.130 3266.820 ;
        RECT 2542.030 3266.760 2542.350 3266.820 ;
        RECT 1890.670 3264.580 1890.990 3264.640 ;
        RECT 1917.810 3264.580 1918.130 3264.640 ;
        RECT 1890.670 3264.440 1918.130 3264.580 ;
        RECT 1890.670 3264.380 1890.990 3264.440 ;
        RECT 1917.810 3264.380 1918.130 3264.440 ;
        RECT 696.970 3264.240 697.290 3264.300 ;
        RECT 2542.030 3264.240 2542.350 3264.300 ;
        RECT 2566.870 3264.240 2567.190 3264.300 ;
        RECT 688.320 3264.100 698.580 3264.240 ;
        RECT 675.810 3263.900 676.130 3263.960 ;
        RECT 688.320 3263.900 688.460 3264.100 ;
        RECT 696.970 3264.040 697.290 3264.100 ;
        RECT 675.810 3263.760 688.460 3263.900 ;
        RECT 698.440 3263.900 698.580 3264.100 ;
        RECT 2542.030 3264.100 2567.190 3264.240 ;
        RECT 2542.030 3264.040 2542.350 3264.100 ;
        RECT 2566.870 3264.040 2567.190 3264.100 ;
        RECT 1292.670 3263.900 1292.990 3263.960 ;
        RECT 1304.185 3263.900 1304.475 3263.945 ;
        RECT 698.440 3263.760 1304.475 3263.900 ;
        RECT 2566.960 3263.900 2567.100 3264.040 ;
        RECT 2594.470 3263.900 2594.790 3263.960 ;
        RECT 2566.960 3263.760 2594.790 3263.900 ;
        RECT 675.810 3263.700 676.130 3263.760 ;
        RECT 1292.670 3263.700 1292.990 3263.760 ;
        RECT 1304.185 3263.715 1304.475 3263.760 ;
        RECT 2594.470 3263.700 2594.790 3263.760 ;
        RECT 1593.985 3254.040 1594.275 3254.085 ;
        RECT 1641.825 3254.040 1642.115 3254.085 ;
        RECT 1593.985 3253.900 1642.115 3254.040 ;
        RECT 1593.985 3253.855 1594.275 3253.900 ;
        RECT 1641.825 3253.855 1642.115 3253.900 ;
        RECT 1690.585 3254.040 1690.875 3254.085 ;
        RECT 1738.425 3254.040 1738.715 3254.085 ;
        RECT 1690.585 3253.900 1738.715 3254.040 ;
        RECT 1690.585 3253.855 1690.875 3253.900 ;
        RECT 1738.425 3253.855 1738.715 3253.900 ;
        RECT 1787.185 3254.040 1787.475 3254.085 ;
        RECT 1835.025 3254.040 1835.315 3254.085 ;
        RECT 1787.185 3253.900 1835.315 3254.040 ;
        RECT 1787.185 3253.855 1787.475 3253.900 ;
        RECT 1835.025 3253.855 1835.315 3253.900 ;
        RECT 2173.585 3254.040 2173.875 3254.085 ;
        RECT 2221.425 3254.040 2221.715 3254.085 ;
        RECT 2173.585 3253.900 2221.715 3254.040 ;
        RECT 2173.585 3253.855 2173.875 3253.900 ;
        RECT 2221.425 3253.855 2221.715 3253.900 ;
        RECT 2270.185 3254.040 2270.475 3254.085 ;
        RECT 2318.025 3254.040 2318.315 3254.085 ;
        RECT 2270.185 3253.900 2318.315 3254.040 ;
        RECT 2270.185 3253.855 2270.475 3253.900 ;
        RECT 2318.025 3253.855 2318.315 3253.900 ;
        RECT 2366.785 3254.040 2367.075 3254.085 ;
        RECT 2414.625 3254.040 2414.915 3254.085 ;
        RECT 2366.785 3253.900 2414.915 3254.040 ;
        RECT 2366.785 3253.855 2367.075 3253.900 ;
        RECT 2414.625 3253.855 2414.915 3253.900 ;
        RECT 2463.385 3254.040 2463.675 3254.085 ;
        RECT 2511.225 3254.040 2511.515 3254.085 ;
        RECT 2463.385 3253.900 2511.515 3254.040 ;
        RECT 2463.385 3253.855 2463.675 3253.900 ;
        RECT 2511.225 3253.855 2511.515 3253.900 ;
        RECT 1400.785 3253.360 1401.075 3253.405 ;
        RECT 1448.625 3253.360 1448.915 3253.405 ;
        RECT 1593.985 3253.360 1594.275 3253.405 ;
        RECT 1690.585 3253.360 1690.875 3253.405 ;
        RECT 1787.185 3253.360 1787.475 3253.405 ;
        RECT 1400.785 3253.220 1448.915 3253.360 ;
        RECT 1400.785 3253.175 1401.075 3253.220 ;
        RECT 1448.625 3253.175 1448.915 3253.220 ;
        RECT 1565.540 3253.220 1594.275 3253.360 ;
        RECT 1559.025 3253.020 1559.315 3253.065 ;
        RECT 1510.800 3252.880 1559.315 3253.020 ;
        RECT 966.085 3252.680 966.375 3252.725 ;
        RECT 1013.925 3252.680 1014.215 3252.725 ;
        RECT 966.085 3252.540 1014.215 3252.680 ;
        RECT 966.085 3252.495 966.375 3252.540 ;
        RECT 1013.925 3252.495 1014.215 3252.540 ;
        RECT 1062.685 3252.680 1062.975 3252.725 ;
        RECT 1110.525 3252.680 1110.815 3252.725 ;
        RECT 1062.685 3252.540 1110.815 3252.680 ;
        RECT 1062.685 3252.495 1062.975 3252.540 ;
        RECT 1110.525 3252.495 1110.815 3252.540 ;
        RECT 1159.285 3252.680 1159.575 3252.725 ;
        RECT 1207.125 3252.680 1207.415 3252.725 ;
        RECT 1159.285 3252.540 1207.415 3252.680 ;
        RECT 1159.285 3252.495 1159.575 3252.540 ;
        RECT 1207.125 3252.495 1207.415 3252.540 ;
        RECT 1255.885 3252.680 1256.175 3252.725 ;
        RECT 1303.725 3252.680 1304.015 3252.725 ;
        RECT 1400.785 3252.680 1401.075 3252.725 ;
        RECT 1510.800 3252.680 1510.940 3252.880 ;
        RECT 1559.025 3252.835 1559.315 3252.880 ;
        RECT 1559.485 3253.020 1559.775 3253.065 ;
        RECT 1565.540 3253.020 1565.680 3253.220 ;
        RECT 1593.985 3253.175 1594.275 3253.220 ;
        RECT 1662.140 3253.220 1690.875 3253.360 ;
        RECT 1559.485 3252.880 1565.680 3253.020 ;
        RECT 1641.825 3253.020 1642.115 3253.065 ;
        RECT 1655.625 3253.020 1655.915 3253.065 ;
        RECT 1641.825 3252.880 1655.915 3253.020 ;
        RECT 1559.485 3252.835 1559.775 3252.880 ;
        RECT 1641.825 3252.835 1642.115 3252.880 ;
        RECT 1655.625 3252.835 1655.915 3252.880 ;
        RECT 1656.085 3253.020 1656.375 3253.065 ;
        RECT 1662.140 3253.020 1662.280 3253.220 ;
        RECT 1690.585 3253.175 1690.875 3253.220 ;
        RECT 1758.740 3253.220 1787.475 3253.360 ;
        RECT 1656.085 3252.880 1662.280 3253.020 ;
        RECT 1738.425 3253.020 1738.715 3253.065 ;
        RECT 1752.225 3253.020 1752.515 3253.065 ;
        RECT 1738.425 3252.880 1752.515 3253.020 ;
        RECT 1656.085 3252.835 1656.375 3252.880 ;
        RECT 1738.425 3252.835 1738.715 3252.880 ;
        RECT 1752.225 3252.835 1752.515 3252.880 ;
        RECT 1752.685 3253.020 1752.975 3253.065 ;
        RECT 1758.740 3253.020 1758.880 3253.220 ;
        RECT 1787.185 3253.175 1787.475 3253.220 ;
        RECT 2125.285 3253.360 2125.575 3253.405 ;
        RECT 2173.585 3253.360 2173.875 3253.405 ;
        RECT 2270.185 3253.360 2270.475 3253.405 ;
        RECT 2366.785 3253.360 2367.075 3253.405 ;
        RECT 2463.385 3253.360 2463.675 3253.405 ;
        RECT 2125.285 3253.220 2173.875 3253.360 ;
        RECT 2125.285 3253.175 2125.575 3253.220 ;
        RECT 2173.585 3253.175 2173.875 3253.220 ;
        RECT 2241.740 3253.220 2270.475 3253.360 ;
        RECT 1752.685 3252.880 1758.880 3253.020 ;
        RECT 1835.025 3253.020 1835.315 3253.065 ;
        RECT 1849.285 3253.020 1849.575 3253.065 ;
        RECT 1835.025 3252.880 1849.575 3253.020 ;
        RECT 1752.685 3252.835 1752.975 3252.880 ;
        RECT 1835.025 3252.835 1835.315 3252.880 ;
        RECT 1849.285 3252.835 1849.575 3252.880 ;
        RECT 1849.745 3253.020 1850.035 3253.065 ;
        RECT 2221.425 3253.020 2221.715 3253.065 ;
        RECT 2235.225 3253.020 2235.515 3253.065 ;
        RECT 1849.745 3252.880 1883.540 3253.020 ;
        RECT 1849.745 3252.835 1850.035 3252.880 ;
        RECT 1255.885 3252.540 1304.015 3252.680 ;
        RECT 1255.885 3252.495 1256.175 3252.540 ;
        RECT 1303.725 3252.495 1304.015 3252.540 ;
        RECT 1372.340 3252.540 1401.075 3252.680 ;
        RECT 1333.150 3252.340 1333.470 3252.400 ;
        RECT 1365.825 3252.340 1366.115 3252.385 ;
        RECT 1317.600 3252.200 1366.115 3252.340 ;
        RECT 1013.925 3251.815 1014.215 3252.045 ;
        RECT 1110.525 3251.815 1110.815 3252.045 ;
        RECT 1207.125 3251.815 1207.415 3252.045 ;
        RECT 1303.725 3252.000 1304.015 3252.045 ;
        RECT 1317.600 3252.000 1317.740 3252.200 ;
        RECT 1333.150 3252.140 1333.470 3252.200 ;
        RECT 1365.825 3252.155 1366.115 3252.200 ;
        RECT 1366.285 3252.340 1366.575 3252.385 ;
        RECT 1372.340 3252.340 1372.480 3252.540 ;
        RECT 1400.785 3252.495 1401.075 3252.540 ;
        RECT 1468.940 3252.540 1510.940 3252.680 ;
        RECT 1883.400 3252.680 1883.540 3252.880 ;
        RECT 2221.425 3252.880 2235.515 3253.020 ;
        RECT 2221.425 3252.835 2221.715 3252.880 ;
        RECT 2235.225 3252.835 2235.515 3252.880 ;
        RECT 2235.685 3253.020 2235.975 3253.065 ;
        RECT 2241.740 3253.020 2241.880 3253.220 ;
        RECT 2270.185 3253.175 2270.475 3253.220 ;
        RECT 2338.340 3253.220 2367.075 3253.360 ;
        RECT 2235.685 3252.880 2241.880 3253.020 ;
        RECT 2318.025 3253.020 2318.315 3253.065 ;
        RECT 2331.825 3253.020 2332.115 3253.065 ;
        RECT 2318.025 3252.880 2332.115 3253.020 ;
        RECT 2235.685 3252.835 2235.975 3252.880 ;
        RECT 2318.025 3252.835 2318.315 3252.880 ;
        RECT 2331.825 3252.835 2332.115 3252.880 ;
        RECT 2332.285 3253.020 2332.575 3253.065 ;
        RECT 2338.340 3253.020 2338.480 3253.220 ;
        RECT 2366.785 3253.175 2367.075 3253.220 ;
        RECT 2434.940 3253.220 2463.675 3253.360 ;
        RECT 2332.285 3252.880 2338.480 3253.020 ;
        RECT 2414.625 3253.020 2414.915 3253.065 ;
        RECT 2428.425 3253.020 2428.715 3253.065 ;
        RECT 2414.625 3252.880 2428.715 3253.020 ;
        RECT 2332.285 3252.835 2332.575 3252.880 ;
        RECT 2414.625 3252.835 2414.915 3252.880 ;
        RECT 2428.425 3252.835 2428.715 3252.880 ;
        RECT 2428.885 3253.020 2429.175 3253.065 ;
        RECT 2434.940 3253.020 2435.080 3253.220 ;
        RECT 2463.385 3253.175 2463.675 3253.220 ;
        RECT 2428.885 3252.880 2435.080 3253.020 ;
        RECT 2511.225 3253.020 2511.515 3253.065 ;
        RECT 2525.485 3253.020 2525.775 3253.065 ;
        RECT 2511.225 3252.880 2525.775 3253.020 ;
        RECT 2428.885 3252.835 2429.175 3252.880 ;
        RECT 2511.225 3252.835 2511.515 3252.880 ;
        RECT 2525.485 3252.835 2525.775 3252.880 ;
        RECT 2525.945 3253.020 2526.235 3253.065 ;
        RECT 2525.945 3252.880 2559.740 3253.020 ;
        RECT 2525.945 3252.835 2526.235 3252.880 ;
        RECT 2028.685 3252.680 2028.975 3252.725 ;
        RECT 2038.790 3252.680 2039.110 3252.740 ;
        RECT 2559.600 3252.680 2559.740 3252.880 ;
        RECT 1883.400 3252.540 1897.340 3252.680 ;
        RECT 1366.285 3252.200 1372.480 3252.340 ;
        RECT 1448.625 3252.340 1448.915 3252.385 ;
        RECT 1462.425 3252.340 1462.715 3252.385 ;
        RECT 1448.625 3252.200 1462.715 3252.340 ;
        RECT 1366.285 3252.155 1366.575 3252.200 ;
        RECT 1448.625 3252.155 1448.915 3252.200 ;
        RECT 1462.425 3252.155 1462.715 3252.200 ;
        RECT 1462.885 3252.340 1463.175 3252.385 ;
        RECT 1468.940 3252.340 1469.080 3252.540 ;
        RECT 1462.885 3252.200 1469.080 3252.340 ;
        RECT 1897.200 3252.340 1897.340 3252.540 ;
        RECT 2028.685 3252.540 2081.340 3252.680 ;
        RECT 2559.600 3252.540 2573.540 3252.680 ;
        RECT 2028.685 3252.495 2028.975 3252.540 ;
        RECT 2038.790 3252.480 2039.110 3252.540 ;
        RECT 1935.750 3252.340 1936.070 3252.400 ;
        RECT 1897.200 3252.200 1936.070 3252.340 ;
        RECT 1462.885 3252.155 1463.175 3252.200 ;
        RECT 1935.750 3252.140 1936.070 3252.200 ;
        RECT 1303.725 3251.860 1317.740 3252.000 ;
        RECT 1303.725 3251.815 1304.015 3251.860 ;
        RECT 966.085 3251.660 966.375 3251.705 ;
        RECT 724.200 3251.520 773.100 3251.660 ;
        RECT 688.230 3251.320 688.550 3251.380 ;
        RECT 724.200 3251.320 724.340 3251.520 ;
      LAYER met1 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met1 ;
        RECT 688.230 3251.180 724.340 3251.320 ;
        RECT 772.960 3251.320 773.100 3251.520 ;
        RECT 820.800 3251.520 869.700 3251.660 ;
        RECT 820.800 3251.320 820.940 3251.520 ;
        RECT 772.960 3251.180 820.940 3251.320 ;
        RECT 869.560 3251.320 869.700 3251.520 ;
        RECT 917.400 3251.520 966.375 3251.660 ;
        RECT 1014.000 3251.660 1014.140 3251.815 ;
        RECT 1062.685 3251.660 1062.975 3251.705 ;
        RECT 1014.000 3251.520 1062.975 3251.660 ;
        RECT 1110.600 3251.660 1110.740 3251.815 ;
        RECT 1159.285 3251.660 1159.575 3251.705 ;
        RECT 1110.600 3251.520 1159.575 3251.660 ;
        RECT 1207.200 3251.660 1207.340 3251.815 ;
        RECT 1255.885 3251.660 1256.175 3251.705 ;
        RECT 1207.200 3251.520 1256.175 3251.660 ;
        RECT 2081.200 3251.660 2081.340 3252.540 ;
        RECT 2573.400 3252.340 2573.540 3252.540 ;
        RECT 2582.050 3252.340 2582.370 3252.400 ;
        RECT 2573.400 3252.200 2582.370 3252.340 ;
        RECT 2582.050 3252.140 2582.370 3252.200 ;
        RECT 2125.285 3251.660 2125.575 3251.705 ;
        RECT 2081.200 3251.520 2125.575 3251.660 ;
        RECT 917.400 3251.320 917.540 3251.520 ;
        RECT 966.085 3251.475 966.375 3251.520 ;
        RECT 1062.685 3251.475 1062.975 3251.520 ;
        RECT 1159.285 3251.475 1159.575 3251.520 ;
        RECT 1255.885 3251.475 1256.175 3251.520 ;
        RECT 2125.285 3251.475 2125.575 3251.520 ;
        RECT 869.560 3251.180 917.540 3251.320 ;
        RECT 688.230 3251.120 688.550 3251.180 ;
      LAYER met1 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met1 ;
        RECT 1459.190 3229.560 1459.510 3229.620 ;
        RECT 1536.930 3229.560 1537.250 3229.620 ;
        RECT 1459.190 3229.420 1537.250 3229.560 ;
        RECT 1459.190 3229.360 1459.510 3229.420 ;
        RECT 1536.930 3229.360 1537.250 3229.420 ;
        RECT 1452.290 3222.420 1452.610 3222.480 ;
        RECT 1535.550 3222.420 1535.870 3222.480 ;
        RECT 1452.290 3222.280 1535.870 3222.420 ;
        RECT 1452.290 3222.220 1452.610 3222.280 ;
        RECT 1535.550 3222.220 1535.870 3222.280 ;
        RECT 1438.490 3215.620 1438.810 3215.680 ;
        RECT 1535.550 3215.620 1535.870 3215.680 ;
        RECT 1438.490 3215.480 1535.870 3215.620 ;
        RECT 1438.490 3215.420 1438.810 3215.480 ;
        RECT 1535.550 3215.420 1535.870 3215.480 ;
        RECT 1431.590 3208.820 1431.910 3208.880 ;
        RECT 1538.310 3208.820 1538.630 3208.880 ;
        RECT 1431.590 3208.680 1538.630 3208.820 ;
        RECT 1431.590 3208.620 1431.910 3208.680 ;
        RECT 1538.310 3208.620 1538.630 3208.680 ;
        RECT 1424.690 3201.680 1425.010 3201.740 ;
        RECT 1538.310 3201.680 1538.630 3201.740 ;
        RECT 1424.690 3201.540 1538.630 3201.680 ;
        RECT 1424.690 3201.480 1425.010 3201.540 ;
        RECT 1538.310 3201.480 1538.630 3201.540 ;
        RECT 1459.650 3188.080 1459.970 3188.140 ;
        RECT 1534.170 3188.080 1534.490 3188.140 ;
        RECT 1459.650 3187.940 1534.490 3188.080 ;
        RECT 1459.650 3187.880 1459.970 3187.940 ;
        RECT 1534.170 3187.880 1534.490 3187.940 ;
        RECT 1352.010 2901.460 1352.330 2901.520 ;
        RECT 1395.710 2901.460 1396.030 2901.520 ;
        RECT 1352.010 2901.320 1396.030 2901.460 ;
        RECT 1352.010 2901.260 1352.330 2901.320 ;
        RECT 1395.710 2901.260 1396.030 2901.320 ;
        RECT 1514.390 2898.400 1514.710 2898.460 ;
        RECT 1538.310 2898.400 1538.630 2898.460 ;
        RECT 1514.390 2898.260 1538.630 2898.400 ;
        RECT 1514.390 2898.200 1514.710 2898.260 ;
        RECT 1538.310 2898.200 1538.630 2898.260 ;
      LAYER met1 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met1 ;
        RECT 1945.870 3250.980 1946.190 3251.040 ;
        RECT 2028.685 3250.980 2028.975 3251.025 ;
        RECT 1945.870 3250.840 2028.975 3250.980 ;
        RECT 1945.870 3250.780 1946.190 3250.840 ;
        RECT 2028.685 3250.795 2028.975 3250.840 ;
      LAYER met1 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met1 ;
        RECT 386.930 2794.360 387.250 2794.420 ;
        RECT 431.550 2794.360 431.870 2794.420 ;
        RECT 433.390 2794.360 433.710 2794.420 ;
        RECT 386.930 2794.220 433.710 2794.360 ;
        RECT 386.930 2794.160 387.250 2794.220 ;
        RECT 431.550 2794.160 431.870 2794.220 ;
        RECT 433.390 2794.160 433.710 2794.220 ;
        RECT 468.810 2794.360 469.130 2794.420 ;
        RECT 686.390 2794.360 686.710 2794.420 ;
        RECT 468.810 2794.220 686.710 2794.360 ;
        RECT 468.810 2794.160 469.130 2794.220 ;
        RECT 686.390 2794.160 686.710 2794.220 ;
        RECT 1738.410 2794.360 1738.730 2794.420 ;
        RECT 1780.270 2794.360 1780.590 2794.420 ;
        RECT 1738.410 2794.220 1780.590 2794.360 ;
        RECT 1738.410 2794.160 1738.730 2794.220 ;
        RECT 1780.270 2794.160 1780.590 2794.220 ;
        RECT 2340.090 2794.360 2340.410 2794.420 ;
        RECT 2382.870 2794.360 2383.190 2794.420 ;
        RECT 2340.090 2794.220 2383.190 2794.360 ;
        RECT 2340.090 2794.160 2340.410 2794.220 ;
        RECT 2382.870 2794.160 2383.190 2794.220 ;
        RECT 330.810 2794.020 331.130 2794.080 ;
        RECT 1001.030 2794.020 1001.350 2794.080 ;
        RECT 330.810 2793.880 1001.350 2794.020 ;
        RECT 330.810 2793.820 331.130 2793.880 ;
        RECT 1001.030 2793.820 1001.350 2793.880 ;
        RECT 1076.470 2794.020 1076.790 2794.080 ;
        RECT 1122.470 2794.020 1122.790 2794.080 ;
        RECT 1076.470 2793.880 1122.790 2794.020 ;
        RECT 1076.470 2793.820 1076.790 2793.880 ;
        RECT 1122.470 2793.820 1122.790 2793.880 ;
        RECT 1432.050 2794.020 1432.370 2794.080 ;
        RECT 2268.330 2794.020 2268.650 2794.080 ;
        RECT 2287.190 2794.020 2287.510 2794.080 ;
        RECT 2332.730 2794.020 2333.050 2794.080 ;
        RECT 2377.350 2794.020 2377.670 2794.080 ;
        RECT 1432.050 2793.880 2276.840 2794.020 ;
        RECT 1432.050 2793.820 1432.370 2793.880 ;
        RECT 2268.330 2793.820 2268.650 2793.880 ;
        RECT 374.970 2793.680 375.290 2793.740 ;
        RECT 420.970 2793.680 421.290 2793.740 ;
        RECT 466.510 2793.680 466.830 2793.740 ;
        RECT 513.890 2793.680 514.210 2793.740 ;
        RECT 374.970 2793.540 514.210 2793.680 ;
        RECT 374.970 2793.480 375.290 2793.540 ;
        RECT 420.970 2793.480 421.290 2793.540 ;
        RECT 466.510 2793.480 466.830 2793.540 ;
        RECT 513.890 2793.480 514.210 2793.540 ;
        RECT 514.365 2793.680 514.655 2793.725 ;
        RECT 531.370 2793.680 531.690 2793.740 ;
        RECT 514.365 2793.540 531.690 2793.680 ;
        RECT 514.365 2793.495 514.655 2793.540 ;
        RECT 531.370 2793.480 531.690 2793.540 ;
        RECT 536.430 2793.680 536.750 2793.740 ;
        RECT 707.090 2793.680 707.410 2793.740 ;
        RECT 536.430 2793.540 707.410 2793.680 ;
        RECT 536.430 2793.480 536.750 2793.540 ;
        RECT 707.090 2793.480 707.410 2793.540 ;
        RECT 1093.950 2793.680 1094.270 2793.740 ;
        RECT 1139.950 2793.680 1140.270 2793.740 ;
        RECT 1186.870 2793.680 1187.190 2793.740 ;
        RECT 1093.950 2793.540 1187.190 2793.680 ;
        RECT 1093.950 2793.480 1094.270 2793.540 ;
        RECT 1139.950 2793.480 1140.270 2793.540 ;
        RECT 1186.870 2793.480 1187.190 2793.540 ;
        RECT 1432.510 2793.680 1432.830 2793.740 ;
        RECT 2273.850 2793.680 2274.170 2793.740 ;
        RECT 1432.510 2793.540 2274.170 2793.680 ;
        RECT 1432.510 2793.480 1432.830 2793.540 ;
        RECT 2273.850 2793.480 2274.170 2793.540 ;
        RECT 392.450 2793.340 392.770 2793.400 ;
        RECT 439.370 2793.340 439.690 2793.400 ;
        RECT 485.830 2793.340 486.150 2793.400 ;
        RECT 392.450 2793.200 486.150 2793.340 ;
        RECT 392.450 2793.140 392.770 2793.200 ;
        RECT 439.370 2793.140 439.690 2793.200 ;
        RECT 485.830 2793.140 486.150 2793.200 ;
        RECT 486.305 2793.340 486.595 2793.385 ;
        RECT 497.330 2793.340 497.650 2793.400 ;
        RECT 486.305 2793.200 497.650 2793.340 ;
        RECT 486.305 2793.155 486.595 2793.200 ;
        RECT 497.330 2793.140 497.650 2793.200 ;
        RECT 498.725 2793.340 499.015 2793.385 ;
        RECT 509.765 2793.340 510.055 2793.385 ;
        RECT 498.725 2793.200 510.055 2793.340 ;
        RECT 498.725 2793.155 499.015 2793.200 ;
        RECT 509.765 2793.155 510.055 2793.200 ;
        RECT 510.210 2793.340 510.530 2793.400 ;
        RECT 700.190 2793.340 700.510 2793.400 ;
        RECT 510.210 2793.200 700.510 2793.340 ;
        RECT 510.210 2793.140 510.530 2793.200 ;
        RECT 700.190 2793.140 700.510 2793.200 ;
        RECT 1110.970 2793.340 1111.290 2793.400 ;
        RECT 1159.270 2793.340 1159.590 2793.400 ;
        RECT 1110.970 2793.200 1159.590 2793.340 ;
        RECT 1110.970 2793.140 1111.290 2793.200 ;
        RECT 1159.270 2793.140 1159.590 2793.200 ;
        RECT 1631.690 2793.340 1632.010 2793.400 ;
        RECT 1677.230 2793.340 1677.550 2793.400 ;
        RECT 1721.390 2793.340 1721.710 2793.400 ;
        RECT 1766.470 2793.340 1766.790 2793.400 ;
        RECT 1631.690 2793.200 1766.790 2793.340 ;
        RECT 1631.690 2793.140 1632.010 2793.200 ;
        RECT 1677.230 2793.140 1677.550 2793.200 ;
        RECT 1721.390 2793.140 1721.710 2793.200 ;
        RECT 1766.470 2793.140 1766.790 2793.200 ;
        RECT 379.570 2793.000 379.890 2793.060 ;
        RECT 426.950 2793.000 427.270 2793.060 ;
        RECT 379.570 2792.860 427.270 2793.000 ;
        RECT 379.570 2792.800 379.890 2792.860 ;
        RECT 426.950 2792.800 427.270 2792.860 ;
        RECT 433.390 2793.000 433.710 2793.060 ;
        RECT 478.470 2793.000 478.790 2793.060 ;
        RECT 499.185 2793.000 499.475 2793.045 ;
        RECT 520.790 2793.000 521.110 2793.060 ;
        RECT 433.390 2792.860 499.475 2793.000 ;
        RECT 433.390 2792.800 433.710 2792.860 ;
        RECT 478.470 2792.800 478.790 2792.860 ;
        RECT 499.185 2792.815 499.475 2792.860 ;
        RECT 499.720 2792.860 521.110 2793.000 ;
        RECT 397.050 2792.660 397.370 2792.720 ;
        RECT 444.430 2792.660 444.750 2792.720 ;
        RECT 491.810 2792.660 492.130 2792.720 ;
        RECT 499.720 2792.660 499.860 2792.860 ;
        RECT 520.790 2792.800 521.110 2792.860 ;
        RECT 542.410 2793.000 542.730 2793.060 ;
        RECT 741.590 2793.000 741.910 2793.060 ;
        RECT 542.410 2792.860 741.910 2793.000 ;
        RECT 542.410 2792.800 542.730 2792.860 ;
        RECT 741.590 2792.800 741.910 2792.860 ;
        RECT 1087.510 2793.000 1087.830 2793.060 ;
        RECT 1129.370 2793.000 1129.690 2793.060 ;
        RECT 1173.070 2793.000 1173.390 2793.060 ;
        RECT 1087.510 2792.860 1173.390 2793.000 ;
        RECT 1087.510 2792.800 1087.830 2792.860 ;
        RECT 1129.370 2792.800 1129.690 2792.860 ;
        RECT 1173.070 2792.800 1173.390 2792.860 ;
        RECT 1680.450 2793.000 1680.770 2793.060 ;
        RECT 1683.210 2793.000 1683.530 2793.060 ;
        RECT 1730.130 2793.000 1730.450 2793.060 ;
        RECT 1773.370 2793.000 1773.690 2793.060 ;
        RECT 1680.450 2792.860 1773.690 2793.000 ;
        RECT 2276.700 2793.000 2276.840 2793.880 ;
        RECT 2287.190 2793.880 2388.620 2794.020 ;
        RECT 2287.190 2793.820 2287.510 2793.880 ;
        RECT 2332.730 2793.820 2333.050 2793.880 ;
        RECT 2377.350 2793.820 2377.670 2793.880 ;
        RECT 2294.090 2793.680 2294.410 2793.740 ;
        RECT 2340.090 2793.680 2340.410 2793.740 ;
        RECT 2294.090 2793.540 2340.410 2793.680 ;
        RECT 2294.090 2793.480 2294.410 2793.540 ;
        RECT 2340.090 2793.480 2340.410 2793.540 ;
        RECT 2340.550 2793.680 2340.870 2793.740 ;
        RECT 2343.770 2793.680 2344.090 2793.740 ;
        RECT 2387.930 2793.680 2388.250 2793.740 ;
        RECT 2340.550 2793.540 2388.250 2793.680 ;
        RECT 2340.550 2793.480 2340.870 2793.540 ;
        RECT 2343.770 2793.480 2344.090 2793.540 ;
        RECT 2387.930 2793.480 2388.250 2793.540 ;
        RECT 2280.290 2793.340 2280.610 2793.400 ;
        RECT 2326.290 2793.340 2326.610 2793.400 ;
        RECT 2374.130 2793.340 2374.450 2793.400 ;
        RECT 2280.290 2793.200 2374.450 2793.340 ;
        RECT 2388.480 2793.340 2388.620 2793.880 ;
        RECT 2421.970 2793.340 2422.290 2793.400 ;
        RECT 2388.480 2793.200 2422.290 2793.340 ;
        RECT 2280.290 2793.140 2280.610 2793.200 ;
        RECT 2326.290 2793.140 2326.610 2793.200 ;
        RECT 2374.130 2793.140 2374.450 2793.200 ;
        RECT 2421.970 2793.140 2422.290 2793.200 ;
        RECT 2315.250 2793.000 2315.570 2793.060 ;
        RECT 2360.790 2793.000 2361.110 2793.060 ;
        RECT 2408.170 2793.000 2408.490 2793.060 ;
        RECT 2276.700 2792.860 2408.490 2793.000 ;
        RECT 1680.450 2792.800 1680.770 2792.860 ;
        RECT 1683.210 2792.800 1683.530 2792.860 ;
        RECT 1730.130 2792.800 1730.450 2792.860 ;
        RECT 1773.370 2792.800 1773.690 2792.860 ;
        RECT 2315.250 2792.800 2315.570 2792.860 ;
        RECT 2360.790 2792.800 2361.110 2792.860 ;
        RECT 2408.170 2792.800 2408.490 2792.860 ;
        RECT 397.050 2792.520 492.130 2792.660 ;
        RECT 397.050 2792.460 397.370 2792.520 ;
        RECT 444.430 2792.460 444.750 2792.520 ;
        RECT 491.810 2792.460 492.130 2792.520 ;
        RECT 492.360 2792.520 499.860 2792.660 ;
        RECT 500.090 2792.660 500.410 2792.720 ;
        RECT 524.010 2792.660 524.330 2792.720 ;
        RECT 720.890 2792.660 721.210 2792.720 ;
        RECT 500.090 2792.520 521.480 2792.660 ;
        RECT 403.950 2792.320 404.270 2792.380 ;
        RECT 449.030 2792.320 449.350 2792.380 ;
        RECT 469.285 2792.320 469.575 2792.365 ;
        RECT 403.950 2792.180 469.575 2792.320 ;
        RECT 403.950 2792.120 404.270 2792.180 ;
        RECT 449.030 2792.120 449.350 2792.180 ;
        RECT 469.285 2792.135 469.575 2792.180 ;
        RECT 473.870 2792.320 474.190 2792.380 ;
        RECT 492.360 2792.320 492.500 2792.520 ;
        RECT 500.090 2792.460 500.410 2792.520 ;
        RECT 473.870 2792.180 492.500 2792.320 ;
        RECT 521.340 2792.320 521.480 2792.520 ;
        RECT 524.010 2792.520 721.210 2792.660 ;
        RECT 524.010 2792.460 524.330 2792.520 ;
        RECT 720.890 2792.460 721.210 2792.520 ;
        RECT 1042.430 2792.660 1042.750 2792.720 ;
        RECT 1087.970 2792.660 1088.290 2792.720 ;
        RECT 1135.810 2792.660 1136.130 2792.720 ;
        RECT 1179.970 2792.660 1180.290 2792.720 ;
        RECT 1042.430 2792.520 1180.290 2792.660 ;
        RECT 1042.430 2792.460 1042.750 2792.520 ;
        RECT 1087.970 2792.460 1088.290 2792.520 ;
        RECT 1135.810 2792.460 1136.130 2792.520 ;
        RECT 1179.970 2792.460 1180.290 2792.520 ;
        RECT 1652.390 2792.660 1652.710 2792.720 ;
        RECT 1699.310 2792.660 1699.630 2792.720 ;
        RECT 1748.530 2792.660 1748.850 2792.720 ;
        RECT 1790.850 2792.660 1791.170 2792.720 ;
        RECT 1652.390 2792.520 1791.170 2792.660 ;
        RECT 1652.390 2792.460 1652.710 2792.520 ;
        RECT 1699.310 2792.460 1699.630 2792.520 ;
        RECT 1748.530 2792.460 1748.850 2792.520 ;
        RECT 1790.850 2792.460 1791.170 2792.520 ;
        RECT 2266.490 2792.660 2266.810 2792.720 ;
        RECT 2308.350 2792.660 2308.670 2792.720 ;
        RECT 2356.650 2792.660 2356.970 2792.720 ;
        RECT 2401.730 2792.660 2402.050 2792.720 ;
        RECT 2266.490 2792.520 2402.050 2792.660 ;
        RECT 2266.490 2792.460 2266.810 2792.520 ;
        RECT 2308.350 2792.460 2308.670 2792.520 ;
        RECT 2356.650 2792.460 2356.970 2792.520 ;
        RECT 2401.730 2792.460 2402.050 2792.520 ;
        RECT 700.650 2792.320 700.970 2792.380 ;
        RECT 521.340 2792.180 700.970 2792.320 ;
        RECT 473.870 2792.120 474.190 2792.180 ;
        RECT 700.650 2792.120 700.970 2792.180 ;
        RECT 1065.890 2792.320 1066.210 2792.380 ;
        RECT 1110.970 2792.320 1111.290 2792.380 ;
        RECT 1065.890 2792.180 1111.290 2792.320 ;
        RECT 1065.890 2792.120 1066.210 2792.180 ;
        RECT 1110.970 2792.120 1111.290 2792.180 ;
        RECT 1646.410 2792.320 1646.730 2792.380 ;
        RECT 1695.170 2792.320 1695.490 2792.380 ;
        RECT 1741.170 2792.320 1741.490 2792.380 ;
        RECT 1787.170 2792.320 1787.490 2792.380 ;
        RECT 1646.410 2792.180 1787.490 2792.320 ;
        RECT 1646.410 2792.120 1646.730 2792.180 ;
        RECT 1695.170 2792.120 1695.490 2792.180 ;
        RECT 1741.170 2792.120 1741.490 2792.180 ;
        RECT 1787.170 2792.120 1787.490 2792.180 ;
        RECT 2273.850 2792.320 2274.170 2792.380 ;
        RECT 2321.230 2792.320 2321.550 2792.380 ;
        RECT 2367.230 2792.320 2367.550 2792.380 ;
        RECT 2415.070 2792.320 2415.390 2792.380 ;
        RECT 2273.850 2792.180 2415.390 2792.320 ;
        RECT 2273.850 2792.120 2274.170 2792.180 ;
        RECT 2321.230 2792.120 2321.550 2792.180 ;
        RECT 2367.230 2792.120 2367.550 2792.180 ;
        RECT 2415.070 2792.120 2415.390 2792.180 ;
        RECT 368.530 2791.980 368.850 2792.040 ;
        RECT 414.530 2791.980 414.850 2792.040 ;
        RECT 462.370 2791.980 462.690 2792.040 ;
        RECT 465.590 2791.980 465.910 2792.040 ;
        RECT 368.530 2791.840 465.910 2791.980 ;
        RECT 368.530 2791.780 368.850 2791.840 ;
        RECT 414.530 2791.780 414.850 2791.840 ;
        RECT 462.370 2791.780 462.690 2791.840 ;
        RECT 465.590 2791.780 465.910 2791.840 ;
        RECT 489.050 2791.980 489.370 2792.040 ;
        RECT 693.290 2791.980 693.610 2792.040 ;
        RECT 489.050 2791.840 693.610 2791.980 ;
        RECT 489.050 2791.780 489.370 2791.840 ;
        RECT 693.290 2791.780 693.610 2791.840 ;
        RECT 1042.905 2791.980 1043.195 2792.025 ;
        RECT 1053.010 2791.980 1053.330 2792.040 ;
        RECT 1100.390 2791.980 1100.710 2792.040 ;
        RECT 1147.310 2791.980 1147.630 2792.040 ;
        RECT 1628.485 2791.980 1628.775 2792.025 ;
        RECT 1670.330 2791.980 1670.650 2792.040 ;
        RECT 1676.310 2791.980 1676.630 2792.040 ;
        RECT 1042.905 2791.840 1166.860 2791.980 ;
        RECT 1042.905 2791.795 1043.195 2791.840 ;
        RECT 1053.010 2791.780 1053.330 2791.840 ;
        RECT 1100.390 2791.780 1100.710 2791.840 ;
        RECT 1147.310 2791.780 1147.630 2791.840 ;
        RECT 407.170 2791.640 407.490 2791.700 ;
        RECT 409.930 2791.640 410.250 2791.700 ;
        RECT 455.470 2791.640 455.790 2791.700 ;
        RECT 407.170 2791.500 455.790 2791.640 ;
        RECT 407.170 2791.440 407.490 2791.500 ;
        RECT 409.930 2791.440 410.250 2791.500 ;
        RECT 455.470 2791.440 455.790 2791.500 ;
        RECT 460.990 2791.640 461.310 2791.700 ;
        RECT 687.310 2791.640 687.630 2791.700 ;
        RECT 460.990 2791.500 687.630 2791.640 ;
        RECT 460.990 2791.440 461.310 2791.500 ;
        RECT 687.310 2791.440 687.630 2791.500 ;
        RECT 1055.770 2791.640 1056.090 2791.700 ;
        RECT 1058.990 2791.640 1059.310 2791.700 ;
        RECT 1105.450 2791.640 1105.770 2791.700 ;
        RECT 1152.370 2791.640 1152.690 2791.700 ;
        RECT 1055.770 2791.500 1152.690 2791.640 ;
        RECT 1055.770 2791.440 1056.090 2791.500 ;
        RECT 1058.990 2791.440 1059.310 2791.500 ;
        RECT 1105.450 2791.440 1105.770 2791.500 ;
        RECT 1152.370 2791.440 1152.690 2791.500 ;
        RECT 371.290 2791.300 371.610 2791.360 ;
        RECT 686.850 2791.300 687.170 2791.360 ;
        RECT 371.290 2791.160 687.170 2791.300 ;
        RECT 371.290 2791.100 371.610 2791.160 ;
        RECT 686.850 2791.100 687.170 2791.160 ;
        RECT 1034.610 2791.300 1034.930 2791.360 ;
        RECT 1076.470 2791.300 1076.790 2791.360 ;
        RECT 1034.610 2791.160 1076.790 2791.300 ;
        RECT 1034.610 2791.100 1034.930 2791.160 ;
        RECT 1076.470 2791.100 1076.790 2791.160 ;
        RECT 1122.470 2791.300 1122.790 2791.360 ;
        RECT 1166.170 2791.300 1166.490 2791.360 ;
        RECT 1122.470 2791.160 1166.490 2791.300 ;
        RECT 1166.720 2791.300 1166.860 2791.840 ;
        RECT 1628.485 2791.840 1676.630 2791.980 ;
        RECT 1628.485 2791.795 1628.775 2791.840 ;
        RECT 1670.330 2791.780 1670.650 2791.840 ;
        RECT 1676.310 2791.780 1676.630 2791.840 ;
        RECT 1687.810 2791.980 1688.130 2792.040 ;
        RECT 1738.410 2791.980 1738.730 2792.040 ;
        RECT 1687.810 2791.840 1738.730 2791.980 ;
        RECT 1687.810 2791.780 1688.130 2791.840 ;
        RECT 1738.410 2791.780 1738.730 2791.840 ;
        RECT 1762.790 2791.980 1763.110 2792.040 ;
        RECT 2381.030 2791.980 2381.350 2792.040 ;
        RECT 1762.790 2791.840 2381.350 2791.980 ;
        RECT 1762.790 2791.780 1763.110 2791.840 ;
        RECT 2381.030 2791.780 2381.350 2791.840 ;
        RECT 2382.870 2791.980 2383.190 2792.040 ;
        RECT 2428.870 2791.980 2429.190 2792.040 ;
        RECT 2382.870 2791.840 2429.190 2791.980 ;
        RECT 2382.870 2791.780 2383.190 2791.840 ;
        RECT 2428.870 2791.780 2429.190 2791.840 ;
        RECT 1665.730 2791.640 1666.050 2791.700 ;
        RECT 1712.650 2791.640 1712.970 2791.700 ;
        RECT 1742.090 2791.640 1742.410 2791.700 ;
        RECT 1657.080 2791.500 1742.410 2791.640 ;
        RECT 1193.770 2791.300 1194.090 2791.360 ;
        RECT 1166.720 2791.160 1194.090 2791.300 ;
        RECT 1122.470 2791.100 1122.790 2791.160 ;
        RECT 1166.170 2791.100 1166.490 2791.160 ;
        RECT 1193.770 2791.100 1194.090 2791.160 ;
        RECT 362.550 2790.960 362.870 2791.020 ;
        RECT 407.170 2790.960 407.490 2791.020 ;
        RECT 362.550 2790.820 407.490 2790.960 ;
        RECT 362.550 2790.760 362.870 2790.820 ;
        RECT 407.170 2790.760 407.490 2790.820 ;
        RECT 419.130 2790.960 419.450 2791.020 ;
        RECT 748.490 2790.960 748.810 2791.020 ;
        RECT 419.130 2790.820 748.810 2790.960 ;
        RECT 419.130 2790.760 419.450 2790.820 ;
        RECT 748.490 2790.760 748.810 2790.820 ;
        RECT 1018.970 2790.960 1019.290 2791.020 ;
        RECT 1065.890 2790.960 1066.210 2791.020 ;
        RECT 1018.970 2790.820 1066.210 2790.960 ;
        RECT 1018.970 2790.760 1019.290 2790.820 ;
        RECT 1065.890 2790.760 1066.210 2790.820 ;
        RECT 384.170 2790.620 384.490 2790.680 ;
        RECT 727.790 2790.620 728.110 2790.680 ;
        RECT 384.170 2790.480 728.110 2790.620 ;
        RECT 384.170 2790.420 384.490 2790.480 ;
        RECT 727.790 2790.420 728.110 2790.480 ;
        RECT 1076.010 2790.620 1076.330 2790.680 ;
        RECT 1110.985 2790.620 1111.275 2790.665 ;
        RECT 1076.010 2790.480 1111.275 2790.620 ;
        RECT 1076.010 2790.420 1076.330 2790.480 ;
        RECT 1110.985 2790.435 1111.275 2790.480 ;
        RECT 1425.610 2790.620 1425.930 2790.680 ;
        RECT 1642.270 2790.620 1642.590 2790.680 ;
        RECT 1425.610 2790.480 1642.590 2790.620 ;
        RECT 1425.610 2790.420 1425.930 2790.480 ;
        RECT 1642.270 2790.420 1642.590 2790.480 ;
        RECT 406.250 2790.280 406.570 2790.340 ;
        RECT 762.750 2790.280 763.070 2790.340 ;
        RECT 406.250 2790.140 763.070 2790.280 ;
        RECT 406.250 2790.080 406.570 2790.140 ;
        RECT 762.750 2790.080 763.070 2790.140 ;
        RECT 1158.825 2790.280 1159.115 2790.325 ;
        RECT 1159.270 2790.280 1159.590 2790.340 ;
        RECT 1158.825 2790.140 1159.590 2790.280 ;
        RECT 1158.825 2790.095 1159.115 2790.140 ;
        RECT 1159.270 2790.080 1159.590 2790.140 ;
        RECT 1562.690 2790.280 1563.010 2790.340 ;
        RECT 1614.670 2790.280 1614.990 2790.340 ;
        RECT 1562.690 2790.140 1614.990 2790.280 ;
        RECT 1562.690 2790.080 1563.010 2790.140 ;
        RECT 1614.670 2790.080 1614.990 2790.140 ;
        RECT 1617.890 2790.280 1618.210 2790.340 ;
        RECT 1657.080 2790.280 1657.220 2791.500 ;
        RECT 1665.730 2791.440 1666.050 2791.500 ;
        RECT 1712.650 2791.440 1712.970 2791.500 ;
        RECT 1742.090 2791.440 1742.410 2791.500 ;
        RECT 1763.250 2791.640 1763.570 2791.700 ;
        RECT 2387.470 2791.640 2387.790 2791.700 ;
        RECT 1763.250 2791.500 2387.790 2791.640 ;
        RECT 1763.250 2791.440 1763.570 2791.500 ;
        RECT 2387.470 2791.440 2387.790 2791.500 ;
        RECT 2387.930 2791.640 2388.250 2791.700 ;
        RECT 2435.770 2791.640 2436.090 2791.700 ;
        RECT 2387.930 2791.500 2436.090 2791.640 ;
        RECT 2387.930 2791.440 2388.250 2791.500 ;
        RECT 2435.770 2791.440 2436.090 2791.500 ;
        RECT 1658.830 2791.300 1659.150 2791.360 ;
        RECT 1706.210 2791.300 1706.530 2791.360 ;
        RECT 1752.670 2791.300 1752.990 2791.360 ;
        RECT 1617.890 2790.140 1657.220 2790.280 ;
        RECT 1657.540 2791.160 1752.990 2791.300 ;
        RECT 1617.890 2790.080 1618.210 2790.140 ;
        RECT 396.590 2789.940 396.910 2790.000 ;
        RECT 762.290 2789.940 762.610 2790.000 ;
        RECT 396.590 2789.800 762.610 2789.940 ;
        RECT 396.590 2789.740 396.910 2789.800 ;
        RECT 762.290 2789.740 762.610 2789.800 ;
        RECT 1548.890 2789.940 1549.210 2790.000 ;
        RECT 1607.770 2789.940 1608.090 2790.000 ;
        RECT 1548.890 2789.800 1608.090 2789.940 ;
        RECT 1548.890 2789.740 1549.210 2789.800 ;
        RECT 1607.770 2789.740 1608.090 2789.800 ;
        RECT 1610.990 2789.940 1611.310 2790.000 ;
        RECT 1657.540 2789.940 1657.680 2791.160 ;
        RECT 1658.830 2791.100 1659.150 2791.160 ;
        RECT 1706.210 2791.100 1706.530 2791.160 ;
        RECT 1752.670 2791.100 1752.990 2791.160 ;
        RECT 1769.690 2791.300 1770.010 2791.360 ;
        RECT 2394.370 2791.300 2394.690 2791.360 ;
        RECT 1769.690 2791.160 2394.690 2791.300 ;
        RECT 1769.690 2791.100 1770.010 2791.160 ;
        RECT 2394.370 2791.100 2394.690 2791.160 ;
        RECT 2394.830 2791.300 2395.150 2791.360 ;
        RECT 2442.670 2791.300 2442.990 2791.360 ;
        RECT 2394.830 2791.160 2442.990 2791.300 ;
        RECT 2394.830 2791.100 2395.150 2791.160 ;
        RECT 2442.670 2791.100 2442.990 2791.160 ;
        RECT 1676.310 2790.960 1676.630 2791.020 ;
        RECT 1718.170 2790.960 1718.490 2791.020 ;
        RECT 1760.030 2790.960 1760.350 2791.020 ;
        RECT 1676.310 2790.820 1760.350 2790.960 ;
        RECT 1676.310 2790.760 1676.630 2790.820 ;
        RECT 1718.170 2790.760 1718.490 2790.820 ;
        RECT 1760.030 2790.760 1760.350 2790.820 ;
        RECT 1770.150 2790.960 1770.470 2791.020 ;
        RECT 2401.730 2790.960 2402.050 2791.020 ;
        RECT 1770.150 2790.820 2402.050 2790.960 ;
        RECT 1770.150 2790.760 1770.470 2790.820 ;
        RECT 2401.730 2790.760 2402.050 2790.820 ;
        RECT 1783.490 2790.620 1783.810 2790.680 ;
        RECT 2415.070 2790.620 2415.390 2790.680 ;
        RECT 1783.490 2790.480 2415.390 2790.620 ;
        RECT 1783.490 2790.420 1783.810 2790.480 ;
        RECT 2415.070 2790.420 2415.390 2790.480 ;
        RECT 1776.590 2790.280 1776.910 2790.340 ;
        RECT 2408.170 2790.280 2408.490 2790.340 ;
        RECT 1776.590 2790.140 2408.490 2790.280 ;
        RECT 1776.590 2790.080 1776.910 2790.140 ;
        RECT 2408.170 2790.080 2408.490 2790.140 ;
        RECT 1610.990 2789.800 1657.680 2789.940 ;
        RECT 1783.950 2789.940 1784.270 2790.000 ;
        RECT 2421.970 2789.940 2422.290 2790.000 ;
        RECT 1783.950 2789.800 2422.290 2789.940 ;
        RECT 1610.990 2789.740 1611.310 2789.800 ;
        RECT 1783.950 2789.740 1784.270 2789.800 ;
        RECT 2421.970 2789.740 2422.290 2789.800 ;
        RECT 469.285 2789.600 469.575 2789.645 ;
        RECT 485.385 2789.600 485.675 2789.645 ;
        RECT 469.285 2789.460 485.675 2789.600 ;
        RECT 469.285 2789.415 469.575 2789.460 ;
        RECT 485.385 2789.415 485.675 2789.460 ;
        RECT 485.830 2789.600 486.150 2789.660 ;
        RECT 498.725 2789.600 499.015 2789.645 ;
        RECT 485.830 2789.460 499.015 2789.600 ;
        RECT 485.830 2789.400 486.150 2789.460 ;
        RECT 498.725 2789.415 499.015 2789.460 ;
        RECT 499.185 2789.600 499.475 2789.645 ;
        RECT 527.690 2789.600 528.010 2789.660 ;
        RECT 499.185 2789.460 528.010 2789.600 ;
        RECT 499.185 2789.415 499.475 2789.460 ;
        RECT 527.690 2789.400 528.010 2789.460 ;
        RECT 648.210 2789.600 648.530 2789.660 ;
        RECT 1042.905 2789.600 1043.195 2789.645 ;
        RECT 648.210 2789.460 1043.195 2789.600 ;
        RECT 648.210 2789.400 648.530 2789.460 ;
        RECT 1042.905 2789.415 1043.195 2789.460 ;
        RECT 1110.985 2789.600 1111.275 2789.645 ;
        RECT 1117.870 2789.600 1118.190 2789.660 ;
        RECT 1158.825 2789.600 1159.115 2789.645 ;
        RECT 1110.985 2789.460 1159.115 2789.600 ;
        RECT 1110.985 2789.415 1111.275 2789.460 ;
        RECT 1117.870 2789.400 1118.190 2789.460 ;
        RECT 1158.825 2789.415 1159.115 2789.460 ;
        RECT 1432.970 2789.600 1433.290 2789.660 ;
        RECT 1649.170 2789.600 1649.490 2789.660 ;
        RECT 1432.970 2789.460 1649.490 2789.600 ;
        RECT 1432.970 2789.400 1433.290 2789.460 ;
        RECT 1649.170 2789.400 1649.490 2789.460 ;
        RECT 1777.050 2789.600 1777.370 2789.660 ;
        RECT 2415.070 2789.600 2415.390 2789.660 ;
        RECT 1777.050 2789.460 2415.390 2789.600 ;
        RECT 1777.050 2789.400 1777.370 2789.460 ;
        RECT 2415.070 2789.400 2415.390 2789.460 ;
        RECT 445.810 2789.260 446.130 2789.320 ;
        RECT 469.745 2789.260 470.035 2789.305 ;
        RECT 445.810 2789.120 470.035 2789.260 ;
        RECT 445.810 2789.060 446.130 2789.120 ;
        RECT 469.745 2789.075 470.035 2789.120 ;
        RECT 491.365 2789.260 491.655 2789.305 ;
        RECT 531.385 2789.260 531.675 2789.305 ;
        RECT 627.065 2789.260 627.355 2789.305 ;
        RECT 491.365 2789.120 531.675 2789.260 ;
        RECT 491.365 2789.075 491.655 2789.120 ;
        RECT 531.385 2789.075 531.675 2789.120 ;
        RECT 606.440 2789.120 627.355 2789.260 ;
        RECT 465.590 2788.920 465.910 2788.980 ;
        RECT 504.230 2788.920 504.550 2788.980 ;
        RECT 465.590 2788.780 504.550 2788.920 ;
        RECT 465.590 2788.720 465.910 2788.780 ;
        RECT 504.230 2788.720 504.550 2788.780 ;
        RECT 579.225 2788.920 579.515 2788.965 ;
        RECT 606.440 2788.920 606.580 2789.120 ;
        RECT 627.065 2789.075 627.355 2789.120 ;
        RECT 627.510 2789.260 627.830 2789.320 ;
        RECT 1042.430 2789.260 1042.750 2789.320 ;
        RECT 627.510 2789.120 1042.750 2789.260 ;
        RECT 627.510 2789.060 627.830 2789.120 ;
        RECT 1042.430 2789.060 1042.750 2789.120 ;
        RECT 1624.790 2789.260 1625.110 2789.320 ;
        RECT 1628.485 2789.260 1628.775 2789.305 ;
        RECT 1624.790 2789.120 1628.775 2789.260 ;
        RECT 1624.790 2789.060 1625.110 2789.120 ;
        RECT 1628.485 2789.075 1628.775 2789.120 ;
        RECT 1790.390 2789.260 1790.710 2789.320 ;
        RECT 2428.870 2789.260 2429.190 2789.320 ;
        RECT 1790.390 2789.120 2429.190 2789.260 ;
        RECT 1790.390 2789.060 1790.710 2789.120 ;
        RECT 2428.870 2789.060 2429.190 2789.120 ;
        RECT 579.225 2788.780 606.580 2788.920 ;
        RECT 606.810 2788.920 607.130 2788.980 ;
        RECT 1034.610 2788.920 1034.930 2788.980 ;
        RECT 606.810 2788.780 1034.930 2788.920 ;
        RECT 579.225 2788.735 579.515 2788.780 ;
        RECT 606.810 2788.720 607.130 2788.780 ;
        RECT 1034.610 2788.720 1034.930 2788.780 ;
        RECT 1045.190 2788.920 1045.510 2788.980 ;
        RECT 1093.950 2788.920 1094.270 2788.980 ;
        RECT 1045.190 2788.780 1094.270 2788.920 ;
        RECT 1045.190 2788.720 1045.510 2788.780 ;
        RECT 1093.950 2788.720 1094.270 2788.780 ;
        RECT 1438.950 2788.920 1439.270 2788.980 ;
        RECT 1656.070 2788.920 1656.390 2788.980 ;
        RECT 1438.950 2788.780 1656.390 2788.920 ;
        RECT 1438.950 2788.720 1439.270 2788.780 ;
        RECT 1656.070 2788.720 1656.390 2788.780 ;
        RECT 1790.850 2788.920 1791.170 2788.980 ;
        RECT 2435.770 2788.920 2436.090 2788.980 ;
        RECT 1790.850 2788.780 2436.090 2788.920 ;
        RECT 1790.850 2788.720 1791.170 2788.780 ;
        RECT 2435.770 2788.720 2436.090 2788.780 ;
        RECT 426.950 2788.580 427.270 2788.640 ;
        RECT 473.870 2788.580 474.190 2788.640 ;
        RECT 426.950 2788.440 474.190 2788.580 ;
        RECT 426.950 2788.380 427.270 2788.440 ;
        RECT 473.870 2788.380 474.190 2788.440 ;
        RECT 474.345 2788.580 474.635 2788.625 ;
        RECT 491.365 2788.580 491.655 2788.625 ;
        RECT 474.345 2788.440 491.655 2788.580 ;
        RECT 474.345 2788.395 474.635 2788.440 ;
        RECT 491.365 2788.395 491.655 2788.440 ;
        RECT 491.810 2788.580 492.130 2788.640 ;
        RECT 541.490 2788.580 541.810 2788.640 ;
        RECT 491.810 2788.440 541.810 2788.580 ;
        RECT 491.810 2788.380 492.130 2788.440 ;
        RECT 541.490 2788.380 541.810 2788.440 ;
        RECT 586.110 2788.580 586.430 2788.640 ;
        RECT 1018.970 2788.580 1019.290 2788.640 ;
        RECT 586.110 2788.440 1019.290 2788.580 ;
        RECT 586.110 2788.380 586.430 2788.440 ;
        RECT 1018.970 2788.380 1019.290 2788.440 ;
        RECT 1024.490 2788.580 1024.810 2788.640 ;
        RECT 1070.030 2788.580 1070.350 2788.640 ;
        RECT 1076.010 2788.580 1076.330 2788.640 ;
        RECT 1024.490 2788.440 1076.330 2788.580 ;
        RECT 1024.490 2788.380 1024.810 2788.440 ;
        RECT 1070.030 2788.380 1070.350 2788.440 ;
        RECT 1076.010 2788.380 1076.330 2788.440 ;
        RECT 1425.150 2788.580 1425.470 2788.640 ;
        RECT 2249.470 2788.580 2249.790 2788.640 ;
        RECT 1425.150 2788.440 2249.790 2788.580 ;
        RECT 1425.150 2788.380 1425.470 2788.440 ;
        RECT 2249.470 2788.380 2249.790 2788.440 ;
        RECT 2301.910 2788.580 2302.230 2788.640 ;
        RECT 2340.550 2788.580 2340.870 2788.640 ;
        RECT 2301.910 2788.440 2340.870 2788.580 ;
        RECT 2301.910 2788.380 2302.230 2788.440 ;
        RECT 2340.550 2788.380 2340.870 2788.440 ;
        RECT 2374.130 2788.580 2374.450 2788.640 ;
        RECT 2415.070 2788.580 2415.390 2788.640 ;
        RECT 2374.130 2788.440 2415.390 2788.580 ;
        RECT 2374.130 2788.380 2374.450 2788.440 ;
        RECT 2415.070 2788.380 2415.390 2788.440 ;
        RECT 455.470 2788.240 455.790 2788.300 ;
        RECT 500.090 2788.240 500.410 2788.300 ;
        RECT 455.470 2788.100 500.410 2788.240 ;
        RECT 455.470 2788.040 455.790 2788.100 ;
        RECT 500.090 2788.040 500.410 2788.100 ;
        RECT 501.930 2788.240 502.250 2788.300 ;
        RECT 542.410 2788.240 542.730 2788.300 ;
        RECT 501.930 2788.100 542.730 2788.240 ;
        RECT 501.930 2788.040 502.250 2788.100 ;
        RECT 542.410 2788.040 542.730 2788.100 ;
        RECT 1010.690 2788.240 1011.010 2788.300 ;
        RECT 1055.770 2788.240 1056.090 2788.300 ;
        RECT 1010.690 2788.100 1056.090 2788.240 ;
        RECT 1010.690 2788.040 1011.010 2788.100 ;
        RECT 1055.770 2788.040 1056.090 2788.100 ;
        RECT 1576.490 2788.240 1576.810 2788.300 ;
        RECT 1621.570 2788.240 1621.890 2788.300 ;
        RECT 1576.490 2788.100 1621.890 2788.240 ;
        RECT 1576.490 2788.040 1576.810 2788.100 ;
        RECT 1621.570 2788.040 1621.890 2788.100 ;
        RECT 1638.590 2788.240 1638.910 2788.300 ;
        RECT 1680.450 2788.240 1680.770 2788.300 ;
        RECT 1638.590 2788.100 1680.770 2788.240 ;
        RECT 1638.590 2788.040 1638.910 2788.100 ;
        RECT 1680.450 2788.040 1680.770 2788.100 ;
        RECT 2300.990 2788.240 2301.310 2788.300 ;
        RECT 2304.210 2788.240 2304.530 2788.300 ;
        RECT 2350.210 2788.240 2350.530 2788.300 ;
        RECT 2394.830 2788.240 2395.150 2788.300 ;
        RECT 2300.990 2788.100 2395.150 2788.240 ;
        RECT 2300.990 2788.040 2301.310 2788.100 ;
        RECT 2304.210 2788.040 2304.530 2788.100 ;
        RECT 2350.210 2788.040 2350.530 2788.100 ;
        RECT 2394.830 2788.040 2395.150 2788.100 ;
        RECT 337.250 2787.900 337.570 2787.960 ;
        RECT 641.325 2787.900 641.615 2787.945 ;
        RECT 337.250 2787.760 641.615 2787.900 ;
        RECT 337.250 2787.700 337.570 2787.760 ;
        RECT 641.325 2787.715 641.615 2787.760 ;
        RECT 641.785 2787.900 642.075 2787.945 ;
        RECT 1007.470 2787.900 1007.790 2787.960 ;
        RECT 641.785 2787.760 1007.790 2787.900 ;
        RECT 641.785 2787.715 642.075 2787.760 ;
        RECT 1007.470 2787.700 1007.790 2787.760 ;
        RECT 1038.290 2787.900 1038.610 2787.960 ;
        RECT 1087.510 2787.900 1087.830 2787.960 ;
        RECT 1038.290 2787.760 1087.830 2787.900 ;
        RECT 1038.290 2787.700 1038.610 2787.760 ;
        RECT 1087.510 2787.700 1087.830 2787.760 ;
        RECT 1541.990 2787.900 1542.310 2787.960 ;
        RECT 1581.550 2787.900 1581.870 2787.960 ;
        RECT 1541.990 2787.760 1581.870 2787.900 ;
        RECT 1541.990 2787.700 1542.310 2787.760 ;
        RECT 1581.550 2787.700 1581.870 2787.760 ;
        RECT 1645.490 2787.900 1645.810 2787.960 ;
        RECT 1687.810 2787.900 1688.130 2787.960 ;
        RECT 1645.490 2787.760 1688.130 2787.900 ;
        RECT 1645.490 2787.700 1645.810 2787.760 ;
        RECT 1687.810 2787.700 1688.130 2787.760 ;
        RECT 2321.690 2787.900 2322.010 2787.960 ;
        RECT 2442.670 2787.900 2442.990 2787.960 ;
        RECT 2321.690 2787.760 2442.990 2787.900 ;
        RECT 2321.690 2787.700 2322.010 2787.760 ;
        RECT 2442.670 2787.700 2442.990 2787.760 ;
        RECT 531.385 2787.560 531.675 2787.605 ;
        RECT 579.225 2787.560 579.515 2787.605 ;
        RECT 531.385 2787.420 579.515 2787.560 ;
        RECT 531.385 2787.375 531.675 2787.420 ;
        RECT 579.225 2787.375 579.515 2787.420 ;
        RECT 627.065 2787.560 627.355 2787.605 ;
        RECT 627.985 2787.560 628.275 2787.605 ;
        RECT 627.065 2787.420 628.275 2787.560 ;
        RECT 627.065 2787.375 627.355 2787.420 ;
        RECT 627.985 2787.375 628.275 2787.420 ;
        RECT 627.985 2784.500 628.275 2784.545 ;
        RECT 658.790 2784.500 659.110 2784.560 ;
        RECT 627.985 2784.360 659.110 2784.500 ;
        RECT 627.985 2784.315 628.275 2784.360 ;
        RECT 658.790 2784.300 659.110 2784.360 ;
        RECT 482.610 2725.340 482.930 2725.400 ;
        RECT 948.130 2725.340 948.450 2725.400 ;
        RECT 482.610 2725.200 948.450 2725.340 ;
        RECT 482.610 2725.140 482.930 2725.200 ;
        RECT 948.130 2725.140 948.450 2725.200 ;
        RECT 470.650 2725.000 470.970 2725.060 ;
        RECT 942.150 2725.000 942.470 2725.060 ;
        RECT 470.650 2724.860 942.470 2725.000 ;
        RECT 470.650 2724.800 470.970 2724.860 ;
        RECT 942.150 2724.800 942.470 2724.860 ;
        RECT 510.210 2724.660 510.530 2724.720 ;
        RECT 989.530 2724.660 989.850 2724.720 ;
        RECT 510.210 2724.520 989.850 2724.660 ;
        RECT 510.210 2724.460 510.530 2724.520 ;
        RECT 989.530 2724.460 989.850 2724.520 ;
        RECT 460.530 2724.320 460.850 2724.380 ;
        RECT 942.610 2724.320 942.930 2724.380 ;
        RECT 460.530 2724.180 942.930 2724.320 ;
        RECT 460.530 2724.120 460.850 2724.180 ;
        RECT 942.610 2724.120 942.930 2724.180 ;
        RECT 449.950 2723.980 450.270 2724.040 ;
        RECT 943.070 2723.980 943.390 2724.040 ;
        RECT 449.950 2723.840 943.390 2723.980 ;
        RECT 449.950 2723.780 450.270 2723.840 ;
        RECT 943.070 2723.780 943.390 2723.840 ;
        RECT 530.910 2723.640 531.230 2723.700 ;
        RECT 1030.930 2723.640 1031.250 2723.700 ;
        RECT 530.910 2723.500 1031.250 2723.640 ;
        RECT 530.910 2723.440 531.230 2723.500 ;
        RECT 1030.930 2723.440 1031.250 2723.500 ;
        RECT 439.830 2723.300 440.150 2723.360 ;
        RECT 943.530 2723.300 943.850 2723.360 ;
        RECT 439.830 2723.160 943.850 2723.300 ;
        RECT 439.830 2723.100 440.150 2723.160 ;
        RECT 943.530 2723.100 943.850 2723.160 ;
        RECT 551.610 2722.960 551.930 2723.020 ;
        RECT 1062.210 2722.960 1062.530 2723.020 ;
        RECT 551.610 2722.820 1062.530 2722.960 ;
        RECT 551.610 2722.760 551.930 2722.820 ;
        RECT 1062.210 2722.760 1062.530 2722.820 ;
        RECT 429.250 2722.620 429.570 2722.680 ;
        RECT 943.990 2722.620 944.310 2722.680 ;
        RECT 429.250 2722.480 944.310 2722.620 ;
        RECT 429.250 2722.420 429.570 2722.480 ;
        RECT 943.990 2722.420 944.310 2722.480 ;
        RECT 419.130 2722.280 419.450 2722.340 ;
        RECT 944.450 2722.280 944.770 2722.340 ;
        RECT 419.130 2722.140 944.770 2722.280 ;
        RECT 419.130 2722.080 419.450 2722.140 ;
        RECT 944.450 2722.080 944.770 2722.140 ;
        RECT 408.550 2721.940 408.870 2722.000 ;
        RECT 979.870 2721.940 980.190 2722.000 ;
        RECT 408.550 2721.800 980.190 2721.940 ;
        RECT 408.550 2721.740 408.870 2721.800 ;
        RECT 979.870 2721.740 980.190 2721.800 ;
        RECT 433.850 2721.600 434.170 2721.660 ;
        RECT 865.330 2721.600 865.650 2721.660 ;
        RECT 433.850 2721.460 865.650 2721.600 ;
        RECT 433.850 2721.400 434.170 2721.460 ;
        RECT 865.330 2721.400 865.650 2721.460 ;
        RECT 441.210 2721.260 441.530 2721.320 ;
        RECT 875.450 2721.260 875.770 2721.320 ;
        RECT 441.210 2721.120 875.770 2721.260 ;
        RECT 441.210 2721.060 441.530 2721.120 ;
        RECT 875.450 2721.060 875.770 2721.120 ;
        RECT 427.410 2720.920 427.730 2720.980 ;
        RECT 844.170 2720.920 844.490 2720.980 ;
        RECT 427.410 2720.780 844.490 2720.920 ;
        RECT 427.410 2720.720 427.730 2720.780 ;
        RECT 844.170 2720.720 844.490 2720.780 ;
        RECT 434.310 2720.580 434.630 2720.640 ;
        RECT 854.750 2720.580 855.070 2720.640 ;
        RECT 434.310 2720.440 855.070 2720.580 ;
        RECT 434.310 2720.380 434.630 2720.440 ;
        RECT 854.750 2720.380 855.070 2720.440 ;
        RECT 413.610 2720.240 413.930 2720.300 ;
        RECT 823.470 2720.240 823.790 2720.300 ;
        RECT 413.610 2720.100 823.790 2720.240 ;
        RECT 413.610 2720.040 413.930 2720.100 ;
        RECT 823.470 2720.040 823.790 2720.100 ;
        RECT 365.310 2719.900 365.630 2719.960 ;
        RECT 740.670 2719.900 740.990 2719.960 ;
        RECT 365.310 2719.760 740.990 2719.900 ;
        RECT 365.310 2719.700 365.630 2719.760 ;
        RECT 740.670 2719.700 740.990 2719.760 ;
        RECT 289.410 2719.560 289.730 2719.620 ;
        RECT 564.030 2719.560 564.350 2719.620 ;
        RECT 289.410 2719.420 564.350 2719.560 ;
        RECT 289.410 2719.360 289.730 2719.420 ;
        RECT 564.030 2719.360 564.350 2719.420 ;
        RECT 288.950 2719.220 289.270 2719.280 ;
        RECT 553.910 2719.220 554.230 2719.280 ;
        RECT 288.950 2719.080 554.230 2719.220 ;
        RECT 288.950 2719.020 289.270 2719.080 ;
        RECT 553.910 2719.020 554.230 2719.080 ;
        RECT 1103.610 2718.680 1103.930 2718.940 ;
        RECT 358.410 2718.540 358.730 2718.600 ;
        RECT 377.270 2718.540 377.590 2718.600 ;
        RECT 358.410 2718.400 377.590 2718.540 ;
        RECT 358.410 2718.340 358.730 2718.400 ;
        RECT 377.270 2718.340 377.590 2718.400 ;
        RECT 379.110 2718.540 379.430 2718.600 ;
        RECT 727.345 2718.540 727.635 2718.585 ;
        RECT 379.110 2718.400 727.635 2718.540 ;
        RECT 379.110 2718.340 379.430 2718.400 ;
        RECT 727.345 2718.355 727.635 2718.400 ;
        RECT 727.790 2718.540 728.110 2718.600 ;
        RECT 762.305 2718.540 762.595 2718.585 ;
        RECT 727.790 2718.400 762.595 2718.540 ;
        RECT 727.790 2718.340 728.110 2718.400 ;
        RECT 762.305 2718.355 762.595 2718.400 ;
        RECT 762.750 2718.540 763.070 2718.600 ;
        RECT 813.350 2718.540 813.670 2718.600 ;
        RECT 762.750 2718.400 813.670 2718.540 ;
        RECT 762.750 2718.340 763.070 2718.400 ;
        RECT 813.350 2718.340 813.670 2718.400 ;
        RECT 1027.710 2718.540 1028.030 2718.600 ;
        RECT 1093.490 2718.540 1093.810 2718.600 ;
        RECT 1027.710 2718.400 1093.810 2718.540 ;
        RECT 1027.710 2718.340 1028.030 2718.400 ;
        RECT 1093.490 2718.340 1093.810 2718.400 ;
        RECT 1102.690 2718.540 1103.010 2718.600 ;
        RECT 1103.700 2718.540 1103.840 2718.680 ;
        RECT 1102.690 2718.400 1103.840 2718.540 ;
        RECT 1145.010 2718.540 1145.330 2718.600 ;
        RECT 1300.950 2718.540 1301.270 2718.600 ;
        RECT 1145.010 2718.400 1301.270 2718.540 ;
        RECT 1102.690 2718.340 1103.010 2718.400 ;
        RECT 1145.010 2718.340 1145.330 2718.400 ;
        RECT 1300.950 2718.340 1301.270 2718.400 ;
        RECT 351.510 2718.200 351.830 2718.260 ;
        RECT 367.150 2718.200 367.470 2718.260 ;
        RECT 351.510 2718.060 367.470 2718.200 ;
        RECT 351.510 2718.000 351.830 2718.060 ;
        RECT 367.150 2718.000 367.470 2718.060 ;
        RECT 392.910 2718.200 393.230 2718.260 ;
        RECT 782.070 2718.200 782.390 2718.260 ;
        RECT 392.910 2718.060 782.390 2718.200 ;
        RECT 392.910 2718.000 393.230 2718.060 ;
        RECT 782.070 2718.000 782.390 2718.060 ;
        RECT 1034.610 2718.200 1034.930 2718.260 ;
        RECT 1103.610 2718.200 1103.930 2718.260 ;
        RECT 1034.610 2718.060 1103.930 2718.200 ;
        RECT 1034.610 2718.000 1034.930 2718.060 ;
        RECT 1103.610 2718.000 1103.930 2718.060 ;
        RECT 1138.110 2718.200 1138.430 2718.260 ;
        RECT 1290.370 2718.200 1290.690 2718.260 ;
        RECT 1138.110 2718.060 1290.690 2718.200 ;
        RECT 1138.110 2718.000 1138.430 2718.060 ;
        RECT 1290.370 2718.000 1290.690 2718.060 ;
        RECT 305.050 2717.860 305.370 2717.920 ;
        RECT 310.110 2717.860 310.430 2717.920 ;
        RECT 305.050 2717.720 310.430 2717.860 ;
        RECT 305.050 2717.660 305.370 2717.720 ;
        RECT 310.110 2717.660 310.430 2717.720 ;
        RECT 325.750 2717.860 326.070 2717.920 ;
        RECT 330.810 2717.860 331.130 2717.920 ;
        RECT 325.750 2717.720 331.130 2717.860 ;
        RECT 325.750 2717.660 326.070 2717.720 ;
        RECT 330.810 2717.660 331.130 2717.720 ;
        RECT 351.050 2717.860 351.370 2717.920 ;
        RECT 356.570 2717.860 356.890 2717.920 ;
        RECT 351.050 2717.720 356.890 2717.860 ;
        RECT 351.050 2717.660 351.370 2717.720 ;
        RECT 356.570 2717.660 356.890 2717.720 ;
        RECT 399.350 2717.860 399.670 2717.920 ;
        RECT 761.845 2717.860 762.135 2717.905 ;
        RECT 399.350 2717.720 762.135 2717.860 ;
        RECT 399.350 2717.660 399.670 2717.720 ;
        RECT 761.845 2717.675 762.135 2717.720 ;
        RECT 762.290 2717.860 762.610 2717.920 ;
        RECT 792.650 2717.860 792.970 2717.920 ;
        RECT 762.290 2717.720 792.970 2717.860 ;
        RECT 762.290 2717.660 762.610 2717.720 ;
        RECT 792.650 2717.660 792.970 2717.720 ;
        RECT 1041.510 2717.860 1041.830 2717.920 ;
        RECT 1114.190 2717.860 1114.510 2717.920 ;
        RECT 1041.510 2717.720 1114.510 2717.860 ;
        RECT 1041.510 2717.660 1041.830 2717.720 ;
        RECT 1114.190 2717.660 1114.510 2717.720 ;
        RECT 1151.910 2717.860 1152.230 2717.920 ;
        RECT 1311.070 2717.860 1311.390 2717.920 ;
        RECT 1151.910 2717.720 1311.390 2717.860 ;
        RECT 1151.910 2717.660 1152.230 2717.720 ;
        RECT 1311.070 2717.660 1311.390 2717.720 ;
        RECT 287.110 2717.520 287.430 2717.580 ;
        RECT 512.510 2717.520 512.830 2717.580 ;
        RECT 287.110 2717.380 512.830 2717.520 ;
        RECT 287.110 2717.320 287.430 2717.380 ;
        RECT 512.510 2717.320 512.830 2717.380 ;
        RECT 636.710 2717.520 637.030 2717.580 ;
        RECT 1045.190 2717.520 1045.510 2717.580 ;
        RECT 636.710 2717.380 1045.510 2717.520 ;
        RECT 636.710 2717.320 637.030 2717.380 ;
        RECT 1045.190 2717.320 1045.510 2717.380 ;
        RECT 1048.410 2717.520 1048.730 2717.580 ;
        RECT 1124.310 2717.520 1124.630 2717.580 ;
        RECT 1048.410 2717.380 1124.630 2717.520 ;
        RECT 1048.410 2717.320 1048.730 2717.380 ;
        RECT 1124.310 2717.320 1124.630 2717.380 ;
        RECT 1158.810 2717.520 1159.130 2717.580 ;
        RECT 1321.650 2717.520 1321.970 2717.580 ;
        RECT 1158.810 2717.380 1321.970 2717.520 ;
        RECT 1158.810 2717.320 1159.130 2717.380 ;
        RECT 1321.650 2717.320 1321.970 2717.380 ;
        RECT 287.570 2717.180 287.890 2717.240 ;
        RECT 522.630 2717.180 522.950 2717.240 ;
        RECT 287.570 2717.040 522.950 2717.180 ;
        RECT 287.570 2716.980 287.890 2717.040 ;
        RECT 522.630 2716.980 522.950 2717.040 ;
        RECT 616.010 2717.180 616.330 2717.240 ;
        RECT 1038.290 2717.180 1038.610 2717.240 ;
        RECT 616.010 2717.040 1038.610 2717.180 ;
        RECT 616.010 2716.980 616.330 2717.040 ;
        RECT 1038.290 2716.980 1038.610 2717.040 ;
        RECT 1055.310 2717.180 1055.630 2717.240 ;
        RECT 1134.890 2717.180 1135.210 2717.240 ;
        RECT 1055.310 2717.040 1135.210 2717.180 ;
        RECT 1055.310 2716.980 1055.630 2717.040 ;
        RECT 1134.890 2716.980 1135.210 2717.040 ;
        RECT 1165.710 2717.180 1166.030 2717.240 ;
        RECT 1332.230 2717.180 1332.550 2717.240 ;
        RECT 1165.710 2717.040 1332.550 2717.180 ;
        RECT 1165.710 2716.980 1166.030 2717.040 ;
        RECT 1332.230 2716.980 1332.550 2717.040 ;
        RECT 288.030 2716.840 288.350 2716.900 ;
        RECT 533.210 2716.840 533.530 2716.900 ;
        RECT 288.030 2716.700 533.530 2716.840 ;
        RECT 288.030 2716.640 288.350 2716.700 ;
        RECT 533.210 2716.640 533.530 2716.700 ;
        RECT 595.310 2716.840 595.630 2716.900 ;
        RECT 1024.490 2716.840 1024.810 2716.900 ;
        RECT 595.310 2716.700 1024.810 2716.840 ;
        RECT 595.310 2716.640 595.630 2716.700 ;
        RECT 1024.490 2716.640 1024.810 2716.700 ;
        RECT 1061.750 2716.840 1062.070 2716.900 ;
        RECT 1155.590 2716.840 1155.910 2716.900 ;
        RECT 1061.750 2716.700 1155.910 2716.840 ;
        RECT 1061.750 2716.640 1062.070 2716.700 ;
        RECT 1155.590 2716.640 1155.910 2716.700 ;
        RECT 1165.250 2716.840 1165.570 2716.900 ;
        RECT 1342.350 2716.840 1342.670 2716.900 ;
        RECT 1165.250 2716.700 1342.670 2716.840 ;
        RECT 1165.250 2716.640 1165.570 2716.700 ;
        RECT 1342.350 2716.640 1342.670 2716.700 ;
        RECT 455.010 2716.500 455.330 2716.560 ;
        RECT 896.150 2716.500 896.470 2716.560 ;
        RECT 455.010 2716.360 896.470 2716.500 ;
        RECT 455.010 2716.300 455.330 2716.360 ;
        RECT 896.150 2716.300 896.470 2716.360 ;
        RECT 1076.010 2716.500 1076.330 2716.560 ;
        RECT 1176.290 2716.500 1176.610 2716.560 ;
        RECT 1076.010 2716.360 1176.610 2716.500 ;
        RECT 1076.010 2716.300 1076.330 2716.360 ;
        RECT 1176.290 2716.300 1176.610 2716.360 ;
        RECT 1179.510 2716.500 1179.830 2716.560 ;
        RECT 1363.050 2716.500 1363.370 2716.560 ;
        RECT 1179.510 2716.360 1363.370 2716.500 ;
        RECT 1179.510 2716.300 1179.830 2716.360 ;
        RECT 1363.050 2716.300 1363.370 2716.360 ;
        RECT 288.490 2716.160 288.810 2716.220 ;
        RECT 543.330 2716.160 543.650 2716.220 ;
        RECT 288.490 2716.020 543.650 2716.160 ;
        RECT 288.490 2715.960 288.810 2716.020 ;
        RECT 543.330 2715.960 543.650 2716.020 ;
        RECT 574.610 2716.160 574.930 2716.220 ;
        RECT 1010.690 2716.160 1011.010 2716.220 ;
        RECT 574.610 2716.020 1011.010 2716.160 ;
        RECT 574.610 2715.960 574.930 2716.020 ;
        RECT 1010.690 2715.960 1011.010 2716.020 ;
        RECT 1082.450 2716.160 1082.770 2716.220 ;
        RECT 1083.845 2716.160 1084.135 2716.205 ;
        RECT 1145.470 2716.160 1145.790 2716.220 ;
        RECT 1082.450 2716.020 1083.600 2716.160 ;
        RECT 1082.450 2715.960 1082.770 2716.020 ;
        RECT 468.350 2715.820 468.670 2715.880 ;
        RECT 916.850 2715.820 917.170 2715.880 ;
        RECT 468.350 2715.680 917.170 2715.820 ;
        RECT 468.350 2715.620 468.670 2715.680 ;
        RECT 916.850 2715.620 917.170 2715.680 ;
        RECT 1020.810 2715.820 1021.130 2715.880 ;
        RECT 1082.910 2715.820 1083.230 2715.880 ;
        RECT 1020.810 2715.680 1083.230 2715.820 ;
        RECT 1083.460 2715.820 1083.600 2716.020 ;
        RECT 1083.845 2716.020 1145.790 2716.160 ;
        RECT 1083.845 2715.975 1084.135 2716.020 ;
        RECT 1145.470 2715.960 1145.790 2716.020 ;
        RECT 1172.610 2716.160 1172.930 2716.220 ;
        RECT 1352.930 2716.160 1353.250 2716.220 ;
        RECT 1172.610 2716.020 1353.250 2716.160 ;
        RECT 1172.610 2715.960 1172.930 2716.020 ;
        RECT 1352.930 2715.960 1353.250 2716.020 ;
        RECT 1186.870 2715.820 1187.190 2715.880 ;
        RECT 1083.460 2715.680 1187.190 2715.820 ;
        RECT 1020.810 2715.620 1021.130 2715.680 ;
        RECT 1082.910 2715.620 1083.230 2715.680 ;
        RECT 1186.870 2715.620 1187.190 2715.680 ;
        RECT 1193.310 2715.820 1193.630 2715.880 ;
        RECT 1383.750 2715.820 1384.070 2715.880 ;
        RECT 1193.310 2715.680 1384.070 2715.820 ;
        RECT 1193.310 2715.620 1193.630 2715.680 ;
        RECT 1383.750 2715.620 1384.070 2715.680 ;
        RECT 286.190 2715.480 286.510 2715.540 ;
        RECT 398.430 2715.480 398.750 2715.540 ;
        RECT 286.190 2715.340 398.750 2715.480 ;
        RECT 286.190 2715.280 286.510 2715.340 ;
        RECT 398.430 2715.280 398.750 2715.340 ;
        RECT 475.250 2715.480 475.570 2715.540 ;
        RECT 937.550 2715.480 937.870 2715.540 ;
        RECT 475.250 2715.340 937.870 2715.480 ;
        RECT 475.250 2715.280 475.570 2715.340 ;
        RECT 937.550 2715.280 937.870 2715.340 ;
        RECT 1069.110 2715.480 1069.430 2715.540 ;
        RECT 1166.170 2715.480 1166.490 2715.540 ;
        RECT 1069.110 2715.340 1166.490 2715.480 ;
        RECT 1069.110 2715.280 1069.430 2715.340 ;
        RECT 1166.170 2715.280 1166.490 2715.340 ;
        RECT 1186.410 2715.480 1186.730 2715.540 ;
        RECT 1373.630 2715.480 1373.950 2715.540 ;
        RECT 1186.410 2715.340 1373.950 2715.480 ;
        RECT 1186.410 2715.280 1186.730 2715.340 ;
        RECT 1373.630 2715.280 1373.950 2715.340 ;
        RECT 337.710 2715.140 338.030 2715.200 ;
        RECT 491.810 2715.140 492.130 2715.200 ;
        RECT 337.710 2715.000 492.130 2715.140 ;
        RECT 337.710 2714.940 338.030 2715.000 ;
        RECT 491.810 2714.940 492.130 2715.000 ;
        RECT 496.410 2715.140 496.730 2715.200 ;
        RECT 968.830 2715.140 969.150 2715.200 ;
        RECT 496.410 2715.000 969.150 2715.140 ;
        RECT 496.410 2714.940 496.730 2715.000 ;
        RECT 968.830 2714.940 969.150 2715.000 ;
        RECT 1013.910 2715.140 1014.230 2715.200 ;
        RECT 1072.790 2715.140 1073.110 2715.200 ;
        RECT 1013.910 2715.000 1073.110 2715.140 ;
        RECT 1013.910 2714.940 1014.230 2715.000 ;
        RECT 1072.790 2714.940 1073.110 2715.000 ;
        RECT 1089.810 2715.140 1090.130 2715.200 ;
        RECT 1196.990 2715.140 1197.310 2715.200 ;
        RECT 1089.810 2715.000 1197.310 2715.140 ;
        RECT 1089.810 2714.940 1090.130 2715.000 ;
        RECT 1196.990 2714.940 1197.310 2715.000 ;
        RECT 1200.210 2715.140 1200.530 2715.200 ;
        RECT 1394.330 2715.140 1394.650 2715.200 ;
        RECT 1200.210 2715.000 1394.650 2715.140 ;
        RECT 1200.210 2714.940 1200.530 2715.000 ;
        RECT 1394.330 2714.940 1394.650 2715.000 ;
        RECT 286.650 2714.800 286.970 2714.860 ;
        RECT 501.930 2714.800 502.250 2714.860 ;
        RECT 286.650 2714.660 502.250 2714.800 ;
        RECT 286.650 2714.600 286.970 2714.660 ;
        RECT 501.930 2714.600 502.250 2714.660 ;
        RECT 541.490 2714.800 541.810 2714.860 ;
        RECT 719.970 2714.800 720.290 2714.860 ;
        RECT 541.490 2714.660 720.290 2714.800 ;
        RECT 541.490 2714.600 541.810 2714.660 ;
        RECT 719.970 2714.600 720.290 2714.660 ;
        RECT 720.890 2714.800 721.210 2714.860 ;
        RECT 1020.810 2714.800 1021.130 2714.860 ;
        RECT 720.890 2714.660 1021.130 2714.800 ;
        RECT 720.890 2714.600 721.210 2714.660 ;
        RECT 1020.810 2714.600 1021.130 2714.660 ;
        RECT 1054.850 2714.800 1055.170 2714.860 ;
        RECT 1083.845 2714.800 1084.135 2714.845 ;
        RECT 1054.850 2714.660 1084.135 2714.800 ;
        RECT 1054.850 2714.600 1055.170 2714.660 ;
        RECT 1083.845 2714.615 1084.135 2714.660 ;
        RECT 1130.750 2714.800 1131.070 2714.860 ;
        RECT 1280.250 2714.800 1280.570 2714.860 ;
        RECT 1130.750 2714.660 1280.570 2714.800 ;
        RECT 1130.750 2714.600 1131.070 2714.660 ;
        RECT 1280.250 2714.600 1280.570 2714.660 ;
        RECT 527.690 2714.460 528.010 2714.520 ;
        RECT 699.270 2714.460 699.590 2714.520 ;
        RECT 527.690 2714.320 699.590 2714.460 ;
        RECT 527.690 2714.260 528.010 2714.320 ;
        RECT 699.270 2714.260 699.590 2714.320 ;
        RECT 700.650 2714.460 700.970 2714.520 ;
        RECT 979.410 2714.460 979.730 2714.520 ;
        RECT 700.650 2714.320 979.730 2714.460 ;
        RECT 700.650 2714.260 700.970 2714.320 ;
        RECT 979.410 2714.260 979.730 2714.320 ;
        RECT 1131.210 2714.460 1131.530 2714.520 ;
        RECT 1269.670 2714.460 1269.990 2714.520 ;
        RECT 1131.210 2714.320 1269.990 2714.460 ;
        RECT 1131.210 2714.260 1131.530 2714.320 ;
        RECT 1269.670 2714.260 1269.990 2714.320 ;
        RECT 513.890 2714.120 514.210 2714.180 ;
        RECT 678.570 2714.120 678.890 2714.180 ;
        RECT 513.890 2713.980 678.890 2714.120 ;
        RECT 513.890 2713.920 514.210 2713.980 ;
        RECT 678.570 2713.920 678.890 2713.980 ;
        RECT 686.390 2714.120 686.710 2714.180 ;
        RECT 693.290 2714.120 693.610 2714.180 ;
        RECT 958.710 2714.120 959.030 2714.180 ;
        RECT 686.390 2713.980 689.380 2714.120 ;
        RECT 686.390 2713.920 686.710 2713.980 ;
        RECT 520.790 2713.780 521.110 2713.840 ;
        RECT 688.690 2713.780 689.010 2713.840 ;
        RECT 520.790 2713.640 689.010 2713.780 ;
        RECT 689.240 2713.780 689.380 2713.980 ;
        RECT 693.290 2713.980 959.030 2714.120 ;
        RECT 693.290 2713.920 693.610 2713.980 ;
        RECT 958.710 2713.920 959.030 2713.980 ;
        RECT 1117.410 2714.120 1117.730 2714.180 ;
        RECT 1248.970 2714.120 1249.290 2714.180 ;
        RECT 1117.410 2713.980 1249.290 2714.120 ;
        RECT 1117.410 2713.920 1117.730 2713.980 ;
        RECT 1248.970 2713.920 1249.290 2713.980 ;
        RECT 927.430 2713.780 927.750 2713.840 ;
        RECT 689.240 2713.640 927.750 2713.780 ;
        RECT 520.790 2713.580 521.110 2713.640 ;
        RECT 688.690 2713.580 689.010 2713.640 ;
        RECT 927.430 2713.580 927.750 2713.640 ;
        RECT 1123.390 2713.780 1123.710 2713.840 ;
        RECT 1259.550 2713.780 1259.870 2713.840 ;
        RECT 1123.390 2713.640 1259.870 2713.780 ;
        RECT 1123.390 2713.580 1123.710 2713.640 ;
        RECT 1259.550 2713.580 1259.870 2713.640 ;
        RECT 500.090 2713.440 500.410 2713.500 ;
        RECT 657.410 2713.440 657.730 2713.500 ;
        RECT 500.090 2713.300 657.730 2713.440 ;
        RECT 500.090 2713.240 500.410 2713.300 ;
        RECT 657.410 2713.240 657.730 2713.300 ;
        RECT 658.790 2713.440 659.110 2713.500 ;
        RECT 886.030 2713.440 886.350 2713.500 ;
        RECT 658.790 2713.300 886.350 2713.440 ;
        RECT 658.790 2713.240 659.110 2713.300 ;
        RECT 886.030 2713.240 886.350 2713.300 ;
        RECT 1102.690 2713.440 1103.010 2713.500 ;
        RECT 1228.270 2713.440 1228.590 2713.500 ;
        RECT 1102.690 2713.300 1228.590 2713.440 ;
        RECT 1102.690 2713.240 1103.010 2713.300 ;
        RECT 1228.270 2713.240 1228.590 2713.300 ;
        RECT 506.990 2713.100 507.310 2713.160 ;
        RECT 667.990 2713.100 668.310 2713.160 ;
        RECT 506.990 2712.960 668.310 2713.100 ;
        RECT 506.990 2712.900 507.310 2712.960 ;
        RECT 667.990 2712.900 668.310 2712.960 ;
        RECT 687.310 2713.100 687.630 2713.160 ;
        RECT 906.730 2713.100 907.050 2713.160 ;
        RECT 687.310 2712.960 907.050 2713.100 ;
        RECT 687.310 2712.900 687.630 2712.960 ;
        RECT 906.730 2712.900 907.050 2712.960 ;
        RECT 1110.510 2713.100 1110.830 2713.160 ;
        RECT 1238.850 2713.100 1239.170 2713.160 ;
        RECT 1110.510 2712.960 1239.170 2713.100 ;
        RECT 1110.510 2712.900 1110.830 2712.960 ;
        RECT 1238.850 2712.900 1239.170 2712.960 ;
        RECT 542.410 2712.760 542.730 2712.820 ;
        RECT 730.090 2712.760 730.410 2712.820 ;
        RECT 761.370 2712.760 761.690 2712.820 ;
        RECT 542.410 2712.620 730.410 2712.760 ;
        RECT 542.410 2712.560 542.730 2712.620 ;
        RECT 730.090 2712.560 730.410 2712.620 ;
        RECT 734.780 2712.620 761.690 2712.760 ;
        RECT 534.590 2712.420 534.910 2712.480 ;
        RECT 709.390 2712.420 709.710 2712.480 ;
        RECT 534.590 2712.280 709.710 2712.420 ;
        RECT 534.590 2712.220 534.910 2712.280 ;
        RECT 709.390 2712.220 709.710 2712.280 ;
        RECT 727.345 2712.420 727.635 2712.465 ;
        RECT 734.780 2712.420 734.920 2712.620 ;
        RECT 761.370 2712.560 761.690 2712.620 ;
        RECT 762.305 2712.760 762.595 2712.805 ;
        RECT 771.950 2712.760 772.270 2712.820 ;
        RECT 834.050 2712.760 834.370 2712.820 ;
        RECT 762.305 2712.620 772.270 2712.760 ;
        RECT 762.305 2712.575 762.595 2712.620 ;
        RECT 771.950 2712.560 772.270 2712.620 ;
        RECT 783.080 2712.620 834.370 2712.760 ;
        RECT 727.345 2712.280 734.920 2712.420 ;
        RECT 748.490 2712.420 748.810 2712.480 ;
        RECT 783.080 2712.420 783.220 2712.620 ;
        RECT 834.050 2712.560 834.370 2712.620 ;
        RECT 1089.350 2712.760 1089.670 2712.820 ;
        RECT 1207.570 2712.760 1207.890 2712.820 ;
        RECT 1089.350 2712.620 1207.890 2712.760 ;
        RECT 1089.350 2712.560 1089.670 2712.620 ;
        RECT 1207.570 2712.560 1207.890 2712.620 ;
        RECT 748.490 2712.280 783.220 2712.420 ;
        RECT 1096.710 2712.420 1097.030 2712.480 ;
        RECT 1217.690 2712.420 1218.010 2712.480 ;
        RECT 1096.710 2712.280 1218.010 2712.420 ;
        RECT 727.345 2712.235 727.635 2712.280 ;
        RECT 748.490 2712.220 748.810 2712.280 ;
        RECT 1096.710 2712.220 1097.030 2712.280 ;
        RECT 1217.690 2712.220 1218.010 2712.280 ;
        RECT 686.850 2712.080 687.170 2712.140 ;
        RECT 750.790 2712.080 751.110 2712.140 ;
        RECT 686.850 2711.940 751.110 2712.080 ;
        RECT 686.850 2711.880 687.170 2711.940 ;
        RECT 750.790 2711.880 751.110 2711.940 ;
        RECT 761.845 2712.080 762.135 2712.125 ;
        RECT 802.770 2712.080 803.090 2712.140 ;
        RECT 761.845 2711.940 803.090 2712.080 ;
        RECT 761.845 2711.895 762.135 2711.940 ;
        RECT 802.770 2711.880 803.090 2711.940 ;
      LAYER met1 ;
        RECT 300.070 1604.460 1395.190 2695.780 ;
      LAYER met1 ;
        RECT 1411.350 2691.680 1411.670 2691.740 ;
        RECT 1835.470 2691.680 1835.790 2691.740 ;
        RECT 1411.350 2691.540 1835.790 2691.680 ;
        RECT 1411.350 2691.480 1411.670 2691.540 ;
        RECT 1835.470 2691.480 1835.790 2691.540 ;
        RECT 1414.110 2691.340 1414.430 2691.400 ;
        RECT 1842.370 2691.340 1842.690 2691.400 ;
        RECT 1414.110 2691.200 1842.690 2691.340 ;
        RECT 1414.110 2691.140 1414.430 2691.200 ;
        RECT 1842.370 2691.140 1842.690 2691.200 ;
        RECT 1414.110 2684.200 1414.430 2684.260 ;
        RECT 1849.270 2684.200 1849.590 2684.260 ;
        RECT 1414.110 2684.060 1849.590 2684.200 ;
        RECT 1414.110 2684.000 1414.430 2684.060 ;
        RECT 1849.270 2684.000 1849.590 2684.060 ;
        RECT 1414.110 2677.400 1414.430 2677.460 ;
        RECT 1856.170 2677.400 1856.490 2677.460 ;
        RECT 1414.110 2677.260 1856.490 2677.400 ;
        RECT 1414.110 2677.200 1414.430 2677.260 ;
        RECT 1856.170 2677.200 1856.490 2677.260 ;
        RECT 1408.590 2670.940 1408.910 2671.000 ;
        RECT 1863.070 2670.940 1863.390 2671.000 ;
        RECT 1408.590 2670.800 1863.390 2670.940 ;
        RECT 1408.590 2670.740 1408.910 2670.800 ;
        RECT 1863.070 2670.740 1863.390 2670.800 ;
        RECT 1410.430 2670.600 1410.750 2670.660 ;
        RECT 1869.970 2670.600 1870.290 2670.660 ;
        RECT 1410.430 2670.460 1870.290 2670.600 ;
        RECT 1410.430 2670.400 1410.750 2670.460 ;
        RECT 1869.970 2670.400 1870.290 2670.460 ;
        RECT 1410.430 2663.800 1410.750 2663.860 ;
        RECT 1876.870 2663.800 1877.190 2663.860 ;
        RECT 1410.430 2663.660 1877.190 2663.800 ;
        RECT 1410.430 2663.600 1410.750 2663.660 ;
        RECT 1876.870 2663.600 1877.190 2663.660 ;
        RECT 1411.350 2657.000 1411.670 2657.060 ;
        RECT 1877.330 2657.000 1877.650 2657.060 ;
        RECT 1411.350 2656.860 1877.650 2657.000 ;
        RECT 1411.350 2656.800 1411.670 2656.860 ;
        RECT 1877.330 2656.800 1877.650 2656.860 ;
        RECT 1414.110 2656.660 1414.430 2656.720 ;
        RECT 1883.770 2656.660 1884.090 2656.720 ;
        RECT 1414.110 2656.520 1884.090 2656.660 ;
        RECT 1414.110 2656.460 1414.430 2656.520 ;
        RECT 1883.770 2656.460 1884.090 2656.520 ;
        RECT 1414.110 2649.860 1414.430 2649.920 ;
        RECT 1891.130 2649.860 1891.450 2649.920 ;
        RECT 1414.110 2649.720 1891.450 2649.860 ;
        RECT 1414.110 2649.660 1414.430 2649.720 ;
        RECT 1891.130 2649.660 1891.450 2649.720 ;
        RECT 1414.110 2643.060 1414.430 2643.120 ;
        RECT 1898.030 2643.060 1898.350 2643.120 ;
        RECT 1414.110 2642.920 1898.350 2643.060 ;
        RECT 1414.110 2642.860 1414.430 2642.920 ;
        RECT 1898.030 2642.860 1898.350 2642.920 ;
        RECT 1414.110 2636.260 1414.430 2636.320 ;
        RECT 1880.090 2636.260 1880.410 2636.320 ;
        RECT 1414.110 2636.120 1880.410 2636.260 ;
        RECT 1414.110 2636.060 1414.430 2636.120 ;
        RECT 1880.090 2636.060 1880.410 2636.120 ;
        RECT 1411.350 2635.920 1411.670 2635.980 ;
        RECT 1904.930 2635.920 1905.250 2635.980 ;
        RECT 1411.350 2635.780 1905.250 2635.920 ;
        RECT 1411.350 2635.720 1411.670 2635.780 ;
        RECT 1904.930 2635.720 1905.250 2635.780 ;
        RECT 1409.510 2629.120 1409.830 2629.180 ;
        RECT 1873.190 2629.120 1873.510 2629.180 ;
        RECT 1409.510 2628.980 1873.510 2629.120 ;
        RECT 1409.510 2628.920 1409.830 2628.980 ;
        RECT 1873.190 2628.920 1873.510 2628.980 ;
        RECT 1414.110 2622.320 1414.430 2622.380 ;
        RECT 1859.390 2622.320 1859.710 2622.380 ;
        RECT 1414.110 2622.180 1859.710 2622.320 ;
        RECT 1414.110 2622.120 1414.430 2622.180 ;
        RECT 1859.390 2622.120 1859.710 2622.180 ;
        RECT 1414.110 2615.520 1414.430 2615.580 ;
        RECT 1770.610 2615.520 1770.930 2615.580 ;
        RECT 1414.110 2615.380 1770.930 2615.520 ;
        RECT 1414.110 2615.320 1414.430 2615.380 ;
        RECT 1770.610 2615.320 1770.930 2615.380 ;
        RECT 1411.810 2615.180 1412.130 2615.240 ;
        RECT 1838.690 2615.180 1839.010 2615.240 ;
        RECT 1411.810 2615.040 1839.010 2615.180 ;
        RECT 1411.810 2614.980 1412.130 2615.040 ;
        RECT 1838.690 2614.980 1839.010 2615.040 ;
        RECT 1414.110 2608.380 1414.430 2608.440 ;
        RECT 1939.430 2608.380 1939.750 2608.440 ;
        RECT 1414.110 2608.240 1939.750 2608.380 ;
        RECT 1414.110 2608.180 1414.430 2608.240 ;
        RECT 1939.430 2608.180 1939.750 2608.240 ;
        RECT 1414.110 2601.580 1414.430 2601.640 ;
        RECT 1953.230 2601.580 1953.550 2601.640 ;
        RECT 1414.110 2601.440 1953.550 2601.580 ;
        RECT 1414.110 2601.380 1414.430 2601.440 ;
        RECT 1953.230 2601.380 1953.550 2601.440 ;
        RECT 1408.590 2595.460 1408.910 2595.520 ;
        RECT 1418.710 2595.460 1419.030 2595.520 ;
        RECT 1408.590 2595.320 1419.030 2595.460 ;
        RECT 1408.590 2595.260 1408.910 2595.320 ;
        RECT 1418.710 2595.260 1419.030 2595.320 ;
        RECT 1410.430 2587.640 1410.750 2587.700 ;
        RECT 1960.130 2587.640 1960.450 2587.700 ;
        RECT 1410.430 2587.500 1960.450 2587.640 ;
        RECT 1410.430 2587.440 1410.750 2587.500 ;
        RECT 1960.130 2587.440 1960.450 2587.500 ;
        RECT 1411.350 2581.180 1411.670 2581.240 ;
        RECT 1935.290 2581.180 1935.610 2581.240 ;
        RECT 1411.350 2581.040 1935.610 2581.180 ;
        RECT 1411.350 2580.980 1411.670 2581.040 ;
        RECT 1935.290 2580.980 1935.610 2581.040 ;
        RECT 1414.110 2580.840 1414.430 2580.900 ;
        RECT 2097.670 2580.840 2097.990 2580.900 ;
        RECT 1414.110 2580.700 2097.990 2580.840 ;
        RECT 1414.110 2580.640 1414.430 2580.700 ;
        RECT 2097.670 2580.640 2097.990 2580.700 ;
        RECT 1414.110 2574.040 1414.430 2574.100 ;
        RECT 1928.390 2574.040 1928.710 2574.100 ;
        RECT 1414.110 2573.900 1928.710 2574.040 ;
        RECT 1414.110 2573.840 1414.430 2573.900 ;
        RECT 1928.390 2573.840 1928.710 2573.900 ;
        RECT 1411.350 2566.900 1411.670 2566.960 ;
        RECT 2098.130 2566.900 2098.450 2566.960 ;
        RECT 1411.350 2566.760 2098.450 2566.900 ;
        RECT 1411.350 2566.700 1411.670 2566.760 ;
        RECT 2098.130 2566.700 2098.450 2566.760 ;
        RECT 1413.650 2560.440 1413.970 2560.500 ;
        RECT 1928.850 2560.440 1929.170 2560.500 ;
        RECT 1413.650 2560.300 1929.170 2560.440 ;
        RECT 1413.650 2560.240 1413.970 2560.300 ;
        RECT 1928.850 2560.240 1929.170 2560.300 ;
        RECT 1414.110 2560.100 1414.430 2560.160 ;
        RECT 2098.590 2560.100 2098.910 2560.160 ;
        RECT 1414.110 2559.960 2098.910 2560.100 ;
        RECT 1414.110 2559.900 1414.430 2559.960 ;
        RECT 2098.590 2559.900 2098.910 2559.960 ;
        RECT 1408.590 2553.300 1408.910 2553.360 ;
        RECT 1921.490 2553.300 1921.810 2553.360 ;
        RECT 1408.590 2553.160 1921.810 2553.300 ;
        RECT 1408.590 2553.100 1408.910 2553.160 ;
        RECT 1921.490 2553.100 1921.810 2553.160 ;
        RECT 1411.350 2546.500 1411.670 2546.560 ;
        RECT 2099.050 2546.500 2099.370 2546.560 ;
        RECT 1411.350 2546.360 2099.370 2546.500 ;
        RECT 1411.350 2546.300 1411.670 2546.360 ;
        RECT 2099.050 2546.300 2099.370 2546.360 ;
        RECT 1412.730 2539.700 1413.050 2539.760 ;
        RECT 1914.590 2539.700 1914.910 2539.760 ;
        RECT 1412.730 2539.560 1914.910 2539.700 ;
        RECT 1412.730 2539.500 1413.050 2539.560 ;
        RECT 1914.590 2539.500 1914.910 2539.560 ;
        RECT 1414.110 2539.360 1414.430 2539.420 ;
        RECT 2099.510 2539.360 2099.830 2539.420 ;
        RECT 1414.110 2539.220 2099.830 2539.360 ;
        RECT 1414.110 2539.160 1414.430 2539.220 ;
        RECT 2099.510 2539.160 2099.830 2539.220 ;
        RECT 1410.430 2532.560 1410.750 2532.620 ;
        RECT 1915.050 2532.560 1915.370 2532.620 ;
        RECT 1410.430 2532.420 1915.370 2532.560 ;
        RECT 1410.430 2532.360 1410.750 2532.420 ;
        RECT 1915.050 2532.360 1915.370 2532.420 ;
        RECT 1414.110 2526.100 1414.430 2526.160 ;
        RECT 1915.510 2526.100 1915.830 2526.160 ;
        RECT 1414.110 2525.960 1915.830 2526.100 ;
        RECT 1414.110 2525.900 1414.430 2525.960 ;
        RECT 1915.510 2525.900 1915.830 2525.960 ;
        RECT 1413.650 2525.760 1413.970 2525.820 ;
        RECT 2099.970 2525.760 2100.290 2525.820 ;
        RECT 1413.650 2525.620 2100.290 2525.760 ;
        RECT 1413.650 2525.560 1413.970 2525.620 ;
        RECT 2099.970 2525.560 2100.290 2525.620 ;
        RECT 1414.110 2518.620 1414.430 2518.680 ;
        RECT 2100.430 2518.620 2100.750 2518.680 ;
        RECT 1414.110 2518.480 2100.750 2518.620 ;
        RECT 1414.110 2518.420 1414.430 2518.480 ;
        RECT 2100.430 2518.420 2100.750 2518.480 ;
        RECT 1414.110 2511.820 1414.430 2511.880 ;
        RECT 1915.970 2511.820 1916.290 2511.880 ;
        RECT 1414.110 2511.680 1916.290 2511.820 ;
        RECT 1414.110 2511.620 1414.430 2511.680 ;
        RECT 1915.970 2511.620 1916.290 2511.680 ;
        RECT 1414.110 2505.360 1414.430 2505.420 ;
        RECT 1893.890 2505.360 1894.210 2505.420 ;
        RECT 1414.110 2505.220 1894.210 2505.360 ;
        RECT 1414.110 2505.160 1414.430 2505.220 ;
        RECT 1893.890 2505.160 1894.210 2505.220 ;
        RECT 1411.350 2505.020 1411.670 2505.080 ;
        RECT 2052.590 2505.020 2052.910 2505.080 ;
        RECT 1411.350 2504.880 2052.910 2505.020 ;
        RECT 1411.350 2504.820 1411.670 2504.880 ;
        RECT 2052.590 2504.820 2052.910 2504.880 ;
        RECT 1414.110 2491.080 1414.430 2491.140 ;
        RECT 1419.630 2491.080 1419.950 2491.140 ;
        RECT 1414.110 2490.940 1419.950 2491.080 ;
        RECT 1414.110 2490.880 1414.430 2490.940 ;
        RECT 1419.630 2490.880 1419.950 2490.940 ;
        RECT 1414.110 2484.280 1414.430 2484.340 ;
        RECT 2081.570 2484.280 2081.890 2484.340 ;
        RECT 1414.110 2484.140 2081.890 2484.280 ;
        RECT 1414.110 2484.080 1414.430 2484.140 ;
        RECT 2081.570 2484.080 2081.890 2484.140 ;
        RECT 1409.510 2477.480 1409.830 2477.540 ;
        RECT 2494.190 2477.480 2494.510 2477.540 ;
        RECT 1409.510 2477.340 2494.510 2477.480 ;
        RECT 1409.510 2477.280 1409.830 2477.340 ;
        RECT 2494.190 2477.280 2494.510 2477.340 ;
        RECT 1414.110 2470.340 1414.430 2470.400 ;
        RECT 2480.390 2470.340 2480.710 2470.400 ;
        RECT 1414.110 2470.200 2480.710 2470.340 ;
        RECT 1414.110 2470.140 1414.430 2470.200 ;
        RECT 2480.390 2470.140 2480.710 2470.200 ;
        RECT 1414.110 2463.880 1414.430 2463.940 ;
        RECT 2459.690 2463.880 2460.010 2463.940 ;
        RECT 1414.110 2463.740 2460.010 2463.880 ;
        RECT 1414.110 2463.680 1414.430 2463.740 ;
        RECT 2459.690 2463.680 2460.010 2463.740 ;
        RECT 1411.810 2463.540 1412.130 2463.600 ;
        RECT 2466.590 2463.540 2466.910 2463.600 ;
        RECT 1411.810 2463.400 2466.910 2463.540 ;
        RECT 1411.810 2463.340 1412.130 2463.400 ;
        RECT 2466.590 2463.340 2466.910 2463.400 ;
        RECT 1414.110 2456.740 1414.430 2456.800 ;
        RECT 2445.890 2456.740 2446.210 2456.800 ;
        RECT 1414.110 2456.600 2446.210 2456.740 ;
        RECT 1414.110 2456.540 1414.430 2456.600 ;
        RECT 2445.890 2456.540 2446.210 2456.600 ;
        RECT 1414.110 2449.940 1414.430 2450.000 ;
        RECT 2418.290 2449.940 2418.610 2450.000 ;
        RECT 1414.110 2449.800 2418.610 2449.940 ;
        RECT 1414.110 2449.740 1414.430 2449.800 ;
        RECT 2418.290 2449.740 2418.610 2449.800 ;
        RECT 1411.350 2449.600 1411.670 2449.660 ;
        RECT 2425.190 2449.600 2425.510 2449.660 ;
        RECT 1411.350 2449.460 2425.510 2449.600 ;
        RECT 1411.350 2449.400 1411.670 2449.460 ;
        RECT 2425.190 2449.400 2425.510 2449.460 ;
        RECT 1411.350 2442.800 1411.670 2442.860 ;
        RECT 2411.390 2442.800 2411.710 2442.860 ;
        RECT 1411.350 2442.660 2411.710 2442.800 ;
        RECT 1411.350 2442.600 1411.670 2442.660 ;
        RECT 2411.390 2442.600 2411.710 2442.660 ;
        RECT 1414.110 2436.000 1414.430 2436.060 ;
        RECT 2404.490 2436.000 2404.810 2436.060 ;
        RECT 1414.110 2435.860 2404.810 2436.000 ;
        RECT 1414.110 2435.800 1414.430 2435.860 ;
        RECT 2404.490 2435.800 2404.810 2435.860 ;
        RECT 1414.110 2429.540 1414.430 2429.600 ;
        RECT 2328.590 2429.540 2328.910 2429.600 ;
        RECT 1414.110 2429.400 2328.910 2429.540 ;
        RECT 1414.110 2429.340 1414.430 2429.400 ;
        RECT 2328.590 2429.340 2328.910 2429.400 ;
        RECT 1411.350 2429.200 1411.670 2429.260 ;
        RECT 2335.490 2429.200 2335.810 2429.260 ;
        RECT 1411.350 2429.060 2335.810 2429.200 ;
        RECT 1411.350 2429.000 1411.670 2429.060 ;
        RECT 2335.490 2429.000 2335.810 2429.060 ;
        RECT 1408.590 2422.060 1408.910 2422.120 ;
        RECT 2245.790 2422.060 2246.110 2422.120 ;
        RECT 1408.590 2421.920 2246.110 2422.060 ;
        RECT 1408.590 2421.860 1408.910 2421.920 ;
        RECT 2245.790 2421.860 2246.110 2421.920 ;
        RECT 1411.350 2415.260 1411.670 2415.320 ;
        RECT 2231.990 2415.260 2232.310 2415.320 ;
        RECT 1411.350 2415.120 2232.310 2415.260 ;
        RECT 1411.350 2415.060 1411.670 2415.120 ;
        RECT 2231.990 2415.060 2232.310 2415.120 ;
        RECT 1414.110 2408.800 1414.430 2408.860 ;
        RECT 2211.290 2408.800 2211.610 2408.860 ;
        RECT 1414.110 2408.660 2211.610 2408.800 ;
        RECT 1414.110 2408.600 1414.430 2408.660 ;
        RECT 2211.290 2408.600 2211.610 2408.660 ;
        RECT 1412.730 2408.460 1413.050 2408.520 ;
        RECT 2225.090 2408.460 2225.410 2408.520 ;
        RECT 1412.730 2408.320 2225.410 2408.460 ;
        RECT 1412.730 2408.260 1413.050 2408.320 ;
        RECT 2225.090 2408.260 2225.410 2408.320 ;
        RECT 1410.430 2401.320 1410.750 2401.380 ;
        RECT 2176.790 2401.320 2177.110 2401.380 ;
        RECT 1410.430 2401.180 2177.110 2401.320 ;
        RECT 1410.430 2401.120 1410.750 2401.180 ;
        RECT 2176.790 2401.120 2177.110 2401.180 ;
        RECT 1414.110 2394.860 1414.430 2394.920 ;
        RECT 2156.090 2394.860 2156.410 2394.920 ;
        RECT 1414.110 2394.720 2156.410 2394.860 ;
        RECT 1414.110 2394.660 1414.430 2394.720 ;
        RECT 2156.090 2394.660 2156.410 2394.720 ;
        RECT 1413.650 2394.520 1413.970 2394.580 ;
        RECT 2169.890 2394.520 2170.210 2394.580 ;
        RECT 1413.650 2394.380 2170.210 2394.520 ;
        RECT 1413.650 2394.320 1413.970 2394.380 ;
        RECT 2169.890 2394.320 2170.210 2394.380 ;
        RECT 1414.110 2387.720 1414.430 2387.780 ;
        RECT 2149.190 2387.720 2149.510 2387.780 ;
        RECT 1414.110 2387.580 2149.510 2387.720 ;
        RECT 1414.110 2387.520 1414.430 2387.580 ;
        RECT 2149.190 2387.520 2149.510 2387.580 ;
        RECT 1410.430 2380.580 1410.750 2380.640 ;
        RECT 2142.290 2380.580 2142.610 2380.640 ;
        RECT 1410.430 2380.440 2142.610 2380.580 ;
        RECT 1410.430 2380.380 1410.750 2380.440 ;
        RECT 2142.290 2380.380 2142.610 2380.440 ;
        RECT 1414.110 2374.120 1414.430 2374.180 ;
        RECT 2121.590 2374.120 2121.910 2374.180 ;
        RECT 1414.110 2373.980 2121.910 2374.120 ;
        RECT 1414.110 2373.920 1414.430 2373.980 ;
        RECT 2121.590 2373.920 2121.910 2373.980 ;
        RECT 1411.350 2373.780 1411.670 2373.840 ;
        RECT 2135.390 2373.780 2135.710 2373.840 ;
        RECT 1411.350 2373.640 2135.710 2373.780 ;
        RECT 1411.350 2373.580 1411.670 2373.640 ;
        RECT 2135.390 2373.580 2135.710 2373.640 ;
        RECT 1408.590 2366.980 1408.910 2367.040 ;
        RECT 2080.190 2366.980 2080.510 2367.040 ;
        RECT 1408.590 2366.840 2080.510 2366.980 ;
        RECT 1408.590 2366.780 1408.910 2366.840 ;
        RECT 2080.190 2366.780 2080.510 2366.840 ;
        RECT 1410.430 2360.180 1410.750 2360.240 ;
        RECT 2387.930 2360.180 2388.250 2360.240 ;
        RECT 1410.430 2360.040 2388.250 2360.180 ;
        RECT 1410.430 2359.980 1410.750 2360.040 ;
        RECT 2387.930 2359.980 2388.250 2360.040 ;
        RECT 1414.110 2353.380 1414.430 2353.440 ;
        RECT 2045.690 2353.380 2046.010 2353.440 ;
        RECT 1414.110 2353.240 2046.010 2353.380 ;
        RECT 1414.110 2353.180 1414.430 2353.240 ;
        RECT 2045.690 2353.180 2046.010 2353.240 ;
        RECT 1413.650 2353.040 1413.970 2353.100 ;
        RECT 2059.490 2353.040 2059.810 2353.100 ;
        RECT 1413.650 2352.900 2059.810 2353.040 ;
        RECT 1413.650 2352.840 1413.970 2352.900 ;
        RECT 2059.490 2352.840 2059.810 2352.900 ;
        RECT 1409.510 2346.240 1409.830 2346.300 ;
        RECT 2374.130 2346.240 2374.450 2346.300 ;
        RECT 1409.510 2346.100 2374.450 2346.240 ;
        RECT 1409.510 2346.040 1409.830 2346.100 ;
        RECT 2374.130 2346.040 2374.450 2346.100 ;
        RECT 1414.110 2339.440 1414.430 2339.500 ;
        RECT 2367.230 2339.440 2367.550 2339.500 ;
        RECT 1414.110 2339.300 2367.550 2339.440 ;
        RECT 1414.110 2339.240 1414.430 2339.300 ;
        RECT 2367.230 2339.240 2367.550 2339.300 ;
        RECT 1413.650 2332.640 1413.970 2332.700 ;
        RECT 2031.890 2332.640 2032.210 2332.700 ;
        RECT 1413.650 2332.500 2032.210 2332.640 ;
        RECT 1413.650 2332.440 1413.970 2332.500 ;
        RECT 2031.890 2332.440 2032.210 2332.500 ;
        RECT 1414.110 2332.300 1414.430 2332.360 ;
        RECT 2353.430 2332.300 2353.750 2332.360 ;
        RECT 1414.110 2332.160 2353.750 2332.300 ;
        RECT 1414.110 2332.100 1414.430 2332.160 ;
        RECT 2353.430 2332.100 2353.750 2332.160 ;
        RECT 1414.110 2325.500 1414.430 2325.560 ;
        RECT 2238.890 2325.500 2239.210 2325.560 ;
        RECT 1414.110 2325.360 2239.210 2325.500 ;
        RECT 1414.110 2325.300 1414.430 2325.360 ;
        RECT 2238.890 2325.300 2239.210 2325.360 ;
        RECT 1413.650 2319.040 1413.970 2319.100 ;
        RECT 2087.090 2319.040 2087.410 2319.100 ;
        RECT 1413.650 2318.900 2087.410 2319.040 ;
        RECT 1413.650 2318.840 1413.970 2318.900 ;
        RECT 2087.090 2318.840 2087.410 2318.900 ;
        RECT 1414.110 2318.700 1414.430 2318.760 ;
        RECT 2631.730 2318.700 2632.050 2318.760 ;
        RECT 1414.110 2318.560 2632.050 2318.700 ;
        RECT 1414.110 2318.500 1414.430 2318.560 ;
        RECT 2631.730 2318.500 2632.050 2318.560 ;
        RECT 1414.110 2311.900 1414.430 2311.960 ;
        RECT 1418.250 2311.900 1418.570 2311.960 ;
        RECT 1414.110 2311.760 1418.570 2311.900 ;
        RECT 1414.110 2311.700 1414.430 2311.760 ;
        RECT 1418.250 2311.700 1418.570 2311.760 ;
        RECT 1414.110 2304.760 1414.430 2304.820 ;
        RECT 1842.830 2304.760 1843.150 2304.820 ;
        RECT 1414.110 2304.620 1843.150 2304.760 ;
        RECT 1414.110 2304.560 1414.430 2304.620 ;
        RECT 1842.830 2304.560 1843.150 2304.620 ;
        RECT 1413.650 2298.300 1413.970 2298.360 ;
        RECT 1419.170 2298.300 1419.490 2298.360 ;
        RECT 1413.650 2298.160 1419.490 2298.300 ;
        RECT 1413.650 2298.100 1413.970 2298.160 ;
        RECT 1419.170 2298.100 1419.490 2298.160 ;
        RECT 1414.110 2297.960 1414.430 2298.020 ;
        RECT 1849.730 2297.960 1850.050 2298.020 ;
        RECT 1414.110 2297.820 1850.050 2297.960 ;
        RECT 1414.110 2297.760 1414.430 2297.820 ;
        RECT 1849.730 2297.760 1850.050 2297.820 ;
        RECT 1408.590 2291.160 1408.910 2291.220 ;
        RECT 1420.090 2291.160 1420.410 2291.220 ;
        RECT 1408.590 2291.020 1420.410 2291.160 ;
        RECT 1408.590 2290.960 1408.910 2291.020 ;
        RECT 1420.090 2290.960 1420.410 2291.020 ;
        RECT 1410.430 2284.020 1410.750 2284.080 ;
        RECT 1420.550 2284.020 1420.870 2284.080 ;
        RECT 1410.430 2283.880 1420.870 2284.020 ;
        RECT 1410.430 2283.820 1410.750 2283.880 ;
        RECT 1420.550 2283.820 1420.870 2283.880 ;
        RECT 1408.130 2277.560 1408.450 2277.620 ;
        RECT 1421.010 2277.560 1421.330 2277.620 ;
        RECT 1408.130 2277.420 1421.330 2277.560 ;
        RECT 1408.130 2277.360 1408.450 2277.420 ;
        RECT 1421.010 2277.360 1421.330 2277.420 ;
        RECT 1414.110 2277.220 1414.430 2277.280 ;
        RECT 1877.790 2277.220 1878.110 2277.280 ;
        RECT 1414.110 2277.080 1878.110 2277.220 ;
        RECT 1414.110 2277.020 1414.430 2277.080 ;
        RECT 1877.790 2277.020 1878.110 2277.080 ;
        RECT 1410.890 2202.080 1411.210 2202.140 ;
        RECT 1921.950 2202.080 1922.270 2202.140 ;
        RECT 1410.890 2201.940 1922.270 2202.080 ;
        RECT 1410.890 2201.880 1411.210 2201.940 ;
        RECT 1921.950 2201.880 1922.270 2201.940 ;
        RECT 1407.210 2201.400 1407.530 2201.460 ;
        RECT 1935.750 2201.400 1936.070 2201.460 ;
        RECT 1407.210 2201.260 1936.070 2201.400 ;
        RECT 1407.210 2201.200 1407.530 2201.260 ;
        RECT 1935.750 2201.200 1936.070 2201.260 ;
        RECT 1410.890 2194.600 1411.210 2194.660 ;
        RECT 1907.690 2194.600 1908.010 2194.660 ;
        RECT 1410.890 2194.460 1908.010 2194.600 ;
        RECT 1410.890 2194.400 1411.210 2194.460 ;
        RECT 1907.690 2194.400 1908.010 2194.460 ;
        RECT 1410.890 2183.040 1411.210 2183.100 ;
        RECT 1410.520 2182.900 1411.210 2183.040 ;
        RECT 1410.520 2180.660 1410.660 2182.900 ;
        RECT 1410.890 2182.840 1411.210 2182.900 ;
        RECT 1410.890 2181.000 1411.210 2181.060 ;
        RECT 1886.990 2181.000 1887.310 2181.060 ;
        RECT 1410.890 2180.860 1887.310 2181.000 ;
        RECT 1410.890 2180.800 1411.210 2180.860 ;
        RECT 1886.990 2180.800 1887.310 2180.860 ;
        RECT 1900.790 2180.660 1901.110 2180.720 ;
        RECT 1410.520 2180.520 1901.110 2180.660 ;
        RECT 1900.790 2180.460 1901.110 2180.520 ;
        RECT 1410.890 2173.860 1411.210 2173.920 ;
        RECT 1873.650 2173.860 1873.970 2173.920 ;
        RECT 1410.890 2173.720 1873.970 2173.860 ;
        RECT 1410.890 2173.660 1411.210 2173.720 ;
        RECT 1873.650 2173.660 1873.970 2173.720 ;
        RECT 1410.890 2166.720 1411.210 2166.780 ;
        RECT 1866.290 2166.720 1866.610 2166.780 ;
        RECT 1410.890 2166.580 1866.610 2166.720 ;
        RECT 1410.890 2166.520 1411.210 2166.580 ;
        RECT 1866.290 2166.520 1866.610 2166.580 ;
        RECT 1410.445 2157.880 1410.735 2157.925 ;
        RECT 1411.350 2157.880 1411.670 2157.940 ;
        RECT 1410.445 2157.740 1411.670 2157.880 ;
        RECT 1410.445 2157.695 1410.735 2157.740 ;
        RECT 1411.350 2157.680 1411.670 2157.740 ;
        RECT 1411.350 2153.460 1411.670 2153.520 ;
        RECT 1942.190 2153.460 1942.510 2153.520 ;
        RECT 1411.350 2153.320 1942.510 2153.460 ;
        RECT 1411.350 2153.260 1411.670 2153.320 ;
        RECT 1942.190 2153.260 1942.510 2153.320 ;
        RECT 1411.350 2152.780 1411.670 2152.840 ;
        RECT 2321.690 2152.780 2322.010 2152.840 ;
        RECT 1411.350 2152.640 2322.010 2152.780 ;
        RECT 1411.350 2152.580 1411.670 2152.640 ;
        RECT 2321.690 2152.580 2322.010 2152.640 ;
        RECT 1407.210 2145.980 1407.530 2146.040 ;
        RECT 2083.870 2145.980 2084.190 2146.040 ;
        RECT 1407.210 2145.840 2084.190 2145.980 ;
        RECT 1407.210 2145.780 1407.530 2145.840 ;
        RECT 2083.870 2145.780 2084.190 2145.840 ;
        RECT 1411.350 2145.640 1411.670 2145.700 ;
        RECT 1790.850 2145.640 1791.170 2145.700 ;
        RECT 1411.350 2145.500 1791.170 2145.640 ;
        RECT 1411.350 2145.440 1411.670 2145.500 ;
        RECT 1790.850 2145.440 1791.170 2145.500 ;
        RECT 1411.350 2138.840 1411.670 2138.900 ;
        RECT 1790.390 2138.840 1790.710 2138.900 ;
        RECT 1411.350 2138.700 1790.710 2138.840 ;
        RECT 1411.350 2138.640 1411.670 2138.700 ;
        RECT 1790.390 2138.640 1790.710 2138.700 ;
        RECT 1783.950 2138.500 1784.270 2138.560 ;
        RECT 1415.580 2138.360 1784.270 2138.500 ;
        RECT 1415.580 2136.800 1415.720 2138.360 ;
        RECT 1783.950 2138.300 1784.270 2138.360 ;
        RECT 1410.980 2136.660 1415.720 2136.800 ;
        RECT 1410.980 2136.120 1411.120 2136.660 ;
        RECT 1411.350 2136.120 1411.670 2136.180 ;
        RECT 1410.980 2135.980 1411.670 2136.120 ;
        RECT 1411.350 2135.920 1411.670 2135.980 ;
        RECT 1411.350 2132.040 1411.670 2132.100 ;
        RECT 1783.490 2132.040 1783.810 2132.100 ;
        RECT 1411.350 2131.900 1783.810 2132.040 ;
        RECT 1411.350 2131.840 1411.670 2131.900 ;
        RECT 1783.490 2131.840 1783.810 2131.900 ;
        RECT 1411.350 2125.240 1411.670 2125.300 ;
        RECT 1777.050 2125.240 1777.370 2125.300 ;
        RECT 1411.350 2125.100 1777.370 2125.240 ;
        RECT 1411.350 2125.040 1411.670 2125.100 ;
        RECT 1777.050 2125.040 1777.370 2125.100 ;
        RECT 1411.350 2118.100 1411.670 2118.160 ;
        RECT 1776.590 2118.100 1776.910 2118.160 ;
        RECT 1411.350 2117.960 1776.910 2118.100 ;
        RECT 1411.350 2117.900 1411.670 2117.960 ;
        RECT 1776.590 2117.900 1776.910 2117.960 ;
        RECT 1770.150 2117.760 1770.470 2117.820 ;
        RECT 1410.980 2117.620 1770.470 2117.760 ;
        RECT 1410.980 2116.400 1411.120 2117.620 ;
        RECT 1770.150 2117.560 1770.470 2117.620 ;
        RECT 1411.350 2116.400 1411.670 2116.460 ;
        RECT 1410.980 2116.260 1411.670 2116.400 ;
        RECT 1411.350 2116.200 1411.670 2116.260 ;
        RECT 1411.350 2111.300 1411.670 2111.360 ;
        RECT 1769.690 2111.300 1770.010 2111.360 ;
        RECT 1411.350 2111.160 1770.010 2111.300 ;
        RECT 1411.350 2111.100 1411.670 2111.160 ;
        RECT 1769.690 2111.100 1770.010 2111.160 ;
        RECT 1408.130 2106.880 1408.450 2106.940 ;
        RECT 1407.935 2106.740 1408.450 2106.880 ;
        RECT 1408.130 2106.680 1408.450 2106.740 ;
        RECT 1408.130 2106.200 1408.450 2106.260 ;
        RECT 1412.270 2106.200 1412.590 2106.260 ;
        RECT 1408.130 2106.060 1412.590 2106.200 ;
        RECT 1408.130 2106.000 1408.450 2106.060 ;
        RECT 1412.270 2106.000 1412.590 2106.060 ;
        RECT 1412.270 2105.180 1412.590 2105.240 ;
        RECT 1414.110 2105.180 1414.430 2105.240 ;
        RECT 1412.270 2105.040 1414.430 2105.180 ;
        RECT 1412.270 2104.980 1412.590 2105.040 ;
        RECT 1414.110 2104.980 1414.430 2105.040 ;
        RECT 1414.110 2104.500 1414.430 2104.560 ;
        RECT 1763.250 2104.500 1763.570 2104.560 ;
        RECT 1414.110 2104.360 1763.570 2104.500 ;
        RECT 1414.110 2104.300 1414.430 2104.360 ;
        RECT 1763.250 2104.300 1763.570 2104.360 ;
        RECT 1412.730 2097.360 1413.050 2097.420 ;
        RECT 2380.570 2097.360 2380.890 2097.420 ;
        RECT 1412.730 2097.220 2380.890 2097.360 ;
        RECT 1412.730 2097.160 1413.050 2097.220 ;
        RECT 2380.570 2097.160 2380.890 2097.220 ;
        RECT 1414.110 2097.020 1414.430 2097.080 ;
        RECT 1762.790 2097.020 1763.110 2097.080 ;
        RECT 1414.110 2096.880 1763.110 2097.020 ;
        RECT 1414.110 2096.820 1414.430 2096.880 ;
        RECT 1762.790 2096.820 1763.110 2096.880 ;
        RECT 1414.110 2090.560 1414.430 2090.620 ;
        RECT 2373.670 2090.560 2373.990 2090.620 ;
        RECT 1414.110 2090.420 2373.990 2090.560 ;
        RECT 1414.110 2090.360 1414.430 2090.420 ;
        RECT 2373.670 2090.360 2373.990 2090.420 ;
        RECT 1411.350 2088.860 1411.670 2088.920 ;
        RECT 1412.730 2088.860 1413.050 2088.920 ;
        RECT 1411.350 2088.720 1413.050 2088.860 ;
        RECT 1411.350 2088.660 1411.670 2088.720 ;
        RECT 1412.730 2088.660 1413.050 2088.720 ;
        RECT 1410.445 2088.180 1410.735 2088.225 ;
        RECT 1411.350 2088.180 1411.670 2088.240 ;
        RECT 1410.445 2088.040 1411.670 2088.180 ;
        RECT 1410.445 2087.995 1410.735 2088.040 ;
        RECT 1411.350 2087.980 1411.670 2088.040 ;
        RECT 1414.110 2083.760 1414.430 2083.820 ;
        RECT 2366.770 2083.760 2367.090 2083.820 ;
        RECT 1414.110 2083.620 2367.090 2083.760 ;
        RECT 1414.110 2083.560 1414.430 2083.620 ;
        RECT 2366.770 2083.560 2367.090 2083.620 ;
        RECT 1422.850 2082.060 1423.170 2082.120 ;
        RECT 2266.490 2082.060 2266.810 2082.120 ;
        RECT 1422.850 2081.920 2266.810 2082.060 ;
        RECT 1422.850 2081.860 1423.170 2081.920 ;
        RECT 2266.490 2081.860 2266.810 2081.920 ;
        RECT 1431.130 2081.720 1431.450 2081.780 ;
        RECT 2277.070 2081.720 2277.390 2081.780 ;
        RECT 1431.130 2081.580 2277.390 2081.720 ;
        RECT 1431.130 2081.520 1431.450 2081.580 ;
        RECT 2277.070 2081.520 2277.390 2081.580 ;
        RECT 1430.670 2081.380 1430.990 2081.440 ;
        RECT 2283.970 2081.380 2284.290 2081.440 ;
        RECT 1430.670 2081.240 2284.290 2081.380 ;
        RECT 1430.670 2081.180 1430.990 2081.240 ;
        RECT 2283.970 2081.180 2284.290 2081.240 ;
        RECT 1416.410 2081.040 1416.730 2081.100 ;
        RECT 2290.870 2081.040 2291.190 2081.100 ;
        RECT 1416.410 2080.900 2291.190 2081.040 ;
        RECT 1416.410 2080.840 1416.730 2080.900 ;
        RECT 2290.870 2080.840 2291.190 2080.900 ;
        RECT 1415.950 2080.700 1416.270 2080.760 ;
        RECT 2297.770 2080.700 2298.090 2080.760 ;
        RECT 1415.950 2080.560 2298.090 2080.700 ;
        RECT 1415.950 2080.500 1416.270 2080.560 ;
        RECT 2297.770 2080.500 2298.090 2080.560 ;
        RECT 1415.490 2080.360 1415.810 2080.420 ;
        RECT 2305.130 2080.360 2305.450 2080.420 ;
        RECT 1415.490 2080.220 2305.450 2080.360 ;
        RECT 1415.490 2080.160 1415.810 2080.220 ;
        RECT 2305.130 2080.160 2305.450 2080.220 ;
        RECT 1411.350 2077.300 1411.670 2077.360 ;
        RECT 1414.570 2077.300 1414.890 2077.360 ;
        RECT 1411.350 2077.160 1414.890 2077.300 ;
        RECT 1411.350 2077.100 1411.670 2077.160 ;
        RECT 1414.570 2077.100 1414.890 2077.160 ;
        RECT 1414.110 2076.960 1414.430 2077.020 ;
        RECT 2359.870 2076.960 2360.190 2077.020 ;
        RECT 1414.110 2076.820 2360.190 2076.960 ;
        RECT 1414.110 2076.760 1414.430 2076.820 ;
        RECT 2359.870 2076.760 2360.190 2076.820 ;
        RECT 1411.350 2076.620 1411.670 2076.680 ;
        RECT 2352.970 2076.620 2353.290 2076.680 ;
        RECT 1411.350 2076.480 2353.290 2076.620 ;
        RECT 1411.350 2076.420 1411.670 2076.480 ;
        RECT 2352.970 2076.420 2353.290 2076.480 ;
        RECT 1426.990 2076.280 1427.310 2076.340 ;
        RECT 2192.890 2076.280 2193.210 2076.340 ;
        RECT 1426.990 2076.140 2193.210 2076.280 ;
        RECT 1426.990 2076.080 1427.310 2076.140 ;
        RECT 2192.890 2076.080 2193.210 2076.140 ;
        RECT 1426.530 2075.940 1426.850 2076.000 ;
        RECT 2193.350 2075.940 2193.670 2076.000 ;
        RECT 1426.530 2075.800 2193.670 2075.940 ;
        RECT 1426.530 2075.740 1426.850 2075.800 ;
        RECT 2193.350 2075.740 2193.670 2075.800 ;
        RECT 1423.770 2075.600 1424.090 2075.660 ;
        RECT 2190.590 2075.600 2190.910 2075.660 ;
        RECT 1423.770 2075.460 2190.910 2075.600 ;
        RECT 1423.770 2075.400 1424.090 2075.460 ;
        RECT 2190.590 2075.400 2190.910 2075.460 ;
        RECT 1424.230 2075.260 1424.550 2075.320 ;
        RECT 2191.510 2075.260 2191.830 2075.320 ;
        RECT 1424.230 2075.120 2191.830 2075.260 ;
        RECT 1424.230 2075.060 1424.550 2075.120 ;
        RECT 2191.510 2075.060 2191.830 2075.120 ;
        RECT 1423.310 2074.920 1423.630 2074.980 ;
        RECT 2191.050 2074.920 2191.370 2074.980 ;
        RECT 1423.310 2074.780 2191.370 2074.920 ;
        RECT 1423.310 2074.720 1423.630 2074.780 ;
        RECT 2191.050 2074.720 2191.370 2074.780 ;
        RECT 1426.070 2074.580 1426.390 2074.640 ;
        RECT 2228.770 2074.580 2229.090 2074.640 ;
        RECT 1426.070 2074.440 2229.090 2074.580 ;
        RECT 1426.070 2074.380 1426.390 2074.440 ;
        RECT 2228.770 2074.380 2229.090 2074.440 ;
        RECT 1460.110 2074.240 1460.430 2074.300 ;
        RECT 2263.730 2074.240 2264.050 2074.300 ;
        RECT 1460.110 2074.100 2264.050 2074.240 ;
        RECT 1460.110 2074.040 1460.430 2074.100 ;
        RECT 2263.730 2074.040 2264.050 2074.100 ;
        RECT 1415.030 2073.900 1415.350 2073.960 ;
        RECT 2339.630 2073.900 2339.950 2073.960 ;
        RECT 1415.030 2073.760 2339.950 2073.900 ;
        RECT 1415.030 2073.700 1415.350 2073.760 ;
        RECT 2339.630 2073.700 2339.950 2073.760 ;
        RECT 1414.570 2073.560 1414.890 2073.620 ;
        RECT 2346.070 2073.560 2346.390 2073.620 ;
        RECT 1414.570 2073.420 2346.390 2073.560 ;
        RECT 1414.570 2073.360 1414.890 2073.420 ;
        RECT 2346.070 2073.360 2346.390 2073.420 ;
        RECT 1427.450 2073.220 1427.770 2073.280 ;
        RECT 2192.430 2073.220 2192.750 2073.280 ;
        RECT 1427.450 2073.080 2192.750 2073.220 ;
        RECT 1427.450 2073.020 1427.770 2073.080 ;
        RECT 2192.430 2073.020 2192.750 2073.080 ;
        RECT 1427.910 2072.880 1428.230 2072.940 ;
        RECT 2191.970 2072.880 2192.290 2072.940 ;
        RECT 1427.910 2072.740 2192.290 2072.880 ;
        RECT 1427.910 2072.680 1428.230 2072.740 ;
        RECT 2191.970 2072.680 2192.290 2072.740 ;
        RECT 1686.890 2072.540 1687.210 2072.600 ;
        RECT 2270.170 2072.540 2270.490 2072.600 ;
        RECT 1686.890 2072.400 2270.490 2072.540 ;
        RECT 1686.890 2072.340 1687.210 2072.400 ;
        RECT 2270.170 2072.340 2270.490 2072.400 ;
        RECT 1421.930 2072.200 1422.250 2072.260 ;
        RECT 1718.630 2072.200 1718.950 2072.260 ;
        RECT 1421.930 2072.060 1718.950 2072.200 ;
        RECT 1421.930 2072.000 1422.250 2072.060 ;
        RECT 1718.630 2072.000 1718.950 2072.060 ;
        RECT 1422.390 2071.860 1422.710 2071.920 ;
        RECT 1711.270 2071.860 1711.590 2071.920 ;
        RECT 1422.390 2071.720 1711.590 2071.860 ;
        RECT 1422.390 2071.660 1422.710 2071.720 ;
        RECT 1711.270 2071.660 1711.590 2071.720 ;
        RECT 1915.510 2070.160 1915.830 2070.220 ;
        RECT 1922.885 2070.160 1923.175 2070.205 ;
        RECT 1915.510 2070.020 1923.175 2070.160 ;
        RECT 1915.510 2069.960 1915.830 2070.020 ;
        RECT 1922.885 2069.975 1923.175 2070.020 ;
        RECT 1410.890 2069.820 1411.210 2069.880 ;
        RECT 2014.870 2069.820 2015.190 2069.880 ;
        RECT 1410.890 2069.680 2015.190 2069.820 ;
        RECT 1410.890 2069.620 1411.210 2069.680 ;
        RECT 2014.870 2069.620 2015.190 2069.680 ;
        RECT 2238.890 2069.820 2239.210 2069.880 ;
        RECT 2346.990 2069.820 2347.310 2069.880 ;
        RECT 2238.890 2069.680 2347.310 2069.820 ;
        RECT 2238.890 2069.620 2239.210 2069.680 ;
        RECT 2346.990 2069.620 2347.310 2069.680 ;
        RECT 2480.390 2069.820 2480.710 2069.880 ;
        RECT 2525.470 2069.820 2525.790 2069.880 ;
        RECT 2480.390 2069.680 2525.790 2069.820 ;
        RECT 2480.390 2069.620 2480.710 2069.680 ;
        RECT 2525.470 2069.620 2525.790 2069.680 ;
        RECT 1408.145 2069.480 1408.435 2069.525 ;
        RECT 1411.350 2069.480 1411.670 2069.540 ;
        RECT 1408.145 2069.340 1411.670 2069.480 ;
        RECT 1408.145 2069.295 1408.435 2069.340 ;
        RECT 1411.350 2069.280 1411.670 2069.340 ;
        RECT 1417.330 2069.480 1417.650 2069.540 ;
        RECT 1980.370 2069.480 1980.690 2069.540 ;
        RECT 1417.330 2069.340 1980.690 2069.480 ;
        RECT 1417.330 2069.280 1417.650 2069.340 ;
        RECT 1980.370 2069.280 1980.690 2069.340 ;
        RECT 2045.690 2069.480 2046.010 2069.540 ;
        RECT 2380.570 2069.480 2380.890 2069.540 ;
        RECT 2045.690 2069.340 2380.890 2069.480 ;
        RECT 2045.690 2069.280 2046.010 2069.340 ;
        RECT 2380.570 2069.280 2380.890 2069.340 ;
        RECT 2445.890 2069.480 2446.210 2069.540 ;
        RECT 2512.590 2069.480 2512.910 2069.540 ;
        RECT 2445.890 2069.340 2512.910 2069.480 ;
        RECT 2445.890 2069.280 2446.210 2069.340 ;
        RECT 2512.590 2069.280 2512.910 2069.340 ;
        RECT 1408.590 2069.140 1408.910 2069.200 ;
        RECT 1922.425 2069.140 1922.715 2069.185 ;
        RECT 1408.590 2069.000 1922.715 2069.140 ;
        RECT 1408.590 2068.940 1408.910 2069.000 ;
        RECT 1922.425 2068.955 1922.715 2069.000 ;
        RECT 1922.885 2069.140 1923.175 2069.185 ;
        RECT 1932.545 2069.140 1932.835 2069.185 ;
        RECT 1922.885 2069.000 1932.835 2069.140 ;
        RECT 1922.885 2068.955 1923.175 2069.000 ;
        RECT 1932.545 2068.955 1932.835 2069.000 ;
        RECT 1935.750 2069.140 1936.070 2069.200 ;
        RECT 1959.670 2069.140 1959.990 2069.200 ;
        RECT 1935.750 2069.000 1959.990 2069.140 ;
        RECT 1935.750 2068.940 1936.070 2069.000 ;
        RECT 1959.670 2068.940 1959.990 2069.000 ;
        RECT 2059.490 2069.140 2059.810 2069.200 ;
        RECT 2387.470 2069.140 2387.790 2069.200 ;
        RECT 2059.490 2069.000 2387.790 2069.140 ;
        RECT 2059.490 2068.940 2059.810 2069.000 ;
        RECT 2387.470 2068.940 2387.790 2069.000 ;
        RECT 2418.290 2069.140 2418.610 2069.200 ;
        RECT 2497.870 2069.140 2498.190 2069.200 ;
        RECT 2418.290 2069.000 2498.190 2069.140 ;
        RECT 2418.290 2068.940 2418.610 2069.000 ;
        RECT 2497.870 2068.940 2498.190 2069.000 ;
        RECT 1409.510 2068.800 1409.830 2068.860 ;
        RECT 1946.330 2068.800 1946.650 2068.860 ;
        RECT 1409.510 2068.660 1946.650 2068.800 ;
        RECT 1409.510 2068.600 1409.830 2068.660 ;
        RECT 1946.330 2068.600 1946.650 2068.660 ;
        RECT 2031.890 2068.800 2032.210 2068.860 ;
        RECT 2359.870 2068.800 2360.190 2068.860 ;
        RECT 2031.890 2068.660 2360.190 2068.800 ;
        RECT 2031.890 2068.600 2032.210 2068.660 ;
        RECT 2359.870 2068.600 2360.190 2068.660 ;
        RECT 2459.690 2068.800 2460.010 2068.860 ;
        RECT 2518.570 2068.800 2518.890 2068.860 ;
        RECT 2459.690 2068.660 2518.890 2068.800 ;
        RECT 2459.690 2068.600 2460.010 2068.660 ;
        RECT 2518.570 2068.600 2518.890 2068.660 ;
        RECT 1409.970 2068.460 1410.290 2068.520 ;
        RECT 1945.870 2068.460 1946.190 2068.520 ;
        RECT 1409.970 2068.320 1946.190 2068.460 ;
        RECT 1409.970 2068.260 1410.290 2068.320 ;
        RECT 1945.870 2068.260 1946.190 2068.320 ;
        RECT 2080.190 2068.460 2080.510 2068.520 ;
        RECT 2394.370 2068.460 2394.690 2068.520 ;
        RECT 2080.190 2068.320 2394.690 2068.460 ;
        RECT 2080.190 2068.260 2080.510 2068.320 ;
        RECT 2394.370 2068.260 2394.690 2068.320 ;
        RECT 2411.390 2068.460 2411.710 2068.520 ;
        RECT 2491.430 2068.460 2491.750 2068.520 ;
        RECT 2411.390 2068.320 2491.750 2068.460 ;
        RECT 2411.390 2068.260 2411.710 2068.320 ;
        RECT 2491.430 2068.260 2491.750 2068.320 ;
        RECT 2494.190 2068.460 2494.510 2068.520 ;
        RECT 2532.370 2068.460 2532.690 2068.520 ;
        RECT 2494.190 2068.320 2532.690 2068.460 ;
        RECT 2494.190 2068.260 2494.510 2068.320 ;
        RECT 2532.370 2068.260 2532.690 2068.320 ;
        RECT 1409.050 2068.120 1409.370 2068.180 ;
        RECT 1906.785 2068.120 1907.075 2068.165 ;
        RECT 1932.070 2068.120 1932.390 2068.180 ;
        RECT 1409.050 2067.980 1907.075 2068.120 ;
        RECT 1409.050 2067.920 1409.370 2067.980 ;
        RECT 1906.785 2067.935 1907.075 2067.980 ;
        RECT 1907.320 2067.980 1932.390 2068.120 ;
        RECT 1410.430 2067.780 1410.750 2067.840 ;
        RECT 1907.320 2067.780 1907.460 2067.980 ;
        RECT 1932.070 2067.920 1932.390 2067.980 ;
        RECT 1932.545 2068.120 1932.835 2068.165 ;
        RECT 1939.905 2068.120 1940.195 2068.165 ;
        RECT 1932.545 2067.980 1940.195 2068.120 ;
        RECT 1932.545 2067.935 1932.835 2067.980 ;
        RECT 1939.905 2067.935 1940.195 2067.980 ;
        RECT 1942.650 2068.120 1942.970 2068.180 ;
        RECT 2021.770 2068.120 2022.090 2068.180 ;
        RECT 1942.650 2067.980 2022.090 2068.120 ;
        RECT 1942.650 2067.920 1942.970 2067.980 ;
        RECT 2021.770 2067.920 2022.090 2067.980 ;
        RECT 2121.590 2068.120 2121.910 2068.180 ;
        RECT 2402.190 2068.120 2402.510 2068.180 ;
        RECT 2121.590 2067.980 2402.510 2068.120 ;
        RECT 2121.590 2067.920 2121.910 2067.980 ;
        RECT 2402.190 2067.920 2402.510 2067.980 ;
        RECT 2404.490 2068.120 2404.810 2068.180 ;
        RECT 2484.070 2068.120 2484.390 2068.180 ;
        RECT 2404.490 2067.980 2484.390 2068.120 ;
        RECT 2404.490 2067.920 2404.810 2067.980 ;
        RECT 2484.070 2067.920 2484.390 2067.980 ;
        RECT 1410.430 2067.640 1907.460 2067.780 ;
        RECT 1907.690 2067.780 1908.010 2067.840 ;
        RECT 1973.470 2067.780 1973.790 2067.840 ;
        RECT 1907.690 2067.640 1973.790 2067.780 ;
        RECT 1410.430 2067.580 1410.750 2067.640 ;
        RECT 1907.690 2067.580 1908.010 2067.640 ;
        RECT 1973.470 2067.580 1973.790 2067.640 ;
        RECT 2156.090 2067.780 2156.410 2067.840 ;
        RECT 2428.870 2067.780 2429.190 2067.840 ;
        RECT 2156.090 2067.640 2429.190 2067.780 ;
        RECT 2156.090 2067.580 2156.410 2067.640 ;
        RECT 2428.870 2067.580 2429.190 2067.640 ;
        RECT 1413.650 2067.440 1413.970 2067.500 ;
        RECT 1879.645 2067.440 1879.935 2067.485 ;
        RECT 1413.650 2067.300 1879.935 2067.440 ;
        RECT 1413.650 2067.240 1413.970 2067.300 ;
        RECT 1879.645 2067.255 1879.935 2067.300 ;
        RECT 1880.090 2067.440 1880.410 2067.500 ;
        RECT 1911.370 2067.440 1911.690 2067.500 ;
        RECT 1880.090 2067.300 1911.690 2067.440 ;
        RECT 1880.090 2067.240 1880.410 2067.300 ;
        RECT 1911.370 2067.240 1911.690 2067.300 ;
        RECT 1915.970 2067.440 1916.290 2067.500 ;
        RECT 2007.970 2067.440 2008.290 2067.500 ;
        RECT 1915.970 2067.300 2008.290 2067.440 ;
        RECT 1915.970 2067.240 1916.290 2067.300 ;
        RECT 2007.970 2067.240 2008.290 2067.300 ;
        RECT 2142.290 2067.440 2142.610 2067.500 ;
        RECT 2415.070 2067.440 2415.390 2067.500 ;
        RECT 2142.290 2067.300 2415.390 2067.440 ;
        RECT 2142.290 2067.240 2142.610 2067.300 ;
        RECT 2415.070 2067.240 2415.390 2067.300 ;
        RECT 2466.590 2067.440 2466.910 2067.500 ;
        RECT 2519.950 2067.440 2520.270 2067.500 ;
        RECT 2466.590 2067.300 2520.270 2067.440 ;
        RECT 2466.590 2067.240 2466.910 2067.300 ;
        RECT 2519.950 2067.240 2520.270 2067.300 ;
        RECT 1413.190 2067.100 1413.510 2067.160 ;
        RECT 1892.985 2067.100 1893.275 2067.145 ;
        RECT 1413.190 2066.960 1893.275 2067.100 ;
        RECT 1413.190 2066.900 1413.510 2066.960 ;
        RECT 1892.985 2066.915 1893.275 2066.960 ;
        RECT 1894.365 2067.100 1894.655 2067.145 ;
        RECT 1921.965 2067.100 1922.255 2067.145 ;
        RECT 1894.365 2066.960 1922.255 2067.100 ;
        RECT 1894.365 2066.915 1894.655 2066.960 ;
        RECT 1921.965 2066.915 1922.255 2066.960 ;
        RECT 1922.885 2067.100 1923.175 2067.145 ;
        RECT 1987.270 2067.100 1987.590 2067.160 ;
        RECT 1922.885 2066.960 1987.590 2067.100 ;
        RECT 1922.885 2066.915 1923.175 2066.960 ;
        RECT 1987.270 2066.900 1987.590 2066.960 ;
        RECT 2135.390 2067.100 2135.710 2067.160 ;
        RECT 2408.170 2067.100 2408.490 2067.160 ;
        RECT 2135.390 2066.960 2408.490 2067.100 ;
        RECT 2135.390 2066.900 2135.710 2066.960 ;
        RECT 2408.170 2066.900 2408.490 2066.960 ;
        RECT 2425.190 2067.100 2425.510 2067.160 ;
        RECT 2505.230 2067.100 2505.550 2067.160 ;
        RECT 2425.190 2066.960 2505.550 2067.100 ;
        RECT 2425.190 2066.900 2425.510 2066.960 ;
        RECT 2505.230 2066.900 2505.550 2066.960 ;
        RECT 1411.810 2066.760 1412.130 2066.820 ;
        RECT 1910.910 2066.760 1911.230 2066.820 ;
        RECT 1411.810 2066.620 1911.230 2066.760 ;
        RECT 1411.810 2066.560 1412.130 2066.620 ;
        RECT 1910.910 2066.560 1911.230 2066.620 ;
        RECT 1921.505 2066.760 1921.795 2066.805 ;
        RECT 1987.730 2066.760 1988.050 2066.820 ;
        RECT 1921.505 2066.620 1988.050 2066.760 ;
        RECT 1921.505 2066.575 1921.795 2066.620 ;
        RECT 1987.730 2066.560 1988.050 2066.620 ;
        RECT 2149.190 2066.760 2149.510 2066.820 ;
        RECT 2421.970 2066.760 2422.290 2066.820 ;
        RECT 2149.190 2066.620 2422.290 2066.760 ;
        RECT 2149.190 2066.560 2149.510 2066.620 ;
        RECT 2421.970 2066.560 2422.290 2066.620 ;
        RECT 1412.270 2066.420 1412.590 2066.480 ;
        RECT 1911.830 2066.420 1912.150 2066.480 ;
        RECT 1412.270 2066.280 1912.150 2066.420 ;
        RECT 1412.270 2066.220 1412.590 2066.280 ;
        RECT 1911.830 2066.220 1912.150 2066.280 ;
        RECT 1915.050 2066.420 1915.370 2066.480 ;
        RECT 1994.170 2066.420 1994.490 2066.480 ;
        RECT 1915.050 2066.280 1994.490 2066.420 ;
        RECT 1915.050 2066.220 1915.370 2066.280 ;
        RECT 1994.170 2066.220 1994.490 2066.280 ;
        RECT 2176.790 2066.420 2177.110 2066.480 ;
        RECT 2442.670 2066.420 2442.990 2066.480 ;
        RECT 2176.790 2066.280 2442.990 2066.420 ;
        RECT 2176.790 2066.220 2177.110 2066.280 ;
        RECT 2442.670 2066.220 2442.990 2066.280 ;
        RECT 1412.730 2066.080 1413.050 2066.140 ;
        RECT 1887.005 2066.080 1887.295 2066.125 ;
        RECT 1412.730 2065.940 1887.295 2066.080 ;
        RECT 1412.730 2065.880 1413.050 2065.940 ;
        RECT 1887.005 2065.895 1887.295 2065.940 ;
        RECT 1887.465 2066.080 1887.755 2066.125 ;
        RECT 1893.445 2066.080 1893.735 2066.125 ;
        RECT 1887.465 2065.940 1893.735 2066.080 ;
        RECT 1887.465 2065.895 1887.755 2065.940 ;
        RECT 1893.445 2065.895 1893.735 2065.940 ;
        RECT 1893.890 2066.080 1894.210 2066.140 ;
        RECT 1921.490 2066.080 1921.810 2066.140 ;
        RECT 1893.890 2065.940 1921.810 2066.080 ;
        RECT 1893.890 2065.880 1894.210 2065.940 ;
        RECT 1921.490 2065.880 1921.810 2065.940 ;
        RECT 1921.950 2066.080 1922.270 2066.140 ;
        RECT 1966.570 2066.080 1966.890 2066.140 ;
        RECT 1921.950 2065.940 1966.890 2066.080 ;
        RECT 1921.950 2065.880 1922.270 2065.940 ;
        RECT 1966.570 2065.880 1966.890 2065.940 ;
        RECT 2169.890 2066.080 2170.210 2066.140 ;
        RECT 2435.770 2066.080 2436.090 2066.140 ;
        RECT 2169.890 2065.940 2436.090 2066.080 ;
        RECT 2169.890 2065.880 2170.210 2065.940 ;
        RECT 2435.770 2065.880 2436.090 2065.940 ;
        RECT 1413.650 2065.740 1413.970 2065.800 ;
        RECT 1892.985 2065.740 1893.275 2065.785 ;
        RECT 1918.270 2065.740 1918.590 2065.800 ;
        RECT 1413.650 2065.600 1891.360 2065.740 ;
        RECT 1413.650 2065.540 1413.970 2065.600 ;
        RECT 1408.130 2065.400 1408.450 2065.460 ;
        RECT 1890.670 2065.400 1890.990 2065.460 ;
        RECT 1408.130 2065.260 1890.990 2065.400 ;
        RECT 1891.220 2065.400 1891.360 2065.600 ;
        RECT 1892.985 2065.600 1918.590 2065.740 ;
        RECT 1892.985 2065.555 1893.275 2065.600 ;
        RECT 1918.270 2065.540 1918.590 2065.600 ;
        RECT 1922.425 2065.740 1922.715 2065.785 ;
        RECT 1952.770 2065.740 1953.090 2065.800 ;
        RECT 1922.425 2065.600 1953.090 2065.740 ;
        RECT 1922.425 2065.555 1922.715 2065.600 ;
        RECT 1952.770 2065.540 1953.090 2065.600 ;
        RECT 2087.090 2065.740 2087.410 2065.800 ;
        RECT 2340.550 2065.740 2340.870 2065.800 ;
        RECT 2087.090 2065.600 2340.870 2065.740 ;
        RECT 2087.090 2065.540 2087.410 2065.600 ;
        RECT 2340.550 2065.540 2340.870 2065.600 ;
        RECT 1898.030 2065.400 1898.350 2065.460 ;
        RECT 1891.220 2065.260 1898.350 2065.400 ;
        RECT 1408.130 2065.200 1408.450 2065.260 ;
        RECT 1890.670 2065.200 1890.990 2065.260 ;
        RECT 1898.030 2065.200 1898.350 2065.260 ;
        RECT 1900.790 2065.400 1901.110 2065.460 ;
        RECT 1922.885 2065.400 1923.175 2065.445 ;
        RECT 1900.790 2065.260 1923.175 2065.400 ;
        RECT 1900.790 2065.200 1901.110 2065.260 ;
        RECT 1922.885 2065.215 1923.175 2065.260 ;
        RECT 1928.850 2065.400 1929.170 2065.460 ;
        RECT 1980.370 2065.400 1980.690 2065.460 ;
        RECT 1928.850 2065.260 1980.690 2065.400 ;
        RECT 1928.850 2065.200 1929.170 2065.260 ;
        RECT 1980.370 2065.200 1980.690 2065.260 ;
        RECT 2211.290 2065.400 2211.610 2065.460 ;
        RECT 2449.570 2065.400 2449.890 2065.460 ;
        RECT 2211.290 2065.260 2449.890 2065.400 ;
        RECT 2211.290 2065.200 2211.610 2065.260 ;
        RECT 2449.570 2065.200 2449.890 2065.260 ;
        RECT 1411.350 2065.060 1411.670 2065.120 ;
        RECT 1435.270 2065.060 1435.590 2065.120 ;
        RECT 1411.350 2064.920 1435.590 2065.060 ;
        RECT 1411.350 2064.860 1411.670 2064.920 ;
        RECT 1435.270 2064.860 1435.590 2064.920 ;
        RECT 1483.110 2065.060 1483.430 2065.120 ;
        RECT 1531.870 2065.060 1532.190 2065.120 ;
        RECT 1483.110 2064.920 1532.190 2065.060 ;
        RECT 1483.110 2064.860 1483.430 2064.920 ;
        RECT 1531.870 2064.860 1532.190 2064.920 ;
        RECT 1579.710 2065.060 1580.030 2065.120 ;
        RECT 1655.610 2065.060 1655.930 2065.120 ;
        RECT 1579.710 2064.920 1655.930 2065.060 ;
        RECT 1579.710 2064.860 1580.030 2064.920 ;
        RECT 1655.610 2064.860 1655.930 2064.920 ;
        RECT 1676.310 2065.060 1676.630 2065.120 ;
        RECT 1752.210 2065.060 1752.530 2065.120 ;
        RECT 1676.310 2064.920 1752.530 2065.060 ;
        RECT 1676.310 2064.860 1676.630 2064.920 ;
        RECT 1752.210 2064.860 1752.530 2064.920 ;
        RECT 1772.910 2065.060 1773.230 2065.120 ;
        RECT 1821.670 2065.060 1821.990 2065.120 ;
        RECT 1772.910 2064.920 1821.990 2065.060 ;
        RECT 1772.910 2064.860 1773.230 2064.920 ;
        RECT 1821.670 2064.860 1821.990 2064.920 ;
        RECT 1869.525 2065.060 1869.815 2065.105 ;
        RECT 1883.770 2065.060 1884.090 2065.120 ;
        RECT 1869.525 2064.920 1884.090 2065.060 ;
        RECT 1869.525 2064.875 1869.815 2064.920 ;
        RECT 1883.770 2064.860 1884.090 2064.920 ;
        RECT 1887.005 2065.060 1887.295 2065.105 ;
        RECT 1904.470 2065.060 1904.790 2065.120 ;
        RECT 1887.005 2064.920 1904.790 2065.060 ;
        RECT 1887.005 2064.875 1887.295 2064.920 ;
        RECT 1904.470 2064.860 1904.790 2064.920 ;
        RECT 1906.785 2065.060 1907.075 2065.105 ;
        RECT 1938.970 2065.060 1939.290 2065.120 ;
        RECT 1906.785 2064.920 1939.290 2065.060 ;
        RECT 1906.785 2064.875 1907.075 2064.920 ;
        RECT 1938.970 2064.860 1939.290 2064.920 ;
        RECT 1939.445 2065.060 1939.735 2065.105 ;
        RECT 1987.270 2065.060 1987.590 2065.120 ;
        RECT 1939.445 2064.920 1987.590 2065.060 ;
        RECT 1939.445 2064.875 1939.735 2064.920 ;
        RECT 1987.270 2064.860 1987.590 2064.920 ;
        RECT 2225.090 2065.060 2225.410 2065.120 ;
        RECT 2456.470 2065.060 2456.790 2065.120 ;
        RECT 2225.090 2064.920 2456.790 2065.060 ;
        RECT 2225.090 2064.860 2225.410 2064.920 ;
        RECT 2456.470 2064.860 2456.790 2064.920 ;
        RECT 1420.550 2064.720 1420.870 2064.780 ;
        RECT 1869.970 2064.720 1870.290 2064.780 ;
        RECT 1420.550 2064.580 1870.290 2064.720 ;
        RECT 1420.550 2064.520 1420.870 2064.580 ;
        RECT 1869.970 2064.520 1870.290 2064.580 ;
        RECT 1879.645 2064.720 1879.935 2064.765 ;
        RECT 1914.590 2064.720 1914.910 2064.780 ;
        RECT 1921.045 2064.720 1921.335 2064.765 ;
        RECT 1879.645 2064.580 1913.440 2064.720 ;
        RECT 1879.645 2064.535 1879.935 2064.580 ;
        RECT 1421.010 2064.380 1421.330 2064.440 ;
        RECT 1870.890 2064.380 1871.210 2064.440 ;
        RECT 1421.010 2064.240 1871.210 2064.380 ;
        RECT 1421.010 2064.180 1421.330 2064.240 ;
        RECT 1870.890 2064.180 1871.210 2064.240 ;
        RECT 1873.190 2064.380 1873.510 2064.440 ;
        RECT 1911.370 2064.380 1911.690 2064.440 ;
        RECT 1873.190 2064.240 1911.690 2064.380 ;
        RECT 1913.300 2064.380 1913.440 2064.580 ;
        RECT 1914.590 2064.580 1921.335 2064.720 ;
        RECT 1914.590 2064.520 1914.910 2064.580 ;
        RECT 1921.045 2064.535 1921.335 2064.580 ;
        RECT 1921.490 2064.720 1921.810 2064.780 ;
        RECT 2015.790 2064.720 2016.110 2064.780 ;
        RECT 1921.490 2064.580 2016.110 2064.720 ;
        RECT 1921.490 2064.520 1921.810 2064.580 ;
        RECT 2015.790 2064.520 2016.110 2064.580 ;
        RECT 2231.990 2064.720 2232.310 2064.780 ;
        RECT 2456.930 2064.720 2457.250 2064.780 ;
        RECT 2231.990 2064.580 2457.250 2064.720 ;
        RECT 2231.990 2064.520 2232.310 2064.580 ;
        RECT 2456.930 2064.520 2457.250 2064.580 ;
        RECT 1925.170 2064.380 1925.490 2064.440 ;
        RECT 1913.300 2064.240 1925.490 2064.380 ;
        RECT 1873.190 2064.180 1873.510 2064.240 ;
        RECT 1911.370 2064.180 1911.690 2064.240 ;
        RECT 1925.170 2064.180 1925.490 2064.240 ;
        RECT 1928.390 2064.380 1928.710 2064.440 ;
        RECT 1973.470 2064.380 1973.790 2064.440 ;
        RECT 1928.390 2064.240 1973.790 2064.380 ;
        RECT 1928.390 2064.180 1928.710 2064.240 ;
        RECT 1973.470 2064.180 1973.790 2064.240 ;
        RECT 2245.790 2064.380 2246.110 2064.440 ;
        RECT 2463.370 2064.380 2463.690 2064.440 ;
        RECT 2245.790 2064.240 2463.690 2064.380 ;
        RECT 2245.790 2064.180 2246.110 2064.240 ;
        RECT 2463.370 2064.180 2463.690 2064.240 ;
        RECT 1420.090 2064.040 1420.410 2064.100 ;
        RECT 1863.070 2064.040 1863.390 2064.100 ;
        RECT 1420.090 2063.900 1863.390 2064.040 ;
        RECT 1420.090 2063.840 1420.410 2063.900 ;
        RECT 1863.070 2063.840 1863.390 2063.900 ;
        RECT 1866.290 2064.040 1866.610 2064.100 ;
        RECT 2001.070 2064.040 2001.390 2064.100 ;
        RECT 1866.290 2063.900 2001.390 2064.040 ;
        RECT 1866.290 2063.840 1866.610 2063.900 ;
        RECT 2001.070 2063.840 2001.390 2063.900 ;
        RECT 2052.590 2064.040 2052.910 2064.100 ;
        RECT 2587.570 2064.040 2587.890 2064.100 ;
        RECT 2052.590 2063.900 2587.890 2064.040 ;
        RECT 2052.590 2063.840 2052.910 2063.900 ;
        RECT 2587.570 2063.840 2587.890 2063.900 ;
        RECT 1419.170 2063.700 1419.490 2063.760 ;
        RECT 1856.170 2063.700 1856.490 2063.760 ;
        RECT 1419.170 2063.560 1856.490 2063.700 ;
        RECT 1419.170 2063.500 1419.490 2063.560 ;
        RECT 1856.170 2063.500 1856.490 2063.560 ;
        RECT 1856.630 2063.700 1856.950 2063.760 ;
        RECT 1869.525 2063.700 1869.815 2063.745 ;
        RECT 1856.630 2063.560 1869.815 2063.700 ;
        RECT 1856.630 2063.500 1856.950 2063.560 ;
        RECT 1869.525 2063.515 1869.815 2063.560 ;
        RECT 1873.650 2063.700 1873.970 2063.760 ;
        RECT 1886.545 2063.700 1886.835 2063.745 ;
        RECT 1873.650 2063.560 1886.835 2063.700 ;
        RECT 1873.650 2063.500 1873.970 2063.560 ;
        RECT 1886.545 2063.515 1886.835 2063.560 ;
        RECT 1886.990 2063.700 1887.310 2063.760 ;
        RECT 1921.505 2063.700 1921.795 2063.745 ;
        RECT 1886.990 2063.560 1921.795 2063.700 ;
        RECT 1886.990 2063.500 1887.310 2063.560 ;
        RECT 1921.505 2063.515 1921.795 2063.560 ;
        RECT 1921.965 2063.700 1922.255 2063.745 ;
        RECT 1994.170 2063.700 1994.490 2063.760 ;
        RECT 1921.965 2063.560 1994.490 2063.700 ;
        RECT 1921.965 2063.515 1922.255 2063.560 ;
        RECT 1994.170 2063.500 1994.490 2063.560 ;
        RECT 2335.490 2063.700 2335.810 2063.760 ;
        RECT 2478.550 2063.700 2478.870 2063.760 ;
        RECT 2335.490 2063.560 2478.870 2063.700 ;
        RECT 2335.490 2063.500 2335.810 2063.560 ;
        RECT 2478.550 2063.500 2478.870 2063.560 ;
        RECT 1418.250 2063.360 1418.570 2063.420 ;
        RECT 1835.470 2063.360 1835.790 2063.420 ;
        RECT 1418.250 2063.220 1835.790 2063.360 ;
        RECT 1418.250 2063.160 1418.570 2063.220 ;
        RECT 1835.470 2063.160 1835.790 2063.220 ;
        RECT 1838.690 2063.360 1839.010 2063.420 ;
        RECT 1925.170 2063.360 1925.490 2063.420 ;
        RECT 1939.445 2063.360 1939.735 2063.405 ;
        RECT 1838.690 2063.220 1925.490 2063.360 ;
        RECT 1838.690 2063.160 1839.010 2063.220 ;
        RECT 1925.170 2063.160 1925.490 2063.220 ;
        RECT 1925.720 2063.220 1939.735 2063.360 ;
        RECT 1419.630 2063.020 1419.950 2063.080 ;
        RECT 1760.490 2063.020 1760.810 2063.080 ;
        RECT 1419.630 2062.880 1760.810 2063.020 ;
        RECT 1419.630 2062.820 1419.950 2062.880 ;
        RECT 1760.490 2062.820 1760.810 2062.880 ;
        RECT 1921.045 2063.020 1921.335 2063.065 ;
        RECT 1925.720 2063.020 1925.860 2063.220 ;
        RECT 1939.445 2063.175 1939.735 2063.220 ;
        RECT 1939.905 2063.360 1940.195 2063.405 ;
        RECT 2001.070 2063.360 2001.390 2063.420 ;
        RECT 1939.905 2063.220 2001.390 2063.360 ;
        RECT 1939.905 2063.175 1940.195 2063.220 ;
        RECT 2001.070 2063.160 2001.390 2063.220 ;
        RECT 2328.590 2063.360 2328.910 2063.420 ;
        RECT 2470.270 2063.360 2470.590 2063.420 ;
        RECT 2328.590 2063.220 2470.590 2063.360 ;
        RECT 2328.590 2063.160 2328.910 2063.220 ;
        RECT 2470.270 2063.160 2470.590 2063.220 ;
        RECT 1921.045 2062.880 1925.860 2063.020 ;
        RECT 1921.045 2062.835 1921.335 2062.880 ;
        RECT 1418.710 2062.680 1419.030 2062.740 ;
        RECT 1760.030 2062.680 1760.350 2062.740 ;
        RECT 1418.710 2062.540 1760.350 2062.680 ;
        RECT 1418.710 2062.480 1419.030 2062.540 ;
        RECT 1760.030 2062.480 1760.350 2062.540 ;
        RECT 1419.170 2062.340 1419.490 2062.400 ;
        RECT 1766.470 2062.340 1766.790 2062.400 ;
        RECT 1419.170 2062.200 1766.790 2062.340 ;
        RECT 1419.170 2062.140 1419.490 2062.200 ;
        RECT 1766.470 2062.140 1766.790 2062.200 ;
        RECT 1420.090 2062.000 1420.410 2062.060 ;
        RECT 1773.370 2062.000 1773.690 2062.060 ;
        RECT 1420.090 2061.860 1773.690 2062.000 ;
        RECT 1420.090 2061.800 1420.410 2061.860 ;
        RECT 1773.370 2061.800 1773.690 2061.860 ;
        RECT 1420.550 2061.660 1420.870 2061.720 ;
        RECT 1780.730 2061.660 1781.050 2061.720 ;
        RECT 1420.550 2061.520 1781.050 2061.660 ;
        RECT 1420.550 2061.460 1420.870 2061.520 ;
        RECT 1780.730 2061.460 1781.050 2061.520 ;
        RECT 1417.330 2061.320 1417.650 2061.380 ;
        RECT 1787.630 2061.320 1787.950 2061.380 ;
        RECT 1417.330 2061.180 1787.950 2061.320 ;
        RECT 1417.330 2061.120 1417.650 2061.180 ;
        RECT 1787.630 2061.120 1787.950 2061.180 ;
        RECT 1421.010 2060.980 1421.330 2061.040 ;
        RECT 1794.530 2060.980 1794.850 2061.040 ;
        RECT 1421.010 2060.840 1794.850 2060.980 ;
        RECT 1421.010 2060.780 1421.330 2060.840 ;
        RECT 1794.530 2060.780 1794.850 2060.840 ;
        RECT 1715.410 2060.640 1715.730 2060.700 ;
        RECT 2339.170 2060.640 2339.490 2060.700 ;
        RECT 1715.410 2060.500 2339.490 2060.640 ;
        RECT 1715.410 2060.440 1715.730 2060.500 ;
        RECT 2339.170 2060.440 2339.490 2060.500 ;
        RECT 1690.110 2060.300 1690.430 2060.360 ;
        RECT 2318.470 2060.300 2318.790 2060.360 ;
        RECT 1690.110 2060.160 2318.790 2060.300 ;
        RECT 1690.110 2060.100 1690.430 2060.160 ;
        RECT 2318.470 2060.100 2318.790 2060.160 ;
        RECT 1416.870 2059.960 1417.190 2060.020 ;
        RECT 2263.270 2059.960 2263.590 2060.020 ;
        RECT 1416.870 2059.820 2263.590 2059.960 ;
        RECT 1416.870 2059.760 1417.190 2059.820 ;
        RECT 2263.270 2059.760 2263.590 2059.820 ;
        RECT 1462.870 2059.620 1463.190 2059.680 ;
        RECT 2325.370 2059.620 2325.690 2059.680 ;
        RECT 1462.870 2059.480 2325.690 2059.620 ;
        RECT 1462.870 2059.420 1463.190 2059.480 ;
        RECT 2325.370 2059.420 2325.690 2059.480 ;
        RECT 1418.250 2059.280 1418.570 2059.340 ;
        RECT 1753.130 2059.280 1753.450 2059.340 ;
        RECT 1418.250 2059.140 1753.450 2059.280 ;
        RECT 1418.250 2059.080 1418.570 2059.140 ;
        RECT 1753.130 2059.080 1753.450 2059.140 ;
        RECT 1417.790 2058.940 1418.110 2059.000 ;
        RECT 1745.770 2058.940 1746.090 2059.000 ;
        RECT 1417.790 2058.800 1746.090 2058.940 ;
        RECT 1417.790 2058.740 1418.110 2058.800 ;
        RECT 1745.770 2058.740 1746.090 2058.800 ;
        RECT 1434.810 2058.600 1435.130 2058.660 ;
        RECT 1738.870 2058.600 1739.190 2058.660 ;
        RECT 1434.810 2058.460 1739.190 2058.600 ;
        RECT 1434.810 2058.400 1435.130 2058.460 ;
        RECT 1738.870 2058.400 1739.190 2058.460 ;
        RECT 1434.350 2058.260 1434.670 2058.320 ;
        RECT 1731.970 2058.260 1732.290 2058.320 ;
        RECT 1434.350 2058.120 1732.290 2058.260 ;
        RECT 1434.350 2058.060 1434.670 2058.120 ;
        RECT 1731.970 2058.060 1732.290 2058.120 ;
        RECT 1433.430 2057.920 1433.750 2057.980 ;
        RECT 1725.070 2057.920 1725.390 2057.980 ;
        RECT 1433.430 2057.780 1725.390 2057.920 ;
        RECT 1433.430 2057.720 1433.750 2057.780 ;
        RECT 1725.070 2057.720 1725.390 2057.780 ;
        RECT 1433.890 2057.580 1434.210 2057.640 ;
        RECT 1718.170 2057.580 1718.490 2057.640 ;
        RECT 1433.890 2057.440 1718.490 2057.580 ;
        RECT 1433.890 2057.380 1434.210 2057.440 ;
        RECT 1718.170 2057.380 1718.490 2057.440 ;
        RECT 1693.790 2056.560 1694.110 2056.620 ;
        RECT 2028.670 2056.560 2028.990 2056.620 ;
        RECT 1693.790 2056.420 2028.990 2056.560 ;
        RECT 1693.790 2056.360 1694.110 2056.420 ;
        RECT 2028.670 2056.360 2028.990 2056.420 ;
        RECT 1413.650 2056.220 1413.970 2056.280 ;
        RECT 2332.270 2056.220 2332.590 2056.280 ;
        RECT 1413.650 2056.080 2332.590 2056.220 ;
        RECT 1413.650 2056.020 1413.970 2056.080 ;
        RECT 2332.270 2056.020 2332.590 2056.080 ;
        RECT 1414.110 2055.880 1414.430 2055.940 ;
        RECT 1715.410 2055.880 1715.730 2055.940 ;
        RECT 1414.110 2055.740 1715.730 2055.880 ;
        RECT 1414.110 2055.680 1414.430 2055.740 ;
        RECT 1715.410 2055.680 1715.730 2055.740 ;
        RECT 1408.130 2055.540 1408.450 2055.600 ;
        RECT 2193.810 2055.540 2194.130 2055.600 ;
        RECT 1408.130 2055.400 2194.130 2055.540 ;
        RECT 1408.130 2055.340 1408.450 2055.400 ;
        RECT 2193.810 2055.340 2194.130 2055.400 ;
        RECT 1409.970 2055.200 1410.290 2055.260 ;
        RECT 2256.370 2055.200 2256.690 2055.260 ;
        RECT 1409.970 2055.060 2256.690 2055.200 ;
        RECT 1409.970 2055.000 1410.290 2055.060 ;
        RECT 2256.370 2055.000 2256.690 2055.060 ;
        RECT 1410.890 2054.860 1411.210 2054.920 ;
        RECT 2280.290 2054.860 2280.610 2054.920 ;
        RECT 1410.890 2054.720 2280.610 2054.860 ;
        RECT 1410.890 2054.660 1411.210 2054.720 ;
        RECT 2280.290 2054.660 2280.610 2054.720 ;
        RECT 1411.350 2054.520 1411.670 2054.580 ;
        RECT 2287.190 2054.520 2287.510 2054.580 ;
        RECT 1411.350 2054.380 2287.510 2054.520 ;
        RECT 1411.350 2054.320 1411.670 2054.380 ;
        RECT 2287.190 2054.320 2287.510 2054.380 ;
        RECT 1413.190 2054.180 1413.510 2054.240 ;
        RECT 2294.090 2054.180 2294.410 2054.240 ;
        RECT 1413.190 2054.040 2294.410 2054.180 ;
        RECT 1413.190 2053.980 1413.510 2054.040 ;
        RECT 2294.090 2053.980 2294.410 2054.040 ;
        RECT 1412.730 2053.840 1413.050 2053.900 ;
        RECT 2300.990 2053.840 2301.310 2053.900 ;
        RECT 1412.730 2053.700 2301.310 2053.840 ;
        RECT 1412.730 2053.640 1413.050 2053.700 ;
        RECT 2300.990 2053.640 2301.310 2053.700 ;
        RECT 1412.270 2053.500 1412.590 2053.560 ;
        RECT 2301.910 2053.500 2302.230 2053.560 ;
        RECT 1412.270 2053.360 2302.230 2053.500 ;
        RECT 1412.270 2053.300 1412.590 2053.360 ;
        RECT 2301.910 2053.300 2302.230 2053.360 ;
        RECT 1411.810 2053.160 1412.130 2053.220 ;
        RECT 2304.670 2053.160 2304.990 2053.220 ;
        RECT 1411.810 2053.020 2304.990 2053.160 ;
        RECT 1411.810 2052.960 1412.130 2053.020 ;
        RECT 2304.670 2052.960 2304.990 2053.020 ;
        RECT 1414.110 2052.820 1414.430 2052.880 ;
        RECT 2311.570 2052.820 2311.890 2052.880 ;
        RECT 1414.110 2052.680 2311.890 2052.820 ;
        RECT 1414.110 2052.620 1414.430 2052.680 ;
        RECT 2311.570 2052.620 2311.890 2052.680 ;
        RECT 1421.470 2052.480 1421.790 2052.540 ;
        RECT 1704.370 2052.480 1704.690 2052.540 ;
        RECT 1421.470 2052.340 1704.690 2052.480 ;
        RECT 1421.470 2052.280 1421.790 2052.340 ;
        RECT 1704.370 2052.280 1704.690 2052.340 ;
        RECT 1408.590 2049.080 1408.910 2049.140 ;
        RECT 1462.870 2049.080 1463.190 2049.140 ;
        RECT 1408.590 2048.940 1463.190 2049.080 ;
        RECT 1408.590 2048.880 1408.910 2048.940 ;
        RECT 1462.870 2048.880 1463.190 2048.940 ;
        RECT 1408.590 2042.280 1408.910 2042.340 ;
        RECT 1690.110 2042.280 1690.430 2042.340 ;
        RECT 1408.590 2042.140 1690.430 2042.280 ;
        RECT 1408.590 2042.080 1408.910 2042.140 ;
        RECT 1690.110 2042.080 1690.430 2042.140 ;
        RECT 1408.130 2020.180 1408.450 2020.240 ;
        RECT 1416.410 2020.180 1416.730 2020.240 ;
        RECT 1408.130 2020.040 1416.730 2020.180 ;
        RECT 1408.130 2019.980 1408.450 2020.040 ;
        RECT 1416.410 2019.980 1416.730 2020.040 ;
        RECT 1414.110 2011.340 1414.430 2011.400 ;
        RECT 1430.670 2011.340 1430.990 2011.400 ;
        RECT 1414.110 2011.200 1430.990 2011.340 ;
        RECT 1414.110 2011.140 1414.430 2011.200 ;
        RECT 1430.670 2011.140 1430.990 2011.200 ;
        RECT 1414.110 2005.900 1414.430 2005.960 ;
        RECT 1431.130 2005.900 1431.450 2005.960 ;
        RECT 1414.110 2005.760 1431.450 2005.900 ;
        RECT 1414.110 2005.700 1414.430 2005.760 ;
        RECT 1431.130 2005.700 1431.450 2005.760 ;
        RECT 1414.110 2000.800 1414.430 2000.860 ;
        RECT 1686.890 2000.800 1687.210 2000.860 ;
        RECT 1414.110 2000.660 1687.210 2000.800 ;
        RECT 1414.110 2000.600 1414.430 2000.660 ;
        RECT 1686.890 2000.600 1687.210 2000.660 ;
        RECT 1411.350 2000.460 1411.670 2000.520 ;
        RECT 1460.110 2000.460 1460.430 2000.520 ;
        RECT 1411.350 2000.320 1460.430 2000.460 ;
        RECT 1411.350 2000.260 1411.670 2000.320 ;
        RECT 1460.110 2000.260 1460.430 2000.320 ;
        RECT 1408.130 1990.940 1408.450 1991.000 ;
        RECT 1416.870 1990.940 1417.190 1991.000 ;
        RECT 1408.130 1990.800 1417.190 1990.940 ;
        RECT 1408.130 1990.740 1408.450 1990.800 ;
        RECT 1416.870 1990.740 1417.190 1990.800 ;
        RECT 1408.130 1986.180 1408.450 1986.240 ;
        RECT 1421.010 1986.180 1421.330 1986.240 ;
        RECT 1408.130 1986.040 1421.330 1986.180 ;
        RECT 1408.130 1985.980 1408.450 1986.040 ;
        RECT 1421.010 1985.980 1421.330 1986.040 ;
        RECT 1408.130 1982.440 1408.450 1982.500 ;
        RECT 1417.330 1982.440 1417.650 1982.500 ;
        RECT 1408.130 1982.300 1417.650 1982.440 ;
        RECT 1408.130 1982.240 1408.450 1982.300 ;
        RECT 1417.330 1982.240 1417.650 1982.300 ;
        RECT 1410.890 1980.060 1411.210 1980.120 ;
        RECT 1410.695 1979.920 1411.210 1980.060 ;
        RECT 1410.890 1979.860 1411.210 1979.920 ;
        RECT 1408.130 1979.040 1408.450 1979.100 ;
        RECT 1420.550 1979.040 1420.870 1979.100 ;
        RECT 1408.130 1978.900 1420.870 1979.040 ;
        RECT 1408.130 1978.840 1408.450 1978.900 ;
        RECT 1420.550 1978.840 1420.870 1978.900 ;
        RECT 1408.130 1971.900 1408.450 1971.960 ;
        RECT 1420.090 1971.900 1420.410 1971.960 ;
        RECT 1408.130 1971.760 1420.410 1971.900 ;
        RECT 1408.130 1971.700 1408.450 1971.760 ;
        RECT 1420.090 1971.700 1420.410 1971.760 ;
        RECT 1408.130 1966.120 1408.450 1966.180 ;
        RECT 1419.170 1966.120 1419.490 1966.180 ;
        RECT 1408.130 1965.980 1419.490 1966.120 ;
        RECT 1408.130 1965.920 1408.450 1965.980 ;
        RECT 1419.170 1965.920 1419.490 1965.980 ;
        RECT 1408.130 1960.340 1408.450 1960.400 ;
        RECT 1419.630 1960.340 1419.950 1960.400 ;
        RECT 1408.130 1960.200 1419.950 1960.340 ;
        RECT 1408.130 1960.140 1408.450 1960.200 ;
        RECT 1419.630 1960.140 1419.950 1960.200 ;
        RECT 1408.130 1958.300 1408.450 1958.360 ;
        RECT 1418.710 1958.300 1419.030 1958.360 ;
        RECT 1408.130 1958.160 1419.030 1958.300 ;
        RECT 1408.130 1958.100 1408.450 1958.160 ;
        RECT 1418.710 1958.100 1419.030 1958.160 ;
        RECT 1408.130 1950.820 1408.450 1950.880 ;
        RECT 1418.250 1950.820 1418.570 1950.880 ;
        RECT 1408.130 1950.680 1418.570 1950.820 ;
        RECT 1408.130 1950.620 1408.450 1950.680 ;
        RECT 1418.250 1950.620 1418.570 1950.680 ;
        RECT 1408.130 1945.380 1408.450 1945.440 ;
        RECT 1417.790 1945.380 1418.110 1945.440 ;
        RECT 1408.130 1945.240 1418.110 1945.380 ;
        RECT 1408.130 1945.180 1408.450 1945.240 ;
        RECT 1417.790 1945.180 1418.110 1945.240 ;
        RECT 1408.130 1941.640 1408.450 1941.700 ;
        RECT 1434.810 1941.640 1435.130 1941.700 ;
        RECT 1408.130 1941.500 1435.130 1941.640 ;
        RECT 1408.130 1941.440 1408.450 1941.500 ;
        RECT 1434.810 1941.440 1435.130 1941.500 ;
        RECT 1408.130 1935.520 1408.450 1935.580 ;
        RECT 1434.350 1935.520 1434.670 1935.580 ;
        RECT 1408.130 1935.380 1434.670 1935.520 ;
        RECT 1408.130 1935.320 1408.450 1935.380 ;
        RECT 1434.350 1935.320 1434.670 1935.380 ;
        RECT 1410.905 1932.120 1411.195 1932.165 ;
        RECT 1411.350 1932.120 1411.670 1932.180 ;
        RECT 1410.905 1931.980 1411.670 1932.120 ;
        RECT 1410.905 1931.935 1411.195 1931.980 ;
        RECT 1411.350 1931.920 1411.670 1931.980 ;
        RECT 1408.130 1930.420 1408.450 1930.480 ;
        RECT 1433.430 1930.420 1433.750 1930.480 ;
        RECT 1408.130 1930.280 1433.750 1930.420 ;
        RECT 1408.130 1930.220 1408.450 1930.280 ;
        RECT 1433.430 1930.220 1433.750 1930.280 ;
        RECT 1408.130 1926.340 1408.450 1926.400 ;
        RECT 1433.890 1926.340 1434.210 1926.400 ;
        RECT 1408.130 1926.200 1434.210 1926.340 ;
        RECT 1408.130 1926.140 1408.450 1926.200 ;
        RECT 1433.890 1926.140 1434.210 1926.200 ;
        RECT 1408.130 1920.220 1408.450 1920.280 ;
        RECT 1421.930 1920.220 1422.250 1920.280 ;
        RECT 1408.130 1920.080 1422.250 1920.220 ;
        RECT 1408.130 1920.020 1408.450 1920.080 ;
        RECT 1421.930 1920.020 1422.250 1920.080 ;
        RECT 1408.130 1916.480 1408.450 1916.540 ;
        RECT 1422.390 1916.480 1422.710 1916.540 ;
        RECT 1408.130 1916.340 1422.710 1916.480 ;
        RECT 1408.130 1916.280 1408.450 1916.340 ;
        RECT 1422.390 1916.280 1422.710 1916.340 ;
        RECT 1409.050 1911.040 1409.370 1911.100 ;
        RECT 1697.470 1911.040 1697.790 1911.100 ;
        RECT 1409.050 1910.900 1697.790 1911.040 ;
        RECT 1409.050 1910.840 1409.370 1910.900 ;
        RECT 1697.470 1910.840 1697.790 1910.900 ;
        RECT 1408.130 1910.700 1408.450 1910.760 ;
        RECT 1421.470 1910.700 1421.790 1910.760 ;
        RECT 1408.130 1910.560 1421.790 1910.700 ;
        RECT 1408.130 1910.500 1408.450 1910.560 ;
        RECT 1421.470 1910.500 1421.790 1910.560 ;
        RECT 1408.130 1904.240 1408.450 1904.300 ;
        RECT 1690.570 1904.240 1690.890 1904.300 ;
        RECT 1408.130 1904.100 1690.890 1904.240 ;
        RECT 1408.130 1904.040 1408.450 1904.100 ;
        RECT 1690.570 1904.040 1690.890 1904.100 ;
        RECT 1408.130 1897.440 1408.450 1897.500 ;
        RECT 1684.130 1897.440 1684.450 1897.500 ;
        RECT 1408.130 1897.300 1684.450 1897.440 ;
        RECT 1408.130 1897.240 1408.450 1897.300 ;
        RECT 1684.130 1897.240 1684.450 1897.300 ;
        RECT 1408.130 1890.640 1408.450 1890.700 ;
        RECT 1683.670 1890.640 1683.990 1890.700 ;
        RECT 1408.130 1890.500 1683.990 1890.640 ;
        RECT 1408.130 1890.440 1408.450 1890.500 ;
        RECT 1683.670 1890.440 1683.990 1890.500 ;
        RECT 1409.050 1890.300 1409.370 1890.360 ;
        RECT 1676.770 1890.300 1677.090 1890.360 ;
        RECT 1409.050 1890.160 1677.090 1890.300 ;
        RECT 1409.050 1890.100 1409.370 1890.160 ;
        RECT 1676.770 1890.100 1677.090 1890.160 ;
        RECT 1408.130 1883.500 1408.450 1883.560 ;
        RECT 1669.870 1883.500 1670.190 1883.560 ;
        RECT 1408.130 1883.360 1670.190 1883.500 ;
        RECT 1408.130 1883.300 1408.450 1883.360 ;
        RECT 1669.870 1883.300 1670.190 1883.360 ;
        RECT 1408.130 1876.700 1408.450 1876.760 ;
        RECT 1662.970 1876.700 1663.290 1876.760 ;
        RECT 1408.130 1876.560 1663.290 1876.700 ;
        RECT 1408.130 1876.500 1408.450 1876.560 ;
        RECT 1662.970 1876.500 1663.290 1876.560 ;
        RECT 1409.050 1869.900 1409.370 1869.960 ;
        RECT 1649.630 1869.900 1649.950 1869.960 ;
        RECT 1409.050 1869.760 1649.950 1869.900 ;
        RECT 1409.050 1869.700 1409.370 1869.760 ;
        RECT 1649.630 1869.700 1649.950 1869.760 ;
        RECT 1408.130 1865.820 1408.450 1865.880 ;
        RECT 1438.950 1865.820 1439.270 1865.880 ;
        RECT 1408.130 1865.680 1439.270 1865.820 ;
        RECT 1408.130 1865.620 1408.450 1865.680 ;
        RECT 1438.950 1865.620 1439.270 1865.680 ;
        RECT 1408.130 1859.700 1408.450 1859.760 ;
        RECT 1432.970 1859.700 1433.290 1859.760 ;
        RECT 1408.130 1859.560 1433.290 1859.700 ;
        RECT 1408.130 1859.500 1408.450 1859.560 ;
        RECT 1432.970 1859.500 1433.290 1859.560 ;
        RECT 1409.050 1855.960 1409.370 1856.020 ;
        RECT 1635.370 1855.960 1635.690 1856.020 ;
        RECT 1409.050 1855.820 1635.690 1855.960 ;
        RECT 1409.050 1855.760 1409.370 1855.820 ;
        RECT 1635.370 1855.760 1635.690 1855.820 ;
        RECT 1408.130 1854.940 1408.450 1855.000 ;
        RECT 1425.610 1854.940 1425.930 1855.000 ;
        RECT 1408.130 1854.800 1425.930 1854.940 ;
        RECT 1408.130 1854.740 1408.450 1854.800 ;
        RECT 1425.610 1854.740 1425.930 1854.800 ;
        RECT 1411.350 1849.500 1411.670 1849.560 ;
        RECT 1411.155 1849.360 1411.670 1849.500 ;
        RECT 1411.350 1849.300 1411.670 1849.360 ;
        RECT 1408.130 1849.160 1408.450 1849.220 ;
        RECT 1628.470 1849.160 1628.790 1849.220 ;
        RECT 1408.130 1849.020 1628.790 1849.160 ;
        RECT 1408.130 1848.960 1408.450 1849.020 ;
        RECT 1628.470 1848.960 1628.790 1849.020 ;
        RECT 1408.130 1842.360 1408.450 1842.420 ;
        RECT 1576.490 1842.360 1576.810 1842.420 ;
        RECT 1408.130 1842.220 1576.810 1842.360 ;
        RECT 1408.130 1842.160 1408.450 1842.220 ;
        RECT 1576.490 1842.160 1576.810 1842.220 ;
        RECT 1410.890 1835.900 1411.210 1835.960 ;
        RECT 1411.365 1835.900 1411.655 1835.945 ;
        RECT 1410.890 1835.760 1411.655 1835.900 ;
        RECT 1410.890 1835.700 1411.210 1835.760 ;
        RECT 1411.365 1835.715 1411.655 1835.760 ;
        RECT 1410.430 1835.020 1410.750 1835.280 ;
        RECT 1422.390 1835.220 1422.710 1835.280 ;
        RECT 1562.690 1835.220 1563.010 1835.280 ;
        RECT 1422.390 1835.080 1563.010 1835.220 ;
        RECT 1422.390 1835.020 1422.710 1835.080 ;
        RECT 1562.690 1835.020 1563.010 1835.080 ;
        RECT 1410.520 1834.585 1410.660 1835.020 ;
        RECT 1425.610 1834.880 1425.930 1834.940 ;
        RECT 1548.890 1834.880 1549.210 1834.940 ;
        RECT 1425.610 1834.740 1549.210 1834.880 ;
        RECT 1425.610 1834.680 1425.930 1834.740 ;
        RECT 1548.890 1834.680 1549.210 1834.740 ;
        RECT 1410.445 1834.355 1410.735 1834.585 ;
        RECT 1408.130 1828.420 1408.450 1828.480 ;
        RECT 1652.390 1828.420 1652.710 1828.480 ;
        RECT 1408.130 1828.280 1652.710 1828.420 ;
        RECT 1408.130 1828.220 1408.450 1828.280 ;
        RECT 1652.390 1828.220 1652.710 1828.280 ;
        RECT 1411.350 1825.020 1411.670 1825.080 ;
        RECT 1413.650 1825.020 1413.970 1825.080 ;
        RECT 1411.350 1824.880 1413.970 1825.020 ;
        RECT 1411.350 1824.820 1411.670 1824.880 ;
        RECT 1413.650 1824.820 1413.970 1824.880 ;
        RECT 1408.130 1821.620 1408.450 1821.680 ;
        RECT 1646.410 1821.620 1646.730 1821.680 ;
        RECT 1408.130 1821.480 1646.730 1821.620 ;
        RECT 1408.130 1821.420 1408.450 1821.480 ;
        RECT 1646.410 1821.420 1646.730 1821.480 ;
        RECT 1408.130 1814.480 1408.450 1814.540 ;
        RECT 1645.490 1814.480 1645.810 1814.540 ;
        RECT 1408.130 1814.340 1645.810 1814.480 ;
        RECT 1408.130 1814.280 1408.450 1814.340 ;
        RECT 1645.490 1814.280 1645.810 1814.340 ;
        RECT 1409.050 1814.140 1409.370 1814.200 ;
        RECT 1638.590 1814.140 1638.910 1814.200 ;
        RECT 1409.050 1814.000 1638.910 1814.140 ;
        RECT 1409.050 1813.940 1409.370 1814.000 ;
        RECT 1638.590 1813.940 1638.910 1814.000 ;
        RECT 1408.130 1807.680 1408.450 1807.740 ;
        RECT 1631.690 1807.680 1632.010 1807.740 ;
        RECT 1408.130 1807.540 1632.010 1807.680 ;
        RECT 1408.130 1807.480 1408.450 1807.540 ;
        RECT 1631.690 1807.480 1632.010 1807.540 ;
        RECT 1408.130 1800.880 1408.450 1800.940 ;
        RECT 1624.790 1800.880 1625.110 1800.940 ;
        RECT 1408.130 1800.740 1625.110 1800.880 ;
        RECT 1408.130 1800.680 1408.450 1800.740 ;
        RECT 1624.790 1800.680 1625.110 1800.740 ;
        RECT 1409.050 1800.540 1409.370 1800.600 ;
        RECT 1617.890 1800.540 1618.210 1800.600 ;
        RECT 1409.050 1800.400 1618.210 1800.540 ;
        RECT 1409.050 1800.340 1409.370 1800.400 ;
        RECT 1617.890 1800.340 1618.210 1800.400 ;
        RECT 1408.130 1793.740 1408.450 1793.800 ;
        RECT 1610.990 1793.740 1611.310 1793.800 ;
        RECT 1408.130 1793.600 1611.310 1793.740 ;
        RECT 1408.130 1793.540 1408.450 1793.600 ;
        RECT 1610.990 1793.540 1611.310 1793.600 ;
        RECT 1410.445 1787.280 1410.735 1787.325 ;
        RECT 1410.890 1787.280 1411.210 1787.340 ;
        RECT 1410.445 1787.140 1411.210 1787.280 ;
        RECT 1410.445 1787.095 1410.735 1787.140 ;
        RECT 1410.890 1787.080 1411.210 1787.140 ;
        RECT 1408.130 1759.060 1408.450 1759.120 ;
        RECT 1432.510 1759.060 1432.830 1759.120 ;
        RECT 1408.130 1758.920 1432.830 1759.060 ;
        RECT 1408.130 1758.860 1408.450 1758.920 ;
        RECT 1432.510 1758.860 1432.830 1758.920 ;
        RECT 1408.130 1754.640 1408.450 1754.700 ;
        RECT 1432.050 1754.640 1432.370 1754.700 ;
        RECT 1408.130 1754.500 1432.370 1754.640 ;
        RECT 1408.130 1754.440 1408.450 1754.500 ;
        RECT 1432.050 1754.440 1432.370 1754.500 ;
        RECT 1408.130 1751.580 1408.450 1751.640 ;
        RECT 1422.850 1751.580 1423.170 1751.640 ;
        RECT 1408.130 1751.440 1423.170 1751.580 ;
        RECT 1408.130 1751.380 1408.450 1751.440 ;
        RECT 1422.850 1751.380 1423.170 1751.440 ;
        RECT 1408.130 1745.460 1408.450 1745.520 ;
        RECT 1459.190 1745.460 1459.510 1745.520 ;
        RECT 1408.130 1745.320 1459.510 1745.460 ;
        RECT 1408.130 1745.260 1408.450 1745.320 ;
        RECT 1459.190 1745.260 1459.510 1745.320 ;
        RECT 1408.130 1738.660 1408.450 1738.720 ;
        RECT 1452.290 1738.660 1452.610 1738.720 ;
        RECT 1408.130 1738.520 1452.610 1738.660 ;
        RECT 1408.130 1738.460 1408.450 1738.520 ;
        RECT 1452.290 1738.460 1452.610 1738.520 ;
        RECT 1408.130 1733.900 1408.450 1733.960 ;
        RECT 1438.490 1733.900 1438.810 1733.960 ;
        RECT 1408.130 1733.760 1438.810 1733.900 ;
        RECT 1408.130 1733.700 1408.450 1733.760 ;
        RECT 1438.490 1733.700 1438.810 1733.760 ;
        RECT 1408.130 1728.460 1408.450 1728.520 ;
        RECT 1431.590 1728.460 1431.910 1728.520 ;
        RECT 1408.130 1728.320 1431.910 1728.460 ;
        RECT 1408.130 1728.260 1408.450 1728.320 ;
        RECT 1431.590 1728.260 1431.910 1728.320 ;
        RECT 1408.130 1724.380 1408.450 1724.440 ;
        RECT 1424.690 1724.380 1425.010 1724.440 ;
        RECT 1408.130 1724.240 1425.010 1724.380 ;
        RECT 1408.130 1724.180 1408.450 1724.240 ;
        RECT 1424.690 1724.180 1425.010 1724.240 ;
        RECT 1408.130 1717.920 1408.450 1717.980 ;
        RECT 1535.090 1717.920 1535.410 1717.980 ;
        RECT 1408.130 1717.780 1535.410 1717.920 ;
        RECT 1408.130 1717.720 1408.450 1717.780 ;
        RECT 1535.090 1717.720 1535.410 1717.780 ;
        RECT 1409.050 1717.580 1409.370 1717.640 ;
        RECT 1459.650 1717.580 1459.970 1717.640 ;
        RECT 1409.050 1717.440 1459.970 1717.580 ;
        RECT 1409.050 1717.380 1409.370 1717.440 ;
        RECT 1459.650 1717.380 1459.970 1717.440 ;
        RECT 1408.130 1711.120 1408.450 1711.180 ;
        RECT 1541.990 1711.120 1542.310 1711.180 ;
        RECT 1408.130 1710.980 1542.310 1711.120 ;
        RECT 1408.130 1710.920 1408.450 1710.980 ;
        RECT 1541.990 1710.920 1542.310 1710.980 ;
        RECT 1411.350 1704.320 1411.670 1704.380 ;
        RECT 1412.270 1704.320 1412.590 1704.380 ;
        RECT 1411.350 1704.180 1412.590 1704.320 ;
        RECT 1411.350 1704.120 1411.670 1704.180 ;
        RECT 1412.270 1704.120 1412.590 1704.180 ;
        RECT 1408.130 1703.980 1408.450 1704.040 ;
        RECT 1423.770 1703.980 1424.090 1704.040 ;
        RECT 1408.130 1703.840 1424.090 1703.980 ;
        RECT 1408.130 1703.780 1408.450 1703.840 ;
        RECT 1423.770 1703.780 1424.090 1703.840 ;
        RECT 1408.590 1703.300 1408.910 1703.360 ;
        RECT 1423.310 1703.300 1423.630 1703.360 ;
        RECT 1408.590 1703.160 1423.630 1703.300 ;
        RECT 1408.590 1703.100 1408.910 1703.160 ;
        RECT 1423.310 1703.100 1423.630 1703.160 ;
        RECT 1408.130 1694.120 1408.450 1694.180 ;
        RECT 1424.230 1694.120 1424.550 1694.180 ;
        RECT 1408.130 1693.980 1424.550 1694.120 ;
        RECT 1408.130 1693.920 1408.450 1693.980 ;
        RECT 1424.230 1693.920 1424.550 1693.980 ;
        RECT 1411.825 1690.380 1412.115 1690.425 ;
        RECT 1412.270 1690.380 1412.590 1690.440 ;
        RECT 1411.825 1690.240 1412.590 1690.380 ;
        RECT 1411.825 1690.195 1412.115 1690.240 ;
        RECT 1412.270 1690.180 1412.590 1690.240 ;
        RECT 1408.130 1689.700 1408.450 1689.760 ;
        RECT 1427.910 1689.700 1428.230 1689.760 ;
        RECT 1408.130 1689.560 1428.230 1689.700 ;
        RECT 1408.130 1689.500 1408.450 1689.560 ;
        RECT 1427.910 1689.500 1428.230 1689.560 ;
        RECT 1408.590 1683.580 1408.910 1683.640 ;
        RECT 1426.990 1683.580 1427.310 1683.640 ;
        RECT 1408.590 1683.440 1427.310 1683.580 ;
        RECT 1408.590 1683.380 1408.910 1683.440 ;
        RECT 1426.990 1683.380 1427.310 1683.440 ;
        RECT 1408.130 1682.900 1408.450 1682.960 ;
        RECT 1427.450 1682.900 1427.770 1682.960 ;
        RECT 1408.130 1682.760 1427.770 1682.900 ;
        RECT 1408.130 1682.700 1408.450 1682.760 ;
        RECT 1427.450 1682.700 1427.770 1682.760 ;
        RECT 1408.130 1673.040 1408.450 1673.100 ;
        RECT 1426.530 1673.040 1426.850 1673.100 ;
        RECT 1408.130 1672.900 1426.850 1673.040 ;
        RECT 1408.130 1672.840 1408.450 1672.900 ;
        RECT 1426.530 1672.840 1426.850 1672.900 ;
        RECT 1408.590 1669.640 1408.910 1669.700 ;
        RECT 1514.390 1669.640 1514.710 1669.700 ;
        RECT 1408.590 1669.500 1514.710 1669.640 ;
        RECT 1408.590 1669.440 1408.910 1669.500 ;
        RECT 1514.390 1669.440 1514.710 1669.500 ;
        RECT 1408.130 1668.280 1408.450 1668.340 ;
        RECT 1426.070 1668.280 1426.390 1668.340 ;
        RECT 1408.130 1668.140 1426.390 1668.280 ;
        RECT 1408.130 1668.080 1408.450 1668.140 ;
        RECT 1426.070 1668.080 1426.390 1668.140 ;
        RECT 1408.130 1656.040 1408.450 1656.100 ;
        RECT 1601.330 1656.040 1601.650 1656.100 ;
        RECT 1408.130 1655.900 1601.650 1656.040 ;
        RECT 1408.130 1655.840 1408.450 1655.900 ;
        RECT 1601.330 1655.840 1601.650 1655.900 ;
        RECT 1407.670 1648.900 1407.990 1648.960 ;
        RECT 1600.870 1648.900 1601.190 1648.960 ;
        RECT 1407.670 1648.760 1601.190 1648.900 ;
        RECT 1407.670 1648.700 1407.990 1648.760 ;
        RECT 1600.870 1648.700 1601.190 1648.760 ;
        RECT 1408.130 1648.560 1408.450 1648.620 ;
        RECT 1593.970 1648.560 1594.290 1648.620 ;
        RECT 1408.130 1648.420 1594.290 1648.560 ;
        RECT 1408.130 1648.360 1408.450 1648.420 ;
        RECT 1593.970 1648.360 1594.290 1648.420 ;
        RECT 1411.810 1642.440 1412.130 1642.500 ;
        RECT 1411.615 1642.300 1412.130 1642.440 ;
        RECT 1411.810 1642.240 1412.130 1642.300 ;
        RECT 1407.670 1642.100 1407.990 1642.160 ;
        RECT 1587.070 1642.100 1587.390 1642.160 ;
        RECT 1407.670 1641.960 1587.390 1642.100 ;
        RECT 1407.670 1641.900 1407.990 1641.960 ;
        RECT 1587.070 1641.900 1587.390 1641.960 ;
        RECT 1407.670 1627.820 1407.990 1627.880 ;
        RECT 1425.150 1627.820 1425.470 1627.880 ;
        RECT 1407.670 1627.680 1425.470 1627.820 ;
        RECT 1407.670 1627.620 1407.990 1627.680 ;
        RECT 1425.150 1627.620 1425.470 1627.680 ;
        RECT 1414.110 1607.760 1414.430 1607.820 ;
        RECT 1693.790 1607.760 1694.110 1607.820 ;
        RECT 1414.110 1607.620 1694.110 1607.760 ;
        RECT 1414.110 1607.560 1414.430 1607.620 ;
        RECT 1693.790 1607.560 1694.110 1607.620 ;
      LAYER met1 ;
        RECT 1705.000 1605.000 2081.480 2051.235 ;
        RECT 2255.000 1605.000 2631.480 2051.235 ;
        RECT 1550.070 404.460 2645.190 1495.780 ;
      LAYER via ;
        RECT 1318.000 3266.760 1318.260 3267.020 ;
        RECT 1890.700 3266.760 1890.960 3267.020 ;
        RECT 1917.840 3266.760 1918.100 3267.020 ;
        RECT 2542.060 3266.760 2542.320 3267.020 ;
        RECT 1890.700 3264.380 1890.960 3264.640 ;
        RECT 1917.840 3264.380 1918.100 3264.640 ;
        RECT 675.840 3263.700 676.100 3263.960 ;
        RECT 697.000 3264.040 697.260 3264.300 ;
        RECT 2542.060 3264.040 2542.320 3264.300 ;
        RECT 2566.900 3264.040 2567.160 3264.300 ;
        RECT 1292.700 3263.700 1292.960 3263.960 ;
        RECT 2594.500 3263.700 2594.760 3263.960 ;
        RECT 1333.180 3252.140 1333.440 3252.400 ;
        RECT 2038.820 3252.480 2039.080 3252.740 ;
        RECT 1935.780 3252.140 1936.040 3252.400 ;
        RECT 688.260 3251.120 688.520 3251.380 ;
        RECT 2582.080 3252.140 2582.340 3252.400 ;
        RECT 1459.220 3229.360 1459.480 3229.620 ;
        RECT 1536.960 3229.360 1537.220 3229.620 ;
        RECT 1452.320 3222.220 1452.580 3222.480 ;
        RECT 1535.580 3222.220 1535.840 3222.480 ;
        RECT 1438.520 3215.420 1438.780 3215.680 ;
        RECT 1535.580 3215.420 1535.840 3215.680 ;
        RECT 1431.620 3208.620 1431.880 3208.880 ;
        RECT 1538.340 3208.620 1538.600 3208.880 ;
        RECT 1424.720 3201.480 1424.980 3201.740 ;
        RECT 1538.340 3201.480 1538.600 3201.740 ;
        RECT 1459.680 3187.880 1459.940 3188.140 ;
        RECT 1534.200 3187.880 1534.460 3188.140 ;
        RECT 1352.040 2901.260 1352.300 2901.520 ;
        RECT 1395.740 2901.260 1396.000 2901.520 ;
        RECT 1514.420 2898.200 1514.680 2898.460 ;
        RECT 1538.340 2898.200 1538.600 2898.460 ;
        RECT 1945.900 3250.780 1946.160 3251.040 ;
        RECT 386.960 2794.160 387.220 2794.420 ;
        RECT 431.580 2794.160 431.840 2794.420 ;
        RECT 433.420 2794.160 433.680 2794.420 ;
        RECT 468.840 2794.160 469.100 2794.420 ;
        RECT 686.420 2794.160 686.680 2794.420 ;
        RECT 1738.440 2794.160 1738.700 2794.420 ;
        RECT 1780.300 2794.160 1780.560 2794.420 ;
        RECT 2340.120 2794.160 2340.380 2794.420 ;
        RECT 2382.900 2794.160 2383.160 2794.420 ;
        RECT 330.840 2793.820 331.100 2794.080 ;
        RECT 1001.060 2793.820 1001.320 2794.080 ;
        RECT 1076.500 2793.820 1076.760 2794.080 ;
        RECT 1122.500 2793.820 1122.760 2794.080 ;
        RECT 1432.080 2793.820 1432.340 2794.080 ;
        RECT 2268.360 2793.820 2268.620 2794.080 ;
        RECT 375.000 2793.480 375.260 2793.740 ;
        RECT 421.000 2793.480 421.260 2793.740 ;
        RECT 466.540 2793.480 466.800 2793.740 ;
        RECT 513.920 2793.480 514.180 2793.740 ;
        RECT 531.400 2793.480 531.660 2793.740 ;
        RECT 536.460 2793.480 536.720 2793.740 ;
        RECT 707.120 2793.480 707.380 2793.740 ;
        RECT 1093.980 2793.480 1094.240 2793.740 ;
        RECT 1139.980 2793.480 1140.240 2793.740 ;
        RECT 1186.900 2793.480 1187.160 2793.740 ;
        RECT 1432.540 2793.480 1432.800 2793.740 ;
        RECT 2273.880 2793.480 2274.140 2793.740 ;
        RECT 392.480 2793.140 392.740 2793.400 ;
        RECT 439.400 2793.140 439.660 2793.400 ;
        RECT 485.860 2793.140 486.120 2793.400 ;
        RECT 497.360 2793.140 497.620 2793.400 ;
        RECT 510.240 2793.140 510.500 2793.400 ;
        RECT 700.220 2793.140 700.480 2793.400 ;
        RECT 1111.000 2793.140 1111.260 2793.400 ;
        RECT 1159.300 2793.140 1159.560 2793.400 ;
        RECT 1631.720 2793.140 1631.980 2793.400 ;
        RECT 1677.260 2793.140 1677.520 2793.400 ;
        RECT 1721.420 2793.140 1721.680 2793.400 ;
        RECT 1766.500 2793.140 1766.760 2793.400 ;
        RECT 379.600 2792.800 379.860 2793.060 ;
        RECT 426.980 2792.800 427.240 2793.060 ;
        RECT 433.420 2792.800 433.680 2793.060 ;
        RECT 478.500 2792.800 478.760 2793.060 ;
        RECT 397.080 2792.460 397.340 2792.720 ;
        RECT 444.460 2792.460 444.720 2792.720 ;
        RECT 491.840 2792.460 492.100 2792.720 ;
        RECT 520.820 2792.800 521.080 2793.060 ;
        RECT 542.440 2792.800 542.700 2793.060 ;
        RECT 741.620 2792.800 741.880 2793.060 ;
        RECT 1087.540 2792.800 1087.800 2793.060 ;
        RECT 1129.400 2792.800 1129.660 2793.060 ;
        RECT 1173.100 2792.800 1173.360 2793.060 ;
        RECT 1680.480 2792.800 1680.740 2793.060 ;
        RECT 1683.240 2792.800 1683.500 2793.060 ;
        RECT 1730.160 2792.800 1730.420 2793.060 ;
        RECT 1773.400 2792.800 1773.660 2793.060 ;
        RECT 2287.220 2793.820 2287.480 2794.080 ;
        RECT 2332.760 2793.820 2333.020 2794.080 ;
        RECT 2377.380 2793.820 2377.640 2794.080 ;
        RECT 2294.120 2793.480 2294.380 2793.740 ;
        RECT 2340.120 2793.480 2340.380 2793.740 ;
        RECT 2340.580 2793.480 2340.840 2793.740 ;
        RECT 2343.800 2793.480 2344.060 2793.740 ;
        RECT 2387.960 2793.480 2388.220 2793.740 ;
        RECT 2280.320 2793.140 2280.580 2793.400 ;
        RECT 2326.320 2793.140 2326.580 2793.400 ;
        RECT 2374.160 2793.140 2374.420 2793.400 ;
        RECT 2422.000 2793.140 2422.260 2793.400 ;
        RECT 2315.280 2792.800 2315.540 2793.060 ;
        RECT 2360.820 2792.800 2361.080 2793.060 ;
        RECT 2408.200 2792.800 2408.460 2793.060 ;
        RECT 403.980 2792.120 404.240 2792.380 ;
        RECT 449.060 2792.120 449.320 2792.380 ;
        RECT 473.900 2792.120 474.160 2792.380 ;
        RECT 500.120 2792.460 500.380 2792.720 ;
        RECT 524.040 2792.460 524.300 2792.720 ;
        RECT 720.920 2792.460 721.180 2792.720 ;
        RECT 1042.460 2792.460 1042.720 2792.720 ;
        RECT 1088.000 2792.460 1088.260 2792.720 ;
        RECT 1135.840 2792.460 1136.100 2792.720 ;
        RECT 1180.000 2792.460 1180.260 2792.720 ;
        RECT 1652.420 2792.460 1652.680 2792.720 ;
        RECT 1699.340 2792.460 1699.600 2792.720 ;
        RECT 1748.560 2792.460 1748.820 2792.720 ;
        RECT 1790.880 2792.460 1791.140 2792.720 ;
        RECT 2266.520 2792.460 2266.780 2792.720 ;
        RECT 2308.380 2792.460 2308.640 2792.720 ;
        RECT 2356.680 2792.460 2356.940 2792.720 ;
        RECT 2401.760 2792.460 2402.020 2792.720 ;
        RECT 700.680 2792.120 700.940 2792.380 ;
        RECT 1065.920 2792.120 1066.180 2792.380 ;
        RECT 1111.000 2792.120 1111.260 2792.380 ;
        RECT 1646.440 2792.120 1646.700 2792.380 ;
        RECT 1695.200 2792.120 1695.460 2792.380 ;
        RECT 1741.200 2792.120 1741.460 2792.380 ;
        RECT 1787.200 2792.120 1787.460 2792.380 ;
        RECT 2273.880 2792.120 2274.140 2792.380 ;
        RECT 2321.260 2792.120 2321.520 2792.380 ;
        RECT 2367.260 2792.120 2367.520 2792.380 ;
        RECT 2415.100 2792.120 2415.360 2792.380 ;
        RECT 368.560 2791.780 368.820 2792.040 ;
        RECT 414.560 2791.780 414.820 2792.040 ;
        RECT 462.400 2791.780 462.660 2792.040 ;
        RECT 465.620 2791.780 465.880 2792.040 ;
        RECT 489.080 2791.780 489.340 2792.040 ;
        RECT 693.320 2791.780 693.580 2792.040 ;
        RECT 1053.040 2791.780 1053.300 2792.040 ;
        RECT 1100.420 2791.780 1100.680 2792.040 ;
        RECT 1147.340 2791.780 1147.600 2792.040 ;
        RECT 407.200 2791.440 407.460 2791.700 ;
        RECT 409.960 2791.440 410.220 2791.700 ;
        RECT 455.500 2791.440 455.760 2791.700 ;
        RECT 461.020 2791.440 461.280 2791.700 ;
        RECT 687.340 2791.440 687.600 2791.700 ;
        RECT 1055.800 2791.440 1056.060 2791.700 ;
        RECT 1059.020 2791.440 1059.280 2791.700 ;
        RECT 1105.480 2791.440 1105.740 2791.700 ;
        RECT 1152.400 2791.440 1152.660 2791.700 ;
        RECT 371.320 2791.100 371.580 2791.360 ;
        RECT 686.880 2791.100 687.140 2791.360 ;
        RECT 1034.640 2791.100 1034.900 2791.360 ;
        RECT 1076.500 2791.100 1076.760 2791.360 ;
        RECT 1122.500 2791.100 1122.760 2791.360 ;
        RECT 1166.200 2791.100 1166.460 2791.360 ;
        RECT 1670.360 2791.780 1670.620 2792.040 ;
        RECT 1676.340 2791.780 1676.600 2792.040 ;
        RECT 1687.840 2791.780 1688.100 2792.040 ;
        RECT 1738.440 2791.780 1738.700 2792.040 ;
        RECT 1762.820 2791.780 1763.080 2792.040 ;
        RECT 2381.060 2791.780 2381.320 2792.040 ;
        RECT 2382.900 2791.780 2383.160 2792.040 ;
        RECT 2428.900 2791.780 2429.160 2792.040 ;
        RECT 1193.800 2791.100 1194.060 2791.360 ;
        RECT 362.580 2790.760 362.840 2791.020 ;
        RECT 407.200 2790.760 407.460 2791.020 ;
        RECT 419.160 2790.760 419.420 2791.020 ;
        RECT 748.520 2790.760 748.780 2791.020 ;
        RECT 1019.000 2790.760 1019.260 2791.020 ;
        RECT 1065.920 2790.760 1066.180 2791.020 ;
        RECT 384.200 2790.420 384.460 2790.680 ;
        RECT 727.820 2790.420 728.080 2790.680 ;
        RECT 1076.040 2790.420 1076.300 2790.680 ;
        RECT 1425.640 2790.420 1425.900 2790.680 ;
        RECT 1642.300 2790.420 1642.560 2790.680 ;
        RECT 406.280 2790.080 406.540 2790.340 ;
        RECT 762.780 2790.080 763.040 2790.340 ;
        RECT 1159.300 2790.080 1159.560 2790.340 ;
        RECT 1562.720 2790.080 1562.980 2790.340 ;
        RECT 1614.700 2790.080 1614.960 2790.340 ;
        RECT 1617.920 2790.080 1618.180 2790.340 ;
        RECT 1665.760 2791.440 1666.020 2791.700 ;
        RECT 1712.680 2791.440 1712.940 2791.700 ;
        RECT 1742.120 2791.440 1742.380 2791.700 ;
        RECT 1763.280 2791.440 1763.540 2791.700 ;
        RECT 2387.500 2791.440 2387.760 2791.700 ;
        RECT 2387.960 2791.440 2388.220 2791.700 ;
        RECT 2435.800 2791.440 2436.060 2791.700 ;
        RECT 396.620 2789.740 396.880 2790.000 ;
        RECT 762.320 2789.740 762.580 2790.000 ;
        RECT 1548.920 2789.740 1549.180 2790.000 ;
        RECT 1607.800 2789.740 1608.060 2790.000 ;
        RECT 1611.020 2789.740 1611.280 2790.000 ;
        RECT 1658.860 2791.100 1659.120 2791.360 ;
        RECT 1706.240 2791.100 1706.500 2791.360 ;
        RECT 1752.700 2791.100 1752.960 2791.360 ;
        RECT 1769.720 2791.100 1769.980 2791.360 ;
        RECT 2394.400 2791.100 2394.660 2791.360 ;
        RECT 2394.860 2791.100 2395.120 2791.360 ;
        RECT 2442.700 2791.100 2442.960 2791.360 ;
        RECT 1676.340 2790.760 1676.600 2791.020 ;
        RECT 1718.200 2790.760 1718.460 2791.020 ;
        RECT 1760.060 2790.760 1760.320 2791.020 ;
        RECT 1770.180 2790.760 1770.440 2791.020 ;
        RECT 2401.760 2790.760 2402.020 2791.020 ;
        RECT 1783.520 2790.420 1783.780 2790.680 ;
        RECT 2415.100 2790.420 2415.360 2790.680 ;
        RECT 1776.620 2790.080 1776.880 2790.340 ;
        RECT 2408.200 2790.080 2408.460 2790.340 ;
        RECT 1783.980 2789.740 1784.240 2790.000 ;
        RECT 2422.000 2789.740 2422.260 2790.000 ;
        RECT 485.860 2789.400 486.120 2789.660 ;
        RECT 527.720 2789.400 527.980 2789.660 ;
        RECT 648.240 2789.400 648.500 2789.660 ;
        RECT 1117.900 2789.400 1118.160 2789.660 ;
        RECT 1433.000 2789.400 1433.260 2789.660 ;
        RECT 1649.200 2789.400 1649.460 2789.660 ;
        RECT 1777.080 2789.400 1777.340 2789.660 ;
        RECT 2415.100 2789.400 2415.360 2789.660 ;
        RECT 445.840 2789.060 446.100 2789.320 ;
        RECT 465.620 2788.720 465.880 2788.980 ;
        RECT 504.260 2788.720 504.520 2788.980 ;
        RECT 627.540 2789.060 627.800 2789.320 ;
        RECT 1042.460 2789.060 1042.720 2789.320 ;
        RECT 1624.820 2789.060 1625.080 2789.320 ;
        RECT 1790.420 2789.060 1790.680 2789.320 ;
        RECT 2428.900 2789.060 2429.160 2789.320 ;
        RECT 606.840 2788.720 607.100 2788.980 ;
        RECT 1034.640 2788.720 1034.900 2788.980 ;
        RECT 1045.220 2788.720 1045.480 2788.980 ;
        RECT 1093.980 2788.720 1094.240 2788.980 ;
        RECT 1438.980 2788.720 1439.240 2788.980 ;
        RECT 1656.100 2788.720 1656.360 2788.980 ;
        RECT 1790.880 2788.720 1791.140 2788.980 ;
        RECT 2435.800 2788.720 2436.060 2788.980 ;
        RECT 426.980 2788.380 427.240 2788.640 ;
        RECT 473.900 2788.380 474.160 2788.640 ;
        RECT 491.840 2788.380 492.100 2788.640 ;
        RECT 541.520 2788.380 541.780 2788.640 ;
        RECT 586.140 2788.380 586.400 2788.640 ;
        RECT 1019.000 2788.380 1019.260 2788.640 ;
        RECT 1024.520 2788.380 1024.780 2788.640 ;
        RECT 1070.060 2788.380 1070.320 2788.640 ;
        RECT 1076.040 2788.380 1076.300 2788.640 ;
        RECT 1425.180 2788.380 1425.440 2788.640 ;
        RECT 2249.500 2788.380 2249.760 2788.640 ;
        RECT 2301.940 2788.380 2302.200 2788.640 ;
        RECT 2340.580 2788.380 2340.840 2788.640 ;
        RECT 2374.160 2788.380 2374.420 2788.640 ;
        RECT 2415.100 2788.380 2415.360 2788.640 ;
        RECT 455.500 2788.040 455.760 2788.300 ;
        RECT 500.120 2788.040 500.380 2788.300 ;
        RECT 501.960 2788.040 502.220 2788.300 ;
        RECT 542.440 2788.040 542.700 2788.300 ;
        RECT 1010.720 2788.040 1010.980 2788.300 ;
        RECT 1055.800 2788.040 1056.060 2788.300 ;
        RECT 1576.520 2788.040 1576.780 2788.300 ;
        RECT 1621.600 2788.040 1621.860 2788.300 ;
        RECT 1638.620 2788.040 1638.880 2788.300 ;
        RECT 1680.480 2788.040 1680.740 2788.300 ;
        RECT 2301.020 2788.040 2301.280 2788.300 ;
        RECT 2304.240 2788.040 2304.500 2788.300 ;
        RECT 2350.240 2788.040 2350.500 2788.300 ;
        RECT 2394.860 2788.040 2395.120 2788.300 ;
        RECT 337.280 2787.700 337.540 2787.960 ;
        RECT 1007.500 2787.700 1007.760 2787.960 ;
        RECT 1038.320 2787.700 1038.580 2787.960 ;
        RECT 1087.540 2787.700 1087.800 2787.960 ;
        RECT 1542.020 2787.700 1542.280 2787.960 ;
        RECT 1581.580 2787.700 1581.840 2787.960 ;
        RECT 1645.520 2787.700 1645.780 2787.960 ;
        RECT 1687.840 2787.700 1688.100 2787.960 ;
        RECT 2321.720 2787.700 2321.980 2787.960 ;
        RECT 2442.700 2787.700 2442.960 2787.960 ;
        RECT 658.820 2784.300 659.080 2784.560 ;
        RECT 482.640 2725.140 482.900 2725.400 ;
        RECT 948.160 2725.140 948.420 2725.400 ;
        RECT 470.680 2724.800 470.940 2725.060 ;
        RECT 942.180 2724.800 942.440 2725.060 ;
        RECT 510.240 2724.460 510.500 2724.720 ;
        RECT 989.560 2724.460 989.820 2724.720 ;
        RECT 460.560 2724.120 460.820 2724.380 ;
        RECT 942.640 2724.120 942.900 2724.380 ;
        RECT 449.980 2723.780 450.240 2724.040 ;
        RECT 943.100 2723.780 943.360 2724.040 ;
        RECT 530.940 2723.440 531.200 2723.700 ;
        RECT 1030.960 2723.440 1031.220 2723.700 ;
        RECT 439.860 2723.100 440.120 2723.360 ;
        RECT 943.560 2723.100 943.820 2723.360 ;
        RECT 551.640 2722.760 551.900 2723.020 ;
        RECT 1062.240 2722.760 1062.500 2723.020 ;
        RECT 429.280 2722.420 429.540 2722.680 ;
        RECT 944.020 2722.420 944.280 2722.680 ;
        RECT 419.160 2722.080 419.420 2722.340 ;
        RECT 944.480 2722.080 944.740 2722.340 ;
        RECT 408.580 2721.740 408.840 2722.000 ;
        RECT 979.900 2721.740 980.160 2722.000 ;
        RECT 433.880 2721.400 434.140 2721.660 ;
        RECT 865.360 2721.400 865.620 2721.660 ;
        RECT 441.240 2721.060 441.500 2721.320 ;
        RECT 875.480 2721.060 875.740 2721.320 ;
        RECT 427.440 2720.720 427.700 2720.980 ;
        RECT 844.200 2720.720 844.460 2720.980 ;
        RECT 434.340 2720.380 434.600 2720.640 ;
        RECT 854.780 2720.380 855.040 2720.640 ;
        RECT 413.640 2720.040 413.900 2720.300 ;
        RECT 823.500 2720.040 823.760 2720.300 ;
        RECT 365.340 2719.700 365.600 2719.960 ;
        RECT 740.700 2719.700 740.960 2719.960 ;
        RECT 289.440 2719.360 289.700 2719.620 ;
        RECT 564.060 2719.360 564.320 2719.620 ;
        RECT 288.980 2719.020 289.240 2719.280 ;
        RECT 553.940 2719.020 554.200 2719.280 ;
        RECT 1103.640 2718.680 1103.900 2718.940 ;
        RECT 358.440 2718.340 358.700 2718.600 ;
        RECT 377.300 2718.340 377.560 2718.600 ;
        RECT 379.140 2718.340 379.400 2718.600 ;
        RECT 727.820 2718.340 728.080 2718.600 ;
        RECT 762.780 2718.340 763.040 2718.600 ;
        RECT 813.380 2718.340 813.640 2718.600 ;
        RECT 1027.740 2718.340 1028.000 2718.600 ;
        RECT 1093.520 2718.340 1093.780 2718.600 ;
        RECT 1102.720 2718.340 1102.980 2718.600 ;
        RECT 1145.040 2718.340 1145.300 2718.600 ;
        RECT 1300.980 2718.340 1301.240 2718.600 ;
        RECT 351.540 2718.000 351.800 2718.260 ;
        RECT 367.180 2718.000 367.440 2718.260 ;
        RECT 392.940 2718.000 393.200 2718.260 ;
        RECT 782.100 2718.000 782.360 2718.260 ;
        RECT 1034.640 2718.000 1034.900 2718.260 ;
        RECT 1103.640 2718.000 1103.900 2718.260 ;
        RECT 1138.140 2718.000 1138.400 2718.260 ;
        RECT 1290.400 2718.000 1290.660 2718.260 ;
        RECT 305.080 2717.660 305.340 2717.920 ;
        RECT 310.140 2717.660 310.400 2717.920 ;
        RECT 325.780 2717.660 326.040 2717.920 ;
        RECT 330.840 2717.660 331.100 2717.920 ;
        RECT 351.080 2717.660 351.340 2717.920 ;
        RECT 356.600 2717.660 356.860 2717.920 ;
        RECT 399.380 2717.660 399.640 2717.920 ;
        RECT 762.320 2717.660 762.580 2717.920 ;
        RECT 792.680 2717.660 792.940 2717.920 ;
        RECT 1041.540 2717.660 1041.800 2717.920 ;
        RECT 1114.220 2717.660 1114.480 2717.920 ;
        RECT 1151.940 2717.660 1152.200 2717.920 ;
        RECT 1311.100 2717.660 1311.360 2717.920 ;
        RECT 287.140 2717.320 287.400 2717.580 ;
        RECT 512.540 2717.320 512.800 2717.580 ;
        RECT 636.740 2717.320 637.000 2717.580 ;
        RECT 1045.220 2717.320 1045.480 2717.580 ;
        RECT 1048.440 2717.320 1048.700 2717.580 ;
        RECT 1124.340 2717.320 1124.600 2717.580 ;
        RECT 1158.840 2717.320 1159.100 2717.580 ;
        RECT 1321.680 2717.320 1321.940 2717.580 ;
        RECT 287.600 2716.980 287.860 2717.240 ;
        RECT 522.660 2716.980 522.920 2717.240 ;
        RECT 616.040 2716.980 616.300 2717.240 ;
        RECT 1038.320 2716.980 1038.580 2717.240 ;
        RECT 1055.340 2716.980 1055.600 2717.240 ;
        RECT 1134.920 2716.980 1135.180 2717.240 ;
        RECT 1165.740 2716.980 1166.000 2717.240 ;
        RECT 1332.260 2716.980 1332.520 2717.240 ;
        RECT 288.060 2716.640 288.320 2716.900 ;
        RECT 533.240 2716.640 533.500 2716.900 ;
        RECT 595.340 2716.640 595.600 2716.900 ;
        RECT 1024.520 2716.640 1024.780 2716.900 ;
        RECT 1061.780 2716.640 1062.040 2716.900 ;
        RECT 1155.620 2716.640 1155.880 2716.900 ;
        RECT 1165.280 2716.640 1165.540 2716.900 ;
        RECT 1342.380 2716.640 1342.640 2716.900 ;
        RECT 455.040 2716.300 455.300 2716.560 ;
        RECT 896.180 2716.300 896.440 2716.560 ;
        RECT 1076.040 2716.300 1076.300 2716.560 ;
        RECT 1176.320 2716.300 1176.580 2716.560 ;
        RECT 1179.540 2716.300 1179.800 2716.560 ;
        RECT 1363.080 2716.300 1363.340 2716.560 ;
        RECT 288.520 2715.960 288.780 2716.220 ;
        RECT 543.360 2715.960 543.620 2716.220 ;
        RECT 574.640 2715.960 574.900 2716.220 ;
        RECT 1010.720 2715.960 1010.980 2716.220 ;
        RECT 1082.480 2715.960 1082.740 2716.220 ;
        RECT 468.380 2715.620 468.640 2715.880 ;
        RECT 916.880 2715.620 917.140 2715.880 ;
        RECT 1020.840 2715.620 1021.100 2715.880 ;
        RECT 1082.940 2715.620 1083.200 2715.880 ;
        RECT 1145.500 2715.960 1145.760 2716.220 ;
        RECT 1172.640 2715.960 1172.900 2716.220 ;
        RECT 1352.960 2715.960 1353.220 2716.220 ;
        RECT 1186.900 2715.620 1187.160 2715.880 ;
        RECT 1193.340 2715.620 1193.600 2715.880 ;
        RECT 1383.780 2715.620 1384.040 2715.880 ;
        RECT 286.220 2715.280 286.480 2715.540 ;
        RECT 398.460 2715.280 398.720 2715.540 ;
        RECT 475.280 2715.280 475.540 2715.540 ;
        RECT 937.580 2715.280 937.840 2715.540 ;
        RECT 1069.140 2715.280 1069.400 2715.540 ;
        RECT 1166.200 2715.280 1166.460 2715.540 ;
        RECT 1186.440 2715.280 1186.700 2715.540 ;
        RECT 1373.660 2715.280 1373.920 2715.540 ;
        RECT 337.740 2714.940 338.000 2715.200 ;
        RECT 491.840 2714.940 492.100 2715.200 ;
        RECT 496.440 2714.940 496.700 2715.200 ;
        RECT 968.860 2714.940 969.120 2715.200 ;
        RECT 1013.940 2714.940 1014.200 2715.200 ;
        RECT 1072.820 2714.940 1073.080 2715.200 ;
        RECT 1089.840 2714.940 1090.100 2715.200 ;
        RECT 1197.020 2714.940 1197.280 2715.200 ;
        RECT 1200.240 2714.940 1200.500 2715.200 ;
        RECT 1394.360 2714.940 1394.620 2715.200 ;
        RECT 286.680 2714.600 286.940 2714.860 ;
        RECT 501.960 2714.600 502.220 2714.860 ;
        RECT 541.520 2714.600 541.780 2714.860 ;
        RECT 720.000 2714.600 720.260 2714.860 ;
        RECT 720.920 2714.600 721.180 2714.860 ;
        RECT 1020.840 2714.600 1021.100 2714.860 ;
        RECT 1054.880 2714.600 1055.140 2714.860 ;
        RECT 1130.780 2714.600 1131.040 2714.860 ;
        RECT 1280.280 2714.600 1280.540 2714.860 ;
        RECT 527.720 2714.260 527.980 2714.520 ;
        RECT 699.300 2714.260 699.560 2714.520 ;
        RECT 700.680 2714.260 700.940 2714.520 ;
        RECT 979.440 2714.260 979.700 2714.520 ;
        RECT 1131.240 2714.260 1131.500 2714.520 ;
        RECT 1269.700 2714.260 1269.960 2714.520 ;
        RECT 513.920 2713.920 514.180 2714.180 ;
        RECT 678.600 2713.920 678.860 2714.180 ;
        RECT 686.420 2713.920 686.680 2714.180 ;
        RECT 520.820 2713.580 521.080 2713.840 ;
        RECT 688.720 2713.580 688.980 2713.840 ;
        RECT 693.320 2713.920 693.580 2714.180 ;
        RECT 958.740 2713.920 959.000 2714.180 ;
        RECT 1117.440 2713.920 1117.700 2714.180 ;
        RECT 1249.000 2713.920 1249.260 2714.180 ;
        RECT 927.460 2713.580 927.720 2713.840 ;
        RECT 1123.420 2713.580 1123.680 2713.840 ;
        RECT 1259.580 2713.580 1259.840 2713.840 ;
        RECT 500.120 2713.240 500.380 2713.500 ;
        RECT 657.440 2713.240 657.700 2713.500 ;
        RECT 658.820 2713.240 659.080 2713.500 ;
        RECT 886.060 2713.240 886.320 2713.500 ;
        RECT 1102.720 2713.240 1102.980 2713.500 ;
        RECT 1228.300 2713.240 1228.560 2713.500 ;
        RECT 507.020 2712.900 507.280 2713.160 ;
        RECT 668.020 2712.900 668.280 2713.160 ;
        RECT 687.340 2712.900 687.600 2713.160 ;
        RECT 906.760 2712.900 907.020 2713.160 ;
        RECT 1110.540 2712.900 1110.800 2713.160 ;
        RECT 1238.880 2712.900 1239.140 2713.160 ;
        RECT 542.440 2712.560 542.700 2712.820 ;
        RECT 730.120 2712.560 730.380 2712.820 ;
        RECT 534.620 2712.220 534.880 2712.480 ;
        RECT 709.420 2712.220 709.680 2712.480 ;
        RECT 761.400 2712.560 761.660 2712.820 ;
        RECT 771.980 2712.560 772.240 2712.820 ;
        RECT 748.520 2712.220 748.780 2712.480 ;
        RECT 834.080 2712.560 834.340 2712.820 ;
        RECT 1089.380 2712.560 1089.640 2712.820 ;
        RECT 1207.600 2712.560 1207.860 2712.820 ;
        RECT 1096.740 2712.220 1097.000 2712.480 ;
        RECT 1217.720 2712.220 1217.980 2712.480 ;
        RECT 686.880 2711.880 687.140 2712.140 ;
        RECT 750.820 2711.880 751.080 2712.140 ;
        RECT 802.800 2711.880 803.060 2712.140 ;
        RECT 1411.380 2691.480 1411.640 2691.740 ;
        RECT 1835.500 2691.480 1835.760 2691.740 ;
        RECT 1414.140 2691.140 1414.400 2691.400 ;
        RECT 1842.400 2691.140 1842.660 2691.400 ;
        RECT 1414.140 2684.000 1414.400 2684.260 ;
        RECT 1849.300 2684.000 1849.560 2684.260 ;
        RECT 1414.140 2677.200 1414.400 2677.460 ;
        RECT 1856.200 2677.200 1856.460 2677.460 ;
        RECT 1408.620 2670.740 1408.880 2671.000 ;
        RECT 1863.100 2670.740 1863.360 2671.000 ;
        RECT 1410.460 2670.400 1410.720 2670.660 ;
        RECT 1870.000 2670.400 1870.260 2670.660 ;
        RECT 1410.460 2663.600 1410.720 2663.860 ;
        RECT 1876.900 2663.600 1877.160 2663.860 ;
        RECT 1411.380 2656.800 1411.640 2657.060 ;
        RECT 1877.360 2656.800 1877.620 2657.060 ;
        RECT 1414.140 2656.460 1414.400 2656.720 ;
        RECT 1883.800 2656.460 1884.060 2656.720 ;
        RECT 1414.140 2649.660 1414.400 2649.920 ;
        RECT 1891.160 2649.660 1891.420 2649.920 ;
        RECT 1414.140 2642.860 1414.400 2643.120 ;
        RECT 1898.060 2642.860 1898.320 2643.120 ;
        RECT 1414.140 2636.060 1414.400 2636.320 ;
        RECT 1880.120 2636.060 1880.380 2636.320 ;
        RECT 1411.380 2635.720 1411.640 2635.980 ;
        RECT 1904.960 2635.720 1905.220 2635.980 ;
        RECT 1409.540 2628.920 1409.800 2629.180 ;
        RECT 1873.220 2628.920 1873.480 2629.180 ;
        RECT 1414.140 2622.120 1414.400 2622.380 ;
        RECT 1859.420 2622.120 1859.680 2622.380 ;
        RECT 1414.140 2615.320 1414.400 2615.580 ;
        RECT 1770.640 2615.320 1770.900 2615.580 ;
        RECT 1411.840 2614.980 1412.100 2615.240 ;
        RECT 1838.720 2614.980 1838.980 2615.240 ;
        RECT 1414.140 2608.180 1414.400 2608.440 ;
        RECT 1939.460 2608.180 1939.720 2608.440 ;
        RECT 1414.140 2601.380 1414.400 2601.640 ;
        RECT 1953.260 2601.380 1953.520 2601.640 ;
        RECT 1408.620 2595.260 1408.880 2595.520 ;
        RECT 1418.740 2595.260 1419.000 2595.520 ;
        RECT 1410.460 2587.440 1410.720 2587.700 ;
        RECT 1960.160 2587.440 1960.420 2587.700 ;
        RECT 1411.380 2580.980 1411.640 2581.240 ;
        RECT 1935.320 2580.980 1935.580 2581.240 ;
        RECT 1414.140 2580.640 1414.400 2580.900 ;
        RECT 2097.700 2580.640 2097.960 2580.900 ;
        RECT 1414.140 2573.840 1414.400 2574.100 ;
        RECT 1928.420 2573.840 1928.680 2574.100 ;
        RECT 1411.380 2566.700 1411.640 2566.960 ;
        RECT 2098.160 2566.700 2098.420 2566.960 ;
        RECT 1413.680 2560.240 1413.940 2560.500 ;
        RECT 1928.880 2560.240 1929.140 2560.500 ;
        RECT 1414.140 2559.900 1414.400 2560.160 ;
        RECT 2098.620 2559.900 2098.880 2560.160 ;
        RECT 1408.620 2553.100 1408.880 2553.360 ;
        RECT 1921.520 2553.100 1921.780 2553.360 ;
        RECT 1411.380 2546.300 1411.640 2546.560 ;
        RECT 2099.080 2546.300 2099.340 2546.560 ;
        RECT 1412.760 2539.500 1413.020 2539.760 ;
        RECT 1914.620 2539.500 1914.880 2539.760 ;
        RECT 1414.140 2539.160 1414.400 2539.420 ;
        RECT 2099.540 2539.160 2099.800 2539.420 ;
        RECT 1410.460 2532.360 1410.720 2532.620 ;
        RECT 1915.080 2532.360 1915.340 2532.620 ;
        RECT 1414.140 2525.900 1414.400 2526.160 ;
        RECT 1915.540 2525.900 1915.800 2526.160 ;
        RECT 1413.680 2525.560 1413.940 2525.820 ;
        RECT 2100.000 2525.560 2100.260 2525.820 ;
        RECT 1414.140 2518.420 1414.400 2518.680 ;
        RECT 2100.460 2518.420 2100.720 2518.680 ;
        RECT 1414.140 2511.620 1414.400 2511.880 ;
        RECT 1916.000 2511.620 1916.260 2511.880 ;
        RECT 1414.140 2505.160 1414.400 2505.420 ;
        RECT 1893.920 2505.160 1894.180 2505.420 ;
        RECT 1411.380 2504.820 1411.640 2505.080 ;
        RECT 2052.620 2504.820 2052.880 2505.080 ;
        RECT 1414.140 2490.880 1414.400 2491.140 ;
        RECT 1419.660 2490.880 1419.920 2491.140 ;
        RECT 1414.140 2484.080 1414.400 2484.340 ;
        RECT 2081.600 2484.080 2081.860 2484.340 ;
        RECT 1409.540 2477.280 1409.800 2477.540 ;
        RECT 2494.220 2477.280 2494.480 2477.540 ;
        RECT 1414.140 2470.140 1414.400 2470.400 ;
        RECT 2480.420 2470.140 2480.680 2470.400 ;
        RECT 1414.140 2463.680 1414.400 2463.940 ;
        RECT 2459.720 2463.680 2459.980 2463.940 ;
        RECT 1411.840 2463.340 1412.100 2463.600 ;
        RECT 2466.620 2463.340 2466.880 2463.600 ;
        RECT 1414.140 2456.540 1414.400 2456.800 ;
        RECT 2445.920 2456.540 2446.180 2456.800 ;
        RECT 1414.140 2449.740 1414.400 2450.000 ;
        RECT 2418.320 2449.740 2418.580 2450.000 ;
        RECT 1411.380 2449.400 1411.640 2449.660 ;
        RECT 2425.220 2449.400 2425.480 2449.660 ;
        RECT 1411.380 2442.600 1411.640 2442.860 ;
        RECT 2411.420 2442.600 2411.680 2442.860 ;
        RECT 1414.140 2435.800 1414.400 2436.060 ;
        RECT 2404.520 2435.800 2404.780 2436.060 ;
        RECT 1414.140 2429.340 1414.400 2429.600 ;
        RECT 2328.620 2429.340 2328.880 2429.600 ;
        RECT 1411.380 2429.000 1411.640 2429.260 ;
        RECT 2335.520 2429.000 2335.780 2429.260 ;
        RECT 1408.620 2421.860 1408.880 2422.120 ;
        RECT 2245.820 2421.860 2246.080 2422.120 ;
        RECT 1411.380 2415.060 1411.640 2415.320 ;
        RECT 2232.020 2415.060 2232.280 2415.320 ;
        RECT 1414.140 2408.600 1414.400 2408.860 ;
        RECT 2211.320 2408.600 2211.580 2408.860 ;
        RECT 1412.760 2408.260 1413.020 2408.520 ;
        RECT 2225.120 2408.260 2225.380 2408.520 ;
        RECT 1410.460 2401.120 1410.720 2401.380 ;
        RECT 2176.820 2401.120 2177.080 2401.380 ;
        RECT 1414.140 2394.660 1414.400 2394.920 ;
        RECT 2156.120 2394.660 2156.380 2394.920 ;
        RECT 1413.680 2394.320 1413.940 2394.580 ;
        RECT 2169.920 2394.320 2170.180 2394.580 ;
        RECT 1414.140 2387.520 1414.400 2387.780 ;
        RECT 2149.220 2387.520 2149.480 2387.780 ;
        RECT 1410.460 2380.380 1410.720 2380.640 ;
        RECT 2142.320 2380.380 2142.580 2380.640 ;
        RECT 1414.140 2373.920 1414.400 2374.180 ;
        RECT 2121.620 2373.920 2121.880 2374.180 ;
        RECT 1411.380 2373.580 1411.640 2373.840 ;
        RECT 2135.420 2373.580 2135.680 2373.840 ;
        RECT 1408.620 2366.780 1408.880 2367.040 ;
        RECT 2080.220 2366.780 2080.480 2367.040 ;
        RECT 1410.460 2359.980 1410.720 2360.240 ;
        RECT 2387.960 2359.980 2388.220 2360.240 ;
        RECT 1414.140 2353.180 1414.400 2353.440 ;
        RECT 2045.720 2353.180 2045.980 2353.440 ;
        RECT 1413.680 2352.840 1413.940 2353.100 ;
        RECT 2059.520 2352.840 2059.780 2353.100 ;
        RECT 1409.540 2346.040 1409.800 2346.300 ;
        RECT 2374.160 2346.040 2374.420 2346.300 ;
        RECT 1414.140 2339.240 1414.400 2339.500 ;
        RECT 2367.260 2339.240 2367.520 2339.500 ;
        RECT 1413.680 2332.440 1413.940 2332.700 ;
        RECT 2031.920 2332.440 2032.180 2332.700 ;
        RECT 1414.140 2332.100 1414.400 2332.360 ;
        RECT 2353.460 2332.100 2353.720 2332.360 ;
        RECT 1414.140 2325.300 1414.400 2325.560 ;
        RECT 2238.920 2325.300 2239.180 2325.560 ;
        RECT 1413.680 2318.840 1413.940 2319.100 ;
        RECT 2087.120 2318.840 2087.380 2319.100 ;
        RECT 1414.140 2318.500 1414.400 2318.760 ;
        RECT 2631.760 2318.500 2632.020 2318.760 ;
        RECT 1414.140 2311.700 1414.400 2311.960 ;
        RECT 1418.280 2311.700 1418.540 2311.960 ;
        RECT 1414.140 2304.560 1414.400 2304.820 ;
        RECT 1842.860 2304.560 1843.120 2304.820 ;
        RECT 1413.680 2298.100 1413.940 2298.360 ;
        RECT 1419.200 2298.100 1419.460 2298.360 ;
        RECT 1414.140 2297.760 1414.400 2298.020 ;
        RECT 1849.760 2297.760 1850.020 2298.020 ;
        RECT 1408.620 2290.960 1408.880 2291.220 ;
        RECT 1420.120 2290.960 1420.380 2291.220 ;
        RECT 1410.460 2283.820 1410.720 2284.080 ;
        RECT 1420.580 2283.820 1420.840 2284.080 ;
        RECT 1408.160 2277.360 1408.420 2277.620 ;
        RECT 1421.040 2277.360 1421.300 2277.620 ;
        RECT 1414.140 2277.020 1414.400 2277.280 ;
        RECT 1877.820 2277.020 1878.080 2277.280 ;
        RECT 1410.920 2201.880 1411.180 2202.140 ;
        RECT 1921.980 2201.880 1922.240 2202.140 ;
        RECT 1407.240 2201.200 1407.500 2201.460 ;
        RECT 1935.780 2201.200 1936.040 2201.460 ;
        RECT 1410.920 2194.400 1411.180 2194.660 ;
        RECT 1907.720 2194.400 1907.980 2194.660 ;
        RECT 1410.920 2182.840 1411.180 2183.100 ;
        RECT 1410.920 2180.800 1411.180 2181.060 ;
        RECT 1887.020 2180.800 1887.280 2181.060 ;
        RECT 1900.820 2180.460 1901.080 2180.720 ;
        RECT 1410.920 2173.660 1411.180 2173.920 ;
        RECT 1873.680 2173.660 1873.940 2173.920 ;
        RECT 1410.920 2166.520 1411.180 2166.780 ;
        RECT 1866.320 2166.520 1866.580 2166.780 ;
        RECT 1411.380 2157.680 1411.640 2157.940 ;
        RECT 1411.380 2153.260 1411.640 2153.520 ;
        RECT 1942.220 2153.260 1942.480 2153.520 ;
        RECT 1411.380 2152.580 1411.640 2152.840 ;
        RECT 2321.720 2152.580 2321.980 2152.840 ;
        RECT 1407.240 2145.780 1407.500 2146.040 ;
        RECT 2083.900 2145.780 2084.160 2146.040 ;
        RECT 1411.380 2145.440 1411.640 2145.700 ;
        RECT 1790.880 2145.440 1791.140 2145.700 ;
        RECT 1411.380 2138.640 1411.640 2138.900 ;
        RECT 1790.420 2138.640 1790.680 2138.900 ;
        RECT 1783.980 2138.300 1784.240 2138.560 ;
        RECT 1411.380 2135.920 1411.640 2136.180 ;
        RECT 1411.380 2131.840 1411.640 2132.100 ;
        RECT 1783.520 2131.840 1783.780 2132.100 ;
        RECT 1411.380 2125.040 1411.640 2125.300 ;
        RECT 1777.080 2125.040 1777.340 2125.300 ;
        RECT 1411.380 2117.900 1411.640 2118.160 ;
        RECT 1776.620 2117.900 1776.880 2118.160 ;
        RECT 1770.180 2117.560 1770.440 2117.820 ;
        RECT 1411.380 2116.200 1411.640 2116.460 ;
        RECT 1411.380 2111.100 1411.640 2111.360 ;
        RECT 1769.720 2111.100 1769.980 2111.360 ;
        RECT 1408.160 2106.680 1408.420 2106.940 ;
        RECT 1408.160 2106.000 1408.420 2106.260 ;
        RECT 1412.300 2106.000 1412.560 2106.260 ;
        RECT 1412.300 2104.980 1412.560 2105.240 ;
        RECT 1414.140 2104.980 1414.400 2105.240 ;
        RECT 1414.140 2104.300 1414.400 2104.560 ;
        RECT 1763.280 2104.300 1763.540 2104.560 ;
        RECT 1412.760 2097.160 1413.020 2097.420 ;
        RECT 2380.600 2097.160 2380.860 2097.420 ;
        RECT 1414.140 2096.820 1414.400 2097.080 ;
        RECT 1762.820 2096.820 1763.080 2097.080 ;
        RECT 1414.140 2090.360 1414.400 2090.620 ;
        RECT 2373.700 2090.360 2373.960 2090.620 ;
        RECT 1411.380 2088.660 1411.640 2088.920 ;
        RECT 1412.760 2088.660 1413.020 2088.920 ;
        RECT 1411.380 2087.980 1411.640 2088.240 ;
        RECT 1414.140 2083.560 1414.400 2083.820 ;
        RECT 2366.800 2083.560 2367.060 2083.820 ;
        RECT 1422.880 2081.860 1423.140 2082.120 ;
        RECT 2266.520 2081.860 2266.780 2082.120 ;
        RECT 1431.160 2081.520 1431.420 2081.780 ;
        RECT 2277.100 2081.520 2277.360 2081.780 ;
        RECT 1430.700 2081.180 1430.960 2081.440 ;
        RECT 2284.000 2081.180 2284.260 2081.440 ;
        RECT 1416.440 2080.840 1416.700 2081.100 ;
        RECT 2290.900 2080.840 2291.160 2081.100 ;
        RECT 1415.980 2080.500 1416.240 2080.760 ;
        RECT 2297.800 2080.500 2298.060 2080.760 ;
        RECT 1415.520 2080.160 1415.780 2080.420 ;
        RECT 2305.160 2080.160 2305.420 2080.420 ;
        RECT 1411.380 2077.100 1411.640 2077.360 ;
        RECT 1414.600 2077.100 1414.860 2077.360 ;
        RECT 1414.140 2076.760 1414.400 2077.020 ;
        RECT 2359.900 2076.760 2360.160 2077.020 ;
        RECT 1411.380 2076.420 1411.640 2076.680 ;
        RECT 2353.000 2076.420 2353.260 2076.680 ;
        RECT 1427.020 2076.080 1427.280 2076.340 ;
        RECT 2192.920 2076.080 2193.180 2076.340 ;
        RECT 1426.560 2075.740 1426.820 2076.000 ;
        RECT 2193.380 2075.740 2193.640 2076.000 ;
        RECT 1423.800 2075.400 1424.060 2075.660 ;
        RECT 2190.620 2075.400 2190.880 2075.660 ;
        RECT 1424.260 2075.060 1424.520 2075.320 ;
        RECT 2191.540 2075.060 2191.800 2075.320 ;
        RECT 1423.340 2074.720 1423.600 2074.980 ;
        RECT 2191.080 2074.720 2191.340 2074.980 ;
        RECT 1426.100 2074.380 1426.360 2074.640 ;
        RECT 2228.800 2074.380 2229.060 2074.640 ;
        RECT 1460.140 2074.040 1460.400 2074.300 ;
        RECT 2263.760 2074.040 2264.020 2074.300 ;
        RECT 1415.060 2073.700 1415.320 2073.960 ;
        RECT 2339.660 2073.700 2339.920 2073.960 ;
        RECT 1414.600 2073.360 1414.860 2073.620 ;
        RECT 2346.100 2073.360 2346.360 2073.620 ;
        RECT 1427.480 2073.020 1427.740 2073.280 ;
        RECT 2192.460 2073.020 2192.720 2073.280 ;
        RECT 1427.940 2072.680 1428.200 2072.940 ;
        RECT 2192.000 2072.680 2192.260 2072.940 ;
        RECT 1686.920 2072.340 1687.180 2072.600 ;
        RECT 2270.200 2072.340 2270.460 2072.600 ;
        RECT 1421.960 2072.000 1422.220 2072.260 ;
        RECT 1718.660 2072.000 1718.920 2072.260 ;
        RECT 1422.420 2071.660 1422.680 2071.920 ;
        RECT 1711.300 2071.660 1711.560 2071.920 ;
        RECT 1915.540 2069.960 1915.800 2070.220 ;
        RECT 1410.920 2069.620 1411.180 2069.880 ;
        RECT 2014.900 2069.620 2015.160 2069.880 ;
        RECT 2238.920 2069.620 2239.180 2069.880 ;
        RECT 2347.020 2069.620 2347.280 2069.880 ;
        RECT 2480.420 2069.620 2480.680 2069.880 ;
        RECT 2525.500 2069.620 2525.760 2069.880 ;
        RECT 1411.380 2069.280 1411.640 2069.540 ;
        RECT 1417.360 2069.280 1417.620 2069.540 ;
        RECT 1980.400 2069.280 1980.660 2069.540 ;
        RECT 2045.720 2069.280 2045.980 2069.540 ;
        RECT 2380.600 2069.280 2380.860 2069.540 ;
        RECT 2445.920 2069.280 2446.180 2069.540 ;
        RECT 2512.620 2069.280 2512.880 2069.540 ;
        RECT 1408.620 2068.940 1408.880 2069.200 ;
        RECT 1935.780 2068.940 1936.040 2069.200 ;
        RECT 1959.700 2068.940 1959.960 2069.200 ;
        RECT 2059.520 2068.940 2059.780 2069.200 ;
        RECT 2387.500 2068.940 2387.760 2069.200 ;
        RECT 2418.320 2068.940 2418.580 2069.200 ;
        RECT 2497.900 2068.940 2498.160 2069.200 ;
        RECT 1409.540 2068.600 1409.800 2068.860 ;
        RECT 1946.360 2068.600 1946.620 2068.860 ;
        RECT 2031.920 2068.600 2032.180 2068.860 ;
        RECT 2359.900 2068.600 2360.160 2068.860 ;
        RECT 2459.720 2068.600 2459.980 2068.860 ;
        RECT 2518.600 2068.600 2518.860 2068.860 ;
        RECT 1410.000 2068.260 1410.260 2068.520 ;
        RECT 1945.900 2068.260 1946.160 2068.520 ;
        RECT 2080.220 2068.260 2080.480 2068.520 ;
        RECT 2394.400 2068.260 2394.660 2068.520 ;
        RECT 2411.420 2068.260 2411.680 2068.520 ;
        RECT 2491.460 2068.260 2491.720 2068.520 ;
        RECT 2494.220 2068.260 2494.480 2068.520 ;
        RECT 2532.400 2068.260 2532.660 2068.520 ;
        RECT 1409.080 2067.920 1409.340 2068.180 ;
        RECT 1410.460 2067.580 1410.720 2067.840 ;
        RECT 1932.100 2067.920 1932.360 2068.180 ;
        RECT 1942.680 2067.920 1942.940 2068.180 ;
        RECT 2021.800 2067.920 2022.060 2068.180 ;
        RECT 2121.620 2067.920 2121.880 2068.180 ;
        RECT 2402.220 2067.920 2402.480 2068.180 ;
        RECT 2404.520 2067.920 2404.780 2068.180 ;
        RECT 2484.100 2067.920 2484.360 2068.180 ;
        RECT 1907.720 2067.580 1907.980 2067.840 ;
        RECT 1973.500 2067.580 1973.760 2067.840 ;
        RECT 2156.120 2067.580 2156.380 2067.840 ;
        RECT 2428.900 2067.580 2429.160 2067.840 ;
        RECT 1413.680 2067.240 1413.940 2067.500 ;
        RECT 1880.120 2067.240 1880.380 2067.500 ;
        RECT 1911.400 2067.240 1911.660 2067.500 ;
        RECT 1916.000 2067.240 1916.260 2067.500 ;
        RECT 2008.000 2067.240 2008.260 2067.500 ;
        RECT 2142.320 2067.240 2142.580 2067.500 ;
        RECT 2415.100 2067.240 2415.360 2067.500 ;
        RECT 2466.620 2067.240 2466.880 2067.500 ;
        RECT 2519.980 2067.240 2520.240 2067.500 ;
        RECT 1413.220 2066.900 1413.480 2067.160 ;
        RECT 1987.300 2066.900 1987.560 2067.160 ;
        RECT 2135.420 2066.900 2135.680 2067.160 ;
        RECT 2408.200 2066.900 2408.460 2067.160 ;
        RECT 2425.220 2066.900 2425.480 2067.160 ;
        RECT 2505.260 2066.900 2505.520 2067.160 ;
        RECT 1411.840 2066.560 1412.100 2066.820 ;
        RECT 1910.940 2066.560 1911.200 2066.820 ;
        RECT 1987.760 2066.560 1988.020 2066.820 ;
        RECT 2149.220 2066.560 2149.480 2066.820 ;
        RECT 2422.000 2066.560 2422.260 2066.820 ;
        RECT 1412.300 2066.220 1412.560 2066.480 ;
        RECT 1911.860 2066.220 1912.120 2066.480 ;
        RECT 1915.080 2066.220 1915.340 2066.480 ;
        RECT 1994.200 2066.220 1994.460 2066.480 ;
        RECT 2176.820 2066.220 2177.080 2066.480 ;
        RECT 2442.700 2066.220 2442.960 2066.480 ;
        RECT 1412.760 2065.880 1413.020 2066.140 ;
        RECT 1893.920 2065.880 1894.180 2066.140 ;
        RECT 1921.520 2065.880 1921.780 2066.140 ;
        RECT 1921.980 2065.880 1922.240 2066.140 ;
        RECT 1966.600 2065.880 1966.860 2066.140 ;
        RECT 2169.920 2065.880 2170.180 2066.140 ;
        RECT 2435.800 2065.880 2436.060 2066.140 ;
        RECT 1413.680 2065.540 1413.940 2065.800 ;
        RECT 1408.160 2065.200 1408.420 2065.460 ;
        RECT 1890.700 2065.200 1890.960 2065.460 ;
        RECT 1918.300 2065.540 1918.560 2065.800 ;
        RECT 1952.800 2065.540 1953.060 2065.800 ;
        RECT 2087.120 2065.540 2087.380 2065.800 ;
        RECT 2340.580 2065.540 2340.840 2065.800 ;
        RECT 1898.060 2065.200 1898.320 2065.460 ;
        RECT 1900.820 2065.200 1901.080 2065.460 ;
        RECT 1928.880 2065.200 1929.140 2065.460 ;
        RECT 1980.400 2065.200 1980.660 2065.460 ;
        RECT 2211.320 2065.200 2211.580 2065.460 ;
        RECT 2449.600 2065.200 2449.860 2065.460 ;
        RECT 1411.380 2064.860 1411.640 2065.120 ;
        RECT 1435.300 2064.860 1435.560 2065.120 ;
        RECT 1483.140 2064.860 1483.400 2065.120 ;
        RECT 1531.900 2064.860 1532.160 2065.120 ;
        RECT 1579.740 2064.860 1580.000 2065.120 ;
        RECT 1655.640 2064.860 1655.900 2065.120 ;
        RECT 1676.340 2064.860 1676.600 2065.120 ;
        RECT 1752.240 2064.860 1752.500 2065.120 ;
        RECT 1772.940 2064.860 1773.200 2065.120 ;
        RECT 1821.700 2064.860 1821.960 2065.120 ;
        RECT 1883.800 2064.860 1884.060 2065.120 ;
        RECT 1904.500 2064.860 1904.760 2065.120 ;
        RECT 1939.000 2064.860 1939.260 2065.120 ;
        RECT 1987.300 2064.860 1987.560 2065.120 ;
        RECT 2225.120 2064.860 2225.380 2065.120 ;
        RECT 2456.500 2064.860 2456.760 2065.120 ;
        RECT 1420.580 2064.520 1420.840 2064.780 ;
        RECT 1870.000 2064.520 1870.260 2064.780 ;
        RECT 1421.040 2064.180 1421.300 2064.440 ;
        RECT 1870.920 2064.180 1871.180 2064.440 ;
        RECT 1873.220 2064.180 1873.480 2064.440 ;
        RECT 1911.400 2064.180 1911.660 2064.440 ;
        RECT 1914.620 2064.520 1914.880 2064.780 ;
        RECT 1921.520 2064.520 1921.780 2064.780 ;
        RECT 2015.820 2064.520 2016.080 2064.780 ;
        RECT 2232.020 2064.520 2232.280 2064.780 ;
        RECT 2456.960 2064.520 2457.220 2064.780 ;
        RECT 1925.200 2064.180 1925.460 2064.440 ;
        RECT 1928.420 2064.180 1928.680 2064.440 ;
        RECT 1973.500 2064.180 1973.760 2064.440 ;
        RECT 2245.820 2064.180 2246.080 2064.440 ;
        RECT 2463.400 2064.180 2463.660 2064.440 ;
        RECT 1420.120 2063.840 1420.380 2064.100 ;
        RECT 1863.100 2063.840 1863.360 2064.100 ;
        RECT 1866.320 2063.840 1866.580 2064.100 ;
        RECT 2001.100 2063.840 2001.360 2064.100 ;
        RECT 2052.620 2063.840 2052.880 2064.100 ;
        RECT 2587.600 2063.840 2587.860 2064.100 ;
        RECT 1419.200 2063.500 1419.460 2063.760 ;
        RECT 1856.200 2063.500 1856.460 2063.760 ;
        RECT 1856.660 2063.500 1856.920 2063.760 ;
        RECT 1873.680 2063.500 1873.940 2063.760 ;
        RECT 1887.020 2063.500 1887.280 2063.760 ;
        RECT 1994.200 2063.500 1994.460 2063.760 ;
        RECT 2335.520 2063.500 2335.780 2063.760 ;
        RECT 2478.580 2063.500 2478.840 2063.760 ;
        RECT 1418.280 2063.160 1418.540 2063.420 ;
        RECT 1835.500 2063.160 1835.760 2063.420 ;
        RECT 1838.720 2063.160 1838.980 2063.420 ;
        RECT 1925.200 2063.160 1925.460 2063.420 ;
        RECT 1419.660 2062.820 1419.920 2063.080 ;
        RECT 1760.520 2062.820 1760.780 2063.080 ;
        RECT 2001.100 2063.160 2001.360 2063.420 ;
        RECT 2328.620 2063.160 2328.880 2063.420 ;
        RECT 2470.300 2063.160 2470.560 2063.420 ;
        RECT 1418.740 2062.480 1419.000 2062.740 ;
        RECT 1760.060 2062.480 1760.320 2062.740 ;
        RECT 1419.200 2062.140 1419.460 2062.400 ;
        RECT 1766.500 2062.140 1766.760 2062.400 ;
        RECT 1420.120 2061.800 1420.380 2062.060 ;
        RECT 1773.400 2061.800 1773.660 2062.060 ;
        RECT 1420.580 2061.460 1420.840 2061.720 ;
        RECT 1780.760 2061.460 1781.020 2061.720 ;
        RECT 1417.360 2061.120 1417.620 2061.380 ;
        RECT 1787.660 2061.120 1787.920 2061.380 ;
        RECT 1421.040 2060.780 1421.300 2061.040 ;
        RECT 1794.560 2060.780 1794.820 2061.040 ;
        RECT 1715.440 2060.440 1715.700 2060.700 ;
        RECT 2339.200 2060.440 2339.460 2060.700 ;
        RECT 1690.140 2060.100 1690.400 2060.360 ;
        RECT 2318.500 2060.100 2318.760 2060.360 ;
        RECT 1416.900 2059.760 1417.160 2060.020 ;
        RECT 2263.300 2059.760 2263.560 2060.020 ;
        RECT 1462.900 2059.420 1463.160 2059.680 ;
        RECT 2325.400 2059.420 2325.660 2059.680 ;
        RECT 1418.280 2059.080 1418.540 2059.340 ;
        RECT 1753.160 2059.080 1753.420 2059.340 ;
        RECT 1417.820 2058.740 1418.080 2059.000 ;
        RECT 1745.800 2058.740 1746.060 2059.000 ;
        RECT 1434.840 2058.400 1435.100 2058.660 ;
        RECT 1738.900 2058.400 1739.160 2058.660 ;
        RECT 1434.380 2058.060 1434.640 2058.320 ;
        RECT 1732.000 2058.060 1732.260 2058.320 ;
        RECT 1433.460 2057.720 1433.720 2057.980 ;
        RECT 1725.100 2057.720 1725.360 2057.980 ;
        RECT 1433.920 2057.380 1434.180 2057.640 ;
        RECT 1718.200 2057.380 1718.460 2057.640 ;
        RECT 1693.820 2056.360 1694.080 2056.620 ;
        RECT 2028.700 2056.360 2028.960 2056.620 ;
        RECT 1413.680 2056.020 1413.940 2056.280 ;
        RECT 2332.300 2056.020 2332.560 2056.280 ;
        RECT 1414.140 2055.680 1414.400 2055.940 ;
        RECT 1715.440 2055.680 1715.700 2055.940 ;
        RECT 1408.160 2055.340 1408.420 2055.600 ;
        RECT 2193.840 2055.340 2194.100 2055.600 ;
        RECT 1410.000 2055.000 1410.260 2055.260 ;
        RECT 2256.400 2055.000 2256.660 2055.260 ;
        RECT 1410.920 2054.660 1411.180 2054.920 ;
        RECT 2280.320 2054.660 2280.580 2054.920 ;
        RECT 1411.380 2054.320 1411.640 2054.580 ;
        RECT 2287.220 2054.320 2287.480 2054.580 ;
        RECT 1413.220 2053.980 1413.480 2054.240 ;
        RECT 2294.120 2053.980 2294.380 2054.240 ;
        RECT 1412.760 2053.640 1413.020 2053.900 ;
        RECT 2301.020 2053.640 2301.280 2053.900 ;
        RECT 1412.300 2053.300 1412.560 2053.560 ;
        RECT 2301.940 2053.300 2302.200 2053.560 ;
        RECT 1411.840 2052.960 1412.100 2053.220 ;
        RECT 2304.700 2052.960 2304.960 2053.220 ;
        RECT 1414.140 2052.620 1414.400 2052.880 ;
        RECT 2311.600 2052.620 2311.860 2052.880 ;
        RECT 1421.500 2052.280 1421.760 2052.540 ;
        RECT 1704.400 2052.280 1704.660 2052.540 ;
        RECT 1408.620 2048.880 1408.880 2049.140 ;
        RECT 1462.900 2048.880 1463.160 2049.140 ;
        RECT 1408.620 2042.080 1408.880 2042.340 ;
        RECT 1690.140 2042.080 1690.400 2042.340 ;
        RECT 1408.160 2019.980 1408.420 2020.240 ;
        RECT 1416.440 2019.980 1416.700 2020.240 ;
        RECT 1414.140 2011.140 1414.400 2011.400 ;
        RECT 1430.700 2011.140 1430.960 2011.400 ;
        RECT 1414.140 2005.700 1414.400 2005.960 ;
        RECT 1431.160 2005.700 1431.420 2005.960 ;
        RECT 1414.140 2000.600 1414.400 2000.860 ;
        RECT 1686.920 2000.600 1687.180 2000.860 ;
        RECT 1411.380 2000.260 1411.640 2000.520 ;
        RECT 1460.140 2000.260 1460.400 2000.520 ;
        RECT 1408.160 1990.740 1408.420 1991.000 ;
        RECT 1416.900 1990.740 1417.160 1991.000 ;
        RECT 1408.160 1985.980 1408.420 1986.240 ;
        RECT 1421.040 1985.980 1421.300 1986.240 ;
        RECT 1408.160 1982.240 1408.420 1982.500 ;
        RECT 1417.360 1982.240 1417.620 1982.500 ;
        RECT 1410.920 1979.860 1411.180 1980.120 ;
        RECT 1408.160 1978.840 1408.420 1979.100 ;
        RECT 1420.580 1978.840 1420.840 1979.100 ;
        RECT 1408.160 1971.700 1408.420 1971.960 ;
        RECT 1420.120 1971.700 1420.380 1971.960 ;
        RECT 1408.160 1965.920 1408.420 1966.180 ;
        RECT 1419.200 1965.920 1419.460 1966.180 ;
        RECT 1408.160 1960.140 1408.420 1960.400 ;
        RECT 1419.660 1960.140 1419.920 1960.400 ;
        RECT 1408.160 1958.100 1408.420 1958.360 ;
        RECT 1418.740 1958.100 1419.000 1958.360 ;
        RECT 1408.160 1950.620 1408.420 1950.880 ;
        RECT 1418.280 1950.620 1418.540 1950.880 ;
        RECT 1408.160 1945.180 1408.420 1945.440 ;
        RECT 1417.820 1945.180 1418.080 1945.440 ;
        RECT 1408.160 1941.440 1408.420 1941.700 ;
        RECT 1434.840 1941.440 1435.100 1941.700 ;
        RECT 1408.160 1935.320 1408.420 1935.580 ;
        RECT 1434.380 1935.320 1434.640 1935.580 ;
        RECT 1411.380 1931.920 1411.640 1932.180 ;
        RECT 1408.160 1930.220 1408.420 1930.480 ;
        RECT 1433.460 1930.220 1433.720 1930.480 ;
        RECT 1408.160 1926.140 1408.420 1926.400 ;
        RECT 1433.920 1926.140 1434.180 1926.400 ;
        RECT 1408.160 1920.020 1408.420 1920.280 ;
        RECT 1421.960 1920.020 1422.220 1920.280 ;
        RECT 1408.160 1916.280 1408.420 1916.540 ;
        RECT 1422.420 1916.280 1422.680 1916.540 ;
        RECT 1409.080 1910.840 1409.340 1911.100 ;
        RECT 1697.500 1910.840 1697.760 1911.100 ;
        RECT 1408.160 1910.500 1408.420 1910.760 ;
        RECT 1421.500 1910.500 1421.760 1910.760 ;
        RECT 1408.160 1904.040 1408.420 1904.300 ;
        RECT 1690.600 1904.040 1690.860 1904.300 ;
        RECT 1408.160 1897.240 1408.420 1897.500 ;
        RECT 1684.160 1897.240 1684.420 1897.500 ;
        RECT 1408.160 1890.440 1408.420 1890.700 ;
        RECT 1683.700 1890.440 1683.960 1890.700 ;
        RECT 1409.080 1890.100 1409.340 1890.360 ;
        RECT 1676.800 1890.100 1677.060 1890.360 ;
        RECT 1408.160 1883.300 1408.420 1883.560 ;
        RECT 1669.900 1883.300 1670.160 1883.560 ;
        RECT 1408.160 1876.500 1408.420 1876.760 ;
        RECT 1663.000 1876.500 1663.260 1876.760 ;
        RECT 1409.080 1869.700 1409.340 1869.960 ;
        RECT 1649.660 1869.700 1649.920 1869.960 ;
        RECT 1408.160 1865.620 1408.420 1865.880 ;
        RECT 1438.980 1865.620 1439.240 1865.880 ;
        RECT 1408.160 1859.500 1408.420 1859.760 ;
        RECT 1433.000 1859.500 1433.260 1859.760 ;
        RECT 1409.080 1855.760 1409.340 1856.020 ;
        RECT 1635.400 1855.760 1635.660 1856.020 ;
        RECT 1408.160 1854.740 1408.420 1855.000 ;
        RECT 1425.640 1854.740 1425.900 1855.000 ;
        RECT 1411.380 1849.300 1411.640 1849.560 ;
        RECT 1408.160 1848.960 1408.420 1849.220 ;
        RECT 1628.500 1848.960 1628.760 1849.220 ;
        RECT 1408.160 1842.160 1408.420 1842.420 ;
        RECT 1576.520 1842.160 1576.780 1842.420 ;
        RECT 1410.920 1835.700 1411.180 1835.960 ;
        RECT 1410.460 1835.020 1410.720 1835.280 ;
        RECT 1422.420 1835.020 1422.680 1835.280 ;
        RECT 1562.720 1835.020 1562.980 1835.280 ;
        RECT 1425.640 1834.680 1425.900 1834.940 ;
        RECT 1548.920 1834.680 1549.180 1834.940 ;
        RECT 1408.160 1828.220 1408.420 1828.480 ;
        RECT 1652.420 1828.220 1652.680 1828.480 ;
        RECT 1411.380 1824.820 1411.640 1825.080 ;
        RECT 1413.680 1824.820 1413.940 1825.080 ;
        RECT 1408.160 1821.420 1408.420 1821.680 ;
        RECT 1646.440 1821.420 1646.700 1821.680 ;
        RECT 1408.160 1814.280 1408.420 1814.540 ;
        RECT 1645.520 1814.280 1645.780 1814.540 ;
        RECT 1409.080 1813.940 1409.340 1814.200 ;
        RECT 1638.620 1813.940 1638.880 1814.200 ;
        RECT 1408.160 1807.480 1408.420 1807.740 ;
        RECT 1631.720 1807.480 1631.980 1807.740 ;
        RECT 1408.160 1800.680 1408.420 1800.940 ;
        RECT 1624.820 1800.680 1625.080 1800.940 ;
        RECT 1409.080 1800.340 1409.340 1800.600 ;
        RECT 1617.920 1800.340 1618.180 1800.600 ;
        RECT 1408.160 1793.540 1408.420 1793.800 ;
        RECT 1611.020 1793.540 1611.280 1793.800 ;
        RECT 1410.920 1787.080 1411.180 1787.340 ;
        RECT 1408.160 1758.860 1408.420 1759.120 ;
        RECT 1432.540 1758.860 1432.800 1759.120 ;
        RECT 1408.160 1754.440 1408.420 1754.700 ;
        RECT 1432.080 1754.440 1432.340 1754.700 ;
        RECT 1408.160 1751.380 1408.420 1751.640 ;
        RECT 1422.880 1751.380 1423.140 1751.640 ;
        RECT 1408.160 1745.260 1408.420 1745.520 ;
        RECT 1459.220 1745.260 1459.480 1745.520 ;
        RECT 1408.160 1738.460 1408.420 1738.720 ;
        RECT 1452.320 1738.460 1452.580 1738.720 ;
        RECT 1408.160 1733.700 1408.420 1733.960 ;
        RECT 1438.520 1733.700 1438.780 1733.960 ;
        RECT 1408.160 1728.260 1408.420 1728.520 ;
        RECT 1431.620 1728.260 1431.880 1728.520 ;
        RECT 1408.160 1724.180 1408.420 1724.440 ;
        RECT 1424.720 1724.180 1424.980 1724.440 ;
        RECT 1408.160 1717.720 1408.420 1717.980 ;
        RECT 1535.120 1717.720 1535.380 1717.980 ;
        RECT 1409.080 1717.380 1409.340 1717.640 ;
        RECT 1459.680 1717.380 1459.940 1717.640 ;
        RECT 1408.160 1710.920 1408.420 1711.180 ;
        RECT 1542.020 1710.920 1542.280 1711.180 ;
        RECT 1411.380 1704.120 1411.640 1704.380 ;
        RECT 1412.300 1704.120 1412.560 1704.380 ;
        RECT 1408.160 1703.780 1408.420 1704.040 ;
        RECT 1423.800 1703.780 1424.060 1704.040 ;
        RECT 1408.620 1703.100 1408.880 1703.360 ;
        RECT 1423.340 1703.100 1423.600 1703.360 ;
        RECT 1408.160 1693.920 1408.420 1694.180 ;
        RECT 1424.260 1693.920 1424.520 1694.180 ;
        RECT 1412.300 1690.180 1412.560 1690.440 ;
        RECT 1408.160 1689.500 1408.420 1689.760 ;
        RECT 1427.940 1689.500 1428.200 1689.760 ;
        RECT 1408.620 1683.380 1408.880 1683.640 ;
        RECT 1427.020 1683.380 1427.280 1683.640 ;
        RECT 1408.160 1682.700 1408.420 1682.960 ;
        RECT 1427.480 1682.700 1427.740 1682.960 ;
        RECT 1408.160 1672.840 1408.420 1673.100 ;
        RECT 1426.560 1672.840 1426.820 1673.100 ;
        RECT 1408.620 1669.440 1408.880 1669.700 ;
        RECT 1514.420 1669.440 1514.680 1669.700 ;
        RECT 1408.160 1668.080 1408.420 1668.340 ;
        RECT 1426.100 1668.080 1426.360 1668.340 ;
        RECT 1408.160 1655.840 1408.420 1656.100 ;
        RECT 1601.360 1655.840 1601.620 1656.100 ;
        RECT 1407.700 1648.700 1407.960 1648.960 ;
        RECT 1600.900 1648.700 1601.160 1648.960 ;
        RECT 1408.160 1648.360 1408.420 1648.620 ;
        RECT 1594.000 1648.360 1594.260 1648.620 ;
        RECT 1411.840 1642.240 1412.100 1642.500 ;
        RECT 1407.700 1641.900 1407.960 1642.160 ;
        RECT 1587.100 1641.900 1587.360 1642.160 ;
        RECT 1407.700 1627.620 1407.960 1627.880 ;
        RECT 1425.180 1627.620 1425.440 1627.880 ;
        RECT 1414.140 1607.560 1414.400 1607.820 ;
        RECT 1693.820 1607.560 1694.080 1607.820 ;
      LAYER met2 ;
        RECT 1318.000 3266.730 1318.260 3267.050 ;
        RECT 1890.700 3266.730 1890.960 3267.050 ;
        RECT 1917.840 3266.730 1918.100 3267.050 ;
        RECT 2542.060 3266.730 2542.320 3267.050 ;
        RECT 697.000 3264.010 697.260 3264.330 ;
        RECT 675.840 3263.900 676.100 3263.990 ;
        RECT 675.440 3263.760 676.100 3263.900 ;
        RECT 675.440 3255.685 675.580 3263.760 ;
        RECT 675.840 3263.670 676.100 3263.760 ;
        RECT 675.370 3255.315 675.650 3255.685 ;
        RECT 289.430 3230.155 289.710 3230.525 ;
        RECT 288.970 3224.715 289.250 3225.085 ;
        RECT 288.510 3215.875 288.790 3216.245 ;
        RECT 288.050 3209.755 288.330 3210.125 ;
        RECT 287.590 3201.595 287.870 3201.965 ;
        RECT 287.130 3196.155 287.410 3196.525 ;
        RECT 286.670 3187.995 286.950 3188.365 ;
        RECT 286.210 2898.315 286.490 2898.685 ;
        RECT 286.280 2715.570 286.420 2898.315 ;
        RECT 286.220 2715.250 286.480 2715.570 ;
        RECT 286.740 2714.890 286.880 3187.995 ;
        RECT 287.200 2717.610 287.340 3196.155 ;
        RECT 287.140 2717.290 287.400 2717.610 ;
        RECT 287.660 2717.270 287.800 3201.595 ;
        RECT 287.600 2716.950 287.860 2717.270 ;
        RECT 288.120 2716.930 288.260 3209.755 ;
        RECT 288.060 2716.610 288.320 2716.930 ;
        RECT 288.580 2716.250 288.720 3215.875 ;
        RECT 289.040 2719.310 289.180 3224.715 ;
        RECT 289.500 2719.650 289.640 3230.155 ;
      LAYER met2 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met2 ;
        RECT 688.260 3251.090 688.520 3251.410 ;
        RECT 688.320 3248.600 688.460 3251.090 ;
        RECT 688.250 3248.230 688.530 3248.600 ;
        RECT 697.060 2948.325 697.200 3264.010 ;
        RECT 1292.700 3263.670 1292.960 3263.990 ;
        RECT 1292.760 3258.405 1292.900 3263.670 ;
        RECT 1318.060 3258.405 1318.200 3266.730 ;
        RECT 1890.760 3264.670 1890.900 3266.730 ;
        RECT 1917.900 3264.670 1918.040 3266.730 ;
        RECT 1890.700 3264.525 1890.960 3264.670 ;
        RECT 1917.840 3264.525 1918.100 3264.670 ;
        RECT 2542.120 3264.525 2542.260 3266.730 ;
        RECT 1890.690 3264.155 1890.970 3264.525 ;
        RECT 1917.830 3264.155 1918.110 3264.525 ;
        RECT 2542.050 3264.155 2542.330 3264.525 ;
        RECT 2566.890 3264.155 2567.170 3264.525 ;
        RECT 1917.900 3264.025 1918.040 3264.155 ;
        RECT 2542.060 3264.010 2542.320 3264.155 ;
        RECT 2566.900 3264.010 2567.160 3264.155 ;
        RECT 2542.120 3263.855 2542.260 3264.010 ;
        RECT 2594.500 3263.670 2594.760 3263.990 ;
        RECT 1292.690 3258.035 1292.970 3258.405 ;
        RECT 1317.990 3258.035 1318.270 3258.405 ;
        RECT 2038.820 3252.450 2039.080 3252.770 ;
        RECT 1333.180 3252.110 1333.440 3252.430 ;
        RECT 1935.780 3252.110 1936.040 3252.430 ;
        RECT 941.710 3230.155 941.990 3230.525 ;
        RECT 696.990 2947.955 697.270 2948.325 ;
        RECT 337.730 2794.275 338.010 2794.645 ;
        RECT 344.630 2794.275 344.910 2794.645 ;
        RECT 351.530 2794.275 351.810 2794.645 ;
        RECT 358.430 2794.275 358.710 2794.645 ;
        RECT 362.570 2794.275 362.850 2794.645 ;
        RECT 365.330 2794.275 365.610 2794.645 ;
        RECT 368.550 2794.275 368.830 2794.645 ;
        RECT 371.310 2794.275 371.590 2794.645 ;
        RECT 374.990 2794.275 375.270 2794.645 ;
        RECT 379.130 2794.275 379.410 2794.645 ;
        RECT 384.190 2794.275 384.470 2794.645 ;
        RECT 386.950 2794.275 387.230 2794.645 ;
        RECT 392.930 2794.275 393.210 2794.645 ;
        RECT 396.610 2794.275 396.890 2794.645 ;
        RECT 399.370 2794.275 399.650 2794.645 ;
        RECT 403.970 2794.275 404.250 2794.645 ;
        RECT 406.270 2794.275 406.550 2794.645 ;
        RECT 409.950 2794.275 410.230 2794.645 ;
        RECT 414.550 2794.275 414.830 2794.645 ;
        RECT 419.150 2794.275 419.430 2794.645 ;
        RECT 420.990 2794.275 421.270 2794.645 ;
        RECT 427.430 2794.275 427.710 2794.645 ;
        RECT 431.570 2794.275 431.850 2794.645 ;
        RECT 330.840 2793.790 331.100 2794.110 ;
        RECT 310.130 2791.555 310.410 2791.925 ;
        RECT 289.440 2719.330 289.700 2719.650 ;
        RECT 288.980 2718.990 289.240 2719.310 ;
        RECT 310.200 2717.950 310.340 2791.555 ;
        RECT 317.030 2790.875 317.310 2791.245 ;
        RECT 305.080 2717.630 305.340 2717.950 ;
        RECT 310.140 2717.630 310.400 2717.950 ;
        RECT 288.520 2715.930 288.780 2716.250 ;
        RECT 286.680 2714.570 286.940 2714.890 ;
        RECT 305.140 2700.000 305.280 2717.630 ;
        RECT 317.100 2700.010 317.240 2790.875 ;
        RECT 330.900 2717.950 331.040 2793.790 ;
        RECT 337.280 2787.670 337.540 2787.990 ;
        RECT 325.780 2717.630 326.040 2717.950 ;
        RECT 330.840 2717.630 331.100 2717.950 ;
        RECT 315.330 2700.000 317.240 2700.010 ;
        RECT 305.140 2699.940 305.430 2700.000 ;
        RECT 305.150 2696.000 305.430 2699.940 ;
        RECT 315.270 2699.870 317.240 2700.000 ;
        RECT 325.840 2700.000 325.980 2717.630 ;
        RECT 337.340 2700.010 337.480 2787.670 ;
        RECT 337.800 2715.230 337.940 2794.275 ;
        RECT 337.740 2714.910 338.000 2715.230 ;
        RECT 344.700 2712.250 344.840 2794.275 ;
        RECT 351.070 2792.915 351.350 2793.285 ;
        RECT 351.140 2717.950 351.280 2792.915 ;
        RECT 351.600 2718.290 351.740 2794.275 ;
        RECT 358.500 2718.630 358.640 2794.275 ;
        RECT 362.640 2791.050 362.780 2794.275 ;
        RECT 362.580 2790.730 362.840 2791.050 ;
        RECT 365.400 2719.990 365.540 2794.275 ;
        RECT 368.620 2792.070 368.760 2794.275 ;
        RECT 368.560 2791.750 368.820 2792.070 ;
        RECT 371.380 2791.390 371.520 2794.275 ;
        RECT 375.060 2793.770 375.200 2794.275 ;
        RECT 375.000 2793.450 375.260 2793.770 ;
        RECT 371.320 2791.070 371.580 2791.390 ;
        RECT 365.340 2719.670 365.600 2719.990 ;
        RECT 379.200 2718.630 379.340 2794.275 ;
        RECT 379.590 2792.915 379.870 2793.285 ;
        RECT 379.600 2792.770 379.860 2792.915 ;
        RECT 384.260 2790.710 384.400 2794.275 ;
        RECT 386.960 2794.130 387.220 2794.275 ;
        RECT 392.480 2793.285 392.740 2793.430 ;
        RECT 392.470 2792.915 392.750 2793.285 ;
        RECT 384.200 2790.390 384.460 2790.710 ;
        RECT 358.440 2718.310 358.700 2718.630 ;
        RECT 377.300 2718.310 377.560 2718.630 ;
        RECT 379.140 2718.310 379.400 2718.630 ;
        RECT 351.540 2717.970 351.800 2718.290 ;
        RECT 367.180 2717.970 367.440 2718.290 ;
        RECT 351.080 2717.630 351.340 2717.950 ;
        RECT 356.600 2717.630 356.860 2717.950 ;
        RECT 344.700 2712.110 345.300 2712.250 ;
        RECT 336.030 2700.000 337.480 2700.010 ;
        RECT 325.840 2699.940 326.130 2700.000 ;
        RECT 315.270 2696.000 315.550 2699.870 ;
        RECT 325.850 2696.000 326.130 2699.940 ;
        RECT 335.970 2699.870 337.480 2700.000 ;
        RECT 345.160 2700.010 345.300 2712.110 ;
        RECT 345.160 2700.000 346.610 2700.010 ;
        RECT 356.660 2700.000 356.800 2717.630 ;
        RECT 367.240 2700.000 367.380 2717.970 ;
        RECT 377.360 2700.000 377.500 2718.310 ;
        RECT 393.000 2718.290 393.140 2794.275 ;
        RECT 396.680 2790.030 396.820 2794.275 ;
        RECT 397.070 2792.915 397.350 2793.285 ;
        RECT 397.140 2792.750 397.280 2792.915 ;
        RECT 397.080 2792.430 397.340 2792.750 ;
        RECT 396.620 2789.710 396.880 2790.030 ;
        RECT 392.940 2717.970 393.200 2718.290 ;
        RECT 399.440 2717.950 399.580 2794.275 ;
        RECT 404.040 2792.410 404.180 2794.275 ;
        RECT 403.980 2792.090 404.240 2792.410 ;
        RECT 406.340 2790.370 406.480 2794.275 ;
        RECT 410.020 2791.730 410.160 2794.275 ;
        RECT 414.620 2792.070 414.760 2794.275 ;
        RECT 414.560 2791.750 414.820 2792.070 ;
        RECT 407.200 2791.410 407.460 2791.730 ;
        RECT 409.960 2791.410 410.220 2791.730 ;
        RECT 407.260 2791.050 407.400 2791.410 ;
        RECT 419.220 2791.050 419.360 2794.275 ;
        RECT 421.060 2793.770 421.200 2794.275 ;
        RECT 421.000 2793.450 421.260 2793.770 ;
        RECT 426.970 2792.915 427.250 2793.285 ;
        RECT 426.980 2792.770 427.240 2792.915 ;
        RECT 407.200 2790.730 407.460 2791.050 ;
        RECT 419.160 2790.730 419.420 2791.050 ;
        RECT 406.280 2790.050 406.540 2790.370 ;
        RECT 413.630 2789.515 413.910 2789.885 ;
        RECT 408.580 2721.710 408.840 2722.030 ;
        RECT 399.380 2717.630 399.640 2717.950 ;
        RECT 398.460 2715.250 398.720 2715.570 ;
        RECT 387.870 2714.715 388.150 2715.085 ;
        RECT 387.940 2700.000 388.080 2714.715 ;
        RECT 398.520 2700.000 398.660 2715.250 ;
        RECT 408.640 2700.000 408.780 2721.710 ;
        RECT 413.700 2720.330 413.840 2789.515 ;
        RECT 427.040 2788.670 427.180 2792.770 ;
        RECT 426.980 2788.350 427.240 2788.670 ;
        RECT 419.160 2722.050 419.420 2722.370 ;
        RECT 413.640 2720.010 413.900 2720.330 ;
        RECT 419.220 2700.000 419.360 2722.050 ;
        RECT 427.500 2721.010 427.640 2794.275 ;
        RECT 431.580 2794.130 431.840 2794.275 ;
        RECT 433.420 2794.130 433.680 2794.450 ;
        RECT 433.870 2794.275 434.150 2794.645 ;
        RECT 439.390 2794.275 439.670 2794.645 ;
        RECT 441.230 2794.275 441.510 2794.645 ;
        RECT 444.450 2794.275 444.730 2794.645 ;
        RECT 445.830 2794.275 446.110 2794.645 ;
        RECT 449.050 2794.275 449.330 2794.645 ;
        RECT 455.030 2794.275 455.310 2794.645 ;
        RECT 461.010 2794.275 461.290 2794.645 ;
        RECT 462.390 2794.275 462.670 2794.645 ;
        RECT 466.530 2794.275 466.810 2794.645 ;
        RECT 468.830 2794.275 469.110 2794.645 ;
        RECT 475.270 2794.275 475.550 2794.645 ;
        RECT 478.490 2794.275 478.770 2794.645 ;
        RECT 482.630 2794.275 482.910 2794.645 ;
        RECT 485.850 2794.275 486.130 2794.645 ;
        RECT 489.070 2794.275 489.350 2794.645 ;
        RECT 491.830 2794.275 492.110 2794.645 ;
        RECT 496.430 2794.275 496.710 2794.645 ;
        RECT 500.110 2794.275 500.390 2794.645 ;
        RECT 510.230 2794.275 510.510 2794.645 ;
        RECT 524.030 2794.275 524.310 2794.645 ;
        RECT 536.450 2794.275 536.730 2794.645 ;
        RECT 542.430 2794.275 542.710 2794.645 ;
        RECT 433.480 2793.090 433.620 2794.130 ;
        RECT 433.420 2792.770 433.680 2793.090 ;
        RECT 429.280 2722.390 429.540 2722.710 ;
        RECT 427.440 2720.690 427.700 2721.010 ;
        RECT 429.340 2700.000 429.480 2722.390 ;
        RECT 433.940 2721.690 434.080 2794.275 ;
        RECT 439.460 2793.430 439.600 2794.275 ;
        RECT 434.330 2792.915 434.610 2793.285 ;
        RECT 439.400 2793.110 439.660 2793.430 ;
        RECT 433.880 2721.370 434.140 2721.690 ;
        RECT 434.400 2720.670 434.540 2792.915 ;
        RECT 439.860 2723.070 440.120 2723.390 ;
        RECT 434.340 2720.350 434.600 2720.670 ;
        RECT 439.920 2700.000 440.060 2723.070 ;
        RECT 441.300 2721.350 441.440 2794.275 ;
        RECT 444.520 2792.750 444.660 2794.275 ;
        RECT 444.460 2792.430 444.720 2792.750 ;
        RECT 445.900 2789.350 446.040 2794.275 ;
        RECT 449.120 2792.410 449.260 2794.275 ;
        RECT 449.060 2792.090 449.320 2792.410 ;
        RECT 445.840 2789.030 446.100 2789.350 ;
        RECT 449.980 2723.750 450.240 2724.070 ;
        RECT 441.240 2721.030 441.500 2721.350 ;
        RECT 450.040 2700.000 450.180 2723.750 ;
        RECT 455.100 2716.590 455.240 2794.275 ;
        RECT 455.490 2792.915 455.770 2793.285 ;
        RECT 455.560 2791.730 455.700 2792.915 ;
        RECT 461.080 2791.730 461.220 2794.275 ;
        RECT 462.460 2792.070 462.600 2794.275 ;
        RECT 466.600 2793.770 466.740 2794.275 ;
        RECT 468.840 2794.130 469.100 2794.275 ;
        RECT 466.540 2793.450 466.800 2793.770 ;
        RECT 468.370 2792.915 468.650 2793.285 ;
        RECT 473.890 2792.915 474.170 2793.285 ;
        RECT 462.400 2791.750 462.660 2792.070 ;
        RECT 465.620 2791.750 465.880 2792.070 ;
        RECT 455.500 2791.410 455.760 2791.730 ;
        RECT 461.020 2791.410 461.280 2791.730 ;
        RECT 455.560 2788.330 455.700 2791.410 ;
        RECT 465.680 2789.010 465.820 2791.750 ;
        RECT 465.620 2788.690 465.880 2789.010 ;
        RECT 455.500 2788.010 455.760 2788.330 ;
        RECT 460.560 2724.090 460.820 2724.410 ;
        RECT 455.040 2716.270 455.300 2716.590 ;
        RECT 460.620 2700.000 460.760 2724.090 ;
        RECT 468.440 2715.910 468.580 2792.915 ;
        RECT 473.960 2792.410 474.100 2792.915 ;
        RECT 473.900 2792.090 474.160 2792.410 ;
        RECT 473.960 2788.670 474.100 2792.090 ;
        RECT 473.900 2788.350 474.160 2788.670 ;
        RECT 470.680 2724.770 470.940 2725.090 ;
        RECT 468.380 2715.590 468.640 2715.910 ;
        RECT 470.740 2700.000 470.880 2724.770 ;
        RECT 475.340 2715.570 475.480 2794.275 ;
        RECT 478.560 2793.090 478.700 2794.275 ;
        RECT 478.500 2792.770 478.760 2793.090 ;
        RECT 482.700 2725.430 482.840 2794.275 ;
        RECT 485.920 2793.430 486.060 2794.275 ;
        RECT 485.860 2793.110 486.120 2793.430 ;
        RECT 485.920 2789.690 486.060 2793.110 ;
        RECT 489.140 2792.070 489.280 2794.275 ;
        RECT 491.900 2792.750 492.040 2794.275 ;
        RECT 491.840 2792.430 492.100 2792.750 ;
        RECT 489.080 2791.750 489.340 2792.070 ;
        RECT 485.860 2789.370 486.120 2789.690 ;
        RECT 491.900 2788.670 492.040 2792.430 ;
        RECT 491.840 2788.350 492.100 2788.670 ;
        RECT 482.640 2725.110 482.900 2725.430 ;
        RECT 481.250 2716.075 481.530 2716.445 ;
        RECT 475.280 2715.250 475.540 2715.570 ;
        RECT 481.320 2700.000 481.460 2716.075 ;
        RECT 496.500 2715.230 496.640 2794.275 ;
        RECT 497.360 2793.110 497.620 2793.430 ;
        RECT 497.420 2792.605 497.560 2793.110 ;
        RECT 500.180 2792.750 500.320 2794.275 ;
        RECT 510.300 2793.430 510.440 2794.275 ;
        RECT 513.920 2793.450 514.180 2793.770 ;
        RECT 510.240 2793.110 510.500 2793.430 ;
        RECT 497.350 2792.235 497.630 2792.605 ;
        RECT 500.120 2792.430 500.380 2792.750 ;
        RECT 501.950 2792.235 502.230 2792.605 ;
        RECT 500.110 2788.155 500.390 2788.525 ;
        RECT 502.020 2788.330 502.160 2792.235 ;
        RECT 504.250 2788.835 504.530 2789.205 ;
        RECT 507.010 2788.835 507.290 2789.205 ;
        RECT 504.260 2788.690 504.520 2788.835 ;
        RECT 500.120 2788.010 500.380 2788.155 ;
        RECT 501.960 2788.010 502.220 2788.330 ;
        RECT 491.840 2714.910 492.100 2715.230 ;
        RECT 496.440 2714.910 496.700 2715.230 ;
        RECT 491.900 2700.000 492.040 2714.910 ;
        RECT 500.180 2713.530 500.320 2788.010 ;
        RECT 501.960 2714.570 502.220 2714.890 ;
        RECT 500.120 2713.210 500.380 2713.530 ;
        RECT 502.020 2700.000 502.160 2714.570 ;
        RECT 507.080 2713.190 507.220 2788.835 ;
        RECT 513.980 2787.845 514.120 2793.450 ;
        RECT 520.820 2792.770 521.080 2793.090 ;
        RECT 520.880 2787.845 521.020 2792.770 ;
        RECT 524.100 2792.750 524.240 2794.275 ;
        RECT 536.520 2793.770 536.660 2794.275 ;
        RECT 531.400 2793.450 531.660 2793.770 ;
        RECT 536.460 2793.450 536.720 2793.770 ;
        RECT 531.460 2793.285 531.600 2793.450 ;
        RECT 531.390 2792.915 531.670 2793.285 ;
        RECT 542.500 2793.090 542.640 2794.275 ;
        RECT 686.420 2794.130 686.680 2794.450 ;
        RECT 542.440 2792.770 542.700 2793.090 ;
        RECT 524.040 2792.430 524.300 2792.750 ;
        RECT 542.430 2792.235 542.710 2792.605 ;
        RECT 551.630 2792.235 551.910 2792.605 ;
        RECT 527.720 2789.370 527.980 2789.690 ;
        RECT 541.510 2789.515 541.790 2789.885 ;
        RECT 527.780 2787.845 527.920 2789.370 ;
        RECT 541.580 2788.670 541.720 2789.515 ;
        RECT 534.610 2788.155 534.890 2788.525 ;
        RECT 541.520 2788.350 541.780 2788.670 ;
        RECT 510.230 2787.475 510.510 2787.845 ;
        RECT 513.910 2787.475 514.190 2787.845 ;
        RECT 517.130 2787.475 517.410 2787.845 ;
        RECT 520.810 2787.475 521.090 2787.845 ;
        RECT 527.710 2787.475 527.990 2787.845 ;
        RECT 530.930 2787.475 531.210 2787.845 ;
        RECT 510.300 2724.750 510.440 2787.475 ;
        RECT 510.240 2724.430 510.500 2724.750 ;
        RECT 512.540 2717.290 512.800 2717.610 ;
        RECT 507.020 2712.870 507.280 2713.190 ;
        RECT 512.600 2700.000 512.740 2717.290 ;
        RECT 513.980 2714.210 514.120 2787.475 ;
        RECT 517.200 2715.765 517.340 2787.475 ;
        RECT 517.130 2715.395 517.410 2715.765 ;
        RECT 513.920 2713.890 514.180 2714.210 ;
        RECT 520.880 2713.870 521.020 2787.475 ;
        RECT 522.660 2716.950 522.920 2717.270 ;
        RECT 520.820 2713.550 521.080 2713.870 ;
        RECT 522.720 2700.000 522.860 2716.950 ;
        RECT 527.780 2714.550 527.920 2787.475 ;
        RECT 531.000 2723.730 531.140 2787.475 ;
        RECT 530.940 2723.410 531.200 2723.730 ;
        RECT 533.240 2716.610 533.500 2716.930 ;
        RECT 527.720 2714.230 527.980 2714.550 ;
        RECT 533.300 2700.000 533.440 2716.610 ;
        RECT 534.680 2712.510 534.820 2788.155 ;
        RECT 541.580 2714.890 541.720 2788.350 ;
        RECT 542.500 2788.330 542.640 2792.235 ;
        RECT 542.440 2788.010 542.700 2788.330 ;
        RECT 541.520 2714.570 541.780 2714.890 ;
        RECT 542.500 2712.850 542.640 2788.010 ;
        RECT 551.700 2723.050 551.840 2792.235 ;
        RECT 648.240 2789.370 648.500 2789.690 ;
        RECT 627.540 2789.030 627.800 2789.350 ;
        RECT 606.840 2788.690 607.100 2789.010 ;
        RECT 586.140 2788.350 586.400 2788.670 ;
        RECT 551.640 2722.730 551.900 2723.050 ;
        RECT 564.060 2719.330 564.320 2719.650 ;
        RECT 553.940 2718.990 554.200 2719.310 ;
        RECT 543.360 2715.930 543.620 2716.250 ;
        RECT 542.440 2712.530 542.700 2712.850 ;
        RECT 534.620 2712.190 534.880 2712.510 ;
        RECT 543.420 2700.000 543.560 2715.930 ;
        RECT 554.000 2700.000 554.140 2718.990 ;
        RECT 564.120 2700.000 564.260 2719.330 ;
        RECT 574.640 2715.930 574.900 2716.250 ;
        RECT 574.700 2700.000 574.840 2715.930 ;
        RECT 586.200 2700.010 586.340 2788.350 ;
        RECT 595.340 2716.610 595.600 2716.930 ;
        RECT 585.350 2700.000 586.340 2700.010 ;
        RECT 345.160 2699.870 346.830 2700.000 ;
        RECT 356.660 2699.940 356.950 2700.000 ;
        RECT 367.240 2699.940 367.530 2700.000 ;
        RECT 377.360 2699.940 377.650 2700.000 ;
        RECT 387.940 2699.940 388.230 2700.000 ;
        RECT 398.520 2699.940 398.810 2700.000 ;
        RECT 408.640 2699.940 408.930 2700.000 ;
        RECT 419.220 2699.940 419.510 2700.000 ;
        RECT 429.340 2699.940 429.630 2700.000 ;
        RECT 439.920 2699.940 440.210 2700.000 ;
        RECT 450.040 2699.940 450.330 2700.000 ;
        RECT 460.620 2699.940 460.910 2700.000 ;
        RECT 470.740 2699.940 471.030 2700.000 ;
        RECT 481.320 2699.940 481.610 2700.000 ;
        RECT 491.900 2699.940 492.190 2700.000 ;
        RECT 502.020 2699.940 502.310 2700.000 ;
        RECT 512.600 2699.940 512.890 2700.000 ;
        RECT 522.720 2699.940 523.010 2700.000 ;
        RECT 533.300 2699.940 533.590 2700.000 ;
        RECT 543.420 2699.940 543.710 2700.000 ;
        RECT 554.000 2699.940 554.290 2700.000 ;
        RECT 564.120 2699.940 564.410 2700.000 ;
        RECT 574.700 2699.940 574.990 2700.000 ;
        RECT 335.970 2696.000 336.250 2699.870 ;
        RECT 346.550 2696.000 346.830 2699.870 ;
        RECT 356.670 2696.000 356.950 2699.940 ;
        RECT 367.250 2696.000 367.530 2699.940 ;
        RECT 377.370 2696.000 377.650 2699.940 ;
        RECT 387.950 2696.000 388.230 2699.940 ;
        RECT 398.530 2696.000 398.810 2699.940 ;
        RECT 408.650 2696.000 408.930 2699.940 ;
        RECT 419.230 2696.000 419.510 2699.940 ;
        RECT 429.350 2696.000 429.630 2699.940 ;
        RECT 439.930 2696.000 440.210 2699.940 ;
        RECT 450.050 2696.000 450.330 2699.940 ;
        RECT 460.630 2696.000 460.910 2699.940 ;
        RECT 470.750 2696.000 471.030 2699.940 ;
        RECT 481.330 2696.000 481.610 2699.940 ;
        RECT 491.910 2696.000 492.190 2699.940 ;
        RECT 502.030 2696.000 502.310 2699.940 ;
        RECT 512.610 2696.000 512.890 2699.940 ;
        RECT 522.730 2696.000 523.010 2699.940 ;
        RECT 533.310 2696.000 533.590 2699.940 ;
        RECT 543.430 2696.000 543.710 2699.940 ;
        RECT 554.010 2696.000 554.290 2699.940 ;
        RECT 564.130 2696.000 564.410 2699.940 ;
        RECT 574.710 2696.000 574.990 2699.940 ;
        RECT 585.290 2699.870 586.340 2700.000 ;
        RECT 595.400 2700.000 595.540 2716.610 ;
        RECT 606.900 2700.010 607.040 2788.690 ;
        RECT 616.040 2716.950 616.300 2717.270 ;
        RECT 606.050 2700.000 607.040 2700.010 ;
        RECT 595.400 2699.940 595.690 2700.000 ;
        RECT 585.290 2696.000 585.570 2699.870 ;
        RECT 595.410 2696.000 595.690 2699.940 ;
        RECT 605.990 2699.870 607.040 2700.000 ;
        RECT 616.100 2700.000 616.240 2716.950 ;
        RECT 627.600 2700.010 627.740 2789.030 ;
        RECT 636.740 2717.290 637.000 2717.610 ;
        RECT 626.750 2700.000 627.740 2700.010 ;
        RECT 616.100 2699.940 616.390 2700.000 ;
        RECT 605.990 2696.000 606.270 2699.870 ;
        RECT 616.110 2696.000 616.390 2699.940 ;
        RECT 626.690 2699.870 627.740 2700.000 ;
        RECT 636.800 2700.000 636.940 2717.290 ;
        RECT 648.300 2700.010 648.440 2789.370 ;
        RECT 658.820 2784.270 659.080 2784.590 ;
        RECT 658.880 2713.530 659.020 2784.270 ;
        RECT 686.480 2714.210 686.620 2794.130 ;
        RECT 707.120 2793.450 707.380 2793.770 ;
        RECT 700.220 2793.110 700.480 2793.430 ;
        RECT 693.320 2791.750 693.580 2792.070 ;
        RECT 687.340 2791.410 687.600 2791.730 ;
        RECT 686.880 2791.070 687.140 2791.390 ;
        RECT 678.600 2713.890 678.860 2714.210 ;
        RECT 686.420 2713.890 686.680 2714.210 ;
        RECT 657.440 2713.210 657.700 2713.530 ;
        RECT 658.820 2713.210 659.080 2713.530 ;
        RECT 647.450 2700.000 648.440 2700.010 ;
        RECT 636.800 2699.940 637.090 2700.000 ;
        RECT 626.690 2696.000 626.970 2699.870 ;
        RECT 636.810 2696.000 637.090 2699.940 ;
        RECT 647.390 2699.870 648.440 2700.000 ;
        RECT 657.500 2700.000 657.640 2713.210 ;
        RECT 668.020 2712.870 668.280 2713.190 ;
        RECT 668.080 2700.000 668.220 2712.870 ;
        RECT 678.660 2700.000 678.800 2713.890 ;
        RECT 686.940 2712.170 687.080 2791.070 ;
        RECT 687.400 2713.190 687.540 2791.410 ;
        RECT 693.380 2714.210 693.520 2791.750 ;
        RECT 700.280 2718.485 700.420 2793.110 ;
        RECT 700.680 2792.090 700.940 2792.410 ;
        RECT 700.210 2718.115 700.490 2718.485 ;
        RECT 700.740 2714.550 700.880 2792.090 ;
        RECT 707.180 2717.125 707.320 2793.450 ;
        RECT 741.620 2792.770 741.880 2793.090 ;
        RECT 720.920 2792.430 721.180 2792.750 ;
        RECT 707.110 2716.755 707.390 2717.125 ;
        RECT 720.980 2714.890 721.120 2792.430 ;
        RECT 727.820 2790.390 728.080 2790.710 ;
        RECT 727.880 2718.630 728.020 2790.390 ;
        RECT 740.700 2719.670 740.960 2719.990 ;
        RECT 727.820 2718.310 728.080 2718.630 ;
        RECT 720.000 2714.570 720.260 2714.890 ;
        RECT 720.920 2714.570 721.180 2714.890 ;
        RECT 699.300 2714.230 699.560 2714.550 ;
        RECT 700.680 2714.230 700.940 2714.550 ;
        RECT 693.320 2713.890 693.580 2714.210 ;
        RECT 688.720 2713.550 688.980 2713.870 ;
        RECT 687.340 2712.870 687.600 2713.190 ;
        RECT 686.880 2711.850 687.140 2712.170 ;
        RECT 688.780 2700.000 688.920 2713.550 ;
        RECT 699.360 2700.000 699.500 2714.230 ;
        RECT 709.420 2712.190 709.680 2712.510 ;
        RECT 709.480 2700.000 709.620 2712.190 ;
        RECT 720.060 2700.000 720.200 2714.570 ;
        RECT 730.120 2712.530 730.380 2712.850 ;
        RECT 730.180 2700.000 730.320 2712.530 ;
        RECT 740.760 2700.000 740.900 2719.670 ;
        RECT 741.680 2717.805 741.820 2792.770 ;
        RECT 748.520 2790.730 748.780 2791.050 ;
        RECT 741.610 2717.435 741.890 2717.805 ;
        RECT 748.580 2712.510 748.720 2790.730 ;
        RECT 762.780 2790.050 763.040 2790.370 ;
        RECT 762.320 2789.710 762.580 2790.030 ;
        RECT 762.380 2717.950 762.520 2789.710 ;
        RECT 762.840 2718.630 762.980 2790.050 ;
        RECT 865.360 2721.370 865.620 2721.690 ;
        RECT 844.200 2720.690 844.460 2721.010 ;
        RECT 823.500 2720.010 823.760 2720.330 ;
        RECT 762.780 2718.310 763.040 2718.630 ;
        RECT 813.380 2718.310 813.640 2718.630 ;
        RECT 782.100 2717.970 782.360 2718.290 ;
        RECT 762.320 2717.630 762.580 2717.950 ;
        RECT 761.400 2712.530 761.660 2712.850 ;
        RECT 771.980 2712.530 772.240 2712.850 ;
        RECT 748.520 2712.190 748.780 2712.510 ;
        RECT 750.820 2711.850 751.080 2712.170 ;
        RECT 750.880 2700.000 751.020 2711.850 ;
        RECT 761.460 2700.000 761.600 2712.530 ;
        RECT 772.040 2700.000 772.180 2712.530 ;
        RECT 782.160 2700.000 782.300 2717.970 ;
        RECT 792.680 2717.630 792.940 2717.950 ;
        RECT 792.740 2700.000 792.880 2717.630 ;
        RECT 802.800 2711.850 803.060 2712.170 ;
        RECT 802.860 2700.000 803.000 2711.850 ;
        RECT 813.440 2700.000 813.580 2718.310 ;
        RECT 823.560 2700.000 823.700 2720.010 ;
        RECT 834.080 2712.530 834.340 2712.850 ;
        RECT 834.140 2700.000 834.280 2712.530 ;
        RECT 844.260 2700.000 844.400 2720.690 ;
        RECT 854.780 2720.350 855.040 2720.670 ;
        RECT 854.840 2700.000 854.980 2720.350 ;
        RECT 865.420 2700.000 865.560 2721.370 ;
        RECT 875.480 2721.030 875.740 2721.350 ;
        RECT 875.540 2700.000 875.680 2721.030 ;
        RECT 896.180 2716.270 896.440 2716.590 ;
        RECT 941.780 2716.445 941.920 3230.155 ;
        RECT 942.170 3224.715 942.450 3225.085 ;
        RECT 942.240 2725.090 942.380 3224.715 ;
        RECT 942.630 3215.875 942.910 3216.245 ;
        RECT 942.180 2724.770 942.440 2725.090 ;
        RECT 942.700 2724.410 942.840 3215.875 ;
        RECT 943.090 3209.755 943.370 3210.125 ;
        RECT 942.640 2724.090 942.900 2724.410 ;
        RECT 943.160 2724.070 943.300 3209.755 ;
        RECT 943.550 3201.595 943.830 3201.965 ;
        RECT 943.100 2723.750 943.360 2724.070 ;
        RECT 943.620 2723.390 943.760 3201.595 ;
        RECT 944.010 3196.155 944.290 3196.525 ;
        RECT 943.560 2723.070 943.820 2723.390 ;
        RECT 944.080 2722.710 944.220 3196.155 ;
        RECT 944.470 3187.995 944.750 3188.365 ;
        RECT 944.020 2722.390 944.280 2722.710 ;
        RECT 944.540 2722.370 944.680 3187.995 ;
        RECT 944.930 2898.315 945.210 2898.685 ;
        RECT 944.480 2722.050 944.740 2722.370 ;
        RECT 886.060 2713.210 886.320 2713.530 ;
        RECT 886.120 2700.000 886.260 2713.210 ;
        RECT 896.240 2700.000 896.380 2716.270 ;
        RECT 941.710 2716.075 941.990 2716.445 ;
        RECT 916.880 2715.590 917.140 2715.910 ;
        RECT 906.760 2712.870 907.020 2713.190 ;
        RECT 906.820 2700.000 906.960 2712.870 ;
        RECT 916.940 2700.000 917.080 2715.590 ;
        RECT 937.580 2715.250 937.840 2715.570 ;
        RECT 927.460 2713.550 927.720 2713.870 ;
        RECT 927.520 2700.000 927.660 2713.550 ;
        RECT 937.640 2700.000 937.780 2715.250 ;
        RECT 945.000 2715.085 945.140 2898.315 ;
      LAYER met2 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met2 ;
        RECT 1333.240 3249.565 1333.380 3252.110 ;
        RECT 1333.170 3249.195 1333.450 3249.565 ;
        RECT 1536.950 3230.155 1537.230 3230.525 ;
        RECT 1537.020 3229.650 1537.160 3230.155 ;
        RECT 1459.220 3229.330 1459.480 3229.650 ;
        RECT 1536.960 3229.330 1537.220 3229.650 ;
        RECT 1452.320 3222.190 1452.580 3222.510 ;
        RECT 1438.520 3215.390 1438.780 3215.710 ;
        RECT 1431.620 3208.590 1431.880 3208.910 ;
        RECT 1424.720 3201.450 1424.980 3201.770 ;
        RECT 1345.590 2946.595 1345.870 2946.965 ;
        RECT 1345.660 2936.085 1345.800 2946.595 ;
        RECT 1345.590 2935.715 1345.870 2936.085 ;
        RECT 1352.030 2901.715 1352.310 2902.085 ;
        RECT 1352.100 2901.550 1352.240 2901.715 ;
        RECT 1352.040 2901.230 1352.300 2901.550 ;
        RECT 1395.740 2901.230 1396.000 2901.550 ;
        RECT 1054.870 2799.715 1055.150 2800.085 ;
        RECT 979.890 2794.275 980.170 2794.645 ;
        RECT 1001.050 2794.275 1001.330 2794.645 ;
        RECT 1013.930 2794.275 1014.210 2794.645 ;
        RECT 1018.990 2794.275 1019.270 2794.645 ;
        RECT 1020.830 2794.275 1021.110 2794.645 ;
        RECT 1027.730 2794.275 1028.010 2794.645 ;
        RECT 1034.630 2794.275 1034.910 2794.645 ;
        RECT 1042.450 2794.275 1042.730 2794.645 ;
        RECT 1053.030 2794.275 1053.310 2794.645 ;
        RECT 948.160 2725.110 948.420 2725.430 ;
        RECT 944.930 2714.715 945.210 2715.085 ;
        RECT 948.220 2700.000 948.360 2725.110 ;
        RECT 979.960 2722.030 980.100 2794.275 ;
        RECT 1001.120 2794.110 1001.260 2794.275 ;
        RECT 1001.060 2793.790 1001.320 2794.110 ;
        RECT 1010.710 2792.915 1010.990 2793.285 ;
        RECT 1007.490 2788.155 1007.770 2788.525 ;
        RECT 1010.780 2788.330 1010.920 2792.915 ;
        RECT 1007.560 2787.990 1007.700 2788.155 ;
        RECT 1010.720 2788.010 1010.980 2788.330 ;
        RECT 1007.500 2787.670 1007.760 2787.990 ;
        RECT 989.560 2724.430 989.820 2724.750 ;
        RECT 979.900 2721.710 980.160 2722.030 ;
        RECT 968.860 2714.910 969.120 2715.230 ;
        RECT 958.740 2713.890 959.000 2714.210 ;
        RECT 958.800 2700.000 958.940 2713.890 ;
        RECT 968.920 2700.000 969.060 2714.910 ;
        RECT 979.440 2714.230 979.700 2714.550 ;
        RECT 979.500 2700.000 979.640 2714.230 ;
        RECT 989.620 2700.000 989.760 2724.430 ;
        RECT 1000.130 2718.115 1000.410 2718.485 ;
        RECT 1000.200 2700.000 1000.340 2718.115 ;
        RECT 1010.780 2716.250 1010.920 2788.010 ;
        RECT 1010.720 2715.930 1010.980 2716.250 ;
        RECT 1010.250 2715.395 1010.530 2715.765 ;
        RECT 1010.320 2700.000 1010.460 2715.395 ;
        RECT 1014.000 2715.230 1014.140 2794.275 ;
        RECT 1019.060 2791.050 1019.200 2794.275 ;
        RECT 1019.000 2790.730 1019.260 2791.050 ;
        RECT 1019.060 2788.670 1019.200 2790.730 ;
        RECT 1019.000 2788.350 1019.260 2788.670 ;
        RECT 1020.900 2715.910 1021.040 2794.275 ;
        RECT 1024.510 2792.915 1024.790 2793.285 ;
        RECT 1024.580 2788.670 1024.720 2792.915 ;
        RECT 1024.520 2788.350 1024.780 2788.670 ;
        RECT 1024.580 2716.930 1024.720 2788.350 ;
        RECT 1027.800 2718.630 1027.940 2794.275 ;
        RECT 1034.700 2791.390 1034.840 2794.275 ;
        RECT 1042.520 2792.750 1042.660 2794.275 ;
        RECT 1045.210 2792.915 1045.490 2793.285 ;
        RECT 1042.460 2792.430 1042.720 2792.750 ;
        RECT 1034.640 2791.070 1034.900 2791.390 ;
        RECT 1034.700 2789.010 1034.840 2791.070 ;
        RECT 1042.520 2789.350 1042.660 2792.430 ;
        RECT 1042.460 2789.030 1042.720 2789.350 ;
        RECT 1045.280 2789.010 1045.420 2792.915 ;
        RECT 1053.100 2792.070 1053.240 2794.275 ;
        RECT 1053.040 2791.750 1053.300 2792.070 ;
        RECT 1034.640 2788.690 1034.900 2789.010 ;
        RECT 1045.220 2788.690 1045.480 2789.010 ;
        RECT 1038.310 2788.155 1038.590 2788.525 ;
        RECT 1038.380 2787.990 1038.520 2788.155 ;
        RECT 1034.630 2787.475 1034.910 2787.845 ;
        RECT 1038.320 2787.670 1038.580 2787.990 ;
        RECT 1030.960 2723.410 1031.220 2723.730 ;
        RECT 1027.740 2718.310 1028.000 2718.630 ;
        RECT 1024.520 2716.610 1024.780 2716.930 ;
        RECT 1020.840 2715.590 1021.100 2715.910 ;
        RECT 1013.940 2714.910 1014.200 2715.230 ;
        RECT 1020.840 2714.570 1021.100 2714.890 ;
        RECT 1020.900 2700.000 1021.040 2714.570 ;
        RECT 1031.020 2700.000 1031.160 2723.410 ;
        RECT 1034.700 2718.290 1034.840 2787.475 ;
        RECT 1034.640 2717.970 1034.900 2718.290 ;
        RECT 1038.380 2717.270 1038.520 2787.670 ;
        RECT 1041.530 2787.475 1041.810 2787.845 ;
        RECT 1041.600 2717.950 1041.740 2787.475 ;
        RECT 1041.540 2717.630 1041.800 2717.950 ;
        RECT 1045.280 2717.610 1045.420 2788.690 ;
        RECT 1048.430 2787.475 1048.710 2787.845 ;
        RECT 1048.500 2717.610 1048.640 2787.475 ;
        RECT 1045.220 2717.290 1045.480 2717.610 ;
        RECT 1048.440 2717.290 1048.700 2717.610 ;
        RECT 1052.110 2717.435 1052.390 2717.805 ;
        RECT 1038.320 2716.950 1038.580 2717.270 ;
        RECT 1041.530 2716.755 1041.810 2717.125 ;
        RECT 1041.600 2700.000 1041.740 2716.755 ;
        RECT 1052.180 2700.000 1052.320 2717.435 ;
        RECT 1054.940 2714.890 1055.080 2799.715 ;
        RECT 1059.010 2794.275 1059.290 2794.645 ;
        RECT 1065.910 2794.275 1066.190 2794.645 ;
        RECT 1070.050 2794.275 1070.330 2794.645 ;
        RECT 1076.490 2794.275 1076.770 2794.645 ;
        RECT 1087.530 2794.275 1087.810 2794.645 ;
        RECT 1093.970 2794.275 1094.250 2794.645 ;
        RECT 1100.410 2794.275 1100.690 2794.645 ;
        RECT 1105.470 2794.275 1105.750 2794.645 ;
        RECT 1110.990 2794.275 1111.270 2794.645 ;
        RECT 1122.490 2794.275 1122.770 2794.645 ;
        RECT 1129.390 2794.275 1129.670 2794.645 ;
        RECT 1130.770 2794.275 1131.050 2794.645 ;
        RECT 1135.830 2794.275 1136.110 2794.645 ;
        RECT 1138.130 2794.275 1138.410 2794.645 ;
        RECT 1139.970 2794.275 1140.250 2794.645 ;
        RECT 1145.030 2794.275 1145.310 2794.645 ;
        RECT 1147.330 2794.275 1147.610 2794.645 ;
        RECT 1151.930 2794.275 1152.210 2794.645 ;
        RECT 1158.830 2794.275 1159.110 2794.645 ;
        RECT 1165.270 2794.275 1165.550 2794.645 ;
        RECT 1166.190 2794.275 1166.470 2794.645 ;
        RECT 1172.630 2794.275 1172.910 2794.645 ;
        RECT 1179.530 2794.275 1179.810 2794.645 ;
        RECT 1186.430 2794.275 1186.710 2794.645 ;
        RECT 1200.230 2794.275 1200.510 2794.645 ;
        RECT 1059.080 2791.730 1059.220 2794.275 ;
        RECT 1065.980 2792.410 1066.120 2794.275 ;
        RECT 1065.920 2792.090 1066.180 2792.410 ;
        RECT 1055.800 2791.410 1056.060 2791.730 ;
        RECT 1059.020 2791.410 1059.280 2791.730 ;
        RECT 1055.330 2788.155 1055.610 2788.525 ;
        RECT 1055.860 2788.330 1056.000 2791.410 ;
        RECT 1065.980 2791.050 1066.120 2792.090 ;
        RECT 1065.920 2790.730 1066.180 2791.050 ;
        RECT 1070.120 2788.670 1070.260 2794.275 ;
        RECT 1076.560 2794.110 1076.700 2794.275 ;
        RECT 1076.500 2793.790 1076.760 2794.110 ;
        RECT 1076.560 2791.390 1076.700 2793.790 ;
        RECT 1087.600 2793.090 1087.740 2794.275 ;
        RECT 1087.990 2793.595 1088.270 2793.965 ;
        RECT 1094.040 2793.770 1094.180 2794.275 ;
        RECT 1087.540 2792.770 1087.800 2793.090 ;
        RECT 1076.500 2791.070 1076.760 2791.390 ;
        RECT 1076.040 2790.390 1076.300 2790.710 ;
        RECT 1076.100 2788.670 1076.240 2790.390 ;
        RECT 1070.060 2788.350 1070.320 2788.670 ;
        RECT 1076.040 2788.350 1076.300 2788.670 ;
        RECT 1055.400 2717.270 1055.540 2788.155 ;
        RECT 1055.800 2788.010 1056.060 2788.330 ;
        RECT 1087.600 2787.990 1087.740 2792.770 ;
        RECT 1088.060 2792.750 1088.200 2793.595 ;
        RECT 1093.980 2793.450 1094.240 2793.770 ;
        RECT 1088.000 2792.430 1088.260 2792.750 ;
        RECT 1094.040 2789.010 1094.180 2793.450 ;
        RECT 1100.480 2792.070 1100.620 2794.275 ;
        RECT 1100.420 2791.750 1100.680 2792.070 ;
        RECT 1105.540 2791.730 1105.680 2794.275 ;
        RECT 1111.060 2793.430 1111.200 2794.275 ;
        RECT 1122.560 2794.110 1122.700 2794.275 ;
        RECT 1117.890 2793.595 1118.170 2793.965 ;
        RECT 1122.500 2793.790 1122.760 2794.110 ;
        RECT 1111.000 2793.110 1111.260 2793.430 ;
        RECT 1111.060 2792.410 1111.200 2793.110 ;
        RECT 1111.000 2792.090 1111.260 2792.410 ;
        RECT 1105.480 2791.410 1105.740 2791.730 ;
        RECT 1117.960 2789.690 1118.100 2793.595 ;
        RECT 1122.560 2791.390 1122.700 2793.790 ;
        RECT 1129.460 2793.090 1129.600 2794.275 ;
        RECT 1129.400 2792.770 1129.660 2793.090 ;
        RECT 1122.500 2791.070 1122.760 2791.390 ;
        RECT 1117.900 2789.370 1118.160 2789.690 ;
        RECT 1093.980 2788.690 1094.240 2789.010 ;
        RECT 1089.830 2788.155 1090.110 2788.525 ;
        RECT 1062.230 2787.475 1062.510 2787.845 ;
        RECT 1069.130 2787.475 1069.410 2787.845 ;
        RECT 1076.030 2787.475 1076.310 2787.845 ;
        RECT 1082.930 2787.475 1083.210 2787.845 ;
        RECT 1087.540 2787.670 1087.800 2787.990 ;
        RECT 1089.370 2787.475 1089.650 2787.845 ;
        RECT 1062.300 2727.890 1062.440 2787.475 ;
        RECT 1061.840 2727.750 1062.440 2727.890 ;
        RECT 1055.340 2716.950 1055.600 2717.270 ;
        RECT 1061.840 2716.930 1061.980 2727.750 ;
        RECT 1062.240 2722.730 1062.500 2723.050 ;
        RECT 1061.780 2716.610 1062.040 2716.930 ;
        RECT 1054.880 2714.570 1055.140 2714.890 ;
        RECT 1062.300 2700.000 1062.440 2722.730 ;
        RECT 1069.200 2715.570 1069.340 2787.475 ;
        RECT 1076.100 2716.590 1076.240 2787.475 ;
        RECT 1083.000 2727.890 1083.140 2787.475 ;
        RECT 1082.540 2727.750 1083.140 2727.890 ;
        RECT 1076.040 2716.270 1076.300 2716.590 ;
        RECT 1082.540 2716.250 1082.680 2727.750 ;
        RECT 1082.480 2715.930 1082.740 2716.250 ;
        RECT 1082.940 2715.590 1083.200 2715.910 ;
        RECT 1069.140 2715.250 1069.400 2715.570 ;
        RECT 1072.820 2714.910 1073.080 2715.230 ;
        RECT 1072.880 2700.000 1073.020 2714.910 ;
        RECT 1083.000 2700.000 1083.140 2715.590 ;
        RECT 1089.440 2712.850 1089.580 2787.475 ;
        RECT 1089.900 2715.230 1090.040 2788.155 ;
        RECT 1096.730 2787.475 1097.010 2787.845 ;
        RECT 1103.630 2787.475 1103.910 2787.845 ;
        RECT 1110.530 2787.475 1110.810 2787.845 ;
        RECT 1117.430 2787.475 1117.710 2787.845 ;
        RECT 1124.330 2787.475 1124.610 2787.845 ;
        RECT 1093.520 2718.310 1093.780 2718.630 ;
        RECT 1089.840 2714.910 1090.100 2715.230 ;
        RECT 1089.380 2712.530 1089.640 2712.850 ;
        RECT 1093.580 2700.000 1093.720 2718.310 ;
        RECT 1096.800 2712.510 1096.940 2787.475 ;
        RECT 1103.700 2718.970 1103.840 2787.475 ;
        RECT 1103.640 2718.650 1103.900 2718.970 ;
        RECT 1102.720 2718.310 1102.980 2718.630 ;
        RECT 1102.780 2713.530 1102.920 2718.310 ;
        RECT 1103.640 2717.970 1103.900 2718.290 ;
        RECT 1102.720 2713.210 1102.980 2713.530 ;
        RECT 1096.740 2712.190 1097.000 2712.510 ;
        RECT 1103.700 2700.000 1103.840 2717.970 ;
        RECT 1110.600 2713.190 1110.740 2787.475 ;
        RECT 1114.220 2717.630 1114.480 2717.950 ;
        RECT 1110.540 2712.870 1110.800 2713.190 ;
        RECT 1114.280 2700.000 1114.420 2717.630 ;
        RECT 1117.500 2714.210 1117.640 2787.475 ;
        RECT 1124.400 2726.530 1124.540 2787.475 ;
        RECT 1123.480 2726.390 1124.540 2726.530 ;
        RECT 1117.440 2713.890 1117.700 2714.210 ;
        RECT 1123.480 2713.870 1123.620 2726.390 ;
        RECT 1124.340 2717.290 1124.600 2717.610 ;
        RECT 1123.420 2713.550 1123.680 2713.870 ;
        RECT 1124.400 2700.000 1124.540 2717.290 ;
        RECT 1130.840 2714.890 1130.980 2794.275 ;
        RECT 1131.230 2793.595 1131.510 2793.965 ;
        RECT 1130.780 2714.570 1131.040 2714.890 ;
        RECT 1131.300 2714.550 1131.440 2793.595 ;
        RECT 1135.900 2792.750 1136.040 2794.275 ;
        RECT 1135.840 2792.430 1136.100 2792.750 ;
        RECT 1138.200 2718.290 1138.340 2794.275 ;
        RECT 1140.040 2793.770 1140.180 2794.275 ;
        RECT 1139.980 2793.450 1140.240 2793.770 ;
        RECT 1145.100 2718.630 1145.240 2794.275 ;
        RECT 1147.400 2792.070 1147.540 2794.275 ;
        RECT 1147.340 2791.750 1147.600 2792.070 ;
        RECT 1145.040 2718.310 1145.300 2718.630 ;
        RECT 1138.140 2717.970 1138.400 2718.290 ;
        RECT 1152.000 2717.950 1152.140 2794.275 ;
        RECT 1152.390 2791.555 1152.670 2791.925 ;
        RECT 1152.400 2791.410 1152.660 2791.555 ;
        RECT 1151.940 2717.630 1152.200 2717.950 ;
        RECT 1158.900 2717.610 1159.040 2794.275 ;
        RECT 1159.290 2793.595 1159.570 2793.965 ;
        RECT 1159.360 2793.430 1159.500 2793.595 ;
        RECT 1159.300 2793.110 1159.560 2793.430 ;
        RECT 1159.290 2792.235 1159.570 2792.605 ;
        RECT 1159.360 2790.370 1159.500 2792.235 ;
        RECT 1159.300 2790.050 1159.560 2790.370 ;
        RECT 1158.840 2717.290 1159.100 2717.610 ;
        RECT 1134.920 2716.950 1135.180 2717.270 ;
        RECT 1131.240 2714.230 1131.500 2714.550 ;
        RECT 1134.980 2700.000 1135.120 2716.950 ;
        RECT 1165.340 2716.930 1165.480 2794.275 ;
        RECT 1165.730 2793.595 1166.010 2793.965 ;
        RECT 1165.800 2717.270 1165.940 2793.595 ;
        RECT 1166.260 2791.390 1166.400 2794.275 ;
        RECT 1166.200 2791.070 1166.460 2791.390 ;
        RECT 1165.740 2716.950 1166.000 2717.270 ;
        RECT 1155.620 2716.610 1155.880 2716.930 ;
        RECT 1165.280 2716.610 1165.540 2716.930 ;
        RECT 1145.500 2715.930 1145.760 2716.250 ;
        RECT 1145.560 2700.000 1145.700 2715.930 ;
        RECT 1155.680 2700.000 1155.820 2716.610 ;
        RECT 1172.700 2716.250 1172.840 2794.275 ;
        RECT 1173.090 2793.595 1173.370 2793.965 ;
        RECT 1173.160 2793.090 1173.300 2793.595 ;
        RECT 1173.100 2792.770 1173.360 2793.090 ;
        RECT 1179.600 2716.590 1179.740 2794.275 ;
        RECT 1179.990 2793.595 1180.270 2793.965 ;
        RECT 1180.060 2792.750 1180.200 2793.595 ;
        RECT 1180.000 2792.430 1180.260 2792.750 ;
        RECT 1176.320 2716.270 1176.580 2716.590 ;
        RECT 1179.540 2716.270 1179.800 2716.590 ;
        RECT 1172.640 2715.930 1172.900 2716.250 ;
        RECT 1166.200 2715.250 1166.460 2715.570 ;
        RECT 1166.260 2700.000 1166.400 2715.250 ;
        RECT 1176.380 2700.000 1176.520 2716.270 ;
        RECT 1186.500 2715.570 1186.640 2794.275 ;
        RECT 1186.890 2793.595 1187.170 2793.965 ;
        RECT 1186.900 2793.450 1187.160 2793.595 ;
        RECT 1193.790 2791.555 1194.070 2791.925 ;
        RECT 1193.860 2791.390 1194.000 2791.555 ;
        RECT 1193.800 2791.070 1194.060 2791.390 ;
        RECT 1193.330 2790.195 1193.610 2790.565 ;
        RECT 1193.400 2715.910 1193.540 2790.195 ;
        RECT 1186.900 2715.590 1187.160 2715.910 ;
        RECT 1193.340 2715.590 1193.600 2715.910 ;
        RECT 1186.440 2715.250 1186.700 2715.570 ;
        RECT 1186.960 2700.000 1187.100 2715.590 ;
        RECT 1200.300 2715.230 1200.440 2794.275 ;
        RECT 1300.980 2718.310 1301.240 2718.630 ;
        RECT 1290.400 2717.970 1290.660 2718.290 ;
        RECT 1197.020 2714.910 1197.280 2715.230 ;
        RECT 1200.240 2714.910 1200.500 2715.230 ;
        RECT 1197.080 2700.000 1197.220 2714.910 ;
        RECT 1280.280 2714.570 1280.540 2714.890 ;
        RECT 1269.700 2714.230 1269.960 2714.550 ;
        RECT 1249.000 2713.890 1249.260 2714.210 ;
        RECT 1228.300 2713.210 1228.560 2713.530 ;
        RECT 1207.600 2712.530 1207.860 2712.850 ;
        RECT 1207.660 2700.000 1207.800 2712.530 ;
        RECT 1217.720 2712.190 1217.980 2712.510 ;
        RECT 1217.780 2700.000 1217.920 2712.190 ;
        RECT 1228.360 2700.000 1228.500 2713.210 ;
        RECT 1238.880 2712.870 1239.140 2713.190 ;
        RECT 1238.940 2700.000 1239.080 2712.870 ;
        RECT 1249.060 2700.000 1249.200 2713.890 ;
        RECT 1259.580 2713.550 1259.840 2713.870 ;
        RECT 1259.640 2700.000 1259.780 2713.550 ;
        RECT 1269.760 2700.000 1269.900 2714.230 ;
        RECT 1280.340 2700.000 1280.480 2714.570 ;
        RECT 1290.460 2700.000 1290.600 2717.970 ;
        RECT 1301.040 2700.000 1301.180 2718.310 ;
        RECT 1311.100 2717.630 1311.360 2717.950 ;
        RECT 1311.160 2700.000 1311.300 2717.630 ;
        RECT 1321.680 2717.290 1321.940 2717.610 ;
        RECT 1321.740 2700.000 1321.880 2717.290 ;
        RECT 1332.260 2716.950 1332.520 2717.270 ;
        RECT 1332.320 2700.000 1332.460 2716.950 ;
        RECT 1342.380 2716.610 1342.640 2716.930 ;
        RECT 1342.440 2700.000 1342.580 2716.610 ;
        RECT 1363.080 2716.270 1363.340 2716.590 ;
        RECT 1352.960 2715.930 1353.220 2716.250 ;
        RECT 1353.020 2700.000 1353.160 2715.930 ;
        RECT 1363.140 2700.000 1363.280 2716.270 ;
        RECT 1383.780 2715.590 1384.040 2715.910 ;
        RECT 1373.660 2715.250 1373.920 2715.570 ;
        RECT 1373.720 2700.000 1373.860 2715.250 ;
        RECT 1383.840 2700.000 1383.980 2715.590 ;
        RECT 1394.360 2714.910 1394.620 2715.230 ;
        RECT 1394.420 2700.000 1394.560 2714.910 ;
        RECT 657.500 2699.940 657.790 2700.000 ;
        RECT 668.080 2699.940 668.370 2700.000 ;
        RECT 678.660 2699.940 678.950 2700.000 ;
        RECT 688.780 2699.940 689.070 2700.000 ;
        RECT 699.360 2699.940 699.650 2700.000 ;
        RECT 709.480 2699.940 709.770 2700.000 ;
        RECT 720.060 2699.940 720.350 2700.000 ;
        RECT 730.180 2699.940 730.470 2700.000 ;
        RECT 740.760 2699.940 741.050 2700.000 ;
        RECT 750.880 2699.940 751.170 2700.000 ;
        RECT 761.460 2699.940 761.750 2700.000 ;
        RECT 772.040 2699.940 772.330 2700.000 ;
        RECT 782.160 2699.940 782.450 2700.000 ;
        RECT 792.740 2699.940 793.030 2700.000 ;
        RECT 802.860 2699.940 803.150 2700.000 ;
        RECT 813.440 2699.940 813.730 2700.000 ;
        RECT 823.560 2699.940 823.850 2700.000 ;
        RECT 834.140 2699.940 834.430 2700.000 ;
        RECT 844.260 2699.940 844.550 2700.000 ;
        RECT 854.840 2699.940 855.130 2700.000 ;
        RECT 865.420 2699.940 865.710 2700.000 ;
        RECT 875.540 2699.940 875.830 2700.000 ;
        RECT 886.120 2699.940 886.410 2700.000 ;
        RECT 896.240 2699.940 896.530 2700.000 ;
        RECT 906.820 2699.940 907.110 2700.000 ;
        RECT 916.940 2699.940 917.230 2700.000 ;
        RECT 927.520 2699.940 927.810 2700.000 ;
        RECT 937.640 2699.940 937.930 2700.000 ;
        RECT 948.220 2699.940 948.510 2700.000 ;
        RECT 958.800 2699.940 959.090 2700.000 ;
        RECT 968.920 2699.940 969.210 2700.000 ;
        RECT 979.500 2699.940 979.790 2700.000 ;
        RECT 989.620 2699.940 989.910 2700.000 ;
        RECT 1000.200 2699.940 1000.490 2700.000 ;
        RECT 1010.320 2699.940 1010.610 2700.000 ;
        RECT 1020.900 2699.940 1021.190 2700.000 ;
        RECT 1031.020 2699.940 1031.310 2700.000 ;
        RECT 1041.600 2699.940 1041.890 2700.000 ;
        RECT 1052.180 2699.940 1052.470 2700.000 ;
        RECT 1062.300 2699.940 1062.590 2700.000 ;
        RECT 1072.880 2699.940 1073.170 2700.000 ;
        RECT 1083.000 2699.940 1083.290 2700.000 ;
        RECT 1093.580 2699.940 1093.870 2700.000 ;
        RECT 1103.700 2699.940 1103.990 2700.000 ;
        RECT 1114.280 2699.940 1114.570 2700.000 ;
        RECT 1124.400 2699.940 1124.690 2700.000 ;
        RECT 1134.980 2699.940 1135.270 2700.000 ;
        RECT 1145.560 2699.940 1145.850 2700.000 ;
        RECT 1155.680 2699.940 1155.970 2700.000 ;
        RECT 1166.260 2699.940 1166.550 2700.000 ;
        RECT 1176.380 2699.940 1176.670 2700.000 ;
        RECT 1186.960 2699.940 1187.250 2700.000 ;
        RECT 1197.080 2699.940 1197.370 2700.000 ;
        RECT 1207.660 2699.940 1207.950 2700.000 ;
        RECT 1217.780 2699.940 1218.070 2700.000 ;
        RECT 1228.360 2699.940 1228.650 2700.000 ;
        RECT 1238.940 2699.940 1239.230 2700.000 ;
        RECT 1249.060 2699.940 1249.350 2700.000 ;
        RECT 1259.640 2699.940 1259.930 2700.000 ;
        RECT 1269.760 2699.940 1270.050 2700.000 ;
        RECT 1280.340 2699.940 1280.630 2700.000 ;
        RECT 1290.460 2699.940 1290.750 2700.000 ;
        RECT 1301.040 2699.940 1301.330 2700.000 ;
        RECT 1311.160 2699.940 1311.450 2700.000 ;
        RECT 1321.740 2699.940 1322.030 2700.000 ;
        RECT 1332.320 2699.940 1332.610 2700.000 ;
        RECT 1342.440 2699.940 1342.730 2700.000 ;
        RECT 1353.020 2699.940 1353.310 2700.000 ;
        RECT 1363.140 2699.940 1363.430 2700.000 ;
        RECT 1373.720 2699.940 1374.010 2700.000 ;
        RECT 1383.840 2699.940 1384.130 2700.000 ;
        RECT 1394.420 2699.940 1394.710 2700.000 ;
        RECT 647.390 2696.000 647.670 2699.870 ;
        RECT 657.510 2696.000 657.790 2699.940 ;
        RECT 668.090 2696.000 668.370 2699.940 ;
        RECT 678.670 2696.000 678.950 2699.940 ;
        RECT 688.790 2696.000 689.070 2699.940 ;
        RECT 699.370 2696.000 699.650 2699.940 ;
        RECT 709.490 2696.000 709.770 2699.940 ;
        RECT 720.070 2696.000 720.350 2699.940 ;
        RECT 730.190 2696.000 730.470 2699.940 ;
        RECT 740.770 2696.000 741.050 2699.940 ;
        RECT 750.890 2696.000 751.170 2699.940 ;
        RECT 761.470 2696.000 761.750 2699.940 ;
        RECT 772.050 2696.000 772.330 2699.940 ;
        RECT 782.170 2696.000 782.450 2699.940 ;
        RECT 792.750 2696.000 793.030 2699.940 ;
        RECT 802.870 2696.000 803.150 2699.940 ;
        RECT 813.450 2696.000 813.730 2699.940 ;
        RECT 823.570 2696.000 823.850 2699.940 ;
        RECT 834.150 2696.000 834.430 2699.940 ;
        RECT 844.270 2696.000 844.550 2699.940 ;
        RECT 854.850 2696.000 855.130 2699.940 ;
        RECT 865.430 2696.000 865.710 2699.940 ;
        RECT 875.550 2696.000 875.830 2699.940 ;
        RECT 886.130 2696.000 886.410 2699.940 ;
        RECT 896.250 2696.000 896.530 2699.940 ;
        RECT 906.830 2696.000 907.110 2699.940 ;
        RECT 916.950 2696.000 917.230 2699.940 ;
        RECT 927.530 2696.000 927.810 2699.940 ;
        RECT 937.650 2696.000 937.930 2699.940 ;
        RECT 948.230 2696.000 948.510 2699.940 ;
        RECT 958.810 2696.000 959.090 2699.940 ;
        RECT 968.930 2696.000 969.210 2699.940 ;
        RECT 979.510 2696.000 979.790 2699.940 ;
        RECT 989.630 2696.000 989.910 2699.940 ;
        RECT 1000.210 2696.000 1000.490 2699.940 ;
        RECT 1010.330 2696.000 1010.610 2699.940 ;
        RECT 1020.910 2696.000 1021.190 2699.940 ;
        RECT 1031.030 2696.000 1031.310 2699.940 ;
        RECT 1041.610 2696.000 1041.890 2699.940 ;
        RECT 1052.190 2696.000 1052.470 2699.940 ;
        RECT 1062.310 2696.000 1062.590 2699.940 ;
        RECT 1072.890 2696.000 1073.170 2699.940 ;
        RECT 1083.010 2696.000 1083.290 2699.940 ;
        RECT 1093.590 2696.000 1093.870 2699.940 ;
        RECT 1103.710 2696.000 1103.990 2699.940 ;
        RECT 1114.290 2696.000 1114.570 2699.940 ;
        RECT 1124.410 2696.000 1124.690 2699.940 ;
        RECT 1134.990 2696.000 1135.270 2699.940 ;
        RECT 1145.570 2696.000 1145.850 2699.940 ;
        RECT 1155.690 2696.000 1155.970 2699.940 ;
        RECT 1166.270 2696.000 1166.550 2699.940 ;
        RECT 1176.390 2696.000 1176.670 2699.940 ;
        RECT 1186.970 2696.000 1187.250 2699.940 ;
        RECT 1197.090 2696.000 1197.370 2699.940 ;
        RECT 1207.670 2696.000 1207.950 2699.940 ;
        RECT 1217.790 2696.000 1218.070 2699.940 ;
        RECT 1228.370 2696.000 1228.650 2699.940 ;
        RECT 1238.950 2696.000 1239.230 2699.940 ;
        RECT 1249.070 2696.000 1249.350 2699.940 ;
        RECT 1259.650 2696.000 1259.930 2699.940 ;
        RECT 1269.770 2696.000 1270.050 2699.940 ;
        RECT 1280.350 2696.000 1280.630 2699.940 ;
        RECT 1290.470 2696.000 1290.750 2699.940 ;
        RECT 1301.050 2696.000 1301.330 2699.940 ;
        RECT 1311.170 2696.000 1311.450 2699.940 ;
        RECT 1321.750 2696.000 1322.030 2699.940 ;
        RECT 1332.330 2696.000 1332.610 2699.940 ;
        RECT 1342.450 2696.000 1342.730 2699.940 ;
        RECT 1353.030 2696.000 1353.310 2699.940 ;
        RECT 1363.150 2696.000 1363.430 2699.940 ;
        RECT 1373.730 2696.000 1374.010 2699.940 ;
        RECT 1383.850 2696.000 1384.130 2699.940 ;
        RECT 1394.430 2696.000 1394.710 2699.940 ;
      LAYER met2 ;
        RECT 300.090 2695.720 304.870 2696.000 ;
        RECT 305.710 2695.720 314.990 2696.000 ;
        RECT 315.830 2695.720 325.570 2696.000 ;
        RECT 326.410 2695.720 335.690 2696.000 ;
        RECT 336.530 2695.720 346.270 2696.000 ;
        RECT 347.110 2695.720 356.390 2696.000 ;
        RECT 357.230 2695.720 366.970 2696.000 ;
        RECT 367.810 2695.720 377.090 2696.000 ;
        RECT 377.930 2695.720 387.670 2696.000 ;
        RECT 388.510 2695.720 398.250 2696.000 ;
        RECT 399.090 2695.720 408.370 2696.000 ;
        RECT 409.210 2695.720 418.950 2696.000 ;
        RECT 419.790 2695.720 429.070 2696.000 ;
        RECT 429.910 2695.720 439.650 2696.000 ;
        RECT 440.490 2695.720 449.770 2696.000 ;
        RECT 450.610 2695.720 460.350 2696.000 ;
        RECT 461.190 2695.720 470.470 2696.000 ;
        RECT 471.310 2695.720 481.050 2696.000 ;
        RECT 481.890 2695.720 491.630 2696.000 ;
        RECT 492.470 2695.720 501.750 2696.000 ;
        RECT 502.590 2695.720 512.330 2696.000 ;
        RECT 513.170 2695.720 522.450 2696.000 ;
        RECT 523.290 2695.720 533.030 2696.000 ;
        RECT 533.870 2695.720 543.150 2696.000 ;
        RECT 543.990 2695.720 553.730 2696.000 ;
        RECT 554.570 2695.720 563.850 2696.000 ;
        RECT 564.690 2695.720 574.430 2696.000 ;
        RECT 575.270 2695.720 585.010 2696.000 ;
        RECT 585.850 2695.720 595.130 2696.000 ;
        RECT 595.970 2695.720 605.710 2696.000 ;
        RECT 606.550 2695.720 615.830 2696.000 ;
        RECT 616.670 2695.720 626.410 2696.000 ;
        RECT 627.250 2695.720 636.530 2696.000 ;
        RECT 637.370 2695.720 647.110 2696.000 ;
        RECT 647.950 2695.720 657.230 2696.000 ;
        RECT 658.070 2695.720 667.810 2696.000 ;
        RECT 668.650 2695.720 678.390 2696.000 ;
        RECT 679.230 2695.720 688.510 2696.000 ;
        RECT 689.350 2695.720 699.090 2696.000 ;
        RECT 699.930 2695.720 709.210 2696.000 ;
        RECT 710.050 2695.720 719.790 2696.000 ;
        RECT 720.630 2695.720 729.910 2696.000 ;
        RECT 730.750 2695.720 740.490 2696.000 ;
        RECT 741.330 2695.720 750.610 2696.000 ;
        RECT 751.450 2695.720 761.190 2696.000 ;
        RECT 762.030 2695.720 771.770 2696.000 ;
        RECT 772.610 2695.720 781.890 2696.000 ;
        RECT 782.730 2695.720 792.470 2696.000 ;
        RECT 793.310 2695.720 802.590 2696.000 ;
        RECT 803.430 2695.720 813.170 2696.000 ;
        RECT 814.010 2695.720 823.290 2696.000 ;
        RECT 824.130 2695.720 833.870 2696.000 ;
        RECT 834.710 2695.720 843.990 2696.000 ;
        RECT 844.830 2695.720 854.570 2696.000 ;
        RECT 855.410 2695.720 865.150 2696.000 ;
        RECT 865.990 2695.720 875.270 2696.000 ;
        RECT 876.110 2695.720 885.850 2696.000 ;
        RECT 886.690 2695.720 895.970 2696.000 ;
        RECT 896.810 2695.720 906.550 2696.000 ;
        RECT 907.390 2695.720 916.670 2696.000 ;
        RECT 917.510 2695.720 927.250 2696.000 ;
        RECT 928.090 2695.720 937.370 2696.000 ;
        RECT 938.210 2695.720 947.950 2696.000 ;
        RECT 948.790 2695.720 958.530 2696.000 ;
        RECT 959.370 2695.720 968.650 2696.000 ;
        RECT 969.490 2695.720 979.230 2696.000 ;
        RECT 980.070 2695.720 989.350 2696.000 ;
        RECT 990.190 2695.720 999.930 2696.000 ;
        RECT 1000.770 2695.720 1010.050 2696.000 ;
        RECT 1010.890 2695.720 1020.630 2696.000 ;
        RECT 1021.470 2695.720 1030.750 2696.000 ;
        RECT 1031.590 2695.720 1041.330 2696.000 ;
        RECT 1042.170 2695.720 1051.910 2696.000 ;
        RECT 1052.750 2695.720 1062.030 2696.000 ;
        RECT 1062.870 2695.720 1072.610 2696.000 ;
        RECT 1073.450 2695.720 1082.730 2696.000 ;
        RECT 1083.570 2695.720 1093.310 2696.000 ;
        RECT 1094.150 2695.720 1103.430 2696.000 ;
        RECT 1104.270 2695.720 1114.010 2696.000 ;
        RECT 1114.850 2695.720 1124.130 2696.000 ;
        RECT 1124.970 2695.720 1134.710 2696.000 ;
        RECT 1135.550 2695.720 1145.290 2696.000 ;
        RECT 1146.130 2695.720 1155.410 2696.000 ;
        RECT 1156.250 2695.720 1165.990 2696.000 ;
        RECT 1166.830 2695.720 1176.110 2696.000 ;
        RECT 1176.950 2695.720 1186.690 2696.000 ;
        RECT 1187.530 2695.720 1196.810 2696.000 ;
        RECT 1197.650 2695.720 1207.390 2696.000 ;
        RECT 1208.230 2695.720 1217.510 2696.000 ;
        RECT 1218.350 2695.720 1228.090 2696.000 ;
        RECT 1228.930 2695.720 1238.670 2696.000 ;
        RECT 1239.510 2695.720 1248.790 2696.000 ;
        RECT 1249.630 2695.720 1259.370 2696.000 ;
        RECT 1260.210 2695.720 1269.490 2696.000 ;
        RECT 1270.330 2695.720 1280.070 2696.000 ;
        RECT 1280.910 2695.720 1290.190 2696.000 ;
        RECT 1291.030 2695.720 1300.770 2696.000 ;
        RECT 1301.610 2695.720 1310.890 2696.000 ;
        RECT 1311.730 2695.720 1321.470 2696.000 ;
        RECT 1322.310 2695.720 1332.050 2696.000 ;
        RECT 1332.890 2695.720 1342.170 2696.000 ;
        RECT 1343.010 2695.720 1352.750 2696.000 ;
        RECT 1353.590 2695.720 1362.870 2696.000 ;
        RECT 1363.710 2695.720 1373.450 2696.000 ;
        RECT 1374.290 2695.720 1383.570 2696.000 ;
        RECT 1384.410 2695.720 1394.150 2696.000 ;
        RECT 1394.990 2695.720 1395.630 2696.000 ;
        RECT 300.090 1604.280 1395.630 2695.720 ;
      LAYER met2 ;
        RECT 1395.800 1604.530 1395.940 2901.230 ;
        RECT 1407.690 2894.915 1407.970 2895.285 ;
        RECT 1407.230 2204.715 1407.510 2205.085 ;
        RECT 1407.300 2201.490 1407.440 2204.715 ;
        RECT 1407.240 2201.170 1407.500 2201.490 ;
        RECT 1407.230 2149.635 1407.510 2150.005 ;
        RECT 1407.300 2146.070 1407.440 2149.635 ;
        RECT 1407.240 2145.750 1407.500 2146.070 ;
        RECT 1407.760 1649.410 1407.900 2894.915 ;
        RECT 1411.370 2697.035 1411.650 2697.405 ;
        RECT 1411.440 2691.770 1411.580 2697.035 ;
        RECT 1414.130 2692.275 1414.410 2692.645 ;
        RECT 1411.380 2691.450 1411.640 2691.770 ;
        RECT 1414.200 2691.430 1414.340 2692.275 ;
        RECT 1414.140 2691.110 1414.400 2691.430 ;
        RECT 1414.130 2686.835 1414.410 2687.205 ;
        RECT 1414.200 2684.290 1414.340 2686.835 ;
        RECT 1414.140 2683.970 1414.400 2684.290 ;
        RECT 1414.130 2682.075 1414.410 2682.445 ;
        RECT 1414.200 2677.490 1414.340 2682.075 ;
        RECT 1414.140 2677.170 1414.400 2677.490 ;
        RECT 1408.610 2676.635 1408.890 2677.005 ;
        RECT 1408.680 2671.030 1408.820 2676.635 ;
        RECT 1410.450 2671.875 1410.730 2672.245 ;
        RECT 1408.620 2670.710 1408.880 2671.030 ;
        RECT 1410.520 2670.690 1410.660 2671.875 ;
        RECT 1410.460 2670.370 1410.720 2670.690 ;
        RECT 1410.450 2667.115 1410.730 2667.485 ;
        RECT 1410.520 2663.890 1410.660 2667.115 ;
        RECT 1410.460 2663.570 1410.720 2663.890 ;
        RECT 1411.370 2661.675 1411.650 2662.045 ;
        RECT 1411.440 2657.090 1411.580 2661.675 ;
        RECT 1411.380 2656.770 1411.640 2657.090 ;
        RECT 1414.130 2656.915 1414.410 2657.285 ;
        RECT 1414.200 2656.750 1414.340 2656.915 ;
        RECT 1414.140 2656.430 1414.400 2656.750 ;
        RECT 1414.130 2651.475 1414.410 2651.845 ;
        RECT 1414.200 2649.950 1414.340 2651.475 ;
        RECT 1414.140 2649.630 1414.400 2649.950 ;
        RECT 1414.130 2646.715 1414.410 2647.085 ;
        RECT 1414.200 2643.150 1414.340 2646.715 ;
        RECT 1414.140 2642.830 1414.400 2643.150 ;
        RECT 1411.370 2641.275 1411.650 2641.645 ;
        RECT 1411.440 2636.010 1411.580 2641.275 ;
        RECT 1414.130 2636.515 1414.410 2636.885 ;
        RECT 1414.200 2636.350 1414.340 2636.515 ;
        RECT 1414.140 2636.030 1414.400 2636.350 ;
        RECT 1411.380 2635.690 1411.640 2636.010 ;
        RECT 1409.530 2631.755 1409.810 2632.125 ;
        RECT 1409.600 2629.210 1409.740 2631.755 ;
        RECT 1409.540 2628.890 1409.800 2629.210 ;
        RECT 1414.130 2626.315 1414.410 2626.685 ;
        RECT 1414.200 2622.410 1414.340 2626.315 ;
        RECT 1414.140 2622.090 1414.400 2622.410 ;
        RECT 1411.830 2621.555 1412.110 2621.925 ;
        RECT 1411.900 2615.270 1412.040 2621.555 ;
        RECT 1414.130 2616.115 1414.410 2616.485 ;
        RECT 1414.200 2615.610 1414.340 2616.115 ;
        RECT 1414.140 2615.290 1414.400 2615.610 ;
        RECT 1411.840 2614.950 1412.100 2615.270 ;
        RECT 1414.130 2611.355 1414.410 2611.725 ;
        RECT 1414.200 2608.470 1414.340 2611.355 ;
        RECT 1414.140 2608.150 1414.400 2608.470 ;
        RECT 1417.810 2605.915 1418.090 2606.285 ;
        RECT 1414.140 2601.525 1414.400 2601.670 ;
        RECT 1414.130 2601.155 1414.410 2601.525 ;
        RECT 1408.610 2596.395 1408.890 2596.765 ;
        RECT 1408.680 2595.550 1408.820 2596.395 ;
        RECT 1408.620 2595.230 1408.880 2595.550 ;
        RECT 1410.450 2590.955 1410.730 2591.325 ;
        RECT 1410.520 2587.730 1410.660 2590.955 ;
        RECT 1410.460 2587.410 1410.720 2587.730 ;
        RECT 1411.370 2586.195 1411.650 2586.565 ;
        RECT 1411.440 2581.270 1411.580 2586.195 ;
        RECT 1411.380 2580.950 1411.640 2581.270 ;
        RECT 1414.130 2580.755 1414.410 2581.125 ;
        RECT 1414.140 2580.610 1414.400 2580.755 ;
        RECT 1414.130 2575.995 1414.410 2576.365 ;
        RECT 1414.200 2574.130 1414.340 2575.995 ;
        RECT 1414.140 2573.810 1414.400 2574.130 ;
        RECT 1411.370 2571.235 1411.650 2571.605 ;
        RECT 1411.440 2566.990 1411.580 2571.235 ;
        RECT 1411.380 2566.670 1411.640 2566.990 ;
        RECT 1413.670 2565.795 1413.950 2566.165 ;
        RECT 1413.740 2560.530 1413.880 2565.795 ;
        RECT 1414.130 2561.035 1414.410 2561.405 ;
        RECT 1413.680 2560.210 1413.940 2560.530 ;
        RECT 1414.200 2560.190 1414.340 2561.035 ;
        RECT 1414.140 2559.870 1414.400 2560.190 ;
        RECT 1408.610 2555.595 1408.890 2555.965 ;
        RECT 1408.680 2553.390 1408.820 2555.595 ;
        RECT 1408.620 2553.070 1408.880 2553.390 ;
        RECT 1411.370 2550.835 1411.650 2551.205 ;
        RECT 1411.440 2546.590 1411.580 2550.835 ;
        RECT 1411.380 2546.270 1411.640 2546.590 ;
        RECT 1412.750 2545.395 1413.030 2545.765 ;
        RECT 1412.820 2539.790 1412.960 2545.395 ;
        RECT 1414.130 2540.635 1414.410 2541.005 ;
        RECT 1412.760 2539.470 1413.020 2539.790 ;
        RECT 1414.200 2539.450 1414.340 2540.635 ;
        RECT 1414.140 2539.130 1414.400 2539.450 ;
        RECT 1410.450 2535.875 1410.730 2536.245 ;
        RECT 1410.520 2532.650 1410.660 2535.875 ;
        RECT 1410.460 2532.330 1410.720 2532.650 ;
        RECT 1413.670 2530.435 1413.950 2530.805 ;
        RECT 1413.740 2525.850 1413.880 2530.435 ;
        RECT 1414.140 2526.045 1414.400 2526.190 ;
        RECT 1413.680 2525.530 1413.940 2525.850 ;
        RECT 1414.130 2525.675 1414.410 2526.045 ;
        RECT 1414.130 2520.235 1414.410 2520.605 ;
        RECT 1414.200 2518.710 1414.340 2520.235 ;
        RECT 1414.140 2518.390 1414.400 2518.710 ;
        RECT 1414.130 2515.475 1414.410 2515.845 ;
        RECT 1414.200 2511.910 1414.340 2515.475 ;
        RECT 1414.140 2511.590 1414.400 2511.910 ;
        RECT 1411.370 2510.035 1411.650 2510.405 ;
        RECT 1411.440 2505.110 1411.580 2510.035 ;
        RECT 1414.130 2505.275 1414.410 2505.645 ;
        RECT 1414.140 2505.130 1414.400 2505.275 ;
        RECT 1411.380 2504.790 1411.640 2505.110 ;
        RECT 1414.130 2495.075 1414.410 2495.445 ;
        RECT 1414.200 2491.170 1414.340 2495.075 ;
        RECT 1414.140 2490.850 1414.400 2491.170 ;
        RECT 1414.130 2484.875 1414.410 2485.245 ;
        RECT 1414.200 2484.370 1414.340 2484.875 ;
        RECT 1414.140 2484.050 1414.400 2484.370 ;
        RECT 1409.530 2480.115 1409.810 2480.485 ;
        RECT 1409.600 2477.570 1409.740 2480.115 ;
        RECT 1409.540 2477.250 1409.800 2477.570 ;
        RECT 1414.130 2475.355 1414.410 2475.725 ;
        RECT 1414.200 2470.430 1414.340 2475.355 ;
        RECT 1411.830 2469.915 1412.110 2470.285 ;
        RECT 1414.140 2470.110 1414.400 2470.430 ;
        RECT 1411.900 2463.630 1412.040 2469.915 ;
        RECT 1414.130 2465.155 1414.410 2465.525 ;
        RECT 1414.200 2463.970 1414.340 2465.155 ;
        RECT 1414.140 2463.650 1414.400 2463.970 ;
        RECT 1411.840 2463.310 1412.100 2463.630 ;
        RECT 1414.130 2459.715 1414.410 2460.085 ;
        RECT 1414.200 2456.830 1414.340 2459.715 ;
        RECT 1414.140 2456.510 1414.400 2456.830 ;
        RECT 1411.370 2454.955 1411.650 2455.325 ;
        RECT 1411.440 2449.690 1411.580 2454.955 ;
        RECT 1414.140 2449.885 1414.400 2450.030 ;
        RECT 1411.380 2449.370 1411.640 2449.690 ;
        RECT 1414.130 2449.515 1414.410 2449.885 ;
        RECT 1411.370 2444.755 1411.650 2445.125 ;
        RECT 1411.440 2442.890 1411.580 2444.755 ;
        RECT 1411.380 2442.570 1411.640 2442.890 ;
        RECT 1414.130 2439.995 1414.410 2440.365 ;
        RECT 1414.200 2436.090 1414.340 2439.995 ;
        RECT 1414.140 2435.770 1414.400 2436.090 ;
        RECT 1411.370 2434.555 1411.650 2434.925 ;
        RECT 1411.440 2429.290 1411.580 2434.555 ;
        RECT 1414.130 2429.795 1414.410 2430.165 ;
        RECT 1414.200 2429.630 1414.340 2429.795 ;
        RECT 1414.140 2429.310 1414.400 2429.630 ;
        RECT 1411.380 2428.970 1411.640 2429.290 ;
        RECT 1408.610 2424.355 1408.890 2424.725 ;
        RECT 1408.680 2422.150 1408.820 2424.355 ;
        RECT 1408.620 2421.830 1408.880 2422.150 ;
        RECT 1411.370 2419.595 1411.650 2419.965 ;
        RECT 1411.440 2415.350 1411.580 2419.595 ;
        RECT 1411.380 2415.030 1411.640 2415.350 ;
        RECT 1412.750 2414.155 1413.030 2414.525 ;
        RECT 1412.820 2408.550 1412.960 2414.155 ;
        RECT 1414.130 2409.395 1414.410 2409.765 ;
        RECT 1414.200 2408.890 1414.340 2409.395 ;
        RECT 1414.140 2408.570 1414.400 2408.890 ;
        RECT 1412.760 2408.230 1413.020 2408.550 ;
        RECT 1410.450 2404.635 1410.730 2405.005 ;
        RECT 1410.520 2401.410 1410.660 2404.635 ;
        RECT 1410.460 2401.090 1410.720 2401.410 ;
        RECT 1413.670 2399.195 1413.950 2399.565 ;
        RECT 1413.740 2394.610 1413.880 2399.195 ;
        RECT 1414.140 2394.805 1414.400 2394.950 ;
        RECT 1413.680 2394.290 1413.940 2394.610 ;
        RECT 1414.130 2394.435 1414.410 2394.805 ;
        RECT 1414.130 2388.995 1414.410 2389.365 ;
        RECT 1414.200 2387.810 1414.340 2388.995 ;
        RECT 1414.140 2387.490 1414.400 2387.810 ;
        RECT 1410.450 2384.235 1410.730 2384.605 ;
        RECT 1410.520 2380.670 1410.660 2384.235 ;
        RECT 1410.460 2380.350 1410.720 2380.670 ;
        RECT 1411.370 2378.795 1411.650 2379.165 ;
        RECT 1411.440 2373.870 1411.580 2378.795 ;
        RECT 1414.130 2374.035 1414.410 2374.405 ;
        RECT 1414.140 2373.890 1414.400 2374.035 ;
        RECT 1411.380 2373.550 1411.640 2373.870 ;
        RECT 1408.610 2369.275 1408.890 2369.645 ;
        RECT 1408.680 2367.070 1408.820 2369.275 ;
        RECT 1408.620 2366.750 1408.880 2367.070 ;
        RECT 1410.450 2363.835 1410.730 2364.205 ;
        RECT 1410.520 2360.270 1410.660 2363.835 ;
        RECT 1410.460 2359.950 1410.720 2360.270 ;
        RECT 1413.670 2359.075 1413.950 2359.445 ;
        RECT 1413.740 2353.130 1413.880 2359.075 ;
        RECT 1414.130 2353.635 1414.410 2354.005 ;
        RECT 1414.200 2353.470 1414.340 2353.635 ;
        RECT 1414.140 2353.150 1414.400 2353.470 ;
        RECT 1413.680 2352.810 1413.940 2353.130 ;
        RECT 1409.530 2348.875 1409.810 2349.245 ;
        RECT 1409.600 2346.330 1409.740 2348.875 ;
        RECT 1409.540 2346.010 1409.800 2346.330 ;
        RECT 1414.130 2344.115 1414.410 2344.485 ;
        RECT 1414.200 2339.530 1414.340 2344.115 ;
        RECT 1414.140 2339.210 1414.400 2339.530 ;
        RECT 1413.670 2338.675 1413.950 2339.045 ;
        RECT 1413.740 2332.730 1413.880 2338.675 ;
        RECT 1414.130 2333.915 1414.410 2334.285 ;
        RECT 1413.680 2332.410 1413.940 2332.730 ;
        RECT 1414.200 2332.390 1414.340 2333.915 ;
        RECT 1414.140 2332.070 1414.400 2332.390 ;
        RECT 1414.130 2328.475 1414.410 2328.845 ;
        RECT 1414.200 2325.590 1414.340 2328.475 ;
        RECT 1414.140 2325.270 1414.400 2325.590 ;
        RECT 1413.670 2323.715 1413.950 2324.085 ;
        RECT 1413.740 2319.130 1413.880 2323.715 ;
        RECT 1413.680 2318.810 1413.940 2319.130 ;
        RECT 1414.140 2318.645 1414.400 2318.790 ;
        RECT 1414.130 2318.275 1414.410 2318.645 ;
        RECT 1414.130 2313.515 1414.410 2313.885 ;
        RECT 1414.200 2311.990 1414.340 2313.515 ;
        RECT 1414.140 2311.670 1414.400 2311.990 ;
        RECT 1414.130 2308.755 1414.410 2309.125 ;
        RECT 1414.200 2304.850 1414.340 2308.755 ;
        RECT 1414.140 2304.530 1414.400 2304.850 ;
        RECT 1414.130 2303.315 1414.410 2303.685 ;
        RECT 1413.670 2298.555 1413.950 2298.925 ;
        RECT 1413.740 2298.390 1413.880 2298.555 ;
        RECT 1413.680 2298.070 1413.940 2298.390 ;
        RECT 1414.200 2298.050 1414.340 2303.315 ;
        RECT 1414.140 2297.730 1414.400 2298.050 ;
        RECT 1408.610 2293.115 1408.890 2293.485 ;
        RECT 1408.680 2291.250 1408.820 2293.115 ;
        RECT 1408.620 2290.930 1408.880 2291.250 ;
        RECT 1410.450 2288.355 1410.730 2288.725 ;
        RECT 1410.520 2284.110 1410.660 2288.355 ;
        RECT 1410.460 2283.790 1410.720 2284.110 ;
        RECT 1408.150 2282.915 1408.430 2283.285 ;
        RECT 1408.220 2277.650 1408.360 2282.915 ;
        RECT 1414.130 2278.155 1414.410 2278.525 ;
        RECT 1408.160 2277.330 1408.420 2277.650 ;
        RECT 1414.200 2277.310 1414.340 2278.155 ;
        RECT 1414.140 2276.990 1414.400 2277.310 ;
        RECT 1408.150 2273.395 1408.430 2273.765 ;
        RECT 1408.220 2106.970 1408.360 2273.395 ;
        RECT 1412.290 2267.955 1412.570 2268.325 ;
        RECT 1411.370 2263.195 1411.650 2263.565 ;
        RECT 1410.450 2232.595 1410.730 2232.965 ;
        RECT 1409.070 2227.835 1409.350 2228.205 ;
        RECT 1408.610 2212.875 1408.890 2213.245 ;
        RECT 1408.160 2106.650 1408.420 2106.970 ;
        RECT 1408.160 2105.970 1408.420 2106.290 ;
        RECT 1408.220 2065.490 1408.360 2105.970 ;
        RECT 1408.680 2069.230 1408.820 2212.875 ;
        RECT 1408.620 2068.910 1408.880 2069.230 ;
        RECT 1409.140 2068.210 1409.280 2227.835 ;
        RECT 1409.990 2222.395 1410.270 2222.765 ;
        RECT 1409.530 2217.635 1409.810 2218.005 ;
        RECT 1409.600 2068.890 1409.740 2217.635 ;
        RECT 1409.540 2068.570 1409.800 2068.890 ;
        RECT 1410.060 2068.550 1410.200 2222.395 ;
        RECT 1410.000 2068.230 1410.260 2068.550 ;
        RECT 1409.080 2067.890 1409.340 2068.210 ;
        RECT 1410.520 2067.870 1410.660 2232.595 ;
        RECT 1410.910 2202.675 1411.190 2203.045 ;
        RECT 1410.980 2202.170 1411.120 2202.675 ;
        RECT 1410.920 2201.850 1411.180 2202.170 ;
        RECT 1410.910 2197.235 1411.190 2197.605 ;
        RECT 1410.980 2194.690 1411.120 2197.235 ;
        RECT 1410.920 2194.370 1411.180 2194.690 ;
        RECT 1410.910 2187.035 1411.190 2187.405 ;
        RECT 1410.980 2183.130 1411.120 2187.035 ;
        RECT 1410.920 2182.810 1411.180 2183.130 ;
        RECT 1410.910 2182.275 1411.190 2182.645 ;
        RECT 1410.980 2181.090 1411.120 2182.275 ;
        RECT 1410.920 2180.770 1411.180 2181.090 ;
        RECT 1410.910 2177.515 1411.190 2177.885 ;
        RECT 1410.980 2173.950 1411.120 2177.515 ;
        RECT 1410.920 2173.630 1411.180 2173.950 ;
        RECT 1410.910 2172.075 1411.190 2172.445 ;
        RECT 1410.980 2166.810 1411.120 2172.075 ;
        RECT 1410.920 2166.490 1411.180 2166.810 ;
        RECT 1410.910 2161.875 1411.190 2162.245 ;
        RECT 1410.980 2069.910 1411.120 2161.875 ;
        RECT 1411.440 2157.970 1411.580 2263.195 ;
        RECT 1411.830 2257.755 1412.110 2258.125 ;
        RECT 1411.380 2157.650 1411.640 2157.970 ;
        RECT 1411.370 2157.115 1411.650 2157.485 ;
        RECT 1411.440 2153.550 1411.580 2157.115 ;
        RECT 1411.380 2153.230 1411.640 2153.550 ;
        RECT 1411.380 2152.550 1411.640 2152.870 ;
        RECT 1411.440 2147.285 1411.580 2152.550 ;
        RECT 1411.370 2146.915 1411.650 2147.285 ;
        RECT 1411.380 2145.410 1411.640 2145.730 ;
        RECT 1411.440 2142.525 1411.580 2145.410 ;
        RECT 1411.370 2142.155 1411.650 2142.525 ;
        RECT 1411.380 2138.610 1411.640 2138.930 ;
        RECT 1411.440 2137.085 1411.580 2138.610 ;
        RECT 1411.370 2136.715 1411.650 2137.085 ;
        RECT 1411.380 2135.890 1411.640 2136.210 ;
        RECT 1411.440 2135.045 1411.580 2135.890 ;
        RECT 1411.370 2134.675 1411.650 2135.045 ;
        RECT 1411.380 2131.810 1411.640 2132.130 ;
        RECT 1411.440 2126.885 1411.580 2131.810 ;
        RECT 1411.370 2126.515 1411.650 2126.885 ;
        RECT 1411.380 2125.010 1411.640 2125.330 ;
        RECT 1411.440 2122.125 1411.580 2125.010 ;
        RECT 1411.370 2121.755 1411.650 2122.125 ;
        RECT 1411.380 2117.870 1411.640 2118.190 ;
        RECT 1411.440 2117.365 1411.580 2117.870 ;
        RECT 1411.370 2116.995 1411.650 2117.365 ;
        RECT 1411.380 2116.170 1411.640 2116.490 ;
        RECT 1411.440 2111.925 1411.580 2116.170 ;
        RECT 1411.370 2111.555 1411.650 2111.925 ;
        RECT 1411.380 2111.070 1411.640 2111.390 ;
        RECT 1411.440 2107.165 1411.580 2111.070 ;
        RECT 1411.370 2106.795 1411.650 2107.165 ;
        RECT 1411.900 2106.370 1412.040 2257.755 ;
        RECT 1411.440 2106.230 1412.040 2106.370 ;
        RECT 1412.360 2106.290 1412.500 2267.955 ;
        RECT 1412.750 2252.995 1413.030 2253.365 ;
        RECT 1411.440 2088.950 1411.580 2106.230 ;
        RECT 1412.300 2105.970 1412.560 2106.290 ;
        RECT 1412.820 2105.690 1412.960 2252.995 ;
        RECT 1414.130 2248.235 1414.410 2248.605 ;
        RECT 1413.210 2242.795 1413.490 2243.165 ;
        RECT 1411.900 2105.550 1412.960 2105.690 ;
        RECT 1411.380 2088.630 1411.640 2088.950 ;
        RECT 1411.380 2087.950 1411.640 2088.270 ;
        RECT 1411.440 2077.390 1411.580 2087.950 ;
        RECT 1411.380 2077.070 1411.640 2077.390 ;
        RECT 1411.380 2076.390 1411.640 2076.710 ;
        RECT 1411.440 2071.805 1411.580 2076.390 ;
        RECT 1411.370 2071.435 1411.650 2071.805 ;
        RECT 1410.920 2069.590 1411.180 2069.910 ;
        RECT 1411.380 2069.250 1411.640 2069.570 ;
        RECT 1410.460 2067.550 1410.720 2067.870 ;
        RECT 1408.160 2065.170 1408.420 2065.490 ;
        RECT 1411.440 2065.150 1411.580 2069.250 ;
        RECT 1411.900 2066.850 1412.040 2105.550 ;
        RECT 1412.300 2104.950 1412.560 2105.270 ;
        RECT 1411.840 2066.530 1412.100 2066.850 ;
        RECT 1412.360 2066.510 1412.500 2104.950 ;
        RECT 1412.760 2097.130 1413.020 2097.450 ;
        RECT 1412.820 2091.525 1412.960 2097.130 ;
        RECT 1412.750 2091.155 1413.030 2091.525 ;
        RECT 1412.760 2088.630 1413.020 2088.950 ;
        RECT 1412.300 2066.190 1412.560 2066.510 ;
        RECT 1412.820 2066.170 1412.960 2088.630 ;
        RECT 1413.280 2067.190 1413.420 2242.795 ;
        RECT 1413.670 2238.035 1413.950 2238.405 ;
        RECT 1413.740 2067.530 1413.880 2238.035 ;
        RECT 1414.200 2105.270 1414.340 2248.235 ;
        RECT 1417.350 2192.475 1417.630 2192.845 ;
        RECT 1416.890 2167.315 1417.170 2167.685 ;
        RECT 1414.140 2104.950 1414.400 2105.270 ;
        RECT 1414.140 2104.270 1414.400 2104.590 ;
        RECT 1414.200 2101.725 1414.340 2104.270 ;
        RECT 1414.130 2101.355 1414.410 2101.725 ;
        RECT 1414.140 2096.965 1414.400 2097.110 ;
        RECT 1414.130 2096.595 1414.410 2096.965 ;
        RECT 1414.140 2090.330 1414.400 2090.650 ;
        RECT 1414.200 2086.765 1414.340 2090.330 ;
        RECT 1414.130 2086.395 1414.410 2086.765 ;
        RECT 1414.140 2083.530 1414.400 2083.850 ;
        RECT 1414.200 2082.005 1414.340 2083.530 ;
        RECT 1414.130 2081.635 1414.410 2082.005 ;
        RECT 1416.440 2080.810 1416.700 2081.130 ;
        RECT 1415.980 2080.470 1416.240 2080.790 ;
        RECT 1415.520 2080.130 1415.780 2080.450 ;
        RECT 1414.600 2077.070 1414.860 2077.390 ;
        RECT 1414.140 2076.730 1414.400 2077.050 ;
        RECT 1414.200 2076.565 1414.340 2076.730 ;
        RECT 1414.130 2076.195 1414.410 2076.565 ;
        RECT 1414.660 2075.770 1414.800 2077.070 ;
        RECT 1414.200 2075.630 1414.800 2075.770 ;
        RECT 1413.680 2067.210 1413.940 2067.530 ;
        RECT 1413.220 2066.870 1413.480 2067.190 ;
        RECT 1414.200 2066.930 1414.340 2075.630 ;
        RECT 1415.060 2073.670 1415.320 2073.990 ;
        RECT 1414.600 2073.330 1414.860 2073.650 ;
        RECT 1413.740 2066.790 1414.340 2066.930 ;
        RECT 1412.760 2065.850 1413.020 2066.170 ;
        RECT 1413.740 2065.830 1413.880 2066.790 ;
        RECT 1414.130 2066.250 1414.410 2066.365 ;
        RECT 1414.660 2066.250 1414.800 2073.330 ;
        RECT 1414.130 2066.110 1414.800 2066.250 ;
        RECT 1414.130 2065.995 1414.410 2066.110 ;
        RECT 1413.680 2065.510 1413.940 2065.830 ;
        RECT 1411.380 2064.830 1411.640 2065.150 ;
        RECT 1414.130 2061.235 1414.410 2061.605 ;
        RECT 1414.200 2060.810 1414.340 2061.235 ;
        RECT 1415.120 2060.810 1415.260 2073.670 ;
        RECT 1414.200 2060.670 1415.260 2060.810 ;
        RECT 1413.680 2055.990 1413.940 2056.310 ;
        RECT 1408.160 2055.310 1408.420 2055.630 ;
        RECT 1408.220 2034.970 1408.360 2055.310 ;
        RECT 1410.000 2054.970 1410.260 2055.290 ;
        RECT 1408.620 2048.850 1408.880 2049.170 ;
        RECT 1408.680 2046.645 1408.820 2048.850 ;
        RECT 1408.610 2046.275 1408.890 2046.645 ;
        RECT 1408.620 2042.050 1408.880 2042.370 ;
        RECT 1408.680 2041.205 1408.820 2042.050 ;
        RECT 1408.610 2040.835 1408.890 2041.205 ;
        RECT 1408.220 2034.830 1408.820 2034.970 ;
        RECT 1408.160 2019.950 1408.420 2020.270 ;
        RECT 1408.220 2016.045 1408.360 2019.950 ;
        RECT 1408.150 2015.675 1408.430 2016.045 ;
        RECT 1408.160 1990.885 1408.420 1991.030 ;
        RECT 1408.150 1990.515 1408.430 1990.885 ;
        RECT 1408.160 1986.125 1408.420 1986.270 ;
        RECT 1408.150 1985.755 1408.430 1986.125 ;
        RECT 1408.160 1982.210 1408.420 1982.530 ;
        RECT 1408.220 1980.685 1408.360 1982.210 ;
        RECT 1408.150 1980.315 1408.430 1980.685 ;
        RECT 1408.160 1978.810 1408.420 1979.130 ;
        RECT 1408.220 1975.925 1408.360 1978.810 ;
        RECT 1408.150 1975.555 1408.430 1975.925 ;
        RECT 1408.160 1971.670 1408.420 1971.990 ;
        RECT 1408.220 1970.485 1408.360 1971.670 ;
        RECT 1408.150 1970.115 1408.430 1970.485 ;
        RECT 1408.160 1965.890 1408.420 1966.210 ;
        RECT 1408.220 1965.725 1408.360 1965.890 ;
        RECT 1408.150 1965.355 1408.430 1965.725 ;
        RECT 1408.160 1960.285 1408.420 1960.430 ;
        RECT 1408.150 1959.915 1408.430 1960.285 ;
        RECT 1408.160 1958.070 1408.420 1958.390 ;
        RECT 1408.220 1955.525 1408.360 1958.070 ;
        RECT 1408.150 1955.155 1408.430 1955.525 ;
        RECT 1408.160 1950.765 1408.420 1950.910 ;
        RECT 1408.150 1950.395 1408.430 1950.765 ;
        RECT 1408.160 1945.325 1408.420 1945.470 ;
        RECT 1408.150 1944.955 1408.430 1945.325 ;
        RECT 1408.160 1941.410 1408.420 1941.730 ;
        RECT 1408.220 1940.565 1408.360 1941.410 ;
        RECT 1408.150 1940.195 1408.430 1940.565 ;
        RECT 1408.160 1935.290 1408.420 1935.610 ;
        RECT 1408.220 1935.125 1408.360 1935.290 ;
        RECT 1408.150 1934.755 1408.430 1935.125 ;
        RECT 1408.160 1930.365 1408.420 1930.510 ;
        RECT 1408.150 1929.995 1408.430 1930.365 ;
        RECT 1408.160 1926.110 1408.420 1926.430 ;
        RECT 1408.220 1925.605 1408.360 1926.110 ;
        RECT 1408.150 1925.235 1408.430 1925.605 ;
        RECT 1408.160 1920.165 1408.420 1920.310 ;
        RECT 1408.150 1919.795 1408.430 1920.165 ;
        RECT 1408.160 1916.250 1408.420 1916.570 ;
        RECT 1408.220 1915.405 1408.360 1916.250 ;
        RECT 1408.150 1915.035 1408.430 1915.405 ;
        RECT 1408.160 1910.470 1408.420 1910.790 ;
        RECT 1408.220 1909.965 1408.360 1910.470 ;
        RECT 1408.150 1909.595 1408.430 1909.965 ;
        RECT 1408.160 1904.010 1408.420 1904.330 ;
        RECT 1408.220 1899.765 1408.360 1904.010 ;
        RECT 1408.150 1899.395 1408.430 1899.765 ;
        RECT 1408.160 1897.210 1408.420 1897.530 ;
        RECT 1408.220 1895.005 1408.360 1897.210 ;
        RECT 1408.150 1894.635 1408.430 1895.005 ;
        RECT 1408.160 1890.410 1408.420 1890.730 ;
        RECT 1408.220 1890.245 1408.360 1890.410 ;
        RECT 1408.150 1889.875 1408.430 1890.245 ;
        RECT 1408.160 1883.270 1408.420 1883.590 ;
        RECT 1408.220 1880.045 1408.360 1883.270 ;
        RECT 1408.150 1879.675 1408.430 1880.045 ;
        RECT 1408.160 1876.470 1408.420 1876.790 ;
        RECT 1408.220 1874.605 1408.360 1876.470 ;
        RECT 1408.150 1874.235 1408.430 1874.605 ;
        RECT 1408.150 1869.475 1408.430 1869.845 ;
        RECT 1408.220 1865.910 1408.360 1869.475 ;
        RECT 1408.160 1865.590 1408.420 1865.910 ;
        RECT 1408.160 1859.645 1408.420 1859.790 ;
        RECT 1408.150 1859.275 1408.430 1859.645 ;
        RECT 1408.160 1854.885 1408.420 1855.030 ;
        RECT 1408.150 1854.515 1408.430 1854.885 ;
        RECT 1408.160 1848.930 1408.420 1849.250 ;
        RECT 1408.220 1844.685 1408.360 1848.930 ;
        RECT 1408.150 1844.315 1408.430 1844.685 ;
        RECT 1408.160 1842.130 1408.420 1842.450 ;
        RECT 1408.220 1839.245 1408.360 1842.130 ;
        RECT 1408.150 1838.875 1408.430 1839.245 ;
        RECT 1408.160 1828.190 1408.420 1828.510 ;
        RECT 1408.220 1824.285 1408.360 1828.190 ;
        RECT 1408.150 1823.915 1408.430 1824.285 ;
        RECT 1408.160 1821.390 1408.420 1821.710 ;
        RECT 1408.220 1819.525 1408.360 1821.390 ;
        RECT 1408.150 1819.155 1408.430 1819.525 ;
        RECT 1408.160 1814.250 1408.420 1814.570 ;
        RECT 1408.220 1814.085 1408.360 1814.250 ;
        RECT 1408.150 1813.715 1408.430 1814.085 ;
        RECT 1408.160 1807.450 1408.420 1807.770 ;
        RECT 1408.220 1803.885 1408.360 1807.450 ;
        RECT 1408.150 1803.515 1408.430 1803.885 ;
        RECT 1408.160 1800.650 1408.420 1800.970 ;
        RECT 1408.220 1799.125 1408.360 1800.650 ;
        RECT 1408.150 1798.755 1408.430 1799.125 ;
        RECT 1408.160 1793.510 1408.420 1793.830 ;
        RECT 1408.220 1788.925 1408.360 1793.510 ;
        RECT 1408.150 1788.555 1408.430 1788.925 ;
        RECT 1408.160 1759.005 1408.420 1759.150 ;
        RECT 1408.150 1758.635 1408.430 1759.005 ;
        RECT 1408.160 1754.410 1408.420 1754.730 ;
        RECT 1408.220 1753.565 1408.360 1754.410 ;
        RECT 1408.150 1753.195 1408.430 1753.565 ;
        RECT 1408.160 1751.350 1408.420 1751.670 ;
        RECT 1408.220 1748.805 1408.360 1751.350 ;
        RECT 1408.150 1748.435 1408.430 1748.805 ;
        RECT 1408.160 1745.230 1408.420 1745.550 ;
        RECT 1408.220 1743.365 1408.360 1745.230 ;
        RECT 1408.150 1742.995 1408.430 1743.365 ;
        RECT 1408.160 1738.605 1408.420 1738.750 ;
        RECT 1408.150 1738.235 1408.430 1738.605 ;
        RECT 1408.160 1733.670 1408.420 1733.990 ;
        RECT 1408.220 1733.165 1408.360 1733.670 ;
        RECT 1408.150 1732.795 1408.430 1733.165 ;
        RECT 1408.160 1728.405 1408.420 1728.550 ;
        RECT 1408.150 1728.035 1408.430 1728.405 ;
        RECT 1408.160 1724.150 1408.420 1724.470 ;
        RECT 1408.220 1723.645 1408.360 1724.150 ;
        RECT 1408.150 1723.275 1408.430 1723.645 ;
        RECT 1408.150 1717.835 1408.430 1718.205 ;
        RECT 1408.160 1717.690 1408.420 1717.835 ;
        RECT 1408.160 1710.890 1408.420 1711.210 ;
        RECT 1408.220 1708.005 1408.360 1710.890 ;
        RECT 1408.150 1707.635 1408.430 1708.005 ;
        RECT 1408.160 1703.750 1408.420 1704.070 ;
        RECT 1408.680 1703.810 1408.820 2034.830 ;
        RECT 1410.060 2028.850 1410.200 2054.970 ;
        RECT 1410.920 2054.630 1411.180 2054.950 ;
        RECT 1410.980 2029.530 1411.120 2054.630 ;
        RECT 1411.380 2054.290 1411.640 2054.610 ;
        RECT 1411.440 2030.210 1411.580 2054.290 ;
        RECT 1413.220 2053.950 1413.480 2054.270 ;
        RECT 1412.760 2053.610 1413.020 2053.930 ;
        RECT 1412.300 2053.270 1412.560 2053.590 ;
        RECT 1411.840 2052.930 1412.100 2053.250 ;
        RECT 1411.900 2031.005 1412.040 2052.930 ;
        RECT 1412.360 2032.930 1412.500 2053.270 ;
        RECT 1412.820 2033.610 1412.960 2053.610 ;
        RECT 1413.280 2034.290 1413.420 2053.950 ;
        RECT 1413.740 2051.405 1413.880 2055.990 ;
        RECT 1414.130 2055.795 1414.410 2056.165 ;
        RECT 1414.140 2055.650 1414.400 2055.795 ;
        RECT 1414.140 2052.590 1414.400 2052.910 ;
        RECT 1413.670 2051.035 1413.950 2051.405 ;
        RECT 1414.200 2036.445 1414.340 2052.590 ;
        RECT 1414.130 2036.075 1414.410 2036.445 ;
        RECT 1413.280 2034.150 1413.880 2034.290 ;
        RECT 1412.820 2033.470 1413.420 2033.610 ;
        RECT 1412.360 2032.790 1412.960 2032.930 ;
        RECT 1411.830 2030.635 1412.110 2031.005 ;
        RECT 1411.440 2030.070 1412.500 2030.210 ;
        RECT 1410.980 2029.390 1412.040 2029.530 ;
        RECT 1410.060 2028.710 1411.120 2028.850 ;
        RECT 1410.980 1980.150 1411.120 2028.710 ;
        RECT 1411.380 2000.230 1411.640 2000.550 ;
        RECT 1411.440 1995.645 1411.580 2000.230 ;
        RECT 1411.370 1995.275 1411.650 1995.645 ;
        RECT 1410.920 1979.830 1411.180 1980.150 ;
        RECT 1411.380 1931.890 1411.640 1932.210 ;
        RECT 1409.080 1910.810 1409.340 1911.130 ;
        RECT 1409.140 1905.205 1409.280 1910.810 ;
        RECT 1409.070 1904.835 1409.350 1905.205 ;
        RECT 1409.080 1890.070 1409.340 1890.390 ;
        RECT 1409.140 1884.805 1409.280 1890.070 ;
        RECT 1409.070 1884.435 1409.350 1884.805 ;
        RECT 1409.080 1869.670 1409.340 1869.990 ;
        RECT 1409.140 1864.405 1409.280 1869.670 ;
        RECT 1409.070 1864.035 1409.350 1864.405 ;
        RECT 1409.080 1855.730 1409.340 1856.050 ;
        RECT 1409.140 1849.445 1409.280 1855.730 ;
        RECT 1411.440 1849.590 1411.580 1931.890 ;
        RECT 1409.070 1849.075 1409.350 1849.445 ;
        RECT 1411.380 1849.270 1411.640 1849.590 ;
        RECT 1410.920 1835.730 1411.180 1835.990 ;
        RECT 1410.520 1835.670 1411.180 1835.730 ;
        RECT 1410.520 1835.590 1411.120 1835.670 ;
        RECT 1410.520 1835.310 1410.660 1835.590 ;
        RECT 1410.460 1834.990 1410.720 1835.310 ;
        RECT 1411.380 1824.790 1411.640 1825.110 ;
        RECT 1409.080 1813.910 1409.340 1814.230 ;
        RECT 1409.140 1809.325 1409.280 1813.910 ;
        RECT 1409.070 1808.955 1409.350 1809.325 ;
        RECT 1409.080 1800.310 1409.340 1800.630 ;
        RECT 1409.140 1794.365 1409.280 1800.310 ;
        RECT 1409.070 1793.995 1409.350 1794.365 ;
        RECT 1410.920 1787.050 1411.180 1787.370 ;
        RECT 1410.980 1762.970 1411.120 1787.050 ;
        RECT 1411.440 1773.965 1411.580 1824.790 ;
        RECT 1411.370 1773.595 1411.650 1773.965 ;
        RECT 1411.900 1763.765 1412.040 2029.390 ;
        RECT 1412.360 1768.525 1412.500 2030.070 ;
        RECT 1412.820 1778.725 1412.960 2032.790 ;
        RECT 1413.280 1784.165 1413.420 2033.470 ;
        RECT 1413.740 1825.110 1413.880 2034.150 ;
        RECT 1414.130 2026.130 1414.410 2026.245 ;
        RECT 1415.580 2026.130 1415.720 2080.130 ;
        RECT 1414.130 2025.990 1415.720 2026.130 ;
        RECT 1414.130 2025.875 1414.410 2025.990 ;
        RECT 1416.040 2022.050 1416.180 2080.470 ;
        RECT 1414.660 2021.910 1416.180 2022.050 ;
        RECT 1414.130 2021.370 1414.410 2021.485 ;
        RECT 1414.660 2021.370 1414.800 2021.910 ;
        RECT 1414.130 2021.230 1414.800 2021.370 ;
        RECT 1414.130 2021.115 1414.410 2021.230 ;
        RECT 1416.500 2020.270 1416.640 2080.810 ;
        RECT 1416.960 2067.045 1417.100 2167.315 ;
        RECT 1417.420 2069.570 1417.560 2192.475 ;
        RECT 1417.360 2069.250 1417.620 2069.570 ;
        RECT 1417.880 2068.405 1418.020 2605.915 ;
        RECT 1418.740 2595.230 1419.000 2595.550 ;
        RECT 1418.280 2311.670 1418.540 2311.990 ;
        RECT 1417.810 2068.035 1418.090 2068.405 ;
        RECT 1416.890 2066.675 1417.170 2067.045 ;
        RECT 1418.340 2063.450 1418.480 2311.670 ;
        RECT 1418.800 2067.725 1418.940 2595.230 ;
        RECT 1419.660 2490.850 1419.920 2491.170 ;
        RECT 1419.200 2298.070 1419.460 2298.390 ;
        RECT 1418.730 2067.355 1419.010 2067.725 ;
        RECT 1419.260 2063.790 1419.400 2298.070 ;
        RECT 1419.720 2066.365 1419.860 2490.850 ;
        RECT 1420.120 2290.930 1420.380 2291.250 ;
        RECT 1419.650 2065.995 1419.930 2066.365 ;
        RECT 1420.180 2064.130 1420.320 2290.930 ;
        RECT 1420.580 2283.790 1420.840 2284.110 ;
        RECT 1420.640 2064.810 1420.780 2283.790 ;
        RECT 1421.040 2277.330 1421.300 2277.650 ;
        RECT 1420.580 2064.490 1420.840 2064.810 ;
        RECT 1421.100 2064.470 1421.240 2277.330 ;
        RECT 1422.880 2081.830 1423.140 2082.150 ;
        RECT 1421.960 2071.970 1422.220 2072.290 ;
        RECT 1421.040 2064.150 1421.300 2064.470 ;
        RECT 1420.120 2063.810 1420.380 2064.130 ;
        RECT 1419.200 2063.470 1419.460 2063.790 ;
        RECT 1418.280 2063.130 1418.540 2063.450 ;
        RECT 1419.660 2062.790 1419.920 2063.110 ;
        RECT 1418.740 2062.450 1419.000 2062.770 ;
        RECT 1417.360 2061.090 1417.620 2061.410 ;
        RECT 1416.900 2059.730 1417.160 2060.050 ;
        RECT 1416.440 2019.950 1416.700 2020.270 ;
        RECT 1414.140 2011.285 1414.400 2011.430 ;
        RECT 1414.130 2010.915 1414.410 2011.285 ;
        RECT 1414.140 2005.845 1414.400 2005.990 ;
        RECT 1414.130 2005.475 1414.410 2005.845 ;
        RECT 1414.130 2000.715 1414.410 2001.085 ;
        RECT 1414.140 2000.570 1414.400 2000.715 ;
        RECT 1416.960 1991.030 1417.100 2059.730 ;
        RECT 1416.900 1990.710 1417.160 1991.030 ;
        RECT 1417.420 1982.530 1417.560 2061.090 ;
        RECT 1418.280 2059.050 1418.540 2059.370 ;
        RECT 1417.820 2058.710 1418.080 2059.030 ;
        RECT 1417.360 1982.210 1417.620 1982.530 ;
        RECT 1417.880 1945.470 1418.020 2058.710 ;
        RECT 1418.340 1950.910 1418.480 2059.050 ;
        RECT 1418.800 1958.390 1418.940 2062.450 ;
        RECT 1419.200 2062.110 1419.460 2062.430 ;
        RECT 1419.260 1966.210 1419.400 2062.110 ;
        RECT 1419.200 1965.890 1419.460 1966.210 ;
        RECT 1419.720 1960.430 1419.860 2062.790 ;
        RECT 1420.120 2061.770 1420.380 2062.090 ;
        RECT 1420.180 1971.990 1420.320 2061.770 ;
        RECT 1420.580 2061.430 1420.840 2061.750 ;
        RECT 1420.640 1979.130 1420.780 2061.430 ;
        RECT 1421.040 2060.750 1421.300 2061.070 ;
        RECT 1421.100 1986.270 1421.240 2060.750 ;
        RECT 1421.500 2052.250 1421.760 2052.570 ;
        RECT 1421.040 1985.950 1421.300 1986.270 ;
        RECT 1420.580 1978.810 1420.840 1979.130 ;
        RECT 1420.120 1971.670 1420.380 1971.990 ;
        RECT 1419.660 1960.110 1419.920 1960.430 ;
        RECT 1418.740 1958.070 1419.000 1958.390 ;
        RECT 1418.280 1950.590 1418.540 1950.910 ;
        RECT 1417.820 1945.150 1418.080 1945.470 ;
        RECT 1421.560 1910.790 1421.700 2052.250 ;
        RECT 1422.020 1920.310 1422.160 2071.970 ;
        RECT 1422.420 2071.630 1422.680 2071.950 ;
        RECT 1421.960 1919.990 1422.220 1920.310 ;
        RECT 1422.480 1916.570 1422.620 2071.630 ;
        RECT 1422.420 1916.250 1422.680 1916.570 ;
        RECT 1421.500 1910.470 1421.760 1910.790 ;
        RECT 1422.420 1834.990 1422.680 1835.310 ;
        RECT 1422.480 1834.485 1422.620 1834.990 ;
        RECT 1422.410 1834.115 1422.690 1834.485 ;
        RECT 1413.680 1824.790 1413.940 1825.110 ;
        RECT 1413.210 1783.795 1413.490 1784.165 ;
        RECT 1412.750 1778.355 1413.030 1778.725 ;
        RECT 1412.290 1768.155 1412.570 1768.525 ;
        RECT 1411.830 1763.395 1412.110 1763.765 ;
        RECT 1410.980 1762.830 1411.580 1762.970 ;
        RECT 1409.080 1717.350 1409.340 1717.670 ;
        RECT 1409.140 1713.445 1409.280 1717.350 ;
        RECT 1409.070 1713.075 1409.350 1713.445 ;
        RECT 1411.440 1704.410 1411.580 1762.830 ;
        RECT 1422.940 1751.670 1423.080 2081.830 ;
        RECT 1423.800 2075.370 1424.060 2075.690 ;
        RECT 1423.340 2074.690 1423.600 2075.010 ;
        RECT 1422.880 1751.350 1423.140 1751.670 ;
        RECT 1411.380 1704.090 1411.640 1704.410 ;
        RECT 1412.300 1704.090 1412.560 1704.410 ;
        RECT 1408.220 1703.245 1408.360 1703.750 ;
        RECT 1408.680 1703.670 1409.740 1703.810 ;
        RECT 1408.150 1702.875 1408.430 1703.245 ;
        RECT 1408.620 1703.070 1408.880 1703.390 ;
        RECT 1408.680 1698.485 1408.820 1703.070 ;
        RECT 1408.610 1698.115 1408.890 1698.485 ;
        RECT 1408.160 1693.890 1408.420 1694.210 ;
        RECT 1408.220 1693.045 1408.360 1693.890 ;
        RECT 1408.150 1692.675 1408.430 1693.045 ;
        RECT 1408.160 1689.470 1408.420 1689.790 ;
        RECT 1408.220 1688.285 1408.360 1689.470 ;
        RECT 1408.150 1687.915 1408.430 1688.285 ;
        RECT 1408.620 1683.350 1408.880 1683.670 ;
        RECT 1408.160 1682.845 1408.420 1682.990 ;
        RECT 1408.150 1682.475 1408.430 1682.845 ;
        RECT 1408.680 1678.085 1408.820 1683.350 ;
        RECT 1408.610 1677.715 1408.890 1678.085 ;
        RECT 1408.160 1672.810 1408.420 1673.130 ;
        RECT 1408.220 1672.645 1408.360 1672.810 ;
        RECT 1408.150 1672.275 1408.430 1672.645 ;
        RECT 1408.620 1669.410 1408.880 1669.730 ;
        RECT 1408.160 1668.050 1408.420 1668.370 ;
        RECT 1408.220 1667.885 1408.360 1668.050 ;
        RECT 1408.150 1667.515 1408.430 1667.885 ;
        RECT 1408.680 1663.125 1408.820 1669.410 ;
        RECT 1408.610 1662.755 1408.890 1663.125 ;
        RECT 1409.600 1657.685 1409.740 1703.670 ;
        RECT 1412.360 1690.470 1412.500 1704.090 ;
        RECT 1423.400 1703.390 1423.540 2074.690 ;
        RECT 1423.860 1704.070 1424.000 2075.370 ;
        RECT 1424.260 2075.030 1424.520 2075.350 ;
        RECT 1423.800 1703.750 1424.060 1704.070 ;
        RECT 1423.340 1703.070 1423.600 1703.390 ;
        RECT 1424.320 1694.210 1424.460 2075.030 ;
        RECT 1424.780 1724.470 1424.920 3201.450 ;
        RECT 1425.640 2790.390 1425.900 2790.710 ;
        RECT 1425.180 2788.350 1425.440 2788.670 ;
        RECT 1424.720 1724.150 1424.980 1724.470 ;
        RECT 1424.260 1693.890 1424.520 1694.210 ;
        RECT 1412.300 1690.150 1412.560 1690.470 ;
        RECT 1409.530 1657.315 1409.810 1657.685 ;
        RECT 1408.160 1655.810 1408.420 1656.130 ;
        RECT 1408.220 1652.925 1408.360 1655.810 ;
        RECT 1408.150 1652.555 1408.430 1652.925 ;
        RECT 1407.760 1649.270 1408.820 1649.410 ;
        RECT 1407.700 1648.670 1407.960 1648.990 ;
        RECT 1407.760 1647.485 1407.900 1648.670 ;
        RECT 1408.160 1648.330 1408.420 1648.650 ;
        RECT 1407.690 1647.115 1407.970 1647.485 ;
        RECT 1408.220 1642.725 1408.360 1648.330 ;
        RECT 1408.150 1642.355 1408.430 1642.725 ;
        RECT 1407.700 1641.870 1407.960 1642.190 ;
        RECT 1407.760 1637.285 1407.900 1641.870 ;
        RECT 1407.690 1636.915 1407.970 1637.285 ;
        RECT 1407.700 1627.765 1407.960 1627.910 ;
        RECT 1407.690 1627.395 1407.970 1627.765 ;
        RECT 1408.680 1612.125 1408.820 1649.270 ;
        RECT 1411.840 1642.210 1412.100 1642.530 ;
        RECT 1411.900 1632.525 1412.040 1642.210 ;
        RECT 1411.830 1632.155 1412.110 1632.525 ;
        RECT 1425.240 1627.910 1425.380 2788.350 ;
        RECT 1425.700 1855.030 1425.840 2790.390 ;
        RECT 1431.160 2081.490 1431.420 2081.810 ;
        RECT 1430.700 2081.150 1430.960 2081.470 ;
        RECT 1427.020 2076.050 1427.280 2076.370 ;
        RECT 1426.560 2075.710 1426.820 2076.030 ;
        RECT 1426.100 2074.350 1426.360 2074.670 ;
        RECT 1425.640 1854.710 1425.900 1855.030 ;
        RECT 1425.640 1834.650 1425.900 1834.970 ;
        RECT 1425.700 1829.045 1425.840 1834.650 ;
        RECT 1425.630 1828.675 1425.910 1829.045 ;
        RECT 1426.160 1668.370 1426.300 2074.350 ;
        RECT 1426.620 1673.130 1426.760 2075.710 ;
        RECT 1427.080 1683.670 1427.220 2076.050 ;
        RECT 1427.480 2072.990 1427.740 2073.310 ;
        RECT 1427.020 1683.350 1427.280 1683.670 ;
        RECT 1427.540 1682.990 1427.680 2072.990 ;
        RECT 1427.940 2072.650 1428.200 2072.970 ;
        RECT 1428.000 1689.790 1428.140 2072.650 ;
        RECT 1430.760 2011.430 1430.900 2081.150 ;
        RECT 1430.700 2011.110 1430.960 2011.430 ;
        RECT 1431.220 2005.990 1431.360 2081.490 ;
        RECT 1431.160 2005.670 1431.420 2005.990 ;
        RECT 1431.680 1728.550 1431.820 3208.590 ;
        RECT 1432.080 2793.790 1432.340 2794.110 ;
        RECT 1432.140 1754.730 1432.280 2793.790 ;
        RECT 1432.540 2793.450 1432.800 2793.770 ;
        RECT 1432.600 1759.150 1432.740 2793.450 ;
        RECT 1433.000 2789.370 1433.260 2789.690 ;
        RECT 1433.060 1859.790 1433.200 2789.370 ;
        RECT 1435.290 2066.675 1435.570 2067.045 ;
        RECT 1435.360 2065.685 1435.500 2066.675 ;
        RECT 1435.750 2065.995 1436.030 2066.365 ;
        RECT 1435.290 2065.315 1435.570 2065.685 ;
        RECT 1435.300 2065.005 1435.560 2065.150 ;
        RECT 1435.290 2064.635 1435.570 2065.005 ;
        RECT 1435.820 2064.325 1435.960 2065.995 ;
        RECT 1435.750 2063.955 1436.030 2064.325 ;
        RECT 1434.840 2058.370 1435.100 2058.690 ;
        RECT 1434.380 2058.030 1434.640 2058.350 ;
        RECT 1433.460 2057.690 1433.720 2058.010 ;
        RECT 1433.520 1930.510 1433.660 2057.690 ;
        RECT 1433.920 2057.350 1434.180 2057.670 ;
        RECT 1433.460 1930.190 1433.720 1930.510 ;
        RECT 1433.980 1926.430 1434.120 2057.350 ;
        RECT 1434.440 1935.610 1434.580 2058.030 ;
        RECT 1434.900 1941.730 1435.040 2058.370 ;
        RECT 1434.840 1941.410 1435.100 1941.730 ;
        RECT 1434.380 1935.290 1434.640 1935.610 ;
        RECT 1433.920 1926.110 1434.180 1926.430 ;
        RECT 1433.000 1859.470 1433.260 1859.790 ;
        RECT 1432.540 1758.830 1432.800 1759.150 ;
        RECT 1432.080 1754.410 1432.340 1754.730 ;
        RECT 1438.580 1733.990 1438.720 3215.390 ;
        RECT 1438.980 2788.690 1439.240 2789.010 ;
        RECT 1439.040 1865.910 1439.180 2788.690 ;
        RECT 1438.980 1865.590 1439.240 1865.910 ;
        RECT 1452.380 1738.750 1452.520 3222.190 ;
        RECT 1459.280 1745.550 1459.420 3229.330 ;
        RECT 1535.570 3224.715 1535.850 3225.085 ;
        RECT 1535.640 3222.510 1535.780 3224.715 ;
        RECT 1535.580 3222.190 1535.840 3222.510 ;
        RECT 1535.570 3217.235 1535.850 3217.605 ;
        RECT 1535.640 3215.710 1535.780 3217.235 ;
        RECT 1535.580 3215.390 1535.840 3215.710 ;
        RECT 1538.330 3210.435 1538.610 3210.805 ;
        RECT 1538.400 3208.910 1538.540 3210.435 ;
        RECT 1538.340 3208.590 1538.600 3208.910 ;
        RECT 1538.330 3202.275 1538.610 3202.645 ;
        RECT 1538.400 3201.770 1538.540 3202.275 ;
        RECT 1538.340 3201.450 1538.600 3201.770 ;
        RECT 1535.110 3196.155 1535.390 3196.525 ;
        RECT 1534.190 3189.355 1534.470 3189.725 ;
        RECT 1534.260 3188.170 1534.400 3189.355 ;
        RECT 1459.680 3187.850 1459.940 3188.170 ;
        RECT 1534.200 3187.850 1534.460 3188.170 ;
        RECT 1459.220 1745.230 1459.480 1745.550 ;
        RECT 1452.320 1738.430 1452.580 1738.750 ;
        RECT 1438.520 1733.670 1438.780 1733.990 ;
        RECT 1431.620 1728.230 1431.880 1728.550 ;
        RECT 1459.740 1717.670 1459.880 3187.850 ;
        RECT 1514.420 2898.170 1514.680 2898.490 ;
        RECT 1460.140 2074.010 1460.400 2074.330 ;
        RECT 1460.200 2000.550 1460.340 2074.010 ;
        RECT 1483.130 2066.675 1483.410 2067.045 ;
        RECT 1482.670 2065.995 1482.950 2066.365 ;
        RECT 1482.740 2064.325 1482.880 2065.995 ;
        RECT 1483.200 2065.685 1483.340 2066.675 ;
        RECT 1483.130 2065.315 1483.410 2065.685 ;
        RECT 1483.140 2065.005 1483.400 2065.150 ;
        RECT 1483.130 2064.635 1483.410 2065.005 ;
        RECT 1482.670 2063.955 1482.950 2064.325 ;
        RECT 1462.900 2059.390 1463.160 2059.710 ;
        RECT 1462.960 2049.170 1463.100 2059.390 ;
        RECT 1462.900 2048.850 1463.160 2049.170 ;
        RECT 1460.140 2000.230 1460.400 2000.550 ;
        RECT 1459.680 1717.350 1459.940 1717.670 ;
        RECT 1427.940 1689.470 1428.200 1689.790 ;
        RECT 1427.480 1682.670 1427.740 1682.990 ;
        RECT 1426.560 1672.810 1426.820 1673.130 ;
        RECT 1514.480 1669.730 1514.620 2898.170 ;
        RECT 1531.890 2066.675 1532.170 2067.045 ;
        RECT 1531.960 2065.685 1532.100 2066.675 ;
        RECT 1532.350 2065.995 1532.630 2066.365 ;
        RECT 1531.890 2065.315 1532.170 2065.685 ;
        RECT 1531.900 2065.005 1532.160 2065.150 ;
        RECT 1531.890 2064.635 1532.170 2065.005 ;
        RECT 1532.420 2064.325 1532.560 2065.995 ;
        RECT 1532.350 2063.955 1532.630 2064.325 ;
        RECT 1535.180 1718.010 1535.320 3196.155 ;
        RECT 1538.330 2898.995 1538.610 2899.365 ;
        RECT 1538.400 2898.490 1538.540 2898.995 ;
        RECT 1538.340 2898.170 1538.600 2898.490 ;
      LAYER met2 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met2 ;
        RECT 1935.840 3249.565 1935.980 3252.110 ;
        RECT 1945.900 3250.750 1946.160 3251.070 ;
        RECT 1945.960 3249.565 1946.100 3250.750 ;
        RECT 1935.770 3249.195 1936.050 3249.565 ;
        RECT 1945.890 3249.195 1946.170 3249.565 ;
        RECT 1742.110 2796.315 1742.390 2796.685 ;
        RECT 1790.870 2796.315 1791.150 2796.685 ;
        RECT 1587.090 2794.275 1587.370 2794.645 ;
        RECT 1593.990 2794.275 1594.270 2794.645 ;
        RECT 1600.890 2794.275 1601.170 2794.645 ;
        RECT 1628.490 2794.275 1628.770 2794.645 ;
        RECT 1635.390 2794.275 1635.670 2794.645 ;
        RECT 1646.430 2794.275 1646.710 2794.645 ;
        RECT 1649.650 2794.275 1649.930 2794.645 ;
        RECT 1658.850 2794.275 1659.130 2794.645 ;
        RECT 1662.990 2794.275 1663.270 2794.645 ;
        RECT 1669.890 2794.275 1670.170 2794.645 ;
        RECT 1676.790 2794.275 1677.070 2794.645 ;
        RECT 1683.690 2794.275 1683.970 2794.645 ;
        RECT 1687.830 2794.275 1688.110 2794.645 ;
        RECT 1690.590 2794.275 1690.870 2794.645 ;
        RECT 1697.490 2794.275 1697.770 2794.645 ;
        RECT 1704.390 2794.275 1704.670 2794.645 ;
        RECT 1711.290 2794.275 1711.570 2794.645 ;
        RECT 1718.650 2794.275 1718.930 2794.645 ;
        RECT 1721.410 2794.275 1721.690 2794.645 ;
        RECT 1725.090 2794.275 1725.370 2794.645 ;
        RECT 1731.990 2794.275 1732.270 2794.645 ;
        RECT 1562.720 2790.050 1562.980 2790.370 ;
        RECT 1548.920 2789.710 1549.180 2790.030 ;
        RECT 1542.020 2787.670 1542.280 2787.990 ;
        RECT 1535.120 1717.690 1535.380 1718.010 ;
        RECT 1542.080 1711.210 1542.220 2787.670 ;
        RECT 1548.980 1834.970 1549.120 2789.710 ;
        RECT 1562.780 1835.310 1562.920 2790.050 ;
        RECT 1581.570 2788.835 1581.850 2789.205 ;
        RECT 1576.520 2788.010 1576.780 2788.330 ;
        RECT 1576.580 1842.450 1576.720 2788.010 ;
        RECT 1581.640 2787.990 1581.780 2788.835 ;
        RECT 1581.580 2787.670 1581.840 2787.990 ;
        RECT 1579.730 2066.675 1580.010 2067.045 ;
        RECT 1579.270 2065.995 1579.550 2066.365 ;
        RECT 1579.340 2064.325 1579.480 2065.995 ;
        RECT 1579.800 2065.685 1579.940 2066.675 ;
        RECT 1579.730 2065.315 1580.010 2065.685 ;
        RECT 1579.740 2065.005 1580.000 2065.150 ;
        RECT 1579.730 2064.635 1580.010 2065.005 ;
        RECT 1579.270 2063.955 1579.550 2064.325 ;
        RECT 1576.520 1842.130 1576.780 1842.450 ;
        RECT 1562.720 1834.990 1562.980 1835.310 ;
        RECT 1548.920 1834.650 1549.180 1834.970 ;
        RECT 1542.020 1710.890 1542.280 1711.210 ;
        RECT 1514.420 1669.410 1514.680 1669.730 ;
        RECT 1426.100 1668.050 1426.360 1668.370 ;
        RECT 1587.160 1642.190 1587.300 2794.275 ;
        RECT 1594.060 1648.650 1594.200 2794.275 ;
        RECT 1600.960 1648.990 1601.100 2794.275 ;
        RECT 1601.350 2793.595 1601.630 2793.965 ;
        RECT 1611.010 2793.595 1611.290 2793.965 ;
        RECT 1601.420 1656.130 1601.560 2793.595 ;
        RECT 1607.790 2790.195 1608.070 2790.565 ;
        RECT 1607.860 2790.030 1608.000 2790.195 ;
        RECT 1611.080 2790.030 1611.220 2793.595 ;
        RECT 1617.910 2792.915 1618.190 2793.285 ;
        RECT 1624.810 2792.915 1625.090 2793.285 ;
        RECT 1614.690 2790.195 1614.970 2790.565 ;
        RECT 1617.980 2790.370 1618.120 2792.915 ;
        RECT 1614.700 2790.050 1614.960 2790.195 ;
        RECT 1617.920 2790.050 1618.180 2790.370 ;
        RECT 1607.800 2789.710 1608.060 2790.030 ;
        RECT 1611.020 2789.710 1611.280 2790.030 ;
        RECT 1611.080 1793.830 1611.220 2789.710 ;
        RECT 1617.980 1800.630 1618.120 2790.050 ;
        RECT 1624.880 2789.350 1625.020 2792.915 ;
        RECT 1624.820 2789.030 1625.080 2789.350 ;
        RECT 1621.590 2788.155 1621.870 2788.525 ;
        RECT 1621.600 2788.010 1621.860 2788.155 ;
        RECT 1624.880 1800.970 1625.020 2789.030 ;
        RECT 1628.560 1849.250 1628.700 2794.275 ;
        RECT 1631.710 2793.595 1631.990 2793.965 ;
        RECT 1631.780 2793.430 1631.920 2793.595 ;
        RECT 1631.720 2793.110 1631.980 2793.430 ;
        RECT 1628.500 1848.930 1628.760 1849.250 ;
        RECT 1631.780 1807.770 1631.920 2793.110 ;
        RECT 1635.460 1856.050 1635.600 2794.275 ;
        RECT 1642.290 2793.595 1642.570 2793.965 ;
        RECT 1638.610 2792.915 1638.890 2793.285 ;
        RECT 1638.680 2788.330 1638.820 2792.915 ;
        RECT 1642.360 2790.710 1642.500 2793.595 ;
        RECT 1645.510 2792.915 1645.790 2793.285 ;
        RECT 1642.300 2790.390 1642.560 2790.710 ;
        RECT 1638.620 2788.010 1638.880 2788.330 ;
        RECT 1635.400 1855.730 1635.660 1856.050 ;
        RECT 1638.680 1814.230 1638.820 2788.010 ;
        RECT 1645.580 2787.990 1645.720 2792.915 ;
        RECT 1646.500 2792.410 1646.640 2794.275 ;
        RECT 1646.440 2792.090 1646.700 2792.410 ;
        RECT 1645.520 2787.670 1645.780 2787.990 ;
        RECT 1645.580 1814.570 1645.720 2787.670 ;
        RECT 1646.500 1821.710 1646.640 2792.090 ;
        RECT 1649.190 2789.515 1649.470 2789.885 ;
        RECT 1649.200 2789.370 1649.460 2789.515 ;
        RECT 1649.720 1869.990 1649.860 2794.275 ;
        RECT 1652.410 2793.595 1652.690 2793.965 ;
        RECT 1652.480 2792.750 1652.620 2793.595 ;
        RECT 1652.420 2792.430 1652.680 2792.750 ;
        RECT 1649.660 1869.670 1649.920 1869.990 ;
        RECT 1652.480 1828.510 1652.620 2792.430 ;
        RECT 1658.920 2791.390 1659.060 2794.275 ;
        RECT 1658.860 2791.070 1659.120 2791.390 ;
        RECT 1656.090 2788.835 1656.370 2789.205 ;
        RECT 1656.100 2788.690 1656.360 2788.835 ;
        RECT 1655.640 2065.005 1655.900 2065.150 ;
        RECT 1655.630 2064.635 1655.910 2065.005 ;
        RECT 1663.060 1876.790 1663.200 2794.275 ;
        RECT 1665.750 2793.595 1666.030 2793.965 ;
        RECT 1665.820 2791.730 1665.960 2793.595 ;
        RECT 1665.760 2791.410 1666.020 2791.730 ;
        RECT 1669.960 1883.590 1670.100 2794.275 ;
        RECT 1670.350 2793.595 1670.630 2793.965 ;
        RECT 1670.420 2792.070 1670.560 2793.595 ;
        RECT 1670.360 2791.750 1670.620 2792.070 ;
        RECT 1676.340 2791.750 1676.600 2792.070 ;
        RECT 1676.400 2791.050 1676.540 2791.750 ;
        RECT 1676.340 2790.730 1676.600 2791.050 ;
        RECT 1676.330 2066.675 1676.610 2067.045 ;
        RECT 1675.870 2065.995 1676.150 2066.365 ;
        RECT 1675.940 2064.325 1676.080 2065.995 ;
        RECT 1676.400 2065.685 1676.540 2066.675 ;
        RECT 1676.330 2065.315 1676.610 2065.685 ;
        RECT 1676.340 2065.005 1676.600 2065.150 ;
        RECT 1676.330 2064.635 1676.610 2065.005 ;
        RECT 1675.870 2063.955 1676.150 2064.325 ;
        RECT 1676.860 1890.390 1677.000 2794.275 ;
        RECT 1677.250 2793.595 1677.530 2793.965 ;
        RECT 1683.230 2793.595 1683.510 2793.965 ;
        RECT 1677.320 2793.430 1677.460 2793.595 ;
        RECT 1677.260 2793.110 1677.520 2793.430 ;
        RECT 1683.300 2793.090 1683.440 2793.595 ;
        RECT 1680.480 2792.770 1680.740 2793.090 ;
        RECT 1683.240 2792.770 1683.500 2793.090 ;
        RECT 1680.540 2788.330 1680.680 2792.770 ;
        RECT 1680.480 2788.010 1680.740 2788.330 ;
        RECT 1683.760 1890.730 1683.900 2794.275 ;
        RECT 1684.150 2793.595 1684.430 2793.965 ;
        RECT 1684.220 1897.530 1684.360 2793.595 ;
        RECT 1687.900 2792.070 1688.040 2794.275 ;
        RECT 1687.840 2791.750 1688.100 2792.070 ;
        RECT 1687.900 2787.990 1688.040 2791.750 ;
        RECT 1687.840 2787.670 1688.100 2787.990 ;
        RECT 1686.920 2072.310 1687.180 2072.630 ;
        RECT 1686.980 2000.890 1687.120 2072.310 ;
        RECT 1690.140 2060.070 1690.400 2060.390 ;
        RECT 1690.200 2042.370 1690.340 2060.070 ;
        RECT 1690.140 2042.050 1690.400 2042.370 ;
        RECT 1686.920 2000.570 1687.180 2000.890 ;
        RECT 1690.660 1904.330 1690.800 2794.275 ;
        RECT 1695.190 2793.595 1695.470 2793.965 ;
        RECT 1695.260 2792.410 1695.400 2793.595 ;
        RECT 1695.200 2792.090 1695.460 2792.410 ;
        RECT 1693.820 2056.330 1694.080 2056.650 ;
        RECT 1690.600 1904.010 1690.860 1904.330 ;
        RECT 1684.160 1897.210 1684.420 1897.530 ;
        RECT 1683.700 1890.410 1683.960 1890.730 ;
        RECT 1676.800 1890.070 1677.060 1890.390 ;
        RECT 1669.900 1883.270 1670.160 1883.590 ;
        RECT 1663.000 1876.470 1663.260 1876.790 ;
        RECT 1652.420 1828.190 1652.680 1828.510 ;
        RECT 1646.440 1821.390 1646.700 1821.710 ;
        RECT 1645.520 1814.250 1645.780 1814.570 ;
        RECT 1638.620 1813.910 1638.880 1814.230 ;
        RECT 1631.720 1807.450 1631.980 1807.770 ;
        RECT 1624.820 1800.650 1625.080 1800.970 ;
        RECT 1617.920 1800.310 1618.180 1800.630 ;
        RECT 1611.020 1793.510 1611.280 1793.830 ;
        RECT 1601.360 1655.810 1601.620 1656.130 ;
        RECT 1600.900 1648.670 1601.160 1648.990 ;
        RECT 1594.000 1648.330 1594.260 1648.650 ;
        RECT 1587.100 1641.870 1587.360 1642.190 ;
        RECT 1425.180 1627.590 1425.440 1627.910 ;
        RECT 1408.610 1611.755 1408.890 1612.125 ;
        RECT 1693.880 1607.850 1694.020 2056.330 ;
        RECT 1697.560 1911.130 1697.700 2794.275 ;
        RECT 1699.330 2793.595 1699.610 2793.965 ;
        RECT 1699.400 2792.750 1699.540 2793.595 ;
        RECT 1699.340 2792.430 1699.600 2792.750 ;
        RECT 1704.460 2052.570 1704.600 2794.275 ;
        RECT 1706.230 2793.595 1706.510 2793.965 ;
        RECT 1706.300 2791.390 1706.440 2793.595 ;
        RECT 1706.240 2791.070 1706.500 2791.390 ;
        RECT 1711.360 2071.950 1711.500 2794.275 ;
        RECT 1712.670 2793.595 1712.950 2793.965 ;
        RECT 1718.190 2793.595 1718.470 2793.965 ;
        RECT 1712.740 2791.730 1712.880 2793.595 ;
        RECT 1712.680 2791.410 1712.940 2791.730 ;
        RECT 1718.260 2791.050 1718.400 2793.595 ;
        RECT 1718.200 2790.730 1718.460 2791.050 ;
        RECT 1718.190 2788.155 1718.470 2788.525 ;
        RECT 1711.300 2071.630 1711.560 2071.950 ;
        RECT 1715.440 2060.410 1715.700 2060.730 ;
        RECT 1715.500 2055.970 1715.640 2060.410 ;
        RECT 1718.260 2057.670 1718.400 2788.155 ;
        RECT 1718.720 2072.290 1718.860 2794.275 ;
        RECT 1721.480 2793.430 1721.620 2794.275 ;
        RECT 1721.420 2793.110 1721.680 2793.430 ;
        RECT 1718.660 2071.970 1718.920 2072.290 ;
        RECT 1725.160 2058.010 1725.300 2794.275 ;
        RECT 1730.150 2793.595 1730.430 2793.965 ;
        RECT 1730.220 2793.090 1730.360 2793.595 ;
        RECT 1730.160 2792.770 1730.420 2793.090 ;
        RECT 1732.060 2058.350 1732.200 2794.275 ;
        RECT 1738.440 2794.130 1738.700 2794.450 ;
        RECT 1738.890 2794.275 1739.170 2794.645 ;
        RECT 1738.500 2793.965 1738.640 2794.130 ;
        RECT 1738.430 2793.595 1738.710 2793.965 ;
        RECT 1738.500 2792.070 1738.640 2793.595 ;
        RECT 1738.440 2791.750 1738.700 2792.070 ;
        RECT 1738.960 2058.690 1739.100 2794.275 ;
        RECT 1741.190 2793.595 1741.470 2793.965 ;
        RECT 1741.260 2792.410 1741.400 2793.595 ;
        RECT 1741.200 2792.090 1741.460 2792.410 ;
        RECT 1742.180 2791.730 1742.320 2796.315 ;
        RECT 1745.790 2794.275 1746.070 2794.645 ;
        RECT 1760.050 2794.275 1760.330 2794.645 ;
        RECT 1780.290 2794.275 1780.570 2794.645 ;
        RECT 1742.120 2791.410 1742.380 2791.730 ;
        RECT 1745.860 2059.030 1746.000 2794.275 ;
        RECT 1748.550 2793.595 1748.830 2793.965 ;
        RECT 1748.620 2792.750 1748.760 2793.595 ;
        RECT 1748.560 2792.430 1748.820 2792.750 ;
        RECT 1752.690 2792.235 1752.970 2792.605 ;
        RECT 1752.760 2791.390 1752.900 2792.235 ;
        RECT 1752.700 2791.070 1752.960 2791.390 ;
        RECT 1760.120 2791.050 1760.260 2794.275 ;
        RECT 1780.300 2794.130 1780.560 2794.275 ;
        RECT 1766.490 2793.595 1766.770 2793.965 ;
        RECT 1773.390 2793.595 1773.670 2793.965 ;
        RECT 1766.560 2793.430 1766.700 2793.595 ;
        RECT 1766.500 2793.110 1766.760 2793.430 ;
        RECT 1773.460 2793.090 1773.600 2793.595 ;
        RECT 1773.400 2792.770 1773.660 2793.090 ;
        RECT 1790.940 2792.750 1791.080 2796.315 ;
        RECT 1787.190 2792.235 1787.470 2792.605 ;
        RECT 1790.880 2792.430 1791.140 2792.750 ;
        RECT 1787.200 2792.090 1787.460 2792.235 ;
        RECT 1762.820 2791.750 1763.080 2792.070 ;
        RECT 1760.060 2790.730 1760.320 2791.050 ;
        RECT 1760.510 2788.155 1760.790 2788.525 ;
        RECT 1753.150 2787.475 1753.430 2787.845 ;
        RECT 1752.240 2065.005 1752.500 2065.150 ;
        RECT 1752.230 2064.635 1752.510 2065.005 ;
        RECT 1753.220 2059.370 1753.360 2787.475 ;
        RECT 1760.050 2777.275 1760.330 2777.645 ;
        RECT 1760.120 2062.770 1760.260 2777.275 ;
        RECT 1760.580 2063.110 1760.720 2788.155 ;
        RECT 1762.880 2097.110 1763.020 2791.750 ;
        RECT 1763.280 2791.410 1763.540 2791.730 ;
        RECT 1763.340 2104.590 1763.480 2791.410 ;
        RECT 1769.720 2791.070 1769.980 2791.390 ;
        RECT 1766.490 2787.475 1766.770 2787.845 ;
        RECT 1763.280 2104.270 1763.540 2104.590 ;
        RECT 1762.820 2096.790 1763.080 2097.110 ;
        RECT 1760.520 2062.790 1760.780 2063.110 ;
        RECT 1760.060 2062.450 1760.320 2062.770 ;
        RECT 1766.560 2062.430 1766.700 2787.475 ;
        RECT 1769.780 2111.390 1769.920 2791.070 ;
        RECT 1770.180 2790.730 1770.440 2791.050 ;
        RECT 1770.240 2117.850 1770.380 2790.730 ;
        RECT 1783.520 2790.390 1783.780 2790.710 ;
        RECT 1776.620 2790.050 1776.880 2790.370 ;
        RECT 1773.390 2787.475 1773.670 2787.845 ;
        RECT 1770.640 2615.290 1770.900 2615.610 ;
        RECT 1770.180 2117.530 1770.440 2117.850 ;
        RECT 1769.720 2111.070 1769.980 2111.390 ;
        RECT 1770.700 2069.085 1770.840 2615.290 ;
        RECT 1770.630 2068.715 1770.910 2069.085 ;
        RECT 1772.930 2066.675 1773.210 2067.045 ;
        RECT 1772.470 2065.995 1772.750 2066.365 ;
        RECT 1772.540 2064.325 1772.680 2065.995 ;
        RECT 1773.000 2065.685 1773.140 2066.675 ;
        RECT 1772.930 2065.315 1773.210 2065.685 ;
        RECT 1772.940 2065.005 1773.200 2065.150 ;
        RECT 1772.930 2064.635 1773.210 2065.005 ;
        RECT 1772.470 2063.955 1772.750 2064.325 ;
        RECT 1766.500 2062.110 1766.760 2062.430 ;
        RECT 1773.460 2062.090 1773.600 2787.475 ;
        RECT 1776.680 2118.190 1776.820 2790.050 ;
        RECT 1777.080 2789.370 1777.340 2789.690 ;
        RECT 1777.140 2125.330 1777.280 2789.370 ;
        RECT 1780.750 2787.475 1781.030 2787.845 ;
        RECT 1777.080 2125.010 1777.340 2125.330 ;
        RECT 1776.620 2117.870 1776.880 2118.190 ;
        RECT 1773.400 2061.770 1773.660 2062.090 ;
        RECT 1780.820 2061.750 1780.960 2787.475 ;
        RECT 1783.580 2132.130 1783.720 2790.390 ;
        RECT 1783.980 2789.710 1784.240 2790.030 ;
        RECT 1784.040 2138.590 1784.180 2789.710 ;
        RECT 1790.420 2789.030 1790.680 2789.350 ;
        RECT 1787.650 2787.475 1787.930 2787.845 ;
        RECT 1783.980 2138.270 1784.240 2138.590 ;
        RECT 1783.520 2131.810 1783.780 2132.130 ;
        RECT 1780.760 2061.430 1781.020 2061.750 ;
        RECT 1787.720 2061.410 1787.860 2787.475 ;
        RECT 1790.480 2138.930 1790.620 2789.030 ;
        RECT 1790.880 2788.690 1791.140 2789.010 ;
        RECT 1790.940 2145.730 1791.080 2788.690 ;
        RECT 1794.550 2777.275 1794.830 2777.645 ;
        RECT 1790.880 2145.410 1791.140 2145.730 ;
        RECT 1790.420 2138.610 1790.680 2138.930 ;
        RECT 1787.660 2061.090 1787.920 2061.410 ;
        RECT 1794.620 2061.070 1794.760 2777.275 ;
        RECT 1835.500 2691.450 1835.760 2691.770 ;
        RECT 1835.560 2069.765 1835.700 2691.450 ;
        RECT 1842.400 2691.110 1842.660 2691.430 ;
        RECT 1838.720 2614.950 1838.980 2615.270 ;
        RECT 1835.490 2069.395 1835.770 2069.765 ;
        RECT 1821.690 2066.675 1821.970 2067.045 ;
        RECT 1821.760 2065.685 1821.900 2066.675 ;
        RECT 1821.690 2065.315 1821.970 2065.685 ;
        RECT 1821.700 2064.830 1821.960 2065.150 ;
        RECT 1821.760 2064.325 1821.900 2064.830 ;
        RECT 1821.690 2063.955 1821.970 2064.325 ;
        RECT 1835.490 2063.275 1835.770 2063.645 ;
        RECT 1838.780 2063.450 1838.920 2614.950 ;
        RECT 1842.460 2065.685 1842.600 2691.110 ;
        RECT 1849.300 2683.970 1849.560 2684.290 ;
        RECT 1842.860 2304.530 1843.120 2304.850 ;
        RECT 1842.920 2069.765 1843.060 2304.530 ;
        RECT 1842.850 2069.395 1843.130 2069.765 ;
        RECT 1849.360 2065.685 1849.500 2683.970 ;
        RECT 1856.200 2677.170 1856.460 2677.490 ;
        RECT 1849.760 2297.730 1850.020 2298.050 ;
        RECT 1849.820 2069.765 1849.960 2297.730 ;
        RECT 1856.260 2069.765 1856.400 2677.170 ;
        RECT 1863.100 2670.710 1863.360 2671.030 ;
        RECT 1859.420 2622.090 1859.680 2622.410 ;
        RECT 1859.480 2070.445 1859.620 2622.090 ;
        RECT 1859.410 2070.075 1859.690 2070.445 ;
        RECT 1863.160 2069.765 1863.300 2670.710 ;
        RECT 1870.000 2670.370 1870.260 2670.690 ;
        RECT 1866.320 2166.490 1866.580 2166.810 ;
        RECT 1849.750 2069.395 1850.030 2069.765 ;
        RECT 1856.190 2069.395 1856.470 2069.765 ;
        RECT 1863.090 2069.395 1863.370 2069.765 ;
        RECT 1841.470 2065.315 1841.750 2065.685 ;
        RECT 1842.390 2065.315 1842.670 2065.685 ;
        RECT 1849.290 2065.315 1849.570 2065.685 ;
        RECT 1854.810 2065.315 1855.090 2065.685 ;
        RECT 1841.540 2063.645 1841.680 2065.315 ;
        RECT 1854.880 2063.645 1855.020 2065.315 ;
        RECT 1856.650 2063.955 1856.930 2064.325 ;
        RECT 1866.380 2064.130 1866.520 2166.490 ;
        RECT 1869.530 2066.675 1869.810 2067.045 ;
        RECT 1869.600 2065.005 1869.740 2066.675 ;
        RECT 1870.060 2066.365 1870.200 2670.370 ;
        RECT 1876.900 2663.570 1877.160 2663.890 ;
        RECT 1873.220 2628.890 1873.480 2629.210 ;
        RECT 1869.990 2065.995 1870.270 2066.365 ;
        RECT 1869.530 2064.635 1869.810 2065.005 ;
        RECT 1870.000 2064.490 1870.260 2064.810 ;
        RECT 1870.060 2064.325 1870.200 2064.490 ;
        RECT 1873.280 2064.470 1873.420 2628.890 ;
        RECT 1873.680 2173.630 1873.940 2173.950 ;
        RECT 1856.720 2063.790 1856.860 2063.955 ;
        RECT 1863.100 2063.810 1863.360 2064.130 ;
        RECT 1866.320 2063.810 1866.580 2064.130 ;
        RECT 1869.990 2063.955 1870.270 2064.325 ;
        RECT 1870.920 2064.150 1871.180 2064.470 ;
        RECT 1873.220 2064.150 1873.480 2064.470 ;
        RECT 1856.200 2063.645 1856.460 2063.790 ;
        RECT 1835.500 2063.130 1835.760 2063.275 ;
        RECT 1838.720 2063.130 1838.980 2063.450 ;
        RECT 1841.470 2063.275 1841.750 2063.645 ;
        RECT 1854.810 2063.275 1855.090 2063.645 ;
        RECT 1856.190 2063.275 1856.470 2063.645 ;
        RECT 1856.660 2063.470 1856.920 2063.790 ;
        RECT 1863.160 2063.645 1863.300 2063.810 ;
        RECT 1870.980 2063.645 1871.120 2064.150 ;
        RECT 1873.740 2063.790 1873.880 2173.630 ;
        RECT 1876.960 2066.365 1877.100 2663.570 ;
        RECT 1877.360 2656.770 1877.620 2657.090 ;
        RECT 1876.890 2065.995 1877.170 2066.365 ;
        RECT 1877.420 2065.685 1877.560 2656.770 ;
        RECT 1883.800 2656.430 1884.060 2656.750 ;
        RECT 1880.120 2636.030 1880.380 2636.350 ;
        RECT 1877.820 2276.990 1878.080 2277.310 ;
        RECT 1877.880 2066.365 1878.020 2276.990 ;
        RECT 1880.180 2067.530 1880.320 2636.030 ;
        RECT 1880.120 2067.210 1880.380 2067.530 ;
        RECT 1883.860 2066.365 1884.000 2656.430 ;
        RECT 1891.160 2649.630 1891.420 2649.950 ;
        RECT 1887.020 2180.770 1887.280 2181.090 ;
        RECT 1877.810 2065.995 1878.090 2066.365 ;
        RECT 1883.790 2065.995 1884.070 2066.365 ;
        RECT 1877.350 2065.315 1877.630 2065.685 ;
        RECT 1883.800 2064.830 1884.060 2065.150 ;
        RECT 1883.860 2064.325 1884.000 2064.830 ;
        RECT 1883.790 2063.955 1884.070 2064.325 ;
        RECT 1887.080 2063.790 1887.220 2180.770 ;
        RECT 1891.220 2066.365 1891.360 2649.630 ;
        RECT 1898.060 2642.830 1898.320 2643.150 ;
        RECT 1893.920 2505.130 1894.180 2505.450 ;
        RECT 1891.150 2065.995 1891.430 2066.365 ;
        RECT 1893.980 2066.170 1894.120 2505.130 ;
        RECT 1898.120 2069.765 1898.260 2642.830 ;
        RECT 1904.960 2635.690 1905.220 2636.010 ;
        RECT 1900.820 2180.430 1901.080 2180.750 ;
        RECT 1898.050 2069.395 1898.330 2069.765 ;
        RECT 1898.970 2066.675 1899.250 2067.045 ;
        RECT 1893.920 2065.850 1894.180 2066.170 ;
        RECT 1890.700 2065.170 1890.960 2065.490 ;
        RECT 1898.060 2065.170 1898.320 2065.490 ;
        RECT 1890.760 2064.325 1890.900 2065.170 ;
        RECT 1898.120 2064.325 1898.260 2065.170 ;
        RECT 1899.040 2064.325 1899.180 2066.675 ;
        RECT 1900.880 2065.490 1901.020 2180.430 ;
        RECT 1903.110 2068.715 1903.390 2069.085 ;
        RECT 1903.180 2066.365 1903.320 2068.715 ;
        RECT 1905.020 2067.045 1905.160 2635.690 ;
        RECT 1939.460 2608.150 1939.720 2608.470 ;
        RECT 1935.320 2580.950 1935.580 2581.270 ;
        RECT 1928.420 2573.810 1928.680 2574.130 ;
        RECT 1921.520 2553.070 1921.780 2553.390 ;
        RECT 1914.620 2539.470 1914.880 2539.790 ;
        RECT 1907.720 2194.370 1907.980 2194.690 ;
        RECT 1907.780 2067.870 1907.920 2194.370 ;
        RECT 1907.720 2067.550 1907.980 2067.870 ;
        RECT 1911.400 2067.210 1911.660 2067.530 ;
        RECT 1911.460 2067.045 1911.600 2067.210 ;
        RECT 1904.950 2066.675 1905.230 2067.045 ;
        RECT 1910.940 2066.530 1911.200 2066.850 ;
        RECT 1911.390 2066.675 1911.670 2067.045 ;
        RECT 1903.110 2065.995 1903.390 2066.365 ;
        RECT 1911.000 2065.685 1911.140 2066.530 ;
        RECT 1911.860 2066.190 1912.120 2066.510 ;
        RECT 1911.920 2065.685 1912.060 2066.190 ;
        RECT 1900.820 2065.170 1901.080 2065.490 ;
        RECT 1910.930 2065.315 1911.210 2065.685 ;
        RECT 1911.850 2065.315 1912.130 2065.685 ;
        RECT 1904.500 2064.830 1904.760 2065.150 ;
        RECT 1890.690 2063.955 1890.970 2064.325 ;
        RECT 1898.050 2063.955 1898.330 2064.325 ;
        RECT 1898.970 2063.955 1899.250 2064.325 ;
        RECT 1863.090 2063.275 1863.370 2063.645 ;
        RECT 1870.910 2063.275 1871.190 2063.645 ;
        RECT 1873.680 2063.470 1873.940 2063.790 ;
        RECT 1887.020 2063.470 1887.280 2063.790 ;
        RECT 1904.560 2063.645 1904.700 2064.830 ;
        RECT 1914.680 2064.810 1914.820 2539.470 ;
        RECT 1915.080 2532.330 1915.340 2532.650 ;
        RECT 1915.140 2066.510 1915.280 2532.330 ;
        RECT 1915.540 2525.870 1915.800 2526.190 ;
        RECT 1915.600 2070.250 1915.740 2525.870 ;
        RECT 1916.000 2511.590 1916.260 2511.910 ;
        RECT 1915.540 2069.930 1915.800 2070.250 ;
        RECT 1916.060 2067.530 1916.200 2511.590 ;
        RECT 1921.580 2069.085 1921.720 2553.070 ;
        RECT 1921.980 2201.850 1922.240 2202.170 ;
        RECT 1921.510 2068.715 1921.790 2069.085 ;
        RECT 1916.000 2067.210 1916.260 2067.530 ;
        RECT 1915.080 2066.190 1915.340 2066.510 ;
        RECT 1922.040 2066.170 1922.180 2201.850 ;
        RECT 1926.570 2067.355 1926.850 2067.725 ;
        RECT 1921.520 2065.850 1921.780 2066.170 ;
        RECT 1921.980 2065.850 1922.240 2066.170 ;
        RECT 1918.300 2065.510 1918.560 2065.830 ;
        RECT 1914.620 2064.490 1914.880 2064.810 ;
        RECT 1911.400 2064.150 1911.660 2064.470 ;
        RECT 1911.460 2063.645 1911.600 2064.150 ;
        RECT 1918.360 2063.645 1918.500 2065.510 ;
        RECT 1921.580 2064.810 1921.720 2065.850 ;
        RECT 1926.640 2065.685 1926.780 2067.355 ;
        RECT 1925.190 2065.315 1925.470 2065.685 ;
        RECT 1926.570 2065.315 1926.850 2065.685 ;
        RECT 1921.520 2064.490 1921.780 2064.810 ;
        RECT 1925.260 2064.470 1925.400 2065.315 ;
        RECT 1928.480 2064.470 1928.620 2573.810 ;
        RECT 1928.880 2560.210 1929.140 2560.530 ;
        RECT 1928.940 2065.490 1929.080 2560.210 ;
        RECT 1932.100 2067.890 1932.360 2068.210 ;
        RECT 1932.160 2067.725 1932.300 2067.890 ;
        RECT 1932.090 2067.355 1932.370 2067.725 ;
        RECT 1928.880 2065.170 1929.140 2065.490 ;
        RECT 1925.200 2064.150 1925.460 2064.470 ;
        RECT 1928.420 2064.150 1928.680 2064.470 ;
        RECT 1935.380 2063.645 1935.520 2580.950 ;
        RECT 1935.780 2201.170 1936.040 2201.490 ;
        RECT 1935.840 2069.230 1935.980 2201.170 ;
        RECT 1939.520 2069.765 1939.660 2608.150 ;
        RECT 1953.260 2601.350 1953.520 2601.670 ;
        RECT 1942.220 2153.230 1942.480 2153.550 ;
        RECT 1942.280 2096.850 1942.420 2153.230 ;
        RECT 1942.280 2096.710 1942.880 2096.850 ;
        RECT 1939.450 2069.395 1939.730 2069.765 ;
        RECT 1935.780 2068.910 1936.040 2069.230 ;
        RECT 1942.740 2068.210 1942.880 2096.710 ;
        RECT 1953.320 2069.765 1953.460 2601.350 ;
        RECT 1960.160 2587.410 1960.420 2587.730 ;
        RECT 1960.220 2069.765 1960.360 2587.410 ;
        RECT 2031.920 2332.410 2032.180 2332.730 ;
        RECT 2014.900 2069.765 2015.160 2069.910 ;
        RECT 1953.250 2069.395 1953.530 2069.765 ;
        RECT 1960.150 2069.395 1960.430 2069.765 ;
        RECT 1980.400 2069.250 1980.660 2069.570 ;
        RECT 2014.890 2069.395 2015.170 2069.765 ;
        RECT 1959.700 2069.085 1959.960 2069.230 ;
        RECT 1980.460 2069.085 1980.600 2069.250 ;
        RECT 1946.360 2068.570 1946.620 2068.890 ;
        RECT 1959.690 2068.715 1959.970 2069.085 ;
        RECT 1980.390 2068.715 1980.670 2069.085 ;
        RECT 2031.980 2068.890 2032.120 2332.410 ;
        RECT 2038.880 2069.765 2039.020 3252.450 ;
        RECT 2582.080 3252.110 2582.340 3252.430 ;
        RECT 2190.610 3230.155 2190.890 3230.525 ;
        RECT 2097.700 2580.610 2097.960 2580.930 ;
        RECT 2052.620 2504.790 2052.880 2505.110 ;
        RECT 2045.720 2353.150 2045.980 2353.470 ;
        RECT 2038.810 2069.395 2039.090 2069.765 ;
        RECT 2045.780 2069.570 2045.920 2353.150 ;
        RECT 2052.680 2069.765 2052.820 2504.790 ;
        RECT 2081.600 2484.050 2081.860 2484.370 ;
        RECT 2080.220 2366.750 2080.480 2367.070 ;
        RECT 2059.520 2352.810 2059.780 2353.130 ;
        RECT 2045.720 2069.250 2045.980 2069.570 ;
        RECT 2052.610 2069.395 2052.890 2069.765 ;
        RECT 2031.920 2068.570 2032.180 2068.890 ;
        RECT 1945.900 2068.230 1946.160 2068.550 ;
        RECT 1942.680 2067.890 1942.940 2068.210 ;
        RECT 1945.960 2067.725 1946.100 2068.230 ;
        RECT 1945.890 2067.355 1946.170 2067.725 ;
        RECT 1939.000 2064.830 1939.260 2065.150 ;
        RECT 1946.420 2065.005 1946.560 2068.570 ;
        RECT 2021.800 2067.890 2022.060 2068.210 ;
        RECT 1973.500 2067.725 1973.760 2067.870 ;
        RECT 2021.860 2067.725 2022.000 2067.890 ;
        RECT 1946.810 2067.355 1947.090 2067.725 ;
        RECT 1973.490 2067.355 1973.770 2067.725 ;
        RECT 1939.060 2063.645 1939.200 2064.830 ;
        RECT 1945.430 2064.635 1945.710 2065.005 ;
        RECT 1946.350 2064.635 1946.630 2065.005 ;
        RECT 1945.500 2064.210 1945.640 2064.635 ;
        RECT 1946.880 2064.210 1947.020 2067.355 ;
        RECT 2008.000 2067.210 2008.260 2067.530 ;
        RECT 2021.790 2067.355 2022.070 2067.725 ;
        RECT 1987.300 2067.045 1987.560 2067.190 ;
        RECT 2008.060 2067.045 2008.200 2067.210 ;
        RECT 1966.130 2066.675 1966.410 2067.045 ;
        RECT 1987.290 2066.675 1987.570 2067.045 ;
        RECT 1952.800 2065.510 1953.060 2065.830 ;
        RECT 1952.860 2065.005 1953.000 2065.510 ;
        RECT 1952.790 2064.635 1953.070 2065.005 ;
        RECT 1966.200 2064.325 1966.340 2066.675 ;
        RECT 1987.760 2066.530 1988.020 2066.850 ;
        RECT 2007.990 2066.675 2008.270 2067.045 ;
        RECT 1966.600 2065.850 1966.860 2066.170 ;
        RECT 1966.660 2065.005 1966.800 2065.850 ;
        RECT 1987.820 2065.685 1987.960 2066.530 ;
        RECT 1994.200 2066.190 1994.460 2066.510 ;
        RECT 1994.260 2065.685 1994.400 2066.190 ;
        RECT 1980.400 2065.170 1980.660 2065.490 ;
        RECT 1987.750 2065.315 1988.030 2065.685 ;
        RECT 1994.190 2065.315 1994.470 2065.685 ;
        RECT 1980.460 2065.005 1980.600 2065.170 ;
        RECT 1987.300 2065.005 1987.560 2065.150 ;
        RECT 1966.590 2064.635 1966.870 2065.005 ;
        RECT 1980.390 2064.635 1980.670 2065.005 ;
        RECT 1987.290 2064.635 1987.570 2065.005 ;
        RECT 2015.820 2064.490 2016.080 2064.810 ;
        RECT 1973.500 2064.325 1973.760 2064.470 ;
        RECT 2015.880 2064.325 2016.020 2064.490 ;
        RECT 1945.500 2064.070 1947.020 2064.210 ;
        RECT 1966.130 2063.955 1966.410 2064.325 ;
        RECT 1973.490 2063.955 1973.770 2064.325 ;
        RECT 2001.090 2063.955 2001.370 2064.325 ;
        RECT 2015.810 2063.955 2016.090 2064.325 ;
        RECT 2052.680 2064.130 2052.820 2069.395 ;
        RECT 2059.580 2069.230 2059.720 2352.810 ;
        RECT 2059.520 2068.910 2059.780 2069.230 ;
        RECT 2080.280 2068.550 2080.420 2366.750 ;
        RECT 2080.220 2068.230 2080.480 2068.550 ;
        RECT 2001.100 2063.810 2001.360 2063.955 ;
        RECT 2052.620 2063.810 2052.880 2064.130 ;
        RECT 1994.200 2063.645 1994.460 2063.790 ;
        RECT 1904.490 2063.275 1904.770 2063.645 ;
        RECT 1911.390 2063.275 1911.670 2063.645 ;
        RECT 1918.290 2063.275 1918.570 2063.645 ;
        RECT 1925.190 2063.275 1925.470 2063.645 ;
        RECT 1935.310 2063.275 1935.590 2063.645 ;
        RECT 1938.990 2063.275 1939.270 2063.645 ;
        RECT 1994.190 2063.275 1994.470 2063.645 ;
        RECT 2001.090 2063.275 2001.370 2063.645 ;
        RECT 1925.200 2063.130 1925.460 2063.275 ;
        RECT 2001.100 2063.130 2001.360 2063.275 ;
        RECT 1794.560 2060.750 1794.820 2061.070 ;
        RECT 1753.160 2059.050 1753.420 2059.370 ;
        RECT 1745.800 2058.710 1746.060 2059.030 ;
        RECT 1738.900 2058.370 1739.160 2058.690 ;
        RECT 1732.000 2058.030 1732.260 2058.350 ;
        RECT 1725.100 2057.690 1725.360 2058.010 ;
        RECT 1718.200 2057.350 1718.460 2057.670 ;
        RECT 2028.690 2057.155 2028.970 2057.525 ;
        RECT 2028.760 2056.650 2028.900 2057.155 ;
        RECT 2028.700 2056.330 2028.960 2056.650 ;
        RECT 1715.440 2055.650 1715.700 2055.970 ;
        RECT 1704.400 2052.250 1704.660 2052.570 ;
        RECT 1697.500 1910.810 1697.760 1911.130 ;
        RECT 1414.140 1607.530 1414.400 1607.850 ;
        RECT 1693.820 1607.530 1694.080 1607.850 ;
        RECT 1414.200 1607.365 1414.340 1607.530 ;
        RECT 1414.130 1606.995 1414.410 1607.365 ;
      LAYER met2 ;
        RECT 1705.000 1605.000 2081.480 2051.235 ;
      LAYER met2 ;
        RECT 2081.660 1956.770 2081.800 2484.050 ;
        RECT 2087.120 2318.810 2087.380 2319.130 ;
        RECT 2083.900 2145.750 2084.160 2146.070 ;
        RECT 2083.960 1965.045 2084.100 2145.750 ;
        RECT 2087.180 2065.830 2087.320 2318.810 ;
        RECT 2087.120 2065.510 2087.380 2065.830 ;
        RECT 2083.890 1964.675 2084.170 1965.045 ;
        RECT 2082.050 1956.770 2082.330 1956.885 ;
        RECT 2081.660 1956.630 2082.330 1956.770 ;
        RECT 2082.050 1956.515 2082.330 1956.630 ;
        RECT 2097.760 1705.285 2097.900 2580.610 ;
        RECT 2098.160 2566.670 2098.420 2566.990 ;
        RECT 2098.220 1708.685 2098.360 2566.670 ;
        RECT 2098.620 2559.870 2098.880 2560.190 ;
        RECT 2098.680 1718.885 2098.820 2559.870 ;
        RECT 2099.080 2546.270 2099.340 2546.590 ;
        RECT 2099.140 1722.285 2099.280 2546.270 ;
        RECT 2099.540 2539.130 2099.800 2539.450 ;
        RECT 2099.600 1733.165 2099.740 2539.130 ;
        RECT 2100.000 2525.530 2100.260 2525.850 ;
        RECT 2099.530 1732.795 2099.810 1733.165 ;
        RECT 2099.070 1721.915 2099.350 1722.285 ;
        RECT 2098.610 1718.515 2098.890 1718.885 ;
        RECT 2098.150 1708.315 2098.430 1708.685 ;
        RECT 2097.690 1704.915 2097.970 1705.285 ;
        RECT 2097.760 1625.725 2097.900 1704.915 ;
        RECT 2098.220 1629.125 2098.360 1708.315 ;
        RECT 2098.680 1640.685 2098.820 1718.515 ;
        RECT 2099.140 1646.125 2099.280 1721.915 ;
        RECT 2099.600 1654.965 2099.740 1732.795 ;
        RECT 2100.060 1732.485 2100.200 2525.530 ;
        RECT 2100.460 2518.390 2100.720 2518.710 ;
        RECT 2100.520 1746.085 2100.660 2518.390 ;
        RECT 2176.820 2401.090 2177.080 2401.410 ;
        RECT 2156.120 2394.630 2156.380 2394.950 ;
        RECT 2149.220 2387.490 2149.480 2387.810 ;
        RECT 2142.320 2380.350 2142.580 2380.670 ;
        RECT 2121.620 2373.890 2121.880 2374.210 ;
        RECT 2121.680 2068.210 2121.820 2373.890 ;
        RECT 2135.420 2373.550 2135.680 2373.870 ;
        RECT 2121.620 2067.890 2121.880 2068.210 ;
        RECT 2135.480 2067.190 2135.620 2373.550 ;
        RECT 2142.380 2067.530 2142.520 2380.350 ;
        RECT 2142.320 2067.210 2142.580 2067.530 ;
        RECT 2135.420 2066.870 2135.680 2067.190 ;
        RECT 2149.280 2066.850 2149.420 2387.490 ;
        RECT 2156.180 2067.870 2156.320 2394.630 ;
        RECT 2169.920 2394.290 2170.180 2394.610 ;
        RECT 2156.120 2067.550 2156.380 2067.870 ;
        RECT 2149.220 2066.530 2149.480 2066.850 ;
        RECT 2169.980 2066.170 2170.120 2394.290 ;
        RECT 2176.880 2066.510 2177.020 2401.090 ;
        RECT 2190.680 2075.690 2190.820 3230.155 ;
        RECT 2191.070 3224.715 2191.350 3225.085 ;
        RECT 2190.620 2075.370 2190.880 2075.690 ;
        RECT 2191.140 2075.010 2191.280 3224.715 ;
        RECT 2191.530 3215.875 2191.810 3216.245 ;
        RECT 2191.600 2075.350 2191.740 3215.875 ;
        RECT 2191.990 3209.755 2192.270 3210.125 ;
        RECT 2191.540 2075.030 2191.800 2075.350 ;
        RECT 2191.080 2074.690 2191.340 2075.010 ;
        RECT 2192.060 2072.970 2192.200 3209.755 ;
        RECT 2192.450 3201.595 2192.730 3201.965 ;
        RECT 2192.520 2073.310 2192.660 3201.595 ;
        RECT 2192.910 3196.155 2193.190 3196.525 ;
        RECT 2192.980 2076.370 2193.120 3196.155 ;
        RECT 2193.370 3187.995 2193.650 3188.365 ;
        RECT 2192.920 2076.050 2193.180 2076.370 ;
        RECT 2193.440 2076.030 2193.580 3187.995 ;
        RECT 2193.830 2898.315 2194.110 2898.685 ;
        RECT 2193.380 2075.710 2193.640 2076.030 ;
        RECT 2192.460 2072.990 2192.720 2073.310 ;
        RECT 2192.000 2072.650 2192.260 2072.970 ;
        RECT 2176.820 2066.190 2177.080 2066.510 ;
        RECT 2169.920 2065.850 2170.180 2066.170 ;
        RECT 2193.900 2055.630 2194.040 2898.315 ;
      LAYER met2 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met2 ;
        RECT 2582.140 3249.565 2582.280 3252.110 ;
        RECT 2582.070 3249.195 2582.350 3249.565 ;
        RECT 2594.560 2946.965 2594.700 3263.670 ;
        RECT 2594.490 2946.595 2594.770 2946.965 ;
        RECT 2594.560 2938.805 2594.700 2946.595 ;
        RECT 2594.490 2938.435 2594.770 2938.805 ;
        RECT 2228.790 2794.275 2229.070 2794.645 ;
        RECT 2256.390 2794.275 2256.670 2794.645 ;
        RECT 2263.290 2794.275 2263.570 2794.645 ;
        RECT 2268.350 2794.275 2268.630 2794.645 ;
        RECT 2270.190 2794.275 2270.470 2794.645 ;
        RECT 2277.090 2794.275 2277.370 2794.645 ;
        RECT 2283.990 2794.275 2284.270 2794.645 ;
        RECT 2290.890 2794.275 2291.170 2794.645 ;
        RECT 2297.790 2794.275 2298.070 2794.645 ;
        RECT 2305.150 2794.275 2305.430 2794.645 ;
        RECT 2308.370 2794.275 2308.650 2794.645 ;
        RECT 2311.590 2794.275 2311.870 2794.645 ;
        RECT 2318.490 2794.275 2318.770 2794.645 ;
        RECT 2325.390 2794.275 2325.670 2794.645 ;
        RECT 2332.290 2794.275 2332.570 2794.645 ;
        RECT 2339.190 2794.275 2339.470 2794.645 ;
        RECT 2211.320 2408.570 2211.580 2408.890 ;
        RECT 2211.380 2065.490 2211.520 2408.570 ;
        RECT 2225.120 2408.230 2225.380 2408.550 ;
        RECT 2211.320 2065.170 2211.580 2065.490 ;
        RECT 2225.180 2065.150 2225.320 2408.230 ;
        RECT 2228.860 2074.670 2229.000 2794.275 ;
        RECT 2249.490 2788.835 2249.770 2789.205 ;
        RECT 2249.560 2788.670 2249.700 2788.835 ;
        RECT 2249.500 2788.350 2249.760 2788.670 ;
        RECT 2245.820 2421.830 2246.080 2422.150 ;
        RECT 2232.020 2415.030 2232.280 2415.350 ;
        RECT 2228.800 2074.350 2229.060 2074.670 ;
        RECT 2225.120 2064.830 2225.380 2065.150 ;
        RECT 2232.080 2064.810 2232.220 2415.030 ;
        RECT 2238.920 2325.270 2239.180 2325.590 ;
        RECT 2238.980 2069.910 2239.120 2325.270 ;
        RECT 2238.920 2069.590 2239.180 2069.910 ;
        RECT 2232.020 2064.490 2232.280 2064.810 ;
        RECT 2245.880 2064.470 2246.020 2421.830 ;
        RECT 2245.820 2064.150 2246.080 2064.470 ;
        RECT 2193.840 2055.310 2194.100 2055.630 ;
        RECT 2256.460 2055.290 2256.600 2794.275 ;
        RECT 2263.360 2060.050 2263.500 2794.275 ;
        RECT 2268.420 2794.110 2268.560 2794.275 ;
        RECT 2263.750 2793.595 2264.030 2793.965 ;
        RECT 2268.360 2793.790 2268.620 2794.110 ;
        RECT 2263.820 2074.330 2263.960 2793.595 ;
        RECT 2266.510 2792.915 2266.790 2793.285 ;
        RECT 2266.580 2792.750 2266.720 2792.915 ;
        RECT 2266.520 2792.430 2266.780 2792.750 ;
        RECT 2266.580 2082.150 2266.720 2792.430 ;
        RECT 2266.520 2081.830 2266.780 2082.150 ;
        RECT 2263.760 2074.010 2264.020 2074.330 ;
        RECT 2270.260 2072.630 2270.400 2794.275 ;
        RECT 2273.870 2793.595 2274.150 2793.965 ;
        RECT 2273.880 2793.450 2274.140 2793.595 ;
        RECT 2273.940 2792.410 2274.080 2793.450 ;
        RECT 2273.880 2792.090 2274.140 2792.410 ;
        RECT 2277.160 2081.810 2277.300 2794.275 ;
        RECT 2280.310 2793.595 2280.590 2793.965 ;
        RECT 2280.380 2793.430 2280.520 2793.595 ;
        RECT 2280.320 2793.110 2280.580 2793.430 ;
        RECT 2277.100 2081.490 2277.360 2081.810 ;
        RECT 2270.200 2072.310 2270.460 2072.630 ;
        RECT 2263.300 2059.730 2263.560 2060.050 ;
        RECT 2256.400 2054.970 2256.660 2055.290 ;
        RECT 2280.380 2054.950 2280.520 2793.110 ;
        RECT 2284.060 2081.470 2284.200 2794.275 ;
        RECT 2287.280 2794.110 2287.420 2794.265 ;
        RECT 2287.220 2793.965 2287.480 2794.110 ;
        RECT 2287.210 2793.595 2287.490 2793.965 ;
        RECT 2284.000 2081.150 2284.260 2081.470 ;
        RECT 2280.320 2054.630 2280.580 2054.950 ;
        RECT 2287.280 2054.610 2287.420 2793.595 ;
        RECT 2290.960 2081.130 2291.100 2794.275 ;
        RECT 2294.110 2793.595 2294.390 2793.965 ;
        RECT 2294.120 2793.450 2294.380 2793.595 ;
        RECT 2290.900 2080.810 2291.160 2081.130 ;
        RECT 2287.220 2054.290 2287.480 2054.610 ;
        RECT 2294.180 2054.270 2294.320 2793.450 ;
        RECT 2297.860 2080.790 2298.000 2794.275 ;
        RECT 2304.690 2793.595 2304.970 2793.965 ;
        RECT 2301.930 2792.915 2302.210 2793.285 ;
        RECT 2302.000 2788.670 2302.140 2792.915 ;
        RECT 2301.940 2788.350 2302.200 2788.670 ;
        RECT 2301.020 2788.010 2301.280 2788.330 ;
        RECT 2297.800 2080.470 2298.060 2080.790 ;
        RECT 2294.120 2053.950 2294.380 2054.270 ;
        RECT 2301.080 2053.930 2301.220 2788.010 ;
        RECT 2301.020 2053.610 2301.280 2053.930 ;
        RECT 2302.000 2053.590 2302.140 2788.350 ;
        RECT 2304.230 2788.155 2304.510 2788.525 ;
        RECT 2304.240 2788.010 2304.500 2788.155 ;
        RECT 2301.940 2053.270 2302.200 2053.590 ;
        RECT 2304.760 2053.250 2304.900 2793.595 ;
        RECT 2305.220 2080.450 2305.360 2794.275 ;
        RECT 2308.440 2792.750 2308.580 2794.275 ;
        RECT 2308.380 2792.430 2308.640 2792.750 ;
        RECT 2305.160 2080.130 2305.420 2080.450 ;
        RECT 2304.700 2052.930 2304.960 2053.250 ;
        RECT 2311.660 2052.910 2311.800 2794.275 ;
        RECT 2315.270 2793.595 2315.550 2793.965 ;
        RECT 2315.340 2793.090 2315.480 2793.595 ;
        RECT 2315.280 2792.770 2315.540 2793.090 ;
        RECT 2318.560 2060.390 2318.700 2794.275 ;
        RECT 2321.250 2793.595 2321.530 2793.965 ;
        RECT 2321.320 2792.410 2321.460 2793.595 ;
        RECT 2321.260 2792.090 2321.520 2792.410 ;
        RECT 2321.720 2787.670 2321.980 2787.990 ;
        RECT 2321.780 2152.870 2321.920 2787.670 ;
        RECT 2321.720 2152.550 2321.980 2152.870 ;
        RECT 2318.500 2060.070 2318.760 2060.390 ;
        RECT 2325.460 2059.710 2325.600 2794.275 ;
        RECT 2326.310 2793.595 2326.590 2793.965 ;
        RECT 2326.380 2793.430 2326.520 2793.595 ;
        RECT 2326.320 2793.110 2326.580 2793.430 ;
        RECT 2328.620 2429.310 2328.880 2429.630 ;
        RECT 2328.680 2063.450 2328.820 2429.310 ;
        RECT 2328.620 2063.130 2328.880 2063.450 ;
        RECT 2325.400 2059.390 2325.660 2059.710 ;
        RECT 2332.360 2056.310 2332.500 2794.275 ;
        RECT 2332.760 2793.965 2333.020 2794.110 ;
        RECT 2332.750 2793.595 2333.030 2793.965 ;
        RECT 2335.520 2428.970 2335.780 2429.290 ;
        RECT 2335.580 2063.790 2335.720 2428.970 ;
        RECT 2335.520 2063.470 2335.780 2063.790 ;
        RECT 2339.260 2060.730 2339.400 2794.275 ;
        RECT 2340.120 2794.130 2340.380 2794.450 ;
        RECT 2343.790 2794.275 2344.070 2794.645 ;
        RECT 2346.090 2794.275 2346.370 2794.645 ;
        RECT 2352.990 2794.275 2353.270 2794.645 ;
        RECT 2359.890 2794.275 2360.170 2794.645 ;
        RECT 2366.790 2794.275 2367.070 2794.645 ;
        RECT 2373.690 2794.275 2373.970 2794.645 ;
        RECT 2377.370 2794.275 2377.650 2794.645 ;
        RECT 2380.590 2794.275 2380.870 2794.645 ;
        RECT 2382.890 2794.275 2383.170 2794.645 ;
        RECT 2387.950 2794.275 2388.230 2794.645 ;
        RECT 2394.850 2794.275 2395.130 2794.645 ;
        RECT 2401.750 2794.275 2402.030 2794.645 ;
        RECT 2339.650 2793.595 2339.930 2793.965 ;
        RECT 2340.180 2793.770 2340.320 2794.130 ;
        RECT 2343.860 2793.770 2344.000 2794.275 ;
        RECT 2339.720 2073.990 2339.860 2793.595 ;
        RECT 2340.120 2793.450 2340.380 2793.770 ;
        RECT 2340.580 2793.450 2340.840 2793.770 ;
        RECT 2343.800 2793.450 2344.060 2793.770 ;
        RECT 2340.180 2793.285 2340.320 2793.450 ;
        RECT 2340.110 2792.915 2340.390 2793.285 ;
        RECT 2340.640 2788.670 2340.780 2793.450 ;
        RECT 2340.580 2788.350 2340.840 2788.670 ;
        RECT 2339.660 2073.670 2339.920 2073.990 ;
        RECT 2346.160 2073.650 2346.300 2794.275 ;
        RECT 2350.230 2792.915 2350.510 2793.285 ;
        RECT 2350.300 2788.330 2350.440 2792.915 ;
        RECT 2350.240 2788.010 2350.500 2788.330 ;
        RECT 2353.060 2076.710 2353.200 2794.275 ;
        RECT 2356.670 2793.595 2356.950 2793.965 ;
        RECT 2356.740 2792.750 2356.880 2793.595 ;
        RECT 2356.680 2792.430 2356.940 2792.750 ;
        RECT 2353.460 2332.070 2353.720 2332.390 ;
        RECT 2353.000 2076.390 2353.260 2076.710 ;
        RECT 2346.100 2073.330 2346.360 2073.650 ;
        RECT 2347.020 2069.590 2347.280 2069.910 ;
        RECT 2353.520 2069.765 2353.660 2332.070 ;
        RECT 2359.960 2077.050 2360.100 2794.275 ;
        RECT 2360.810 2793.595 2361.090 2793.965 ;
        RECT 2360.880 2793.090 2361.020 2793.595 ;
        RECT 2360.820 2792.770 2361.080 2793.090 ;
        RECT 2366.860 2083.850 2367.000 2794.275 ;
        RECT 2367.250 2793.595 2367.530 2793.965 ;
        RECT 2367.320 2792.410 2367.460 2793.595 ;
        RECT 2367.260 2792.090 2367.520 2792.410 ;
        RECT 2367.260 2339.210 2367.520 2339.530 ;
        RECT 2366.800 2083.530 2367.060 2083.850 ;
        RECT 2359.900 2076.730 2360.160 2077.050 ;
        RECT 2340.580 2065.510 2340.840 2065.830 ;
        RECT 2340.640 2063.645 2340.780 2065.510 ;
        RECT 2347.080 2063.645 2347.220 2069.590 ;
        RECT 2353.450 2069.395 2353.730 2069.765 ;
        RECT 2359.900 2068.570 2360.160 2068.890 ;
        RECT 2359.960 2063.645 2360.100 2068.570 ;
        RECT 2340.570 2063.275 2340.850 2063.645 ;
        RECT 2347.010 2063.275 2347.290 2063.645 ;
        RECT 2359.890 2063.275 2360.170 2063.645 ;
        RECT 2339.200 2060.410 2339.460 2060.730 ;
        RECT 2332.300 2055.990 2332.560 2056.310 ;
        RECT 2311.600 2052.590 2311.860 2052.910 ;
        RECT 2367.320 2052.085 2367.460 2339.210 ;
        RECT 2373.760 2090.650 2373.900 2794.275 ;
        RECT 2377.440 2794.110 2377.580 2794.275 ;
        RECT 2374.150 2793.595 2374.430 2793.965 ;
        RECT 2377.380 2793.790 2377.640 2794.110 ;
        RECT 2374.220 2793.430 2374.360 2793.595 ;
        RECT 2374.160 2793.110 2374.420 2793.430 ;
        RECT 2374.220 2788.670 2374.360 2793.110 ;
        RECT 2374.160 2788.350 2374.420 2788.670 ;
        RECT 2374.160 2346.010 2374.420 2346.330 ;
        RECT 2373.700 2090.330 2373.960 2090.650 ;
        RECT 2374.220 2069.765 2374.360 2346.010 ;
        RECT 2380.660 2097.450 2380.800 2794.275 ;
        RECT 2382.900 2794.130 2383.160 2794.275 ;
        RECT 2381.050 2792.915 2381.330 2793.285 ;
        RECT 2381.120 2792.070 2381.260 2792.915 ;
        RECT 2382.960 2792.070 2383.100 2794.130 ;
        RECT 2388.020 2793.770 2388.160 2794.275 ;
        RECT 2387.960 2793.450 2388.220 2793.770 ;
        RECT 2381.060 2791.750 2381.320 2792.070 ;
        RECT 2382.900 2791.750 2383.160 2792.070 ;
        RECT 2387.490 2791.555 2387.770 2791.925 ;
        RECT 2388.020 2791.730 2388.160 2793.450 ;
        RECT 2394.390 2792.235 2394.670 2792.605 ;
        RECT 2387.500 2791.410 2387.760 2791.555 ;
        RECT 2387.960 2791.410 2388.220 2791.730 ;
        RECT 2394.460 2791.390 2394.600 2792.235 ;
        RECT 2394.920 2791.390 2395.060 2794.275 ;
        RECT 2401.820 2792.750 2401.960 2794.275 ;
        RECT 2421.990 2793.595 2422.270 2793.965 ;
        RECT 2422.060 2793.430 2422.200 2793.595 ;
        RECT 2408.190 2792.915 2408.470 2793.285 ;
        RECT 2422.000 2793.110 2422.260 2793.430 ;
        RECT 2408.200 2792.770 2408.460 2792.915 ;
        RECT 2401.760 2792.430 2402.020 2792.750 ;
        RECT 2408.190 2792.235 2408.470 2792.605 ;
        RECT 2415.090 2792.235 2415.370 2792.605 ;
        RECT 2428.890 2792.235 2429.170 2792.605 ;
        RECT 2435.790 2792.235 2436.070 2792.605 ;
        RECT 2401.750 2791.555 2402.030 2791.925 ;
        RECT 2394.400 2791.070 2394.660 2791.390 ;
        RECT 2394.860 2791.070 2395.120 2791.390 ;
        RECT 2394.920 2788.330 2395.060 2791.070 ;
        RECT 2401.820 2791.050 2401.960 2791.555 ;
        RECT 2401.760 2790.730 2402.020 2791.050 ;
        RECT 2408.260 2790.370 2408.400 2792.235 ;
        RECT 2415.100 2792.090 2415.360 2792.235 ;
        RECT 2428.960 2792.070 2429.100 2792.235 ;
        RECT 2428.900 2791.750 2429.160 2792.070 ;
        RECT 2435.860 2791.730 2436.000 2792.235 ;
        RECT 2435.800 2791.410 2436.060 2791.730 ;
        RECT 2442.690 2791.555 2442.970 2791.925 ;
        RECT 2442.760 2791.390 2442.900 2791.555 ;
        RECT 2415.090 2790.875 2415.370 2791.245 ;
        RECT 2442.700 2791.070 2442.960 2791.390 ;
        RECT 2415.160 2790.710 2415.300 2790.875 ;
        RECT 2415.100 2790.390 2415.360 2790.710 ;
        RECT 2408.200 2790.050 2408.460 2790.370 ;
        RECT 2421.990 2790.195 2422.270 2790.565 ;
        RECT 2422.060 2790.030 2422.200 2790.195 ;
        RECT 2415.090 2789.515 2415.370 2789.885 ;
        RECT 2422.000 2789.710 2422.260 2790.030 ;
        RECT 2428.890 2789.515 2429.170 2789.885 ;
        RECT 2415.100 2789.370 2415.360 2789.515 ;
        RECT 2428.960 2789.350 2429.100 2789.515 ;
        RECT 2415.090 2788.835 2415.370 2789.205 ;
        RECT 2428.900 2789.030 2429.160 2789.350 ;
        RECT 2435.790 2788.835 2436.070 2789.205 ;
        RECT 2415.160 2788.670 2415.300 2788.835 ;
        RECT 2435.800 2788.690 2436.060 2788.835 ;
        RECT 2415.100 2788.350 2415.360 2788.670 ;
        RECT 2394.860 2788.010 2395.120 2788.330 ;
        RECT 2442.690 2788.155 2442.970 2788.525 ;
        RECT 2442.760 2787.990 2442.900 2788.155 ;
        RECT 2442.700 2787.670 2442.960 2787.990 ;
        RECT 2494.220 2477.250 2494.480 2477.570 ;
        RECT 2480.420 2470.110 2480.680 2470.430 ;
        RECT 2459.720 2463.650 2459.980 2463.970 ;
        RECT 2445.920 2456.510 2446.180 2456.830 ;
        RECT 2418.320 2449.710 2418.580 2450.030 ;
        RECT 2411.420 2442.570 2411.680 2442.890 ;
        RECT 2404.520 2435.770 2404.780 2436.090 ;
        RECT 2387.960 2359.950 2388.220 2360.270 ;
        RECT 2380.600 2097.130 2380.860 2097.450 ;
        RECT 2388.020 2069.765 2388.160 2359.950 ;
        RECT 2374.150 2069.395 2374.430 2069.765 ;
        RECT 2380.600 2069.250 2380.860 2069.570 ;
        RECT 2387.950 2069.395 2388.230 2069.765 ;
        RECT 2380.660 2069.085 2380.800 2069.250 ;
        RECT 2387.500 2069.085 2387.760 2069.230 ;
        RECT 2380.590 2068.715 2380.870 2069.085 ;
        RECT 2387.490 2068.715 2387.770 2069.085 ;
        RECT 2394.400 2068.405 2394.660 2068.550 ;
        RECT 2394.390 2068.035 2394.670 2068.405 ;
        RECT 2404.580 2068.210 2404.720 2435.770 ;
        RECT 2411.480 2068.550 2411.620 2442.570 ;
        RECT 2418.380 2069.230 2418.520 2449.710 ;
        RECT 2425.220 2449.370 2425.480 2449.690 ;
        RECT 2418.320 2068.910 2418.580 2069.230 ;
        RECT 2411.420 2068.230 2411.680 2068.550 ;
        RECT 2402.220 2067.890 2402.480 2068.210 ;
        RECT 2404.520 2067.890 2404.780 2068.210 ;
        RECT 2402.280 2067.725 2402.420 2067.890 ;
        RECT 2402.210 2067.355 2402.490 2067.725 ;
        RECT 2415.100 2067.210 2415.360 2067.530 ;
        RECT 2408.200 2067.045 2408.460 2067.190 ;
        RECT 2415.160 2067.045 2415.300 2067.210 ;
        RECT 2425.280 2067.190 2425.420 2449.370 ;
        RECT 2445.980 2069.570 2446.120 2456.510 ;
        RECT 2445.920 2069.250 2446.180 2069.570 ;
        RECT 2459.780 2068.890 2459.920 2463.650 ;
        RECT 2466.620 2463.310 2466.880 2463.630 ;
        RECT 2459.720 2068.570 2459.980 2068.890 ;
        RECT 2428.900 2067.725 2429.160 2067.870 ;
        RECT 2428.890 2067.355 2429.170 2067.725 ;
        RECT 2466.680 2067.530 2466.820 2463.310 ;
        RECT 2480.480 2069.910 2480.620 2470.110 ;
        RECT 2480.420 2069.590 2480.680 2069.910 ;
        RECT 2494.280 2068.550 2494.420 2477.250 ;
        RECT 2631.760 2318.470 2632.020 2318.790 ;
        RECT 2525.500 2069.590 2525.760 2069.910 ;
        RECT 2512.620 2069.250 2512.880 2069.570 ;
        RECT 2497.900 2068.910 2498.160 2069.230 ;
        RECT 2491.460 2068.230 2491.720 2068.550 ;
        RECT 2494.220 2068.230 2494.480 2068.550 ;
        RECT 2484.100 2067.890 2484.360 2068.210 ;
        RECT 2466.620 2067.210 2466.880 2067.530 ;
        RECT 2408.190 2066.675 2408.470 2067.045 ;
        RECT 2415.090 2066.675 2415.370 2067.045 ;
        RECT 2425.220 2066.870 2425.480 2067.190 ;
        RECT 2422.000 2066.530 2422.260 2066.850 ;
        RECT 2422.060 2066.365 2422.200 2066.530 ;
        RECT 2442.700 2066.365 2442.960 2066.510 ;
        RECT 2421.990 2065.995 2422.270 2066.365 ;
        RECT 2435.800 2065.850 2436.060 2066.170 ;
        RECT 2442.690 2065.995 2442.970 2066.365 ;
        RECT 2435.860 2065.685 2436.000 2065.850 ;
        RECT 2435.790 2065.315 2436.070 2065.685 ;
        RECT 2449.600 2065.170 2449.860 2065.490 ;
        RECT 2449.660 2065.005 2449.800 2065.170 ;
        RECT 2456.500 2065.005 2456.760 2065.150 ;
        RECT 2449.590 2064.635 2449.870 2065.005 ;
        RECT 2456.490 2064.635 2456.770 2065.005 ;
        RECT 2456.960 2064.490 2457.220 2064.810 ;
        RECT 2457.020 2063.645 2457.160 2064.490 ;
        RECT 2463.400 2064.150 2463.660 2064.470 ;
        RECT 2463.460 2063.645 2463.600 2064.150 ;
        RECT 2478.580 2063.645 2478.840 2063.790 ;
        RECT 2484.160 2063.645 2484.300 2067.890 ;
        RECT 2491.520 2063.645 2491.660 2068.230 ;
        RECT 2497.960 2063.645 2498.100 2068.910 ;
        RECT 2505.260 2066.870 2505.520 2067.190 ;
        RECT 2505.320 2063.645 2505.460 2066.870 ;
        RECT 2512.680 2063.645 2512.820 2069.250 ;
        RECT 2525.560 2069.085 2525.700 2069.590 ;
        RECT 2518.600 2068.570 2518.860 2068.890 ;
        RECT 2525.490 2068.715 2525.770 2069.085 ;
        RECT 2518.660 2063.645 2518.800 2068.570 ;
        RECT 2532.400 2068.405 2532.660 2068.550 ;
        RECT 2532.390 2068.035 2532.670 2068.405 ;
        RECT 2519.980 2067.210 2520.240 2067.530 ;
        RECT 2520.040 2063.645 2520.180 2067.210 ;
        RECT 2587.600 2063.810 2587.860 2064.130 ;
        RECT 2587.660 2063.645 2587.800 2063.810 ;
        RECT 2456.950 2063.275 2457.230 2063.645 ;
        RECT 2463.390 2063.275 2463.670 2063.645 ;
        RECT 2470.290 2063.275 2470.570 2063.645 ;
        RECT 2478.570 2063.275 2478.850 2063.645 ;
        RECT 2484.090 2063.275 2484.370 2063.645 ;
        RECT 2491.450 2063.275 2491.730 2063.645 ;
        RECT 2497.890 2063.275 2498.170 2063.645 ;
        RECT 2505.250 2063.275 2505.530 2063.645 ;
        RECT 2512.610 2063.275 2512.890 2063.645 ;
        RECT 2518.590 2063.275 2518.870 2063.645 ;
        RECT 2519.970 2063.275 2520.250 2063.645 ;
        RECT 2587.590 2063.275 2587.870 2063.645 ;
        RECT 2470.300 2063.130 2470.560 2063.275 ;
        RECT 2367.250 2051.715 2367.530 2052.085 ;
        RECT 2100.450 1745.715 2100.730 1746.085 ;
        RECT 2099.990 1732.115 2100.270 1732.485 ;
        RECT 2100.060 1660.405 2100.200 1732.115 ;
        RECT 2100.520 1668.565 2100.660 1745.715 ;
        RECT 2100.450 1668.195 2100.730 1668.565 ;
        RECT 2099.990 1660.035 2100.270 1660.405 ;
        RECT 2099.530 1654.595 2099.810 1654.965 ;
        RECT 2099.070 1645.755 2099.350 1646.125 ;
        RECT 2098.610 1640.315 2098.890 1640.685 ;
        RECT 2098.150 1628.755 2098.430 1629.125 ;
        RECT 2097.690 1625.355 2097.970 1625.725 ;
      LAYER met2 ;
        RECT 2255.000 1605.000 2631.480 2051.235 ;
      LAYER met2 ;
        RECT 2631.820 2049.930 2631.960 2318.470 ;
        RECT 2632.210 2049.930 2632.490 2050.045 ;
        RECT 2631.820 2049.790 2632.490 2049.930 ;
        RECT 2632.210 2049.675 2632.490 2049.790 ;
        RECT 1396.650 1604.530 1396.930 1604.645 ;
        RECT 1395.800 1604.390 1396.930 1604.530 ;
      LAYER met2 ;
        RECT 300.090 1602.195 304.410 1604.280 ;
        RECT 305.250 1602.195 314.070 1604.280 ;
        RECT 314.910 1602.195 323.730 1604.280 ;
        RECT 324.570 1602.195 333.390 1604.280 ;
        RECT 334.230 1602.195 343.050 1604.280 ;
        RECT 343.890 1602.195 352.710 1604.280 ;
        RECT 353.550 1602.195 362.370 1604.280 ;
        RECT 363.210 1602.195 372.490 1604.280 ;
        RECT 373.330 1602.195 382.150 1604.280 ;
        RECT 382.990 1602.195 391.810 1604.280 ;
        RECT 392.650 1602.195 401.470 1604.280 ;
        RECT 402.310 1602.195 411.130 1604.280 ;
        RECT 411.970 1602.195 420.790 1604.280 ;
        RECT 421.630 1602.195 430.910 1604.280 ;
        RECT 431.750 1602.195 440.570 1604.280 ;
        RECT 441.410 1602.195 450.230 1604.280 ;
        RECT 451.070 1602.195 459.890 1604.280 ;
        RECT 460.730 1602.195 469.550 1604.280 ;
        RECT 470.390 1602.195 479.210 1604.280 ;
        RECT 480.050 1602.195 489.330 1604.280 ;
        RECT 490.170 1602.195 498.990 1604.280 ;
        RECT 499.830 1602.195 508.650 1604.280 ;
        RECT 509.490 1602.195 518.310 1604.280 ;
        RECT 519.150 1602.195 527.970 1604.280 ;
        RECT 528.810 1602.195 537.630 1604.280 ;
        RECT 538.470 1602.195 547.290 1604.280 ;
        RECT 548.130 1602.195 557.410 1604.280 ;
        RECT 558.250 1602.195 567.070 1604.280 ;
        RECT 567.910 1602.195 576.730 1604.280 ;
        RECT 577.570 1602.195 586.390 1604.280 ;
        RECT 587.230 1602.195 596.050 1604.280 ;
        RECT 596.890 1602.195 605.710 1604.280 ;
        RECT 606.550 1602.195 615.830 1604.280 ;
        RECT 616.670 1602.195 625.490 1604.280 ;
        RECT 626.330 1602.195 635.150 1604.280 ;
        RECT 635.990 1602.195 644.810 1604.280 ;
        RECT 645.650 1602.195 654.470 1604.280 ;
        RECT 655.310 1602.195 664.130 1604.280 ;
        RECT 664.970 1602.195 674.250 1604.280 ;
        RECT 675.090 1602.195 683.910 1604.280 ;
        RECT 684.750 1602.195 693.570 1604.280 ;
        RECT 694.410 1602.195 703.230 1604.280 ;
        RECT 704.070 1602.195 712.890 1604.280 ;
        RECT 713.730 1602.195 722.550 1604.280 ;
        RECT 723.390 1602.195 732.670 1604.280 ;
        RECT 733.510 1602.195 742.330 1604.280 ;
        RECT 743.170 1602.195 751.990 1604.280 ;
        RECT 752.830 1602.195 761.650 1604.280 ;
        RECT 762.490 1602.195 771.310 1604.280 ;
        RECT 772.150 1602.195 780.970 1604.280 ;
        RECT 781.810 1602.195 790.630 1604.280 ;
        RECT 791.470 1602.195 800.750 1604.280 ;
        RECT 801.590 1602.195 810.410 1604.280 ;
        RECT 811.250 1602.195 820.070 1604.280 ;
        RECT 820.910 1602.195 829.730 1604.280 ;
        RECT 830.570 1602.195 839.390 1604.280 ;
        RECT 840.230 1602.195 849.050 1604.280 ;
        RECT 849.890 1602.195 859.170 1604.280 ;
        RECT 860.010 1602.195 868.830 1604.280 ;
        RECT 869.670 1602.195 878.490 1604.280 ;
        RECT 879.330 1602.195 888.150 1604.280 ;
        RECT 888.990 1602.195 897.810 1604.280 ;
        RECT 898.650 1602.195 907.470 1604.280 ;
        RECT 908.310 1602.195 917.590 1604.280 ;
        RECT 918.430 1602.195 927.250 1604.280 ;
        RECT 928.090 1602.195 936.910 1604.280 ;
        RECT 937.750 1602.195 946.570 1604.280 ;
        RECT 947.410 1602.195 956.230 1604.280 ;
        RECT 957.070 1602.195 965.890 1604.280 ;
        RECT 966.730 1602.195 975.550 1604.280 ;
        RECT 976.390 1602.195 985.670 1604.280 ;
        RECT 986.510 1602.195 995.330 1604.280 ;
        RECT 996.170 1602.195 1004.990 1604.280 ;
        RECT 1005.830 1602.195 1014.650 1604.280 ;
        RECT 1015.490 1602.195 1024.310 1604.280 ;
        RECT 1025.150 1602.195 1033.970 1604.280 ;
        RECT 1034.810 1602.195 1044.090 1604.280 ;
        RECT 1044.930 1602.195 1053.750 1604.280 ;
        RECT 1054.590 1602.195 1063.410 1604.280 ;
        RECT 1064.250 1602.195 1073.070 1604.280 ;
        RECT 1073.910 1602.195 1082.730 1604.280 ;
        RECT 1083.570 1602.195 1092.390 1604.280 ;
        RECT 1093.230 1602.195 1102.510 1604.280 ;
        RECT 1103.350 1602.195 1112.170 1604.280 ;
        RECT 1113.010 1602.195 1121.830 1604.280 ;
        RECT 1122.670 1602.195 1131.490 1604.280 ;
        RECT 1132.330 1602.195 1141.150 1604.280 ;
        RECT 1141.990 1602.195 1150.810 1604.280 ;
        RECT 1151.650 1602.195 1160.930 1604.280 ;
        RECT 1161.770 1602.195 1170.590 1604.280 ;
        RECT 1171.430 1602.195 1180.250 1604.280 ;
        RECT 1181.090 1602.195 1189.910 1604.280 ;
        RECT 1190.750 1602.195 1199.570 1604.280 ;
        RECT 1200.410 1602.195 1209.230 1604.280 ;
        RECT 1210.070 1602.195 1218.890 1604.280 ;
        RECT 1219.730 1602.195 1229.010 1604.280 ;
        RECT 1229.850 1602.195 1238.670 1604.280 ;
        RECT 1239.510 1602.195 1248.330 1604.280 ;
        RECT 1249.170 1602.195 1257.990 1604.280 ;
        RECT 1258.830 1602.195 1267.650 1604.280 ;
        RECT 1268.490 1602.195 1277.310 1604.280 ;
        RECT 1278.150 1602.195 1287.430 1604.280 ;
        RECT 1288.270 1602.195 1297.090 1604.280 ;
        RECT 1297.930 1602.195 1306.750 1604.280 ;
        RECT 1307.590 1602.195 1316.410 1604.280 ;
        RECT 1317.250 1602.195 1326.070 1604.280 ;
        RECT 1326.910 1602.195 1335.730 1604.280 ;
        RECT 1336.570 1602.195 1345.850 1604.280 ;
        RECT 1346.690 1602.195 1355.510 1604.280 ;
        RECT 1356.350 1602.195 1365.170 1604.280 ;
        RECT 1366.010 1602.195 1374.830 1604.280 ;
        RECT 1375.670 1602.195 1384.490 1604.280 ;
        RECT 1385.330 1602.195 1394.150 1604.280 ;
        RECT 1394.990 1602.195 1395.630 1604.280 ;
      LAYER met2 ;
        RECT 1396.650 1604.275 1396.930 1604.390 ;
        RECT 1555.150 1496.000 1555.430 1500.000 ;
        RECT 1565.270 1496.000 1565.550 1500.000 ;
        RECT 1575.850 1496.000 1576.130 1500.000 ;
        RECT 1585.970 1496.000 1586.250 1500.000 ;
        RECT 1596.550 1496.000 1596.830 1500.000 ;
        RECT 1606.670 1496.000 1606.950 1500.000 ;
        RECT 1617.250 1496.000 1617.530 1500.000 ;
        RECT 1627.370 1496.000 1627.650 1500.000 ;
        RECT 1637.950 1496.000 1638.230 1500.000 ;
        RECT 1648.530 1496.000 1648.810 1500.000 ;
        RECT 1658.650 1496.000 1658.930 1500.000 ;
        RECT 1669.230 1496.000 1669.510 1500.000 ;
        RECT 1679.350 1496.000 1679.630 1500.000 ;
        RECT 1689.930 1496.000 1690.210 1500.000 ;
        RECT 1700.050 1496.000 1700.330 1500.000 ;
        RECT 1710.630 1496.000 1710.910 1500.000 ;
        RECT 1720.750 1496.000 1721.030 1500.000 ;
        RECT 1731.330 1496.000 1731.610 1500.000 ;
        RECT 1741.910 1496.000 1742.190 1500.000 ;
        RECT 1752.030 1496.000 1752.310 1500.000 ;
        RECT 1762.610 1496.000 1762.890 1500.000 ;
        RECT 1772.730 1496.000 1773.010 1500.000 ;
        RECT 1783.310 1496.000 1783.590 1500.000 ;
        RECT 1793.430 1496.000 1793.710 1500.000 ;
        RECT 1804.010 1496.000 1804.290 1500.000 ;
        RECT 1814.130 1496.000 1814.410 1500.000 ;
        RECT 1824.710 1496.000 1824.990 1500.000 ;
        RECT 1835.290 1496.000 1835.570 1500.000 ;
        RECT 1845.410 1496.000 1845.690 1500.000 ;
        RECT 1855.990 1496.000 1856.270 1500.000 ;
        RECT 1866.110 1496.000 1866.390 1500.000 ;
        RECT 1876.690 1496.000 1876.970 1500.000 ;
        RECT 1886.810 1496.000 1887.090 1500.000 ;
        RECT 1897.390 1496.000 1897.670 1500.000 ;
        RECT 1907.510 1496.000 1907.790 1500.000 ;
        RECT 1918.090 1496.000 1918.370 1500.000 ;
        RECT 1928.670 1496.000 1928.950 1500.000 ;
        RECT 1938.790 1496.000 1939.070 1500.000 ;
        RECT 1949.370 1496.000 1949.650 1500.000 ;
        RECT 1959.490 1496.000 1959.770 1500.000 ;
        RECT 1970.070 1496.000 1970.350 1500.000 ;
        RECT 1980.190 1496.000 1980.470 1500.000 ;
        RECT 1990.770 1496.000 1991.050 1500.000 ;
        RECT 2000.890 1496.000 2001.170 1500.000 ;
        RECT 2011.470 1496.000 2011.750 1500.000 ;
        RECT 2022.050 1496.000 2022.330 1500.000 ;
        RECT 2032.170 1496.000 2032.450 1500.000 ;
        RECT 2042.750 1496.000 2043.030 1500.000 ;
        RECT 2052.870 1496.000 2053.150 1500.000 ;
        RECT 2063.450 1496.000 2063.730 1500.000 ;
        RECT 2073.570 1496.000 2073.850 1500.000 ;
        RECT 2084.150 1496.000 2084.430 1500.000 ;
        RECT 2094.270 1496.000 2094.550 1500.000 ;
        RECT 2104.850 1496.000 2105.130 1500.000 ;
        RECT 2115.430 1496.000 2115.710 1500.000 ;
        RECT 2125.550 1496.000 2125.830 1500.000 ;
        RECT 2136.130 1496.000 2136.410 1500.000 ;
        RECT 2146.250 1496.000 2146.530 1500.000 ;
        RECT 2156.830 1496.000 2157.110 1500.000 ;
        RECT 2166.950 1496.000 2167.230 1500.000 ;
        RECT 2177.530 1496.000 2177.810 1500.000 ;
        RECT 2187.650 1496.000 2187.930 1500.000 ;
        RECT 2198.230 1496.000 2198.510 1500.000 ;
        RECT 2208.810 1496.000 2209.090 1500.000 ;
        RECT 2218.930 1496.000 2219.210 1500.000 ;
        RECT 2229.510 1496.000 2229.790 1500.000 ;
        RECT 2239.630 1496.000 2239.910 1500.000 ;
        RECT 2250.210 1496.000 2250.490 1500.000 ;
        RECT 2260.330 1496.000 2260.610 1500.000 ;
        RECT 2270.910 1496.000 2271.190 1500.000 ;
        RECT 2281.030 1496.000 2281.310 1500.000 ;
        RECT 2291.610 1496.000 2291.890 1500.000 ;
        RECT 2302.190 1496.000 2302.470 1500.000 ;
        RECT 2312.310 1496.000 2312.590 1500.000 ;
        RECT 2322.890 1496.000 2323.170 1500.000 ;
        RECT 2333.010 1496.000 2333.290 1500.000 ;
        RECT 2343.590 1496.000 2343.870 1500.000 ;
        RECT 2353.710 1496.000 2353.990 1500.000 ;
        RECT 2364.290 1496.000 2364.570 1500.000 ;
        RECT 2374.410 1496.000 2374.690 1500.000 ;
        RECT 2384.990 1496.000 2385.270 1500.000 ;
        RECT 2395.570 1496.000 2395.850 1500.000 ;
        RECT 2405.690 1496.000 2405.970 1500.000 ;
        RECT 2416.270 1496.000 2416.550 1500.000 ;
        RECT 2426.390 1496.000 2426.670 1500.000 ;
        RECT 2436.970 1496.000 2437.250 1500.000 ;
        RECT 2447.090 1496.000 2447.370 1500.000 ;
        RECT 2457.670 1496.000 2457.950 1500.000 ;
        RECT 2467.790 1496.000 2468.070 1500.000 ;
        RECT 2478.370 1496.000 2478.650 1500.000 ;
        RECT 2488.950 1496.000 2489.230 1500.000 ;
        RECT 2499.070 1496.000 2499.350 1500.000 ;
        RECT 2509.650 1496.000 2509.930 1500.000 ;
        RECT 2519.770 1496.000 2520.050 1500.000 ;
        RECT 2530.350 1496.000 2530.630 1500.000 ;
        RECT 2540.470 1496.000 2540.750 1500.000 ;
        RECT 2551.050 1496.000 2551.330 1500.000 ;
        RECT 2561.170 1496.000 2561.450 1500.000 ;
        RECT 2571.750 1496.000 2572.030 1500.000 ;
        RECT 2582.330 1496.000 2582.610 1500.000 ;
        RECT 2592.450 1496.000 2592.730 1500.000 ;
        RECT 2603.030 1496.000 2603.310 1500.000 ;
        RECT 2613.150 1496.000 2613.430 1500.000 ;
        RECT 2623.730 1496.000 2624.010 1500.000 ;
        RECT 2633.850 1496.000 2634.130 1500.000 ;
        RECT 2644.430 1496.000 2644.710 1500.000 ;
      LAYER met2 ;
        RECT 1550.090 1495.720 1554.870 1496.000 ;
        RECT 1555.710 1495.720 1564.990 1496.000 ;
        RECT 1565.830 1495.720 1575.570 1496.000 ;
        RECT 1576.410 1495.720 1585.690 1496.000 ;
        RECT 1586.530 1495.720 1596.270 1496.000 ;
        RECT 1597.110 1495.720 1606.390 1496.000 ;
        RECT 1607.230 1495.720 1616.970 1496.000 ;
        RECT 1617.810 1495.720 1627.090 1496.000 ;
        RECT 1627.930 1495.720 1637.670 1496.000 ;
        RECT 1638.510 1495.720 1648.250 1496.000 ;
        RECT 1649.090 1495.720 1658.370 1496.000 ;
        RECT 1659.210 1495.720 1668.950 1496.000 ;
        RECT 1669.790 1495.720 1679.070 1496.000 ;
        RECT 1679.910 1495.720 1689.650 1496.000 ;
        RECT 1690.490 1495.720 1699.770 1496.000 ;
        RECT 1700.610 1495.720 1710.350 1496.000 ;
        RECT 1711.190 1495.720 1720.470 1496.000 ;
        RECT 1721.310 1495.720 1731.050 1496.000 ;
        RECT 1731.890 1495.720 1741.630 1496.000 ;
        RECT 1742.470 1495.720 1751.750 1496.000 ;
        RECT 1752.590 1495.720 1762.330 1496.000 ;
        RECT 1763.170 1495.720 1772.450 1496.000 ;
        RECT 1773.290 1495.720 1783.030 1496.000 ;
        RECT 1783.870 1495.720 1793.150 1496.000 ;
        RECT 1793.990 1495.720 1803.730 1496.000 ;
        RECT 1804.570 1495.720 1813.850 1496.000 ;
        RECT 1814.690 1495.720 1824.430 1496.000 ;
        RECT 1825.270 1495.720 1835.010 1496.000 ;
        RECT 1835.850 1495.720 1845.130 1496.000 ;
        RECT 1845.970 1495.720 1855.710 1496.000 ;
        RECT 1856.550 1495.720 1865.830 1496.000 ;
        RECT 1866.670 1495.720 1876.410 1496.000 ;
        RECT 1877.250 1495.720 1886.530 1496.000 ;
        RECT 1887.370 1495.720 1897.110 1496.000 ;
        RECT 1897.950 1495.720 1907.230 1496.000 ;
        RECT 1908.070 1495.720 1917.810 1496.000 ;
        RECT 1918.650 1495.720 1928.390 1496.000 ;
        RECT 1929.230 1495.720 1938.510 1496.000 ;
        RECT 1939.350 1495.720 1949.090 1496.000 ;
        RECT 1949.930 1495.720 1959.210 1496.000 ;
        RECT 1960.050 1495.720 1969.790 1496.000 ;
        RECT 1970.630 1495.720 1979.910 1496.000 ;
        RECT 1980.750 1495.720 1990.490 1496.000 ;
        RECT 1991.330 1495.720 2000.610 1496.000 ;
        RECT 2001.450 1495.720 2011.190 1496.000 ;
        RECT 2012.030 1495.720 2021.770 1496.000 ;
        RECT 2022.610 1495.720 2031.890 1496.000 ;
        RECT 2032.730 1495.720 2042.470 1496.000 ;
        RECT 2043.310 1495.720 2052.590 1496.000 ;
        RECT 2053.430 1495.720 2063.170 1496.000 ;
        RECT 2064.010 1495.720 2073.290 1496.000 ;
        RECT 2074.130 1495.720 2083.870 1496.000 ;
        RECT 2084.710 1495.720 2093.990 1496.000 ;
        RECT 2094.830 1495.720 2104.570 1496.000 ;
        RECT 2105.410 1495.720 2115.150 1496.000 ;
        RECT 2115.990 1495.720 2125.270 1496.000 ;
        RECT 2126.110 1495.720 2135.850 1496.000 ;
        RECT 2136.690 1495.720 2145.970 1496.000 ;
        RECT 2146.810 1495.720 2156.550 1496.000 ;
        RECT 2157.390 1495.720 2166.670 1496.000 ;
        RECT 2167.510 1495.720 2177.250 1496.000 ;
        RECT 2178.090 1495.720 2187.370 1496.000 ;
        RECT 2188.210 1495.720 2197.950 1496.000 ;
        RECT 2198.790 1495.720 2208.530 1496.000 ;
        RECT 2209.370 1495.720 2218.650 1496.000 ;
        RECT 2219.490 1495.720 2229.230 1496.000 ;
        RECT 2230.070 1495.720 2239.350 1496.000 ;
        RECT 2240.190 1495.720 2249.930 1496.000 ;
        RECT 2250.770 1495.720 2260.050 1496.000 ;
        RECT 2260.890 1495.720 2270.630 1496.000 ;
        RECT 2271.470 1495.720 2280.750 1496.000 ;
        RECT 2281.590 1495.720 2291.330 1496.000 ;
        RECT 2292.170 1495.720 2301.910 1496.000 ;
        RECT 2302.750 1495.720 2312.030 1496.000 ;
        RECT 2312.870 1495.720 2322.610 1496.000 ;
        RECT 2323.450 1495.720 2332.730 1496.000 ;
        RECT 2333.570 1495.720 2343.310 1496.000 ;
        RECT 2344.150 1495.720 2353.430 1496.000 ;
        RECT 2354.270 1495.720 2364.010 1496.000 ;
        RECT 2364.850 1495.720 2374.130 1496.000 ;
        RECT 2374.970 1495.720 2384.710 1496.000 ;
        RECT 2385.550 1495.720 2395.290 1496.000 ;
        RECT 2396.130 1495.720 2405.410 1496.000 ;
        RECT 2406.250 1495.720 2415.990 1496.000 ;
        RECT 2416.830 1495.720 2426.110 1496.000 ;
        RECT 2426.950 1495.720 2436.690 1496.000 ;
        RECT 2437.530 1495.720 2446.810 1496.000 ;
        RECT 2447.650 1495.720 2457.390 1496.000 ;
        RECT 2458.230 1495.720 2467.510 1496.000 ;
        RECT 2468.350 1495.720 2478.090 1496.000 ;
        RECT 2478.930 1495.720 2488.670 1496.000 ;
        RECT 2489.510 1495.720 2498.790 1496.000 ;
        RECT 2499.630 1495.720 2509.370 1496.000 ;
        RECT 2510.210 1495.720 2519.490 1496.000 ;
        RECT 2520.330 1495.720 2530.070 1496.000 ;
        RECT 2530.910 1495.720 2540.190 1496.000 ;
        RECT 2541.030 1495.720 2550.770 1496.000 ;
        RECT 2551.610 1495.720 2560.890 1496.000 ;
        RECT 2561.730 1495.720 2571.470 1496.000 ;
        RECT 2572.310 1495.720 2582.050 1496.000 ;
        RECT 2582.890 1495.720 2592.170 1496.000 ;
        RECT 2593.010 1495.720 2602.750 1496.000 ;
        RECT 2603.590 1495.720 2612.870 1496.000 ;
        RECT 2613.710 1495.720 2623.450 1496.000 ;
        RECT 2624.290 1495.720 2633.570 1496.000 ;
        RECT 2634.410 1495.720 2644.150 1496.000 ;
        RECT 2644.990 1495.720 2645.630 1496.000 ;
        RECT 1550.090 404.280 2645.630 1495.720 ;
        RECT 1550.090 402.195 1554.410 404.280 ;
      LAYER met2 ;
        RECT 1554.690 400.000 1554.970 404.000 ;
      LAYER met2 ;
        RECT 1555.250 402.195 1564.070 404.280 ;
      LAYER met2 ;
        RECT 1564.350 400.000 1564.630 404.000 ;
      LAYER met2 ;
        RECT 1564.910 402.195 1573.730 404.280 ;
      LAYER met2 ;
        RECT 1574.010 400.000 1574.290 404.000 ;
      LAYER met2 ;
        RECT 1574.570 402.195 1583.390 404.280 ;
      LAYER met2 ;
        RECT 1583.670 400.000 1583.950 404.000 ;
      LAYER met2 ;
        RECT 1584.230 402.195 1593.050 404.280 ;
      LAYER met2 ;
        RECT 1593.330 400.000 1593.610 404.000 ;
      LAYER met2 ;
        RECT 1593.890 402.195 1602.710 404.280 ;
      LAYER met2 ;
        RECT 1602.990 400.000 1603.270 404.000 ;
      LAYER met2 ;
        RECT 1603.550 402.195 1612.370 404.280 ;
      LAYER met2 ;
        RECT 1612.650 400.000 1612.930 404.000 ;
      LAYER met2 ;
        RECT 1613.210 402.195 1622.490 404.280 ;
      LAYER met2 ;
        RECT 1622.770 400.000 1623.050 404.000 ;
      LAYER met2 ;
        RECT 1623.330 402.195 1632.150 404.280 ;
      LAYER met2 ;
        RECT 1632.430 400.000 1632.710 404.000 ;
      LAYER met2 ;
        RECT 1632.990 402.195 1641.810 404.280 ;
      LAYER met2 ;
        RECT 1642.090 400.000 1642.370 404.000 ;
      LAYER met2 ;
        RECT 1642.650 402.195 1651.470 404.280 ;
      LAYER met2 ;
        RECT 1651.750 400.000 1652.030 404.000 ;
      LAYER met2 ;
        RECT 1652.310 402.195 1661.130 404.280 ;
      LAYER met2 ;
        RECT 1661.410 400.000 1661.690 404.000 ;
      LAYER met2 ;
        RECT 1661.970 402.195 1670.790 404.280 ;
      LAYER met2 ;
        RECT 1671.070 400.000 1671.350 404.000 ;
      LAYER met2 ;
        RECT 1671.630 402.195 1680.910 404.280 ;
      LAYER met2 ;
        RECT 1681.190 400.000 1681.470 404.000 ;
      LAYER met2 ;
        RECT 1681.750 402.195 1690.570 404.280 ;
      LAYER met2 ;
        RECT 1690.850 400.000 1691.130 404.000 ;
      LAYER met2 ;
        RECT 1691.410 402.195 1700.230 404.280 ;
      LAYER met2 ;
        RECT 1700.510 400.000 1700.790 404.000 ;
      LAYER met2 ;
        RECT 1701.070 402.195 1709.890 404.280 ;
      LAYER met2 ;
        RECT 1710.170 400.000 1710.450 404.000 ;
      LAYER met2 ;
        RECT 1710.730 402.195 1719.550 404.280 ;
      LAYER met2 ;
        RECT 1719.830 400.000 1720.110 404.000 ;
      LAYER met2 ;
        RECT 1720.390 402.195 1729.210 404.280 ;
      LAYER met2 ;
        RECT 1729.490 400.000 1729.770 404.000 ;
      LAYER met2 ;
        RECT 1730.050 402.195 1739.330 404.280 ;
      LAYER met2 ;
        RECT 1739.610 400.000 1739.890 404.000 ;
      LAYER met2 ;
        RECT 1740.170 402.195 1748.990 404.280 ;
      LAYER met2 ;
        RECT 1749.270 400.000 1749.550 404.000 ;
      LAYER met2 ;
        RECT 1749.830 402.195 1758.650 404.280 ;
      LAYER met2 ;
        RECT 1758.930 400.000 1759.210 404.000 ;
      LAYER met2 ;
        RECT 1759.490 402.195 1768.310 404.280 ;
      LAYER met2 ;
        RECT 1768.590 400.000 1768.870 404.000 ;
      LAYER met2 ;
        RECT 1769.150 402.195 1777.970 404.280 ;
      LAYER met2 ;
        RECT 1778.250 400.000 1778.530 404.000 ;
      LAYER met2 ;
        RECT 1778.810 402.195 1787.630 404.280 ;
      LAYER met2 ;
        RECT 1787.910 400.000 1788.190 404.000 ;
      LAYER met2 ;
        RECT 1788.470 402.195 1797.290 404.280 ;
      LAYER met2 ;
        RECT 1797.570 400.000 1797.850 404.000 ;
      LAYER met2 ;
        RECT 1798.130 402.195 1807.410 404.280 ;
      LAYER met2 ;
        RECT 1807.690 400.000 1807.970 404.000 ;
      LAYER met2 ;
        RECT 1808.250 402.195 1817.070 404.280 ;
      LAYER met2 ;
        RECT 1817.350 400.000 1817.630 404.000 ;
      LAYER met2 ;
        RECT 1817.910 402.195 1826.730 404.280 ;
      LAYER met2 ;
        RECT 1827.010 400.000 1827.290 404.000 ;
      LAYER met2 ;
        RECT 1827.570 402.195 1836.390 404.280 ;
      LAYER met2 ;
        RECT 1836.670 400.000 1836.950 404.000 ;
      LAYER met2 ;
        RECT 1837.230 402.195 1846.050 404.280 ;
      LAYER met2 ;
        RECT 1846.330 400.000 1846.610 404.000 ;
      LAYER met2 ;
        RECT 1846.890 402.195 1855.710 404.280 ;
      LAYER met2 ;
        RECT 1855.990 400.000 1856.270 404.000 ;
      LAYER met2 ;
        RECT 1856.550 402.195 1865.830 404.280 ;
      LAYER met2 ;
        RECT 1866.110 400.000 1866.390 404.000 ;
      LAYER met2 ;
        RECT 1866.670 402.195 1875.490 404.280 ;
      LAYER met2 ;
        RECT 1875.770 400.000 1876.050 404.000 ;
      LAYER met2 ;
        RECT 1876.330 402.195 1885.150 404.280 ;
      LAYER met2 ;
        RECT 1885.430 400.000 1885.710 404.000 ;
      LAYER met2 ;
        RECT 1885.990 402.195 1894.810 404.280 ;
      LAYER met2 ;
        RECT 1895.090 400.000 1895.370 404.000 ;
      LAYER met2 ;
        RECT 1895.650 402.195 1904.470 404.280 ;
      LAYER met2 ;
        RECT 1904.750 400.000 1905.030 404.000 ;
      LAYER met2 ;
        RECT 1905.310 402.195 1914.130 404.280 ;
      LAYER met2 ;
        RECT 1914.410 400.000 1914.690 404.000 ;
      LAYER met2 ;
        RECT 1914.970 402.195 1924.250 404.280 ;
      LAYER met2 ;
        RECT 1924.530 400.000 1924.810 404.000 ;
      LAYER met2 ;
        RECT 1925.090 402.195 1933.910 404.280 ;
      LAYER met2 ;
        RECT 1934.190 400.000 1934.470 404.000 ;
      LAYER met2 ;
        RECT 1934.750 402.195 1943.570 404.280 ;
      LAYER met2 ;
        RECT 1943.850 400.000 1944.130 404.000 ;
      LAYER met2 ;
        RECT 1944.410 402.195 1953.230 404.280 ;
      LAYER met2 ;
        RECT 1953.510 400.000 1953.790 404.000 ;
      LAYER met2 ;
        RECT 1954.070 402.195 1962.890 404.280 ;
      LAYER met2 ;
        RECT 1963.170 400.000 1963.450 404.000 ;
      LAYER met2 ;
        RECT 1963.730 402.195 1972.550 404.280 ;
      LAYER met2 ;
        RECT 1972.830 400.000 1973.110 404.000 ;
      LAYER met2 ;
        RECT 1973.390 402.195 1982.670 404.280 ;
      LAYER met2 ;
        RECT 1982.950 400.000 1983.230 404.000 ;
      LAYER met2 ;
        RECT 1983.510 402.195 1992.330 404.280 ;
      LAYER met2 ;
        RECT 1992.610 400.000 1992.890 404.000 ;
      LAYER met2 ;
        RECT 1993.170 402.195 2001.990 404.280 ;
      LAYER met2 ;
        RECT 2002.270 400.000 2002.550 404.000 ;
      LAYER met2 ;
        RECT 2002.830 402.195 2011.650 404.280 ;
      LAYER met2 ;
        RECT 2011.930 400.000 2012.210 404.000 ;
      LAYER met2 ;
        RECT 2012.490 402.195 2021.310 404.280 ;
      LAYER met2 ;
        RECT 2021.590 400.000 2021.870 404.000 ;
      LAYER met2 ;
        RECT 2022.150 402.195 2030.970 404.280 ;
      LAYER met2 ;
        RECT 2031.250 400.000 2031.530 404.000 ;
      LAYER met2 ;
        RECT 2031.810 402.195 2040.630 404.280 ;
      LAYER met2 ;
        RECT 2040.910 400.000 2041.190 404.000 ;
      LAYER met2 ;
        RECT 2041.470 402.195 2050.750 404.280 ;
      LAYER met2 ;
        RECT 2051.030 400.000 2051.310 404.000 ;
      LAYER met2 ;
        RECT 2051.590 402.195 2060.410 404.280 ;
      LAYER met2 ;
        RECT 2060.690 400.000 2060.970 404.000 ;
      LAYER met2 ;
        RECT 2061.250 402.195 2070.070 404.280 ;
      LAYER met2 ;
        RECT 2070.350 400.000 2070.630 404.000 ;
      LAYER met2 ;
        RECT 2070.910 402.195 2079.730 404.280 ;
      LAYER met2 ;
        RECT 2080.010 400.000 2080.290 404.000 ;
      LAYER met2 ;
        RECT 2080.570 402.195 2089.390 404.280 ;
      LAYER met2 ;
        RECT 2089.670 400.000 2089.950 404.000 ;
      LAYER met2 ;
        RECT 2090.230 402.195 2099.050 404.280 ;
      LAYER met2 ;
        RECT 2099.330 400.000 2099.610 404.000 ;
      LAYER met2 ;
        RECT 2099.890 402.195 2109.170 404.280 ;
      LAYER met2 ;
        RECT 2109.450 400.000 2109.730 404.000 ;
      LAYER met2 ;
        RECT 2110.010 402.195 2118.830 404.280 ;
      LAYER met2 ;
        RECT 2119.110 400.000 2119.390 404.000 ;
      LAYER met2 ;
        RECT 2119.670 402.195 2128.490 404.280 ;
      LAYER met2 ;
        RECT 2128.770 400.000 2129.050 404.000 ;
      LAYER met2 ;
        RECT 2129.330 402.195 2138.150 404.280 ;
      LAYER met2 ;
        RECT 2138.430 400.000 2138.710 404.000 ;
      LAYER met2 ;
        RECT 2138.990 402.195 2147.810 404.280 ;
      LAYER met2 ;
        RECT 2148.090 400.000 2148.370 404.000 ;
      LAYER met2 ;
        RECT 2148.650 402.195 2157.470 404.280 ;
      LAYER met2 ;
        RECT 2157.750 400.000 2158.030 404.000 ;
      LAYER met2 ;
        RECT 2158.310 402.195 2167.590 404.280 ;
      LAYER met2 ;
        RECT 2167.870 400.000 2168.150 404.000 ;
      LAYER met2 ;
        RECT 2168.430 402.195 2177.250 404.280 ;
      LAYER met2 ;
        RECT 2177.530 400.000 2177.810 404.000 ;
      LAYER met2 ;
        RECT 2178.090 402.195 2186.910 404.280 ;
      LAYER met2 ;
        RECT 2187.190 400.000 2187.470 404.000 ;
      LAYER met2 ;
        RECT 2187.750 402.195 2196.570 404.280 ;
      LAYER met2 ;
        RECT 2196.850 400.000 2197.130 404.000 ;
      LAYER met2 ;
        RECT 2197.410 402.195 2206.230 404.280 ;
      LAYER met2 ;
        RECT 2206.510 400.000 2206.790 404.000 ;
      LAYER met2 ;
        RECT 2207.070 402.195 2215.890 404.280 ;
      LAYER met2 ;
        RECT 2216.170 400.000 2216.450 404.000 ;
      LAYER met2 ;
        RECT 2216.730 402.195 2225.550 404.280 ;
      LAYER met2 ;
        RECT 2225.830 400.000 2226.110 404.000 ;
      LAYER met2 ;
        RECT 2226.390 402.195 2235.670 404.280 ;
      LAYER met2 ;
        RECT 2235.950 400.000 2236.230 404.000 ;
      LAYER met2 ;
        RECT 2236.510 402.195 2245.330 404.280 ;
      LAYER met2 ;
        RECT 2245.610 400.000 2245.890 404.000 ;
      LAYER met2 ;
        RECT 2246.170 402.195 2254.990 404.280 ;
      LAYER met2 ;
        RECT 2255.270 400.000 2255.550 404.000 ;
      LAYER met2 ;
        RECT 2255.830 402.195 2264.650 404.280 ;
      LAYER met2 ;
        RECT 2264.930 400.000 2265.210 404.000 ;
      LAYER met2 ;
        RECT 2265.490 402.195 2274.310 404.280 ;
      LAYER met2 ;
        RECT 2274.590 400.000 2274.870 404.000 ;
      LAYER met2 ;
        RECT 2275.150 402.195 2283.970 404.280 ;
      LAYER met2 ;
        RECT 2284.250 400.000 2284.530 404.000 ;
      LAYER met2 ;
        RECT 2284.810 402.195 2294.090 404.280 ;
      LAYER met2 ;
        RECT 2294.370 400.000 2294.650 404.000 ;
      LAYER met2 ;
        RECT 2294.930 402.195 2303.750 404.280 ;
      LAYER met2 ;
        RECT 2304.030 400.000 2304.310 404.000 ;
      LAYER met2 ;
        RECT 2304.590 402.195 2313.410 404.280 ;
      LAYER met2 ;
        RECT 2313.690 400.000 2313.970 404.000 ;
      LAYER met2 ;
        RECT 2314.250 402.195 2323.070 404.280 ;
      LAYER met2 ;
        RECT 2323.350 400.000 2323.630 404.000 ;
      LAYER met2 ;
        RECT 2323.910 402.195 2332.730 404.280 ;
      LAYER met2 ;
        RECT 2333.010 400.000 2333.290 404.000 ;
      LAYER met2 ;
        RECT 2333.570 402.195 2342.390 404.280 ;
      LAYER met2 ;
        RECT 2342.670 400.000 2342.950 404.000 ;
      LAYER met2 ;
        RECT 2343.230 402.195 2352.510 404.280 ;
      LAYER met2 ;
        RECT 2352.790 400.000 2353.070 404.000 ;
      LAYER met2 ;
        RECT 2353.350 402.195 2362.170 404.280 ;
      LAYER met2 ;
        RECT 2362.450 400.000 2362.730 404.000 ;
      LAYER met2 ;
        RECT 2363.010 402.195 2371.830 404.280 ;
      LAYER met2 ;
        RECT 2372.110 400.000 2372.390 404.000 ;
      LAYER met2 ;
        RECT 2372.670 402.195 2381.490 404.280 ;
      LAYER met2 ;
        RECT 2381.770 400.000 2382.050 404.000 ;
      LAYER met2 ;
        RECT 2382.330 402.195 2391.150 404.280 ;
      LAYER met2 ;
        RECT 2391.430 400.000 2391.710 404.000 ;
      LAYER met2 ;
        RECT 2391.990 402.195 2400.810 404.280 ;
      LAYER met2 ;
        RECT 2401.090 400.000 2401.370 404.000 ;
      LAYER met2 ;
        RECT 2401.650 402.195 2410.930 404.280 ;
      LAYER met2 ;
        RECT 2411.210 400.000 2411.490 404.000 ;
      LAYER met2 ;
        RECT 2411.770 402.195 2420.590 404.280 ;
      LAYER met2 ;
        RECT 2420.870 400.000 2421.150 404.000 ;
      LAYER met2 ;
        RECT 2421.430 402.195 2430.250 404.280 ;
      LAYER met2 ;
        RECT 2430.530 400.000 2430.810 404.000 ;
      LAYER met2 ;
        RECT 2431.090 402.195 2439.910 404.280 ;
      LAYER met2 ;
        RECT 2440.190 400.000 2440.470 404.000 ;
      LAYER met2 ;
        RECT 2440.750 402.195 2449.570 404.280 ;
      LAYER met2 ;
        RECT 2449.850 400.000 2450.130 404.000 ;
      LAYER met2 ;
        RECT 2450.410 402.195 2459.230 404.280 ;
      LAYER met2 ;
        RECT 2459.510 400.000 2459.790 404.000 ;
      LAYER met2 ;
        RECT 2460.070 402.195 2468.890 404.280 ;
      LAYER met2 ;
        RECT 2469.170 400.000 2469.450 404.000 ;
      LAYER met2 ;
        RECT 2469.730 402.195 2479.010 404.280 ;
      LAYER met2 ;
        RECT 2479.290 400.000 2479.570 404.000 ;
      LAYER met2 ;
        RECT 2479.850 402.195 2488.670 404.280 ;
      LAYER met2 ;
        RECT 2488.950 400.000 2489.230 404.000 ;
      LAYER met2 ;
        RECT 2489.510 402.195 2498.330 404.280 ;
      LAYER met2 ;
        RECT 2498.610 400.000 2498.890 404.000 ;
      LAYER met2 ;
        RECT 2499.170 402.195 2507.990 404.280 ;
      LAYER met2 ;
        RECT 2508.270 400.000 2508.550 404.000 ;
      LAYER met2 ;
        RECT 2508.830 402.195 2517.650 404.280 ;
      LAYER met2 ;
        RECT 2517.930 400.000 2518.210 404.000 ;
      LAYER met2 ;
        RECT 2518.490 402.195 2527.310 404.280 ;
      LAYER met2 ;
        RECT 2527.590 400.000 2527.870 404.000 ;
      LAYER met2 ;
        RECT 2528.150 402.195 2537.430 404.280 ;
      LAYER met2 ;
        RECT 2537.710 400.000 2537.990 404.000 ;
      LAYER met2 ;
        RECT 2538.270 402.195 2547.090 404.280 ;
      LAYER met2 ;
        RECT 2547.370 400.000 2547.650 404.000 ;
      LAYER met2 ;
        RECT 2547.930 402.195 2556.750 404.280 ;
      LAYER met2 ;
        RECT 2557.030 400.000 2557.310 404.000 ;
      LAYER met2 ;
        RECT 2557.590 402.195 2566.410 404.280 ;
      LAYER met2 ;
        RECT 2566.690 400.000 2566.970 404.000 ;
      LAYER met2 ;
        RECT 2567.250 402.195 2576.070 404.280 ;
      LAYER met2 ;
        RECT 2576.350 400.000 2576.630 404.000 ;
      LAYER met2 ;
        RECT 2576.910 402.195 2585.730 404.280 ;
      LAYER met2 ;
        RECT 2586.010 400.000 2586.290 404.000 ;
      LAYER met2 ;
        RECT 2586.570 402.195 2595.850 404.280 ;
      LAYER met2 ;
        RECT 2596.130 400.000 2596.410 404.000 ;
      LAYER met2 ;
        RECT 2596.690 402.195 2605.510 404.280 ;
      LAYER met2 ;
        RECT 2605.790 400.000 2606.070 404.000 ;
      LAYER met2 ;
        RECT 2606.350 402.195 2615.170 404.280 ;
      LAYER met2 ;
        RECT 2615.450 400.000 2615.730 404.000 ;
      LAYER met2 ;
        RECT 2616.010 402.195 2624.830 404.280 ;
      LAYER met2 ;
        RECT 2625.110 400.000 2625.390 404.000 ;
      LAYER met2 ;
        RECT 2625.670 402.195 2634.490 404.280 ;
      LAYER met2 ;
        RECT 2634.770 400.000 2635.050 404.000 ;
      LAYER met2 ;
        RECT 2635.330 402.195 2644.150 404.280 ;
      LAYER met2 ;
        RECT 2644.430 400.000 2644.710 404.000 ;
      LAYER met2 ;
        RECT 2644.990 402.195 2645.630 404.280 ;
      LAYER via2 ;
        RECT 675.370 3255.360 675.650 3255.640 ;
        RECT 289.430 3230.200 289.710 3230.480 ;
        RECT 288.970 3224.760 289.250 3225.040 ;
        RECT 288.510 3215.920 288.790 3216.200 ;
        RECT 288.050 3209.800 288.330 3210.080 ;
        RECT 287.590 3201.640 287.870 3201.920 ;
        RECT 287.130 3196.200 287.410 3196.480 ;
        RECT 286.670 3188.040 286.950 3188.320 ;
        RECT 286.210 2898.360 286.490 2898.640 ;
        RECT 688.250 3248.275 688.530 3248.555 ;
        RECT 1890.690 3264.200 1890.970 3264.480 ;
        RECT 1917.830 3264.200 1918.110 3264.480 ;
        RECT 2542.050 3264.200 2542.330 3264.480 ;
        RECT 2566.890 3264.200 2567.170 3264.480 ;
        RECT 1292.690 3258.080 1292.970 3258.360 ;
        RECT 1317.990 3258.080 1318.270 3258.360 ;
        RECT 941.710 3230.200 941.990 3230.480 ;
        RECT 696.990 2948.000 697.270 2948.280 ;
        RECT 337.730 2794.320 338.010 2794.600 ;
        RECT 344.630 2794.320 344.910 2794.600 ;
        RECT 351.530 2794.320 351.810 2794.600 ;
        RECT 358.430 2794.320 358.710 2794.600 ;
        RECT 362.570 2794.320 362.850 2794.600 ;
        RECT 365.330 2794.320 365.610 2794.600 ;
        RECT 368.550 2794.320 368.830 2794.600 ;
        RECT 371.310 2794.320 371.590 2794.600 ;
        RECT 374.990 2794.320 375.270 2794.600 ;
        RECT 379.130 2794.320 379.410 2794.600 ;
        RECT 384.190 2794.320 384.470 2794.600 ;
        RECT 386.950 2794.320 387.230 2794.600 ;
        RECT 392.930 2794.320 393.210 2794.600 ;
        RECT 396.610 2794.320 396.890 2794.600 ;
        RECT 399.370 2794.320 399.650 2794.600 ;
        RECT 403.970 2794.320 404.250 2794.600 ;
        RECT 406.270 2794.320 406.550 2794.600 ;
        RECT 409.950 2794.320 410.230 2794.600 ;
        RECT 414.550 2794.320 414.830 2794.600 ;
        RECT 419.150 2794.320 419.430 2794.600 ;
        RECT 420.990 2794.320 421.270 2794.600 ;
        RECT 427.430 2794.320 427.710 2794.600 ;
        RECT 431.570 2794.320 431.850 2794.600 ;
        RECT 310.130 2791.600 310.410 2791.880 ;
        RECT 317.030 2790.920 317.310 2791.200 ;
        RECT 351.070 2792.960 351.350 2793.240 ;
        RECT 379.590 2792.960 379.870 2793.240 ;
        RECT 392.470 2792.960 392.750 2793.240 ;
        RECT 397.070 2792.960 397.350 2793.240 ;
        RECT 426.970 2792.960 427.250 2793.240 ;
        RECT 413.630 2789.560 413.910 2789.840 ;
        RECT 387.870 2714.760 388.150 2715.040 ;
        RECT 433.870 2794.320 434.150 2794.600 ;
        RECT 439.390 2794.320 439.670 2794.600 ;
        RECT 441.230 2794.320 441.510 2794.600 ;
        RECT 444.450 2794.320 444.730 2794.600 ;
        RECT 445.830 2794.320 446.110 2794.600 ;
        RECT 449.050 2794.320 449.330 2794.600 ;
        RECT 455.030 2794.320 455.310 2794.600 ;
        RECT 461.010 2794.320 461.290 2794.600 ;
        RECT 462.390 2794.320 462.670 2794.600 ;
        RECT 466.530 2794.320 466.810 2794.600 ;
        RECT 468.830 2794.320 469.110 2794.600 ;
        RECT 475.270 2794.320 475.550 2794.600 ;
        RECT 478.490 2794.320 478.770 2794.600 ;
        RECT 482.630 2794.320 482.910 2794.600 ;
        RECT 485.850 2794.320 486.130 2794.600 ;
        RECT 489.070 2794.320 489.350 2794.600 ;
        RECT 491.830 2794.320 492.110 2794.600 ;
        RECT 496.430 2794.320 496.710 2794.600 ;
        RECT 500.110 2794.320 500.390 2794.600 ;
        RECT 510.230 2794.320 510.510 2794.600 ;
        RECT 524.030 2794.320 524.310 2794.600 ;
        RECT 536.450 2794.320 536.730 2794.600 ;
        RECT 542.430 2794.320 542.710 2794.600 ;
        RECT 434.330 2792.960 434.610 2793.240 ;
        RECT 455.490 2792.960 455.770 2793.240 ;
        RECT 468.370 2792.960 468.650 2793.240 ;
        RECT 473.890 2792.960 474.170 2793.240 ;
        RECT 481.250 2716.120 481.530 2716.400 ;
        RECT 497.350 2792.280 497.630 2792.560 ;
        RECT 501.950 2792.280 502.230 2792.560 ;
        RECT 500.110 2788.200 500.390 2788.480 ;
        RECT 504.250 2788.880 504.530 2789.160 ;
        RECT 507.010 2788.880 507.290 2789.160 ;
        RECT 531.390 2792.960 531.670 2793.240 ;
        RECT 542.430 2792.280 542.710 2792.560 ;
        RECT 551.630 2792.280 551.910 2792.560 ;
        RECT 541.510 2789.560 541.790 2789.840 ;
        RECT 534.610 2788.200 534.890 2788.480 ;
        RECT 510.230 2787.520 510.510 2787.800 ;
        RECT 513.910 2787.520 514.190 2787.800 ;
        RECT 517.130 2787.520 517.410 2787.800 ;
        RECT 520.810 2787.520 521.090 2787.800 ;
        RECT 527.710 2787.520 527.990 2787.800 ;
        RECT 530.930 2787.520 531.210 2787.800 ;
        RECT 517.130 2715.440 517.410 2715.720 ;
        RECT 700.210 2718.160 700.490 2718.440 ;
        RECT 707.110 2716.800 707.390 2717.080 ;
        RECT 741.610 2717.480 741.890 2717.760 ;
        RECT 942.170 3224.760 942.450 3225.040 ;
        RECT 942.630 3215.920 942.910 3216.200 ;
        RECT 943.090 3209.800 943.370 3210.080 ;
        RECT 943.550 3201.640 943.830 3201.920 ;
        RECT 944.010 3196.200 944.290 3196.480 ;
        RECT 944.470 3188.040 944.750 3188.320 ;
        RECT 944.930 2898.360 945.210 2898.640 ;
        RECT 941.710 2716.120 941.990 2716.400 ;
        RECT 1333.170 3249.240 1333.450 3249.520 ;
        RECT 1536.950 3230.200 1537.230 3230.480 ;
        RECT 1345.590 2946.640 1345.870 2946.920 ;
        RECT 1345.590 2935.760 1345.870 2936.040 ;
        RECT 1352.030 2901.760 1352.310 2902.040 ;
        RECT 1054.870 2799.760 1055.150 2800.040 ;
        RECT 979.890 2794.320 980.170 2794.600 ;
        RECT 1001.050 2794.320 1001.330 2794.600 ;
        RECT 1013.930 2794.320 1014.210 2794.600 ;
        RECT 1018.990 2794.320 1019.270 2794.600 ;
        RECT 1020.830 2794.320 1021.110 2794.600 ;
        RECT 1027.730 2794.320 1028.010 2794.600 ;
        RECT 1034.630 2794.320 1034.910 2794.600 ;
        RECT 1042.450 2794.320 1042.730 2794.600 ;
        RECT 1053.030 2794.320 1053.310 2794.600 ;
        RECT 944.930 2714.760 945.210 2715.040 ;
        RECT 1010.710 2792.960 1010.990 2793.240 ;
        RECT 1007.490 2788.200 1007.770 2788.480 ;
        RECT 1000.130 2718.160 1000.410 2718.440 ;
        RECT 1010.250 2715.440 1010.530 2715.720 ;
        RECT 1024.510 2792.960 1024.790 2793.240 ;
        RECT 1045.210 2792.960 1045.490 2793.240 ;
        RECT 1038.310 2788.200 1038.590 2788.480 ;
        RECT 1034.630 2787.520 1034.910 2787.800 ;
        RECT 1041.530 2787.520 1041.810 2787.800 ;
        RECT 1048.430 2787.520 1048.710 2787.800 ;
        RECT 1052.110 2717.480 1052.390 2717.760 ;
        RECT 1041.530 2716.800 1041.810 2717.080 ;
        RECT 1059.010 2794.320 1059.290 2794.600 ;
        RECT 1065.910 2794.320 1066.190 2794.600 ;
        RECT 1070.050 2794.320 1070.330 2794.600 ;
        RECT 1076.490 2794.320 1076.770 2794.600 ;
        RECT 1087.530 2794.320 1087.810 2794.600 ;
        RECT 1093.970 2794.320 1094.250 2794.600 ;
        RECT 1100.410 2794.320 1100.690 2794.600 ;
        RECT 1105.470 2794.320 1105.750 2794.600 ;
        RECT 1110.990 2794.320 1111.270 2794.600 ;
        RECT 1122.490 2794.320 1122.770 2794.600 ;
        RECT 1129.390 2794.320 1129.670 2794.600 ;
        RECT 1130.770 2794.320 1131.050 2794.600 ;
        RECT 1135.830 2794.320 1136.110 2794.600 ;
        RECT 1138.130 2794.320 1138.410 2794.600 ;
        RECT 1139.970 2794.320 1140.250 2794.600 ;
        RECT 1145.030 2794.320 1145.310 2794.600 ;
        RECT 1147.330 2794.320 1147.610 2794.600 ;
        RECT 1151.930 2794.320 1152.210 2794.600 ;
        RECT 1158.830 2794.320 1159.110 2794.600 ;
        RECT 1165.270 2794.320 1165.550 2794.600 ;
        RECT 1166.190 2794.320 1166.470 2794.600 ;
        RECT 1172.630 2794.320 1172.910 2794.600 ;
        RECT 1179.530 2794.320 1179.810 2794.600 ;
        RECT 1186.430 2794.320 1186.710 2794.600 ;
        RECT 1200.230 2794.320 1200.510 2794.600 ;
        RECT 1055.330 2788.200 1055.610 2788.480 ;
        RECT 1087.990 2793.640 1088.270 2793.920 ;
        RECT 1117.890 2793.640 1118.170 2793.920 ;
        RECT 1089.830 2788.200 1090.110 2788.480 ;
        RECT 1062.230 2787.520 1062.510 2787.800 ;
        RECT 1069.130 2787.520 1069.410 2787.800 ;
        RECT 1076.030 2787.520 1076.310 2787.800 ;
        RECT 1082.930 2787.520 1083.210 2787.800 ;
        RECT 1089.370 2787.520 1089.650 2787.800 ;
        RECT 1096.730 2787.520 1097.010 2787.800 ;
        RECT 1103.630 2787.520 1103.910 2787.800 ;
        RECT 1110.530 2787.520 1110.810 2787.800 ;
        RECT 1117.430 2787.520 1117.710 2787.800 ;
        RECT 1124.330 2787.520 1124.610 2787.800 ;
        RECT 1131.230 2793.640 1131.510 2793.920 ;
        RECT 1152.390 2791.600 1152.670 2791.880 ;
        RECT 1159.290 2793.640 1159.570 2793.920 ;
        RECT 1159.290 2792.280 1159.570 2792.560 ;
        RECT 1165.730 2793.640 1166.010 2793.920 ;
        RECT 1173.090 2793.640 1173.370 2793.920 ;
        RECT 1179.990 2793.640 1180.270 2793.920 ;
        RECT 1186.890 2793.640 1187.170 2793.920 ;
        RECT 1193.790 2791.600 1194.070 2791.880 ;
        RECT 1193.330 2790.240 1193.610 2790.520 ;
        RECT 1407.690 2894.960 1407.970 2895.240 ;
        RECT 1407.230 2204.760 1407.510 2205.040 ;
        RECT 1407.230 2149.680 1407.510 2149.960 ;
        RECT 1411.370 2697.080 1411.650 2697.360 ;
        RECT 1414.130 2692.320 1414.410 2692.600 ;
        RECT 1414.130 2686.880 1414.410 2687.160 ;
        RECT 1414.130 2682.120 1414.410 2682.400 ;
        RECT 1408.610 2676.680 1408.890 2676.960 ;
        RECT 1410.450 2671.920 1410.730 2672.200 ;
        RECT 1410.450 2667.160 1410.730 2667.440 ;
        RECT 1411.370 2661.720 1411.650 2662.000 ;
        RECT 1414.130 2656.960 1414.410 2657.240 ;
        RECT 1414.130 2651.520 1414.410 2651.800 ;
        RECT 1414.130 2646.760 1414.410 2647.040 ;
        RECT 1411.370 2641.320 1411.650 2641.600 ;
        RECT 1414.130 2636.560 1414.410 2636.840 ;
        RECT 1409.530 2631.800 1409.810 2632.080 ;
        RECT 1414.130 2626.360 1414.410 2626.640 ;
        RECT 1411.830 2621.600 1412.110 2621.880 ;
        RECT 1414.130 2616.160 1414.410 2616.440 ;
        RECT 1414.130 2611.400 1414.410 2611.680 ;
        RECT 1417.810 2605.960 1418.090 2606.240 ;
        RECT 1414.130 2601.200 1414.410 2601.480 ;
        RECT 1408.610 2596.440 1408.890 2596.720 ;
        RECT 1410.450 2591.000 1410.730 2591.280 ;
        RECT 1411.370 2586.240 1411.650 2586.520 ;
        RECT 1414.130 2580.800 1414.410 2581.080 ;
        RECT 1414.130 2576.040 1414.410 2576.320 ;
        RECT 1411.370 2571.280 1411.650 2571.560 ;
        RECT 1413.670 2565.840 1413.950 2566.120 ;
        RECT 1414.130 2561.080 1414.410 2561.360 ;
        RECT 1408.610 2555.640 1408.890 2555.920 ;
        RECT 1411.370 2550.880 1411.650 2551.160 ;
        RECT 1412.750 2545.440 1413.030 2545.720 ;
        RECT 1414.130 2540.680 1414.410 2540.960 ;
        RECT 1410.450 2535.920 1410.730 2536.200 ;
        RECT 1413.670 2530.480 1413.950 2530.760 ;
        RECT 1414.130 2525.720 1414.410 2526.000 ;
        RECT 1414.130 2520.280 1414.410 2520.560 ;
        RECT 1414.130 2515.520 1414.410 2515.800 ;
        RECT 1411.370 2510.080 1411.650 2510.360 ;
        RECT 1414.130 2505.320 1414.410 2505.600 ;
        RECT 1414.130 2495.120 1414.410 2495.400 ;
        RECT 1414.130 2484.920 1414.410 2485.200 ;
        RECT 1409.530 2480.160 1409.810 2480.440 ;
        RECT 1414.130 2475.400 1414.410 2475.680 ;
        RECT 1411.830 2469.960 1412.110 2470.240 ;
        RECT 1414.130 2465.200 1414.410 2465.480 ;
        RECT 1414.130 2459.760 1414.410 2460.040 ;
        RECT 1411.370 2455.000 1411.650 2455.280 ;
        RECT 1414.130 2449.560 1414.410 2449.840 ;
        RECT 1411.370 2444.800 1411.650 2445.080 ;
        RECT 1414.130 2440.040 1414.410 2440.320 ;
        RECT 1411.370 2434.600 1411.650 2434.880 ;
        RECT 1414.130 2429.840 1414.410 2430.120 ;
        RECT 1408.610 2424.400 1408.890 2424.680 ;
        RECT 1411.370 2419.640 1411.650 2419.920 ;
        RECT 1412.750 2414.200 1413.030 2414.480 ;
        RECT 1414.130 2409.440 1414.410 2409.720 ;
        RECT 1410.450 2404.680 1410.730 2404.960 ;
        RECT 1413.670 2399.240 1413.950 2399.520 ;
        RECT 1414.130 2394.480 1414.410 2394.760 ;
        RECT 1414.130 2389.040 1414.410 2389.320 ;
        RECT 1410.450 2384.280 1410.730 2384.560 ;
        RECT 1411.370 2378.840 1411.650 2379.120 ;
        RECT 1414.130 2374.080 1414.410 2374.360 ;
        RECT 1408.610 2369.320 1408.890 2369.600 ;
        RECT 1410.450 2363.880 1410.730 2364.160 ;
        RECT 1413.670 2359.120 1413.950 2359.400 ;
        RECT 1414.130 2353.680 1414.410 2353.960 ;
        RECT 1409.530 2348.920 1409.810 2349.200 ;
        RECT 1414.130 2344.160 1414.410 2344.440 ;
        RECT 1413.670 2338.720 1413.950 2339.000 ;
        RECT 1414.130 2333.960 1414.410 2334.240 ;
        RECT 1414.130 2328.520 1414.410 2328.800 ;
        RECT 1413.670 2323.760 1413.950 2324.040 ;
        RECT 1414.130 2318.320 1414.410 2318.600 ;
        RECT 1414.130 2313.560 1414.410 2313.840 ;
        RECT 1414.130 2308.800 1414.410 2309.080 ;
        RECT 1414.130 2303.360 1414.410 2303.640 ;
        RECT 1413.670 2298.600 1413.950 2298.880 ;
        RECT 1408.610 2293.160 1408.890 2293.440 ;
        RECT 1410.450 2288.400 1410.730 2288.680 ;
        RECT 1408.150 2282.960 1408.430 2283.240 ;
        RECT 1414.130 2278.200 1414.410 2278.480 ;
        RECT 1408.150 2273.440 1408.430 2273.720 ;
        RECT 1412.290 2268.000 1412.570 2268.280 ;
        RECT 1411.370 2263.240 1411.650 2263.520 ;
        RECT 1410.450 2232.640 1410.730 2232.920 ;
        RECT 1409.070 2227.880 1409.350 2228.160 ;
        RECT 1408.610 2212.920 1408.890 2213.200 ;
        RECT 1409.990 2222.440 1410.270 2222.720 ;
        RECT 1409.530 2217.680 1409.810 2217.960 ;
        RECT 1410.910 2202.720 1411.190 2203.000 ;
        RECT 1410.910 2197.280 1411.190 2197.560 ;
        RECT 1410.910 2187.080 1411.190 2187.360 ;
        RECT 1410.910 2182.320 1411.190 2182.600 ;
        RECT 1410.910 2177.560 1411.190 2177.840 ;
        RECT 1410.910 2172.120 1411.190 2172.400 ;
        RECT 1410.910 2161.920 1411.190 2162.200 ;
        RECT 1411.830 2257.800 1412.110 2258.080 ;
        RECT 1411.370 2157.160 1411.650 2157.440 ;
        RECT 1411.370 2146.960 1411.650 2147.240 ;
        RECT 1411.370 2142.200 1411.650 2142.480 ;
        RECT 1411.370 2136.760 1411.650 2137.040 ;
        RECT 1411.370 2134.720 1411.650 2135.000 ;
        RECT 1411.370 2126.560 1411.650 2126.840 ;
        RECT 1411.370 2121.800 1411.650 2122.080 ;
        RECT 1411.370 2117.040 1411.650 2117.320 ;
        RECT 1411.370 2111.600 1411.650 2111.880 ;
        RECT 1411.370 2106.840 1411.650 2107.120 ;
        RECT 1412.750 2253.040 1413.030 2253.320 ;
        RECT 1414.130 2248.280 1414.410 2248.560 ;
        RECT 1413.210 2242.840 1413.490 2243.120 ;
        RECT 1411.370 2071.480 1411.650 2071.760 ;
        RECT 1412.750 2091.200 1413.030 2091.480 ;
        RECT 1413.670 2238.080 1413.950 2238.360 ;
        RECT 1417.350 2192.520 1417.630 2192.800 ;
        RECT 1416.890 2167.360 1417.170 2167.640 ;
        RECT 1414.130 2101.400 1414.410 2101.680 ;
        RECT 1414.130 2096.640 1414.410 2096.920 ;
        RECT 1414.130 2086.440 1414.410 2086.720 ;
        RECT 1414.130 2081.680 1414.410 2081.960 ;
        RECT 1414.130 2076.240 1414.410 2076.520 ;
        RECT 1414.130 2066.040 1414.410 2066.320 ;
        RECT 1414.130 2061.280 1414.410 2061.560 ;
        RECT 1408.610 2046.320 1408.890 2046.600 ;
        RECT 1408.610 2040.880 1408.890 2041.160 ;
        RECT 1408.150 2015.720 1408.430 2016.000 ;
        RECT 1408.150 1990.560 1408.430 1990.840 ;
        RECT 1408.150 1985.800 1408.430 1986.080 ;
        RECT 1408.150 1980.360 1408.430 1980.640 ;
        RECT 1408.150 1975.600 1408.430 1975.880 ;
        RECT 1408.150 1970.160 1408.430 1970.440 ;
        RECT 1408.150 1965.400 1408.430 1965.680 ;
        RECT 1408.150 1959.960 1408.430 1960.240 ;
        RECT 1408.150 1955.200 1408.430 1955.480 ;
        RECT 1408.150 1950.440 1408.430 1950.720 ;
        RECT 1408.150 1945.000 1408.430 1945.280 ;
        RECT 1408.150 1940.240 1408.430 1940.520 ;
        RECT 1408.150 1934.800 1408.430 1935.080 ;
        RECT 1408.150 1930.040 1408.430 1930.320 ;
        RECT 1408.150 1925.280 1408.430 1925.560 ;
        RECT 1408.150 1919.840 1408.430 1920.120 ;
        RECT 1408.150 1915.080 1408.430 1915.360 ;
        RECT 1408.150 1909.640 1408.430 1909.920 ;
        RECT 1408.150 1899.440 1408.430 1899.720 ;
        RECT 1408.150 1894.680 1408.430 1894.960 ;
        RECT 1408.150 1889.920 1408.430 1890.200 ;
        RECT 1408.150 1879.720 1408.430 1880.000 ;
        RECT 1408.150 1874.280 1408.430 1874.560 ;
        RECT 1408.150 1869.520 1408.430 1869.800 ;
        RECT 1408.150 1859.320 1408.430 1859.600 ;
        RECT 1408.150 1854.560 1408.430 1854.840 ;
        RECT 1408.150 1844.360 1408.430 1844.640 ;
        RECT 1408.150 1838.920 1408.430 1839.200 ;
        RECT 1408.150 1823.960 1408.430 1824.240 ;
        RECT 1408.150 1819.200 1408.430 1819.480 ;
        RECT 1408.150 1813.760 1408.430 1814.040 ;
        RECT 1408.150 1803.560 1408.430 1803.840 ;
        RECT 1408.150 1798.800 1408.430 1799.080 ;
        RECT 1408.150 1788.600 1408.430 1788.880 ;
        RECT 1408.150 1758.680 1408.430 1758.960 ;
        RECT 1408.150 1753.240 1408.430 1753.520 ;
        RECT 1408.150 1748.480 1408.430 1748.760 ;
        RECT 1408.150 1743.040 1408.430 1743.320 ;
        RECT 1408.150 1738.280 1408.430 1738.560 ;
        RECT 1408.150 1732.840 1408.430 1733.120 ;
        RECT 1408.150 1728.080 1408.430 1728.360 ;
        RECT 1408.150 1723.320 1408.430 1723.600 ;
        RECT 1408.150 1717.880 1408.430 1718.160 ;
        RECT 1408.150 1707.680 1408.430 1707.960 ;
        RECT 1414.130 2055.840 1414.410 2056.120 ;
        RECT 1413.670 2051.080 1413.950 2051.360 ;
        RECT 1414.130 2036.120 1414.410 2036.400 ;
        RECT 1411.830 2030.680 1412.110 2030.960 ;
        RECT 1411.370 1995.320 1411.650 1995.600 ;
        RECT 1409.070 1904.880 1409.350 1905.160 ;
        RECT 1409.070 1884.480 1409.350 1884.760 ;
        RECT 1409.070 1864.080 1409.350 1864.360 ;
        RECT 1409.070 1849.120 1409.350 1849.400 ;
        RECT 1409.070 1809.000 1409.350 1809.280 ;
        RECT 1409.070 1794.040 1409.350 1794.320 ;
        RECT 1411.370 1773.640 1411.650 1773.920 ;
        RECT 1414.130 2025.920 1414.410 2026.200 ;
        RECT 1414.130 2021.160 1414.410 2021.440 ;
        RECT 1417.810 2068.080 1418.090 2068.360 ;
        RECT 1416.890 2066.720 1417.170 2067.000 ;
        RECT 1418.730 2067.400 1419.010 2067.680 ;
        RECT 1419.650 2066.040 1419.930 2066.320 ;
        RECT 1414.130 2010.960 1414.410 2011.240 ;
        RECT 1414.130 2005.520 1414.410 2005.800 ;
        RECT 1414.130 2000.760 1414.410 2001.040 ;
        RECT 1422.410 1834.160 1422.690 1834.440 ;
        RECT 1413.210 1783.840 1413.490 1784.120 ;
        RECT 1412.750 1778.400 1413.030 1778.680 ;
        RECT 1412.290 1768.200 1412.570 1768.480 ;
        RECT 1411.830 1763.440 1412.110 1763.720 ;
        RECT 1409.070 1713.120 1409.350 1713.400 ;
        RECT 1408.150 1702.920 1408.430 1703.200 ;
        RECT 1408.610 1698.160 1408.890 1698.440 ;
        RECT 1408.150 1692.720 1408.430 1693.000 ;
        RECT 1408.150 1687.960 1408.430 1688.240 ;
        RECT 1408.150 1682.520 1408.430 1682.800 ;
        RECT 1408.610 1677.760 1408.890 1678.040 ;
        RECT 1408.150 1672.320 1408.430 1672.600 ;
        RECT 1408.150 1667.560 1408.430 1667.840 ;
        RECT 1408.610 1662.800 1408.890 1663.080 ;
        RECT 1409.530 1657.360 1409.810 1657.640 ;
        RECT 1408.150 1652.600 1408.430 1652.880 ;
        RECT 1407.690 1647.160 1407.970 1647.440 ;
        RECT 1408.150 1642.400 1408.430 1642.680 ;
        RECT 1407.690 1636.960 1407.970 1637.240 ;
        RECT 1407.690 1627.440 1407.970 1627.720 ;
        RECT 1411.830 1632.200 1412.110 1632.480 ;
        RECT 1425.630 1828.720 1425.910 1829.000 ;
        RECT 1435.290 2066.720 1435.570 2067.000 ;
        RECT 1435.750 2066.040 1436.030 2066.320 ;
        RECT 1435.290 2065.360 1435.570 2065.640 ;
        RECT 1435.290 2064.680 1435.570 2064.960 ;
        RECT 1435.750 2064.000 1436.030 2064.280 ;
        RECT 1535.570 3224.760 1535.850 3225.040 ;
        RECT 1535.570 3217.280 1535.850 3217.560 ;
        RECT 1538.330 3210.480 1538.610 3210.760 ;
        RECT 1538.330 3202.320 1538.610 3202.600 ;
        RECT 1535.110 3196.200 1535.390 3196.480 ;
        RECT 1534.190 3189.400 1534.470 3189.680 ;
        RECT 1483.130 2066.720 1483.410 2067.000 ;
        RECT 1482.670 2066.040 1482.950 2066.320 ;
        RECT 1483.130 2065.360 1483.410 2065.640 ;
        RECT 1483.130 2064.680 1483.410 2064.960 ;
        RECT 1482.670 2064.000 1482.950 2064.280 ;
        RECT 1531.890 2066.720 1532.170 2067.000 ;
        RECT 1532.350 2066.040 1532.630 2066.320 ;
        RECT 1531.890 2065.360 1532.170 2065.640 ;
        RECT 1531.890 2064.680 1532.170 2064.960 ;
        RECT 1532.350 2064.000 1532.630 2064.280 ;
        RECT 1538.330 2899.040 1538.610 2899.320 ;
        RECT 1935.770 3249.240 1936.050 3249.520 ;
        RECT 1945.890 3249.240 1946.170 3249.520 ;
        RECT 1742.110 2796.360 1742.390 2796.640 ;
        RECT 1790.870 2796.360 1791.150 2796.640 ;
        RECT 1587.090 2794.320 1587.370 2794.600 ;
        RECT 1593.990 2794.320 1594.270 2794.600 ;
        RECT 1600.890 2794.320 1601.170 2794.600 ;
        RECT 1628.490 2794.320 1628.770 2794.600 ;
        RECT 1635.390 2794.320 1635.670 2794.600 ;
        RECT 1646.430 2794.320 1646.710 2794.600 ;
        RECT 1649.650 2794.320 1649.930 2794.600 ;
        RECT 1658.850 2794.320 1659.130 2794.600 ;
        RECT 1662.990 2794.320 1663.270 2794.600 ;
        RECT 1669.890 2794.320 1670.170 2794.600 ;
        RECT 1676.790 2794.320 1677.070 2794.600 ;
        RECT 1683.690 2794.320 1683.970 2794.600 ;
        RECT 1687.830 2794.320 1688.110 2794.600 ;
        RECT 1690.590 2794.320 1690.870 2794.600 ;
        RECT 1697.490 2794.320 1697.770 2794.600 ;
        RECT 1704.390 2794.320 1704.670 2794.600 ;
        RECT 1711.290 2794.320 1711.570 2794.600 ;
        RECT 1718.650 2794.320 1718.930 2794.600 ;
        RECT 1721.410 2794.320 1721.690 2794.600 ;
        RECT 1725.090 2794.320 1725.370 2794.600 ;
        RECT 1731.990 2794.320 1732.270 2794.600 ;
        RECT 1581.570 2788.880 1581.850 2789.160 ;
        RECT 1579.730 2066.720 1580.010 2067.000 ;
        RECT 1579.270 2066.040 1579.550 2066.320 ;
        RECT 1579.730 2065.360 1580.010 2065.640 ;
        RECT 1579.730 2064.680 1580.010 2064.960 ;
        RECT 1579.270 2064.000 1579.550 2064.280 ;
        RECT 1601.350 2793.640 1601.630 2793.920 ;
        RECT 1611.010 2793.640 1611.290 2793.920 ;
        RECT 1607.790 2790.240 1608.070 2790.520 ;
        RECT 1617.910 2792.960 1618.190 2793.240 ;
        RECT 1624.810 2792.960 1625.090 2793.240 ;
        RECT 1614.690 2790.240 1614.970 2790.520 ;
        RECT 1621.590 2788.200 1621.870 2788.480 ;
        RECT 1631.710 2793.640 1631.990 2793.920 ;
        RECT 1642.290 2793.640 1642.570 2793.920 ;
        RECT 1638.610 2792.960 1638.890 2793.240 ;
        RECT 1645.510 2792.960 1645.790 2793.240 ;
        RECT 1649.190 2789.560 1649.470 2789.840 ;
        RECT 1652.410 2793.640 1652.690 2793.920 ;
        RECT 1656.090 2788.880 1656.370 2789.160 ;
        RECT 1655.630 2064.680 1655.910 2064.960 ;
        RECT 1665.750 2793.640 1666.030 2793.920 ;
        RECT 1670.350 2793.640 1670.630 2793.920 ;
        RECT 1676.330 2066.720 1676.610 2067.000 ;
        RECT 1675.870 2066.040 1676.150 2066.320 ;
        RECT 1676.330 2065.360 1676.610 2065.640 ;
        RECT 1676.330 2064.680 1676.610 2064.960 ;
        RECT 1675.870 2064.000 1676.150 2064.280 ;
        RECT 1677.250 2793.640 1677.530 2793.920 ;
        RECT 1683.230 2793.640 1683.510 2793.920 ;
        RECT 1684.150 2793.640 1684.430 2793.920 ;
        RECT 1695.190 2793.640 1695.470 2793.920 ;
        RECT 1408.610 1611.800 1408.890 1612.080 ;
        RECT 1699.330 2793.640 1699.610 2793.920 ;
        RECT 1706.230 2793.640 1706.510 2793.920 ;
        RECT 1712.670 2793.640 1712.950 2793.920 ;
        RECT 1718.190 2793.640 1718.470 2793.920 ;
        RECT 1718.190 2788.200 1718.470 2788.480 ;
        RECT 1730.150 2793.640 1730.430 2793.920 ;
        RECT 1738.890 2794.320 1739.170 2794.600 ;
        RECT 1738.430 2793.640 1738.710 2793.920 ;
        RECT 1741.190 2793.640 1741.470 2793.920 ;
        RECT 1745.790 2794.320 1746.070 2794.600 ;
        RECT 1760.050 2794.320 1760.330 2794.600 ;
        RECT 1780.290 2794.320 1780.570 2794.600 ;
        RECT 1748.550 2793.640 1748.830 2793.920 ;
        RECT 1752.690 2792.280 1752.970 2792.560 ;
        RECT 1766.490 2793.640 1766.770 2793.920 ;
        RECT 1773.390 2793.640 1773.670 2793.920 ;
        RECT 1787.190 2792.280 1787.470 2792.560 ;
        RECT 1760.510 2788.200 1760.790 2788.480 ;
        RECT 1753.150 2787.520 1753.430 2787.800 ;
        RECT 1752.230 2064.680 1752.510 2064.960 ;
        RECT 1760.050 2777.320 1760.330 2777.600 ;
        RECT 1766.490 2787.520 1766.770 2787.800 ;
        RECT 1773.390 2787.520 1773.670 2787.800 ;
        RECT 1770.630 2068.760 1770.910 2069.040 ;
        RECT 1772.930 2066.720 1773.210 2067.000 ;
        RECT 1772.470 2066.040 1772.750 2066.320 ;
        RECT 1772.930 2065.360 1773.210 2065.640 ;
        RECT 1772.930 2064.680 1773.210 2064.960 ;
        RECT 1772.470 2064.000 1772.750 2064.280 ;
        RECT 1780.750 2787.520 1781.030 2787.800 ;
        RECT 1787.650 2787.520 1787.930 2787.800 ;
        RECT 1794.550 2777.320 1794.830 2777.600 ;
        RECT 1835.490 2069.440 1835.770 2069.720 ;
        RECT 1821.690 2066.720 1821.970 2067.000 ;
        RECT 1821.690 2065.360 1821.970 2065.640 ;
        RECT 1821.690 2064.000 1821.970 2064.280 ;
        RECT 1835.490 2063.320 1835.770 2063.600 ;
        RECT 1842.850 2069.440 1843.130 2069.720 ;
        RECT 1859.410 2070.120 1859.690 2070.400 ;
        RECT 1849.750 2069.440 1850.030 2069.720 ;
        RECT 1856.190 2069.440 1856.470 2069.720 ;
        RECT 1863.090 2069.440 1863.370 2069.720 ;
        RECT 1841.470 2065.360 1841.750 2065.640 ;
        RECT 1842.390 2065.360 1842.670 2065.640 ;
        RECT 1849.290 2065.360 1849.570 2065.640 ;
        RECT 1854.810 2065.360 1855.090 2065.640 ;
        RECT 1856.650 2064.000 1856.930 2064.280 ;
        RECT 1869.530 2066.720 1869.810 2067.000 ;
        RECT 1869.990 2066.040 1870.270 2066.320 ;
        RECT 1869.530 2064.680 1869.810 2064.960 ;
        RECT 1869.990 2064.000 1870.270 2064.280 ;
        RECT 1841.470 2063.320 1841.750 2063.600 ;
        RECT 1854.810 2063.320 1855.090 2063.600 ;
        RECT 1856.190 2063.320 1856.470 2063.600 ;
        RECT 1876.890 2066.040 1877.170 2066.320 ;
        RECT 1877.810 2066.040 1878.090 2066.320 ;
        RECT 1883.790 2066.040 1884.070 2066.320 ;
        RECT 1877.350 2065.360 1877.630 2065.640 ;
        RECT 1883.790 2064.000 1884.070 2064.280 ;
        RECT 1891.150 2066.040 1891.430 2066.320 ;
        RECT 1898.050 2069.440 1898.330 2069.720 ;
        RECT 1898.970 2066.720 1899.250 2067.000 ;
        RECT 1903.110 2068.760 1903.390 2069.040 ;
        RECT 1904.950 2066.720 1905.230 2067.000 ;
        RECT 1911.390 2066.720 1911.670 2067.000 ;
        RECT 1903.110 2066.040 1903.390 2066.320 ;
        RECT 1910.930 2065.360 1911.210 2065.640 ;
        RECT 1911.850 2065.360 1912.130 2065.640 ;
        RECT 1890.690 2064.000 1890.970 2064.280 ;
        RECT 1898.050 2064.000 1898.330 2064.280 ;
        RECT 1898.970 2064.000 1899.250 2064.280 ;
        RECT 1863.090 2063.320 1863.370 2063.600 ;
        RECT 1870.910 2063.320 1871.190 2063.600 ;
        RECT 1921.510 2068.760 1921.790 2069.040 ;
        RECT 1926.570 2067.400 1926.850 2067.680 ;
        RECT 1925.190 2065.360 1925.470 2065.640 ;
        RECT 1926.570 2065.360 1926.850 2065.640 ;
        RECT 1932.090 2067.400 1932.370 2067.680 ;
        RECT 1939.450 2069.440 1939.730 2069.720 ;
        RECT 1953.250 2069.440 1953.530 2069.720 ;
        RECT 1960.150 2069.440 1960.430 2069.720 ;
        RECT 2014.890 2069.440 2015.170 2069.720 ;
        RECT 1959.690 2068.760 1959.970 2069.040 ;
        RECT 1980.390 2068.760 1980.670 2069.040 ;
        RECT 2190.610 3230.200 2190.890 3230.480 ;
        RECT 2038.810 2069.440 2039.090 2069.720 ;
        RECT 2052.610 2069.440 2052.890 2069.720 ;
        RECT 1945.890 2067.400 1946.170 2067.680 ;
        RECT 1946.810 2067.400 1947.090 2067.680 ;
        RECT 1973.490 2067.400 1973.770 2067.680 ;
        RECT 1945.430 2064.680 1945.710 2064.960 ;
        RECT 1946.350 2064.680 1946.630 2064.960 ;
        RECT 2021.790 2067.400 2022.070 2067.680 ;
        RECT 1966.130 2066.720 1966.410 2067.000 ;
        RECT 1987.290 2066.720 1987.570 2067.000 ;
        RECT 1952.790 2064.680 1953.070 2064.960 ;
        RECT 2007.990 2066.720 2008.270 2067.000 ;
        RECT 1987.750 2065.360 1988.030 2065.640 ;
        RECT 1994.190 2065.360 1994.470 2065.640 ;
        RECT 1966.590 2064.680 1966.870 2064.960 ;
        RECT 1980.390 2064.680 1980.670 2064.960 ;
        RECT 1987.290 2064.680 1987.570 2064.960 ;
        RECT 1966.130 2064.000 1966.410 2064.280 ;
        RECT 1973.490 2064.000 1973.770 2064.280 ;
        RECT 2001.090 2064.000 2001.370 2064.280 ;
        RECT 2015.810 2064.000 2016.090 2064.280 ;
        RECT 1904.490 2063.320 1904.770 2063.600 ;
        RECT 1911.390 2063.320 1911.670 2063.600 ;
        RECT 1918.290 2063.320 1918.570 2063.600 ;
        RECT 1925.190 2063.320 1925.470 2063.600 ;
        RECT 1935.310 2063.320 1935.590 2063.600 ;
        RECT 1938.990 2063.320 1939.270 2063.600 ;
        RECT 1994.190 2063.320 1994.470 2063.600 ;
        RECT 2001.090 2063.320 2001.370 2063.600 ;
        RECT 2028.690 2057.200 2028.970 2057.480 ;
        RECT 1414.130 1607.040 1414.410 1607.320 ;
        RECT 2083.890 1964.720 2084.170 1965.000 ;
        RECT 2082.050 1956.560 2082.330 1956.840 ;
        RECT 2099.530 1732.840 2099.810 1733.120 ;
        RECT 2099.070 1721.960 2099.350 1722.240 ;
        RECT 2098.610 1718.560 2098.890 1718.840 ;
        RECT 2098.150 1708.360 2098.430 1708.640 ;
        RECT 2097.690 1704.960 2097.970 1705.240 ;
        RECT 2191.070 3224.760 2191.350 3225.040 ;
        RECT 2191.530 3215.920 2191.810 3216.200 ;
        RECT 2191.990 3209.800 2192.270 3210.080 ;
        RECT 2192.450 3201.640 2192.730 3201.920 ;
        RECT 2192.910 3196.200 2193.190 3196.480 ;
        RECT 2193.370 3188.040 2193.650 3188.320 ;
        RECT 2193.830 2898.360 2194.110 2898.640 ;
        RECT 2582.070 3249.240 2582.350 3249.520 ;
        RECT 2594.490 2946.640 2594.770 2946.920 ;
        RECT 2594.490 2938.480 2594.770 2938.760 ;
        RECT 2228.790 2794.320 2229.070 2794.600 ;
        RECT 2256.390 2794.320 2256.670 2794.600 ;
        RECT 2263.290 2794.320 2263.570 2794.600 ;
        RECT 2268.350 2794.320 2268.630 2794.600 ;
        RECT 2270.190 2794.320 2270.470 2794.600 ;
        RECT 2277.090 2794.320 2277.370 2794.600 ;
        RECT 2283.990 2794.320 2284.270 2794.600 ;
        RECT 2290.890 2794.320 2291.170 2794.600 ;
        RECT 2297.790 2794.320 2298.070 2794.600 ;
        RECT 2305.150 2794.320 2305.430 2794.600 ;
        RECT 2308.370 2794.320 2308.650 2794.600 ;
        RECT 2311.590 2794.320 2311.870 2794.600 ;
        RECT 2318.490 2794.320 2318.770 2794.600 ;
        RECT 2325.390 2794.320 2325.670 2794.600 ;
        RECT 2332.290 2794.320 2332.570 2794.600 ;
        RECT 2339.190 2794.320 2339.470 2794.600 ;
        RECT 2249.490 2788.880 2249.770 2789.160 ;
        RECT 2263.750 2793.640 2264.030 2793.920 ;
        RECT 2266.510 2792.960 2266.790 2793.240 ;
        RECT 2273.870 2793.640 2274.150 2793.920 ;
        RECT 2280.310 2793.640 2280.590 2793.920 ;
        RECT 2287.210 2793.640 2287.490 2793.920 ;
        RECT 2294.110 2793.640 2294.390 2793.920 ;
        RECT 2304.690 2793.640 2304.970 2793.920 ;
        RECT 2301.930 2792.960 2302.210 2793.240 ;
        RECT 2304.230 2788.200 2304.510 2788.480 ;
        RECT 2315.270 2793.640 2315.550 2793.920 ;
        RECT 2321.250 2793.640 2321.530 2793.920 ;
        RECT 2326.310 2793.640 2326.590 2793.920 ;
        RECT 2332.750 2793.640 2333.030 2793.920 ;
        RECT 2343.790 2794.320 2344.070 2794.600 ;
        RECT 2346.090 2794.320 2346.370 2794.600 ;
        RECT 2352.990 2794.320 2353.270 2794.600 ;
        RECT 2359.890 2794.320 2360.170 2794.600 ;
        RECT 2366.790 2794.320 2367.070 2794.600 ;
        RECT 2373.690 2794.320 2373.970 2794.600 ;
        RECT 2377.370 2794.320 2377.650 2794.600 ;
        RECT 2380.590 2794.320 2380.870 2794.600 ;
        RECT 2382.890 2794.320 2383.170 2794.600 ;
        RECT 2387.950 2794.320 2388.230 2794.600 ;
        RECT 2394.850 2794.320 2395.130 2794.600 ;
        RECT 2401.750 2794.320 2402.030 2794.600 ;
        RECT 2339.650 2793.640 2339.930 2793.920 ;
        RECT 2340.110 2792.960 2340.390 2793.240 ;
        RECT 2350.230 2792.960 2350.510 2793.240 ;
        RECT 2356.670 2793.640 2356.950 2793.920 ;
        RECT 2360.810 2793.640 2361.090 2793.920 ;
        RECT 2367.250 2793.640 2367.530 2793.920 ;
        RECT 2353.450 2069.440 2353.730 2069.720 ;
        RECT 2340.570 2063.320 2340.850 2063.600 ;
        RECT 2347.010 2063.320 2347.290 2063.600 ;
        RECT 2359.890 2063.320 2360.170 2063.600 ;
        RECT 2374.150 2793.640 2374.430 2793.920 ;
        RECT 2381.050 2792.960 2381.330 2793.240 ;
        RECT 2387.490 2791.600 2387.770 2791.880 ;
        RECT 2394.390 2792.280 2394.670 2792.560 ;
        RECT 2421.990 2793.640 2422.270 2793.920 ;
        RECT 2408.190 2792.960 2408.470 2793.240 ;
        RECT 2408.190 2792.280 2408.470 2792.560 ;
        RECT 2415.090 2792.280 2415.370 2792.560 ;
        RECT 2428.890 2792.280 2429.170 2792.560 ;
        RECT 2435.790 2792.280 2436.070 2792.560 ;
        RECT 2401.750 2791.600 2402.030 2791.880 ;
        RECT 2442.690 2791.600 2442.970 2791.880 ;
        RECT 2415.090 2790.920 2415.370 2791.200 ;
        RECT 2421.990 2790.240 2422.270 2790.520 ;
        RECT 2415.090 2789.560 2415.370 2789.840 ;
        RECT 2428.890 2789.560 2429.170 2789.840 ;
        RECT 2415.090 2788.880 2415.370 2789.160 ;
        RECT 2435.790 2788.880 2436.070 2789.160 ;
        RECT 2442.690 2788.200 2442.970 2788.480 ;
        RECT 2374.150 2069.440 2374.430 2069.720 ;
        RECT 2387.950 2069.440 2388.230 2069.720 ;
        RECT 2380.590 2068.760 2380.870 2069.040 ;
        RECT 2387.490 2068.760 2387.770 2069.040 ;
        RECT 2394.390 2068.080 2394.670 2068.360 ;
        RECT 2402.210 2067.400 2402.490 2067.680 ;
        RECT 2428.890 2067.400 2429.170 2067.680 ;
        RECT 2408.190 2066.720 2408.470 2067.000 ;
        RECT 2415.090 2066.720 2415.370 2067.000 ;
        RECT 2421.990 2066.040 2422.270 2066.320 ;
        RECT 2442.690 2066.040 2442.970 2066.320 ;
        RECT 2435.790 2065.360 2436.070 2065.640 ;
        RECT 2449.590 2064.680 2449.870 2064.960 ;
        RECT 2456.490 2064.680 2456.770 2064.960 ;
        RECT 2525.490 2068.760 2525.770 2069.040 ;
        RECT 2532.390 2068.080 2532.670 2068.360 ;
        RECT 2456.950 2063.320 2457.230 2063.600 ;
        RECT 2463.390 2063.320 2463.670 2063.600 ;
        RECT 2470.290 2063.320 2470.570 2063.600 ;
        RECT 2478.570 2063.320 2478.850 2063.600 ;
        RECT 2484.090 2063.320 2484.370 2063.600 ;
        RECT 2491.450 2063.320 2491.730 2063.600 ;
        RECT 2497.890 2063.320 2498.170 2063.600 ;
        RECT 2505.250 2063.320 2505.530 2063.600 ;
        RECT 2512.610 2063.320 2512.890 2063.600 ;
        RECT 2518.590 2063.320 2518.870 2063.600 ;
        RECT 2519.970 2063.320 2520.250 2063.600 ;
        RECT 2587.590 2063.320 2587.870 2063.600 ;
        RECT 2367.250 2051.760 2367.530 2052.040 ;
        RECT 2100.450 1745.760 2100.730 1746.040 ;
        RECT 2099.990 1732.160 2100.270 1732.440 ;
        RECT 2100.450 1668.240 2100.730 1668.520 ;
        RECT 2099.990 1660.080 2100.270 1660.360 ;
        RECT 2099.530 1654.640 2099.810 1654.920 ;
        RECT 2099.070 1645.800 2099.350 1646.080 ;
        RECT 2098.610 1640.360 2098.890 1640.640 ;
        RECT 2098.150 1628.800 2098.430 1629.080 ;
        RECT 2097.690 1625.400 2097.970 1625.680 ;
        RECT 2632.210 2049.720 2632.490 2050.000 ;
        RECT 1396.650 1604.320 1396.930 1604.600 ;
      LAYER met3 ;
        RECT 1890.665 3264.500 1890.995 3264.505 ;
        RECT 1917.805 3264.500 1918.135 3264.505 ;
        RECT 1890.665 3264.490 1891.250 3264.500 ;
        RECT 1917.550 3264.490 1918.135 3264.500 ;
        RECT 1890.665 3264.190 1891.450 3264.490 ;
        RECT 1917.350 3264.190 1918.135 3264.490 ;
        RECT 1890.665 3264.180 1891.250 3264.190 ;
        RECT 1917.550 3264.180 1918.135 3264.190 ;
        RECT 1890.665 3264.175 1890.995 3264.180 ;
        RECT 1917.805 3264.175 1918.135 3264.180 ;
        RECT 2542.025 3264.500 2542.355 3264.505 ;
        RECT 2566.865 3264.500 2567.195 3264.505 ;
        RECT 2542.025 3264.490 2542.610 3264.500 ;
        RECT 2566.865 3264.490 2567.450 3264.500 ;
        RECT 2542.025 3264.190 2542.810 3264.490 ;
        RECT 2566.865 3264.190 2567.650 3264.490 ;
        RECT 2542.025 3264.180 2542.610 3264.190 ;
        RECT 2566.865 3264.180 2567.450 3264.190 ;
        RECT 2542.025 3264.175 2542.355 3264.180 ;
        RECT 2566.865 3264.175 2567.195 3264.180 ;
        RECT 1292.665 3258.380 1292.995 3258.385 ;
        RECT 1317.965 3258.380 1318.295 3258.385 ;
        RECT 1292.665 3258.370 1293.230 3258.380 ;
        RECT 1317.825 3258.370 1318.295 3258.380 ;
        RECT 1292.665 3258.070 1293.450 3258.370 ;
        RECT 1317.510 3258.070 1318.295 3258.370 ;
        RECT 1292.665 3258.060 1293.230 3258.070 ;
        RECT 1317.825 3258.060 1318.295 3258.070 ;
        RECT 1292.665 3258.055 1292.995 3258.060 ;
        RECT 1317.965 3258.055 1318.295 3258.060 ;
        RECT 646.110 3255.650 646.490 3255.660 ;
        RECT 669.110 3255.650 669.490 3255.660 ;
        RECT 675.345 3255.650 675.675 3255.665 ;
        RECT 646.110 3255.350 675.675 3255.650 ;
        RECT 646.110 3255.340 646.490 3255.350 ;
        RECT 669.110 3255.340 669.490 3255.350 ;
        RECT 675.345 3255.335 675.675 3255.350 ;
        RECT 659.280 3251.235 661.020 3252.140 ;
        RECT 1309.280 3251.235 1311.020 3252.140 ;
        RECT 1909.280 3251.235 1911.020 3252.140 ;
        RECT 2559.280 3251.235 2561.020 3252.140 ;
        RECT 300.000 3232.785 304.600 3233.085 ;
        RECT 289.405 3230.490 289.735 3230.505 ;
        RECT 300.230 3230.490 300.530 3232.785 ;
        RECT 289.405 3230.190 300.530 3230.490 ;
        RECT 289.405 3230.175 289.735 3230.190 ;
        RECT 300.000 3227.145 304.600 3227.445 ;
        RECT 288.945 3225.050 289.275 3225.065 ;
        RECT 300.230 3225.050 300.530 3227.145 ;
        RECT 288.945 3224.750 300.530 3225.050 ;
        RECT 288.945 3224.735 289.275 3224.750 ;
        RECT 300.000 3218.645 304.600 3218.945 ;
        RECT 288.485 3216.210 288.815 3216.225 ;
        RECT 300.230 3216.210 300.530 3218.645 ;
        RECT 288.485 3215.910 300.530 3216.210 ;
        RECT 288.485 3215.895 288.815 3215.910 ;
        RECT 300.000 3213.005 304.600 3213.305 ;
        RECT 288.025 3210.090 288.355 3210.105 ;
        RECT 300.230 3210.090 300.530 3213.005 ;
        RECT 288.025 3209.790 300.530 3210.090 ;
        RECT 288.025 3209.775 288.355 3209.790 ;
        RECT 300.000 3204.505 304.600 3204.805 ;
        RECT 287.565 3201.930 287.895 3201.945 ;
        RECT 300.230 3201.930 300.530 3204.505 ;
        RECT 287.565 3201.630 300.530 3201.930 ;
        RECT 287.565 3201.615 287.895 3201.630 ;
        RECT 300.000 3198.865 304.600 3199.165 ;
        RECT 287.105 3196.490 287.435 3196.505 ;
        RECT 300.230 3196.490 300.530 3198.865 ;
        RECT 287.105 3196.190 300.530 3196.490 ;
        RECT 287.105 3196.175 287.435 3196.190 ;
        RECT 300.000 3190.365 304.600 3190.665 ;
        RECT 286.645 3188.330 286.975 3188.345 ;
        RECT 300.230 3188.330 300.530 3190.365 ;
        RECT 286.645 3188.030 300.530 3188.330 ;
        RECT 286.645 3188.015 286.975 3188.030 ;
        RECT 300.000 2901.125 304.600 2901.425 ;
        RECT 286.185 2898.650 286.515 2898.665 ;
        RECT 300.230 2898.650 300.530 2901.125 ;
        RECT 286.185 2898.350 300.530 2898.650 ;
        RECT 286.185 2898.335 286.515 2898.350 ;
        RECT 302.950 2894.940 303.330 2895.260 ;
        RECT 302.990 2892.925 303.290 2894.940 ;
        RECT 300.000 2892.625 304.600 2892.925 ;
      LAYER met3 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met3 ;
        RECT 688.225 3248.565 688.555 3248.580 ;
        RECT 681.880 3248.265 688.555 3248.565 ;
        RECT 688.225 3248.250 688.555 3248.265 ;
        RECT 950.000 3232.785 954.600 3233.085 ;
        RECT 941.685 3230.490 942.015 3230.505 ;
        RECT 950.670 3230.490 950.970 3232.785 ;
        RECT 941.685 3230.190 950.970 3230.490 ;
        RECT 941.685 3230.175 942.015 3230.190 ;
        RECT 950.000 3227.145 954.600 3227.445 ;
        RECT 942.145 3225.050 942.475 3225.065 ;
        RECT 950.670 3225.050 950.970 3227.145 ;
        RECT 942.145 3224.750 950.970 3225.050 ;
        RECT 942.145 3224.735 942.475 3224.750 ;
        RECT 950.000 3218.645 954.600 3218.945 ;
        RECT 942.605 3216.210 942.935 3216.225 ;
        RECT 950.670 3216.210 950.970 3218.645 ;
        RECT 942.605 3215.910 950.970 3216.210 ;
        RECT 942.605 3215.895 942.935 3215.910 ;
        RECT 950.000 3213.005 954.600 3213.305 ;
        RECT 943.065 3210.090 943.395 3210.105 ;
        RECT 950.670 3210.090 950.970 3213.005 ;
        RECT 943.065 3209.790 950.970 3210.090 ;
        RECT 943.065 3209.775 943.395 3209.790 ;
        RECT 950.000 3204.505 954.600 3204.805 ;
        RECT 943.525 3201.930 943.855 3201.945 ;
        RECT 950.670 3201.930 950.970 3204.505 ;
        RECT 943.525 3201.630 950.970 3201.930 ;
        RECT 943.525 3201.615 943.855 3201.630 ;
        RECT 950.000 3198.865 954.600 3199.165 ;
        RECT 943.985 3196.490 944.315 3196.505 ;
        RECT 950.670 3196.490 950.970 3198.865 ;
        RECT 943.985 3196.190 950.970 3196.490 ;
        RECT 943.985 3196.175 944.315 3196.190 ;
        RECT 950.000 3190.365 954.600 3190.665 ;
        RECT 944.445 3188.330 944.775 3188.345 ;
        RECT 950.670 3188.330 950.970 3190.365 ;
        RECT 944.445 3188.030 950.970 3188.330 ;
        RECT 944.445 3188.015 944.775 3188.030 ;
        RECT 696.965 2948.290 697.295 2948.305 ;
        RECT 684.790 2947.990 697.295 2948.290 ;
        RECT 684.790 2947.210 685.090 2947.990 ;
        RECT 696.965 2947.975 697.295 2947.990 ;
        RECT 681.880 2946.910 686.480 2947.210 ;
        RECT 684.790 2938.710 685.090 2946.910 ;
        RECT 681.880 2938.410 686.480 2938.710 ;
        RECT 684.790 2933.070 685.090 2938.410 ;
        RECT 681.880 2932.770 686.480 2933.070 ;
        RECT 685.710 2924.570 686.010 2932.770 ;
        RECT 681.880 2924.270 686.480 2924.570 ;
        RECT 685.710 2918.930 686.010 2924.270 ;
        RECT 681.880 2918.630 686.480 2918.930 ;
        RECT 685.710 2910.430 686.010 2918.630 ;
        RECT 681.880 2910.130 686.480 2910.430 ;
        RECT 685.710 2904.790 686.010 2910.130 ;
        RECT 681.880 2904.490 686.480 2904.790 ;
        RECT 950.000 2901.125 954.600 2901.425 ;
        RECT 944.905 2898.650 945.235 2898.665 ;
        RECT 950.670 2898.650 950.970 2901.125 ;
        RECT 944.905 2898.350 950.970 2898.650 ;
        RECT 944.905 2898.335 945.235 2898.350 ;
        RECT 944.190 2895.250 944.570 2895.260 ;
        RECT 944.190 2894.950 950.970 2895.250 ;
        RECT 944.190 2894.940 944.570 2894.950 ;
        RECT 950.670 2892.925 950.970 2894.950 ;
        RECT 950.000 2892.625 954.600 2892.925 ;
      LAYER met3 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met3 ;
        RECT 1333.145 3249.530 1333.475 3249.545 ;
        RECT 1333.145 3249.215 1333.690 3249.530 ;
        RECT 1333.390 3248.565 1333.690 3249.215 ;
        RECT 1331.880 3248.265 1336.480 3248.565 ;
        RECT 1550.000 3232.785 1554.600 3233.085 ;
        RECT 1536.925 3230.490 1537.255 3230.505 ;
        RECT 1550.510 3230.490 1550.810 3232.785 ;
        RECT 1536.925 3230.190 1550.810 3230.490 ;
        RECT 1536.925 3230.175 1537.255 3230.190 ;
        RECT 1550.000 3227.145 1554.600 3227.445 ;
        RECT 1535.545 3225.050 1535.875 3225.065 ;
        RECT 1550.510 3225.050 1550.810 3227.145 ;
        RECT 1535.545 3224.750 1550.810 3225.050 ;
        RECT 1535.545 3224.735 1535.875 3224.750 ;
        RECT 1550.000 3218.645 1554.600 3218.945 ;
        RECT 1535.545 3217.570 1535.875 3217.585 ;
        RECT 1550.510 3217.570 1550.810 3218.645 ;
        RECT 1535.545 3217.270 1550.810 3217.570 ;
        RECT 1535.545 3217.255 1535.875 3217.270 ;
        RECT 1550.000 3213.005 1554.600 3213.305 ;
        RECT 1538.305 3210.770 1538.635 3210.785 ;
        RECT 1550.510 3210.770 1550.810 3213.005 ;
        RECT 1538.305 3210.470 1550.810 3210.770 ;
        RECT 1538.305 3210.455 1538.635 3210.470 ;
        RECT 1550.000 3204.505 1554.600 3204.805 ;
        RECT 1538.305 3202.610 1538.635 3202.625 ;
        RECT 1550.510 3202.610 1550.810 3204.505 ;
        RECT 1538.305 3202.310 1550.810 3202.610 ;
        RECT 1538.305 3202.295 1538.635 3202.310 ;
        RECT 1550.000 3198.865 1554.600 3199.165 ;
        RECT 1535.085 3196.490 1535.415 3196.505 ;
        RECT 1550.510 3196.490 1550.810 3198.865 ;
        RECT 1535.085 3196.190 1550.810 3196.490 ;
        RECT 1535.085 3196.175 1535.415 3196.190 ;
        RECT 1550.000 3190.365 1554.600 3190.665 ;
        RECT 1534.165 3189.690 1534.495 3189.705 ;
        RECT 1550.510 3189.690 1550.810 3190.365 ;
        RECT 1534.165 3189.390 1550.810 3189.690 ;
        RECT 1534.165 3189.375 1534.495 3189.390 ;
        RECT 1331.880 2946.930 1336.480 2947.210 ;
        RECT 1345.565 2946.930 1345.895 2946.945 ;
        RECT 1331.880 2946.910 1345.895 2946.930 ;
        RECT 1336.150 2946.630 1345.895 2946.910 ;
        RECT 1345.565 2946.615 1345.895 2946.630 ;
        RECT 1331.880 2938.410 1336.480 2938.710 ;
        RECT 1336.150 2936.050 1336.450 2938.410 ;
        RECT 1345.565 2936.050 1345.895 2936.065 ;
        RECT 1351.750 2936.050 1352.130 2936.060 ;
        RECT 1336.150 2935.750 1352.130 2936.050 ;
        RECT 1336.150 2933.070 1336.450 2935.750 ;
        RECT 1345.565 2935.735 1345.895 2935.750 ;
        RECT 1351.750 2935.740 1352.130 2935.750 ;
        RECT 1331.880 2932.770 1336.480 2933.070 ;
        RECT 1336.150 2924.570 1336.450 2932.770 ;
        RECT 1331.880 2924.270 1336.480 2924.570 ;
        RECT 1336.150 2918.930 1336.450 2924.270 ;
        RECT 1331.880 2918.630 1336.480 2918.930 ;
        RECT 1336.150 2910.430 1336.450 2918.630 ;
        RECT 1331.880 2910.130 1336.480 2910.430 ;
        RECT 1336.150 2904.790 1336.450 2910.130 ;
        RECT 1331.880 2904.490 1336.480 2904.790 ;
        RECT 1336.150 2902.050 1336.450 2904.490 ;
        RECT 1352.005 2902.050 1352.335 2902.065 ;
        RECT 1336.150 2901.750 1352.335 2902.050 ;
        RECT 1352.005 2901.735 1352.335 2901.750 ;
        RECT 1550.000 2901.125 1554.600 2901.425 ;
        RECT 1538.305 2899.330 1538.635 2899.345 ;
        RECT 1550.510 2899.330 1550.810 2901.125 ;
        RECT 1538.305 2899.030 1550.810 2899.330 ;
        RECT 1538.305 2899.015 1538.635 2899.030 ;
        RECT 1407.665 2895.250 1407.995 2895.265 ;
        RECT 1412.470 2895.250 1412.850 2895.260 ;
        RECT 1407.665 2894.950 1412.850 2895.250 ;
        RECT 1407.665 2894.935 1407.995 2894.950 ;
        RECT 1412.470 2894.940 1412.850 2894.950 ;
        RECT 1551.390 2894.940 1551.770 2895.260 ;
        RECT 1551.430 2892.925 1551.730 2894.940 ;
        RECT 1550.000 2892.625 1554.600 2892.925 ;
      LAYER met3 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met3 ;
        RECT 1935.745 3249.530 1936.075 3249.545 ;
        RECT 1945.865 3249.530 1946.195 3249.545 ;
        RECT 1935.340 3249.230 1946.195 3249.530 ;
        RECT 1935.745 3249.215 1936.290 3249.230 ;
        RECT 1945.865 3249.215 1946.195 3249.230 ;
        RECT 1935.990 3248.565 1936.290 3249.215 ;
        RECT 1931.880 3248.265 1936.480 3248.565 ;
        RECT 2200.000 3232.785 2204.600 3233.085 ;
        RECT 2190.585 3230.490 2190.915 3230.505 ;
        RECT 2200.030 3230.490 2200.330 3232.785 ;
        RECT 2190.585 3230.190 2200.330 3230.490 ;
        RECT 2190.585 3230.175 2190.915 3230.190 ;
        RECT 2200.000 3227.145 2204.600 3227.445 ;
        RECT 2191.045 3225.050 2191.375 3225.065 ;
        RECT 2200.030 3225.050 2200.330 3227.145 ;
        RECT 2191.045 3224.750 2200.330 3225.050 ;
        RECT 2191.045 3224.735 2191.375 3224.750 ;
        RECT 2200.000 3218.645 2204.600 3218.945 ;
        RECT 2191.505 3216.210 2191.835 3216.225 ;
        RECT 2200.030 3216.210 2200.330 3218.645 ;
        RECT 2191.505 3215.910 2200.330 3216.210 ;
        RECT 2191.505 3215.895 2191.835 3215.910 ;
        RECT 2200.000 3213.005 2204.600 3213.305 ;
        RECT 2191.965 3210.090 2192.295 3210.105 ;
        RECT 2200.030 3210.090 2200.330 3213.005 ;
        RECT 2191.965 3209.790 2200.330 3210.090 ;
        RECT 2191.965 3209.775 2192.295 3209.790 ;
        RECT 2200.000 3204.505 2204.600 3204.805 ;
        RECT 2192.425 3201.930 2192.755 3201.945 ;
        RECT 2200.030 3201.930 2200.330 3204.505 ;
        RECT 2192.425 3201.630 2200.330 3201.930 ;
        RECT 2192.425 3201.615 2192.755 3201.630 ;
        RECT 2200.000 3198.865 2204.600 3199.165 ;
        RECT 2192.885 3196.490 2193.215 3196.505 ;
        RECT 2200.030 3196.490 2200.330 3198.865 ;
        RECT 2192.885 3196.190 2200.330 3196.490 ;
        RECT 2192.885 3196.175 2193.215 3196.190 ;
        RECT 2200.000 3190.365 2204.600 3190.665 ;
        RECT 2193.345 3188.330 2193.675 3188.345 ;
        RECT 2200.030 3188.330 2200.330 3190.365 ;
        RECT 2193.345 3188.030 2200.330 3188.330 ;
        RECT 2193.345 3188.015 2193.675 3188.030 ;
        RECT 1931.880 2946.910 1936.480 2947.210 ;
        RECT 1935.990 2938.710 1936.290 2946.910 ;
        RECT 1931.880 2938.410 1936.480 2938.710 ;
        RECT 1935.990 2936.050 1936.290 2938.410 ;
        RECT 1937.790 2936.050 1938.170 2936.060 ;
        RECT 1935.990 2935.750 1938.170 2936.050 ;
        RECT 1935.990 2933.070 1936.290 2935.750 ;
        RECT 1937.790 2935.740 1938.170 2935.750 ;
        RECT 1931.880 2932.770 1936.480 2933.070 ;
        RECT 1935.990 2924.570 1936.290 2932.770 ;
        RECT 1931.880 2924.270 1936.480 2924.570 ;
        RECT 1935.990 2918.930 1936.290 2924.270 ;
        RECT 1931.880 2918.630 1936.480 2918.930 ;
        RECT 1935.990 2910.430 1936.290 2918.630 ;
        RECT 1931.880 2910.130 1936.480 2910.430 ;
        RECT 1935.990 2904.790 1936.290 2910.130 ;
        RECT 1931.880 2904.770 1936.480 2904.790 ;
        RECT 1946.070 2904.770 1946.450 2904.780 ;
        RECT 1931.880 2904.490 1946.450 2904.770 ;
        RECT 1935.990 2904.470 1946.450 2904.490 ;
        RECT 1946.070 2904.460 1946.450 2904.470 ;
        RECT 2200.000 2901.125 2204.600 2901.425 ;
        RECT 2193.805 2898.650 2194.135 2898.665 ;
        RECT 2200.030 2898.650 2200.330 2901.125 ;
        RECT 2193.805 2898.350 2200.330 2898.650 ;
        RECT 2193.805 2898.335 2194.135 2898.350 ;
        RECT 2187.110 2895.250 2187.490 2895.260 ;
        RECT 2187.110 2894.950 2200.330 2895.250 ;
        RECT 2187.110 2894.940 2187.490 2894.950 ;
        RECT 2200.030 2892.925 2200.330 2894.950 ;
        RECT 2200.000 2892.625 2204.600 2892.925 ;
      LAYER met3 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met3 ;
        RECT 2582.045 3249.530 2582.375 3249.545 ;
        RECT 2582.045 3249.230 2583.050 3249.530 ;
        RECT 2582.045 3249.215 2582.375 3249.230 ;
        RECT 2582.750 3248.565 2583.050 3249.230 ;
        RECT 2581.880 3248.265 2586.480 3248.565 ;
        RECT 2581.880 2946.930 2586.480 2947.210 ;
        RECT 2594.465 2946.930 2594.795 2946.945 ;
        RECT 2581.880 2946.910 2594.795 2946.930 ;
        RECT 2585.510 2946.630 2594.795 2946.910 ;
        RECT 2594.465 2946.615 2594.795 2946.630 ;
        RECT 2594.465 2938.770 2594.795 2938.785 ;
        RECT 2585.510 2938.710 2594.795 2938.770 ;
        RECT 2581.880 2938.470 2594.795 2938.710 ;
        RECT 2581.880 2938.410 2586.480 2938.470 ;
        RECT 2594.465 2938.455 2594.795 2938.470 ;
        RECT 2585.510 2933.070 2585.810 2938.410 ;
        RECT 2581.880 2932.770 2586.480 2933.070 ;
        RECT 2585.510 2924.570 2585.810 2932.770 ;
        RECT 2581.880 2924.270 2586.480 2924.570 ;
        RECT 2585.510 2918.930 2585.810 2924.270 ;
        RECT 2581.880 2918.630 2586.480 2918.930 ;
        RECT 2585.510 2910.430 2585.810 2918.630 ;
        RECT 2581.880 2910.130 2586.480 2910.430 ;
        RECT 2585.510 2904.790 2585.810 2910.130 ;
        RECT 2581.880 2904.770 2586.480 2904.790 ;
        RECT 2594.670 2904.770 2595.050 2904.780 ;
        RECT 2581.880 2904.490 2595.050 2904.770 ;
        RECT 2585.510 2904.470 2595.050 2904.490 ;
        RECT 2594.670 2904.460 2595.050 2904.470 ;
        RECT 1054.845 2800.050 1055.175 2800.065 ;
        RECT 1055.510 2800.050 1055.890 2800.060 ;
        RECT 1054.845 2799.750 1055.890 2800.050 ;
        RECT 1054.845 2799.735 1055.175 2799.750 ;
        RECT 1055.510 2799.740 1055.890 2799.750 ;
        RECT 1742.085 2796.650 1742.415 2796.665 ;
        RECT 1759.310 2796.650 1759.690 2796.660 ;
        RECT 1742.085 2796.350 1759.690 2796.650 ;
        RECT 1742.085 2796.335 1742.415 2796.350 ;
        RECT 1759.310 2796.340 1759.690 2796.350 ;
        RECT 1790.845 2796.650 1791.175 2796.665 ;
        RECT 1794.270 2796.650 1794.650 2796.660 ;
        RECT 1790.845 2796.350 1794.650 2796.650 ;
        RECT 1790.845 2796.335 1791.175 2796.350 ;
        RECT 1794.270 2796.340 1794.650 2796.350 ;
        RECT 336.990 2794.610 337.370 2794.620 ;
        RECT 337.705 2794.610 338.035 2794.625 ;
        RECT 336.990 2794.310 338.035 2794.610 ;
        RECT 336.990 2794.300 337.370 2794.310 ;
        RECT 337.705 2794.295 338.035 2794.310 ;
        RECT 342.510 2794.610 342.890 2794.620 ;
        RECT 344.605 2794.610 344.935 2794.625 ;
        RECT 342.510 2794.310 344.935 2794.610 ;
        RECT 342.510 2794.300 342.890 2794.310 ;
        RECT 344.605 2794.295 344.935 2794.310 ;
        RECT 350.790 2794.610 351.170 2794.620 ;
        RECT 351.505 2794.610 351.835 2794.625 ;
        RECT 358.405 2794.620 358.735 2794.625 ;
        RECT 350.790 2794.310 351.835 2794.610 ;
        RECT 350.790 2794.300 351.170 2794.310 ;
        RECT 351.505 2794.295 351.835 2794.310 ;
        RECT 358.150 2794.610 358.735 2794.620 ;
        RECT 361.830 2794.610 362.210 2794.620 ;
        RECT 362.545 2794.610 362.875 2794.625 ;
        RECT 358.150 2794.310 358.960 2794.610 ;
        RECT 361.830 2794.310 362.875 2794.610 ;
        RECT 358.150 2794.300 358.735 2794.310 ;
        RECT 361.830 2794.300 362.210 2794.310 ;
        RECT 358.405 2794.295 358.735 2794.300 ;
        RECT 362.545 2794.295 362.875 2794.310 ;
        RECT 364.590 2794.610 364.970 2794.620 ;
        RECT 365.305 2794.610 365.635 2794.625 ;
        RECT 368.525 2794.620 368.855 2794.625 ;
        RECT 371.285 2794.620 371.615 2794.625 ;
        RECT 374.965 2794.620 375.295 2794.625 ;
        RECT 368.270 2794.610 368.855 2794.620 ;
        RECT 371.030 2794.610 371.615 2794.620 ;
        RECT 374.710 2794.610 375.295 2794.620 ;
        RECT 364.590 2794.310 365.635 2794.610 ;
        RECT 368.070 2794.310 368.855 2794.610 ;
        RECT 370.830 2794.310 371.615 2794.610 ;
        RECT 374.510 2794.310 375.295 2794.610 ;
        RECT 364.590 2794.300 364.970 2794.310 ;
        RECT 365.305 2794.295 365.635 2794.310 ;
        RECT 368.270 2794.300 368.855 2794.310 ;
        RECT 371.030 2794.300 371.615 2794.310 ;
        RECT 374.710 2794.300 375.295 2794.310 ;
        RECT 378.390 2794.610 378.770 2794.620 ;
        RECT 379.105 2794.610 379.435 2794.625 ;
        RECT 384.165 2794.620 384.495 2794.625 ;
        RECT 386.925 2794.620 387.255 2794.625 ;
        RECT 383.910 2794.610 384.495 2794.620 ;
        RECT 386.670 2794.610 387.255 2794.620 ;
        RECT 378.390 2794.310 379.435 2794.610 ;
        RECT 383.710 2794.310 384.495 2794.610 ;
        RECT 386.470 2794.310 387.255 2794.610 ;
        RECT 378.390 2794.300 378.770 2794.310 ;
        RECT 368.525 2794.295 368.855 2794.300 ;
        RECT 371.285 2794.295 371.615 2794.300 ;
        RECT 374.965 2794.295 375.295 2794.300 ;
        RECT 379.105 2794.295 379.435 2794.310 ;
        RECT 383.910 2794.300 384.495 2794.310 ;
        RECT 386.670 2794.300 387.255 2794.310 ;
        RECT 390.350 2794.610 390.730 2794.620 ;
        RECT 392.905 2794.610 393.235 2794.625 ;
        RECT 390.350 2794.310 393.235 2794.610 ;
        RECT 390.350 2794.300 390.730 2794.310 ;
        RECT 384.165 2794.295 384.495 2794.300 ;
        RECT 386.925 2794.295 387.255 2794.300 ;
        RECT 392.905 2794.295 393.235 2794.310 ;
        RECT 395.870 2794.610 396.250 2794.620 ;
        RECT 396.585 2794.610 396.915 2794.625 ;
        RECT 399.345 2794.620 399.675 2794.625 ;
        RECT 399.345 2794.610 399.930 2794.620 ;
        RECT 395.870 2794.310 396.915 2794.610 ;
        RECT 399.120 2794.310 399.930 2794.610 ;
        RECT 395.870 2794.300 396.250 2794.310 ;
        RECT 396.585 2794.295 396.915 2794.310 ;
        RECT 399.345 2794.300 399.930 2794.310 ;
        RECT 403.230 2794.610 403.610 2794.620 ;
        RECT 403.945 2794.610 404.275 2794.625 ;
        RECT 406.245 2794.620 406.575 2794.625 ;
        RECT 409.925 2794.620 410.255 2794.625 ;
        RECT 414.525 2794.620 414.855 2794.625 ;
        RECT 419.125 2794.620 419.455 2794.625 ;
        RECT 420.965 2794.620 421.295 2794.625 ;
        RECT 405.990 2794.610 406.575 2794.620 ;
        RECT 409.670 2794.610 410.255 2794.620 ;
        RECT 414.270 2794.610 414.855 2794.620 ;
        RECT 418.870 2794.610 419.455 2794.620 ;
        RECT 403.230 2794.310 404.275 2794.610 ;
        RECT 405.790 2794.310 406.575 2794.610 ;
        RECT 409.470 2794.310 410.255 2794.610 ;
        RECT 414.070 2794.310 414.855 2794.610 ;
        RECT 418.670 2794.310 419.455 2794.610 ;
        RECT 403.230 2794.300 403.610 2794.310 ;
        RECT 399.345 2794.295 399.675 2794.300 ;
        RECT 403.945 2794.295 404.275 2794.310 ;
        RECT 405.990 2794.300 406.575 2794.310 ;
        RECT 409.670 2794.300 410.255 2794.310 ;
        RECT 414.270 2794.300 414.855 2794.310 ;
        RECT 418.870 2794.300 419.455 2794.310 ;
        RECT 420.710 2794.610 421.295 2794.620 ;
        RECT 425.310 2794.610 425.690 2794.620 ;
        RECT 427.405 2794.610 427.735 2794.625 ;
        RECT 420.710 2794.310 421.520 2794.610 ;
        RECT 425.310 2794.310 427.735 2794.610 ;
        RECT 420.710 2794.300 421.295 2794.310 ;
        RECT 425.310 2794.300 425.690 2794.310 ;
        RECT 406.245 2794.295 406.575 2794.300 ;
        RECT 409.925 2794.295 410.255 2794.300 ;
        RECT 414.525 2794.295 414.855 2794.300 ;
        RECT 419.125 2794.295 419.455 2794.300 ;
        RECT 420.965 2794.295 421.295 2794.300 ;
        RECT 427.405 2794.295 427.735 2794.310 ;
        RECT 431.545 2794.620 431.875 2794.625 ;
        RECT 433.845 2794.620 434.175 2794.625 ;
        RECT 439.365 2794.620 439.695 2794.625 ;
        RECT 441.205 2794.620 441.535 2794.625 ;
        RECT 431.545 2794.610 432.130 2794.620 ;
        RECT 433.590 2794.610 434.175 2794.620 ;
        RECT 439.110 2794.610 439.695 2794.620 ;
        RECT 431.545 2794.310 432.330 2794.610 ;
        RECT 433.590 2794.310 434.400 2794.610 ;
        RECT 438.910 2794.310 439.695 2794.610 ;
        RECT 431.545 2794.300 432.130 2794.310 ;
        RECT 433.590 2794.300 434.175 2794.310 ;
        RECT 439.110 2794.300 439.695 2794.310 ;
        RECT 440.950 2794.610 441.535 2794.620 ;
        RECT 444.425 2794.620 444.755 2794.625 ;
        RECT 445.805 2794.620 446.135 2794.625 ;
        RECT 444.425 2794.610 445.010 2794.620 ;
        RECT 445.550 2794.610 446.135 2794.620 ;
        RECT 440.950 2794.310 441.760 2794.610 ;
        RECT 444.200 2794.310 445.010 2794.610 ;
        RECT 445.350 2794.310 446.135 2794.610 ;
        RECT 440.950 2794.300 441.535 2794.310 ;
        RECT 431.545 2794.295 431.875 2794.300 ;
        RECT 433.845 2794.295 434.175 2794.300 ;
        RECT 439.365 2794.295 439.695 2794.300 ;
        RECT 441.205 2794.295 441.535 2794.300 ;
        RECT 444.425 2794.300 445.010 2794.310 ;
        RECT 445.550 2794.300 446.135 2794.310 ;
        RECT 444.425 2794.295 444.755 2794.300 ;
        RECT 445.805 2794.295 446.135 2794.300 ;
        RECT 449.025 2794.620 449.355 2794.625 ;
        RECT 455.005 2794.620 455.335 2794.625 ;
        RECT 449.025 2794.610 449.610 2794.620 ;
        RECT 454.750 2794.610 455.335 2794.620 ;
        RECT 459.350 2794.610 459.730 2794.620 ;
        RECT 460.985 2794.610 461.315 2794.625 ;
        RECT 462.365 2794.620 462.695 2794.625 ;
        RECT 462.110 2794.610 462.695 2794.620 ;
        RECT 449.025 2794.310 449.810 2794.610 ;
        RECT 454.750 2794.310 455.560 2794.610 ;
        RECT 459.350 2794.310 461.315 2794.610 ;
        RECT 461.910 2794.310 462.695 2794.610 ;
        RECT 449.025 2794.300 449.610 2794.310 ;
        RECT 454.750 2794.300 455.335 2794.310 ;
        RECT 459.350 2794.300 459.730 2794.310 ;
        RECT 449.025 2794.295 449.355 2794.300 ;
        RECT 455.005 2794.295 455.335 2794.300 ;
        RECT 460.985 2794.295 461.315 2794.310 ;
        RECT 462.110 2794.300 462.695 2794.310 ;
        RECT 462.365 2794.295 462.695 2794.300 ;
        RECT 466.505 2794.620 466.835 2794.625 ;
        RECT 468.805 2794.620 469.135 2794.625 ;
        RECT 475.245 2794.620 475.575 2794.625 ;
        RECT 466.505 2794.610 467.090 2794.620 ;
        RECT 468.550 2794.610 469.135 2794.620 ;
        RECT 466.505 2794.310 467.290 2794.610 ;
        RECT 468.350 2794.310 469.135 2794.610 ;
        RECT 466.505 2794.300 467.090 2794.310 ;
        RECT 468.550 2794.300 469.135 2794.310 ;
        RECT 474.990 2794.610 475.575 2794.620 ;
        RECT 478.465 2794.620 478.795 2794.625 ;
        RECT 482.605 2794.620 482.935 2794.625 ;
        RECT 478.465 2794.610 479.050 2794.620 ;
        RECT 482.350 2794.610 482.935 2794.620 ;
        RECT 485.110 2794.610 485.490 2794.620 ;
        RECT 485.825 2794.610 486.155 2794.625 ;
        RECT 489.045 2794.620 489.375 2794.625 ;
        RECT 491.805 2794.620 492.135 2794.625 ;
        RECT 488.790 2794.610 489.375 2794.620 ;
        RECT 491.550 2794.610 492.135 2794.620 ;
        RECT 474.990 2794.310 475.800 2794.610 ;
        RECT 478.465 2794.310 479.250 2794.610 ;
        RECT 482.350 2794.310 483.160 2794.610 ;
        RECT 485.110 2794.310 486.155 2794.610 ;
        RECT 488.590 2794.310 489.375 2794.610 ;
        RECT 491.350 2794.310 492.135 2794.610 ;
        RECT 474.990 2794.300 475.575 2794.310 ;
        RECT 466.505 2794.295 466.835 2794.300 ;
        RECT 468.805 2794.295 469.135 2794.300 ;
        RECT 475.245 2794.295 475.575 2794.300 ;
        RECT 478.465 2794.300 479.050 2794.310 ;
        RECT 482.350 2794.300 482.935 2794.310 ;
        RECT 485.110 2794.300 485.490 2794.310 ;
        RECT 478.465 2794.295 478.795 2794.300 ;
        RECT 482.605 2794.295 482.935 2794.300 ;
        RECT 485.825 2794.295 486.155 2794.310 ;
        RECT 488.790 2794.300 489.375 2794.310 ;
        RECT 491.550 2794.300 492.135 2794.310 ;
        RECT 495.230 2794.610 495.610 2794.620 ;
        RECT 496.405 2794.610 496.735 2794.625 ;
        RECT 500.085 2794.620 500.415 2794.625 ;
        RECT 510.205 2794.620 510.535 2794.625 ;
        RECT 524.005 2794.620 524.335 2794.625 ;
        RECT 499.830 2794.610 500.415 2794.620 ;
        RECT 509.950 2794.610 510.535 2794.620 ;
        RECT 523.750 2794.610 524.335 2794.620 ;
        RECT 495.230 2794.310 496.735 2794.610 ;
        RECT 499.630 2794.310 500.415 2794.610 ;
        RECT 509.750 2794.310 510.535 2794.610 ;
        RECT 523.550 2794.310 524.335 2794.610 ;
        RECT 495.230 2794.300 495.610 2794.310 ;
        RECT 489.045 2794.295 489.375 2794.300 ;
        RECT 491.805 2794.295 492.135 2794.300 ;
        RECT 496.405 2794.295 496.735 2794.310 ;
        RECT 499.830 2794.300 500.415 2794.310 ;
        RECT 509.950 2794.300 510.535 2794.310 ;
        RECT 523.750 2794.300 524.335 2794.310 ;
        RECT 535.710 2794.610 536.090 2794.620 ;
        RECT 536.425 2794.610 536.755 2794.625 ;
        RECT 542.405 2794.620 542.735 2794.625 ;
        RECT 542.150 2794.610 542.735 2794.620 ;
        RECT 535.710 2794.310 536.755 2794.610 ;
        RECT 541.950 2794.310 542.735 2794.610 ;
        RECT 535.710 2794.300 536.090 2794.310 ;
        RECT 500.085 2794.295 500.415 2794.300 ;
        RECT 510.205 2794.295 510.535 2794.300 ;
        RECT 524.005 2794.295 524.335 2794.300 ;
        RECT 536.425 2794.295 536.755 2794.310 ;
        RECT 542.150 2794.300 542.735 2794.310 ;
        RECT 542.405 2794.295 542.735 2794.300 ;
        RECT 979.865 2794.610 980.195 2794.625 ;
        RECT 1001.025 2794.620 1001.355 2794.625 ;
        RECT 980.990 2794.610 981.370 2794.620 ;
        RECT 1001.025 2794.610 1001.610 2794.620 ;
        RECT 979.865 2794.310 981.370 2794.610 ;
        RECT 1000.800 2794.310 1001.610 2794.610 ;
        RECT 979.865 2794.295 980.195 2794.310 ;
        RECT 980.990 2794.300 981.370 2794.310 ;
        RECT 1001.025 2794.300 1001.610 2794.310 ;
        RECT 1013.190 2794.610 1013.570 2794.620 ;
        RECT 1013.905 2794.610 1014.235 2794.625 ;
        RECT 1018.965 2794.620 1019.295 2794.625 ;
        RECT 1018.710 2794.610 1019.295 2794.620 ;
        RECT 1013.190 2794.310 1014.235 2794.610 ;
        RECT 1018.510 2794.310 1019.295 2794.610 ;
        RECT 1013.190 2794.300 1013.570 2794.310 ;
        RECT 1001.025 2794.295 1001.355 2794.300 ;
        RECT 1013.905 2794.295 1014.235 2794.310 ;
        RECT 1018.710 2794.300 1019.295 2794.310 ;
        RECT 1019.630 2794.610 1020.010 2794.620 ;
        RECT 1020.805 2794.610 1021.135 2794.625 ;
        RECT 1019.630 2794.310 1021.135 2794.610 ;
        RECT 1019.630 2794.300 1020.010 2794.310 ;
        RECT 1018.965 2794.295 1019.295 2794.300 ;
        RECT 1020.805 2794.295 1021.135 2794.310 ;
        RECT 1026.990 2794.610 1027.370 2794.620 ;
        RECT 1027.705 2794.610 1028.035 2794.625 ;
        RECT 1026.990 2794.310 1028.035 2794.610 ;
        RECT 1026.990 2794.300 1027.370 2794.310 ;
        RECT 1027.705 2794.295 1028.035 2794.310 ;
        RECT 1030.670 2794.610 1031.050 2794.620 ;
        RECT 1034.605 2794.610 1034.935 2794.625 ;
        RECT 1030.670 2794.310 1034.935 2794.610 ;
        RECT 1030.670 2794.300 1031.050 2794.310 ;
        RECT 1034.605 2794.295 1034.935 2794.310 ;
        RECT 1041.710 2794.610 1042.090 2794.620 ;
        RECT 1042.425 2794.610 1042.755 2794.625 ;
        RECT 1053.005 2794.620 1053.335 2794.625 ;
        RECT 1052.750 2794.610 1053.335 2794.620 ;
        RECT 1041.710 2794.310 1042.755 2794.610 ;
        RECT 1052.550 2794.310 1053.335 2794.610 ;
        RECT 1041.710 2794.300 1042.090 2794.310 ;
        RECT 1042.425 2794.295 1042.755 2794.310 ;
        RECT 1052.750 2794.300 1053.335 2794.310 ;
        RECT 1053.005 2794.295 1053.335 2794.300 ;
        RECT 1058.985 2794.620 1059.315 2794.625 ;
        RECT 1065.885 2794.620 1066.215 2794.625 ;
        RECT 1058.985 2794.610 1059.570 2794.620 ;
        RECT 1065.630 2794.610 1066.215 2794.620 ;
        RECT 1058.985 2794.310 1059.770 2794.610 ;
        RECT 1065.430 2794.310 1066.215 2794.610 ;
        RECT 1058.985 2794.300 1059.570 2794.310 ;
        RECT 1065.630 2794.300 1066.215 2794.310 ;
        RECT 1058.985 2794.295 1059.315 2794.300 ;
        RECT 1065.885 2794.295 1066.215 2794.300 ;
        RECT 1070.025 2794.620 1070.355 2794.625 ;
        RECT 1076.465 2794.620 1076.795 2794.625 ;
        RECT 1070.025 2794.610 1070.610 2794.620 ;
        RECT 1076.465 2794.610 1077.050 2794.620 ;
        RECT 1083.110 2794.610 1083.490 2794.620 ;
        RECT 1087.505 2794.610 1087.835 2794.625 ;
        RECT 1070.025 2794.310 1070.810 2794.610 ;
        RECT 1076.465 2794.310 1077.250 2794.610 ;
        RECT 1083.110 2794.310 1087.835 2794.610 ;
        RECT 1070.025 2794.300 1070.610 2794.310 ;
        RECT 1076.465 2794.300 1077.050 2794.310 ;
        RECT 1083.110 2794.300 1083.490 2794.310 ;
        RECT 1070.025 2794.295 1070.355 2794.300 ;
        RECT 1076.465 2794.295 1076.795 2794.300 ;
        RECT 1087.505 2794.295 1087.835 2794.310 ;
        RECT 1093.945 2794.620 1094.275 2794.625 ;
        RECT 1100.385 2794.620 1100.715 2794.625 ;
        RECT 1105.445 2794.620 1105.775 2794.625 ;
        RECT 1093.945 2794.610 1094.530 2794.620 ;
        RECT 1100.385 2794.610 1100.970 2794.620 ;
        RECT 1105.190 2794.610 1105.775 2794.620 ;
        RECT 1093.945 2794.310 1094.730 2794.610 ;
        RECT 1100.385 2794.310 1101.170 2794.610 ;
        RECT 1104.990 2794.310 1105.775 2794.610 ;
        RECT 1093.945 2794.300 1094.530 2794.310 ;
        RECT 1100.385 2794.300 1100.970 2794.310 ;
        RECT 1105.190 2794.300 1105.775 2794.310 ;
        RECT 1093.945 2794.295 1094.275 2794.300 ;
        RECT 1100.385 2794.295 1100.715 2794.300 ;
        RECT 1105.445 2794.295 1105.775 2794.300 ;
        RECT 1110.965 2794.610 1111.295 2794.625 ;
        RECT 1122.465 2794.620 1122.795 2794.625 ;
        RECT 1129.365 2794.620 1129.695 2794.625 ;
        RECT 1111.630 2794.610 1112.010 2794.620 ;
        RECT 1110.965 2794.310 1112.010 2794.610 ;
        RECT 1110.965 2794.295 1111.295 2794.310 ;
        RECT 1111.630 2794.300 1112.010 2794.310 ;
        RECT 1122.465 2794.610 1123.050 2794.620 ;
        RECT 1129.110 2794.610 1129.695 2794.620 ;
        RECT 1130.745 2794.620 1131.075 2794.625 ;
        RECT 1135.805 2794.620 1136.135 2794.625 ;
        RECT 1130.745 2794.610 1131.330 2794.620 ;
        RECT 1135.550 2794.610 1136.135 2794.620 ;
        RECT 1122.465 2794.310 1123.250 2794.610 ;
        RECT 1128.910 2794.310 1129.695 2794.610 ;
        RECT 1130.520 2794.310 1131.330 2794.610 ;
        RECT 1135.350 2794.310 1136.135 2794.610 ;
        RECT 1122.465 2794.300 1123.050 2794.310 ;
        RECT 1129.110 2794.300 1129.695 2794.310 ;
        RECT 1122.465 2794.295 1122.795 2794.300 ;
        RECT 1129.365 2794.295 1129.695 2794.300 ;
        RECT 1130.745 2794.300 1131.330 2794.310 ;
        RECT 1135.550 2794.300 1136.135 2794.310 ;
        RECT 1137.390 2794.610 1137.770 2794.620 ;
        RECT 1138.105 2794.610 1138.435 2794.625 ;
        RECT 1137.390 2794.310 1138.435 2794.610 ;
        RECT 1137.390 2794.300 1137.770 2794.310 ;
        RECT 1130.745 2794.295 1131.075 2794.300 ;
        RECT 1135.805 2794.295 1136.135 2794.300 ;
        RECT 1138.105 2794.295 1138.435 2794.310 ;
        RECT 1139.945 2794.620 1140.275 2794.625 ;
        RECT 1139.945 2794.610 1140.530 2794.620 ;
        RECT 1143.830 2794.610 1144.210 2794.620 ;
        RECT 1145.005 2794.610 1145.335 2794.625 ;
        RECT 1139.945 2794.310 1140.730 2794.610 ;
        RECT 1143.830 2794.310 1145.335 2794.610 ;
        RECT 1139.945 2794.300 1140.530 2794.310 ;
        RECT 1143.830 2794.300 1144.210 2794.310 ;
        RECT 1139.945 2794.295 1140.275 2794.300 ;
        RECT 1145.005 2794.295 1145.335 2794.310 ;
        RECT 1147.305 2794.620 1147.635 2794.625 ;
        RECT 1147.305 2794.610 1147.890 2794.620 ;
        RECT 1151.190 2794.610 1151.570 2794.620 ;
        RECT 1151.905 2794.610 1152.235 2794.625 ;
        RECT 1147.305 2794.310 1148.090 2794.610 ;
        RECT 1151.190 2794.310 1152.235 2794.610 ;
        RECT 1147.305 2794.300 1147.890 2794.310 ;
        RECT 1151.190 2794.300 1151.570 2794.310 ;
        RECT 1147.305 2794.295 1147.635 2794.300 ;
        RECT 1151.905 2794.295 1152.235 2794.310 ;
        RECT 1153.950 2794.610 1154.330 2794.620 ;
        RECT 1158.805 2794.610 1159.135 2794.625 ;
        RECT 1165.245 2794.620 1165.575 2794.625 ;
        RECT 1153.950 2794.310 1159.135 2794.610 ;
        RECT 1153.950 2794.300 1154.330 2794.310 ;
        RECT 1158.805 2794.295 1159.135 2794.310 ;
        RECT 1164.990 2794.610 1165.575 2794.620 ;
        RECT 1166.165 2794.610 1166.495 2794.625 ;
        RECT 1172.605 2794.620 1172.935 2794.625 ;
        RECT 1167.750 2794.610 1168.130 2794.620 ;
        RECT 1164.990 2794.310 1165.800 2794.610 ;
        RECT 1166.165 2794.310 1168.130 2794.610 ;
        RECT 1164.990 2794.300 1165.575 2794.310 ;
        RECT 1165.245 2794.295 1165.575 2794.300 ;
        RECT 1166.165 2794.295 1166.495 2794.310 ;
        RECT 1167.750 2794.300 1168.130 2794.310 ;
        RECT 1172.350 2794.610 1172.935 2794.620 ;
        RECT 1178.790 2794.610 1179.170 2794.620 ;
        RECT 1179.505 2794.610 1179.835 2794.625 ;
        RECT 1186.405 2794.620 1186.735 2794.625 ;
        RECT 1172.350 2794.310 1173.160 2794.610 ;
        RECT 1178.790 2794.310 1179.835 2794.610 ;
        RECT 1172.350 2794.300 1172.935 2794.310 ;
        RECT 1178.790 2794.300 1179.170 2794.310 ;
        RECT 1172.605 2794.295 1172.935 2794.300 ;
        RECT 1179.505 2794.295 1179.835 2794.310 ;
        RECT 1186.150 2794.610 1186.735 2794.620 ;
        RECT 1198.110 2794.610 1198.490 2794.620 ;
        RECT 1200.205 2794.610 1200.535 2794.625 ;
        RECT 1587.065 2794.620 1587.395 2794.625 ;
        RECT 1587.065 2794.610 1587.650 2794.620 ;
        RECT 1186.150 2794.310 1186.960 2794.610 ;
        RECT 1198.110 2794.310 1200.535 2794.610 ;
        RECT 1586.840 2794.310 1587.650 2794.610 ;
        RECT 1186.150 2794.300 1186.735 2794.310 ;
        RECT 1198.110 2794.300 1198.490 2794.310 ;
        RECT 1186.405 2794.295 1186.735 2794.300 ;
        RECT 1200.205 2794.295 1200.535 2794.310 ;
        RECT 1587.065 2794.300 1587.650 2794.310 ;
        RECT 1593.965 2794.610 1594.295 2794.625 ;
        RECT 1600.865 2794.620 1601.195 2794.625 ;
        RECT 1594.630 2794.610 1595.010 2794.620 ;
        RECT 1600.865 2794.610 1601.450 2794.620 ;
        RECT 1593.965 2794.310 1595.010 2794.610 ;
        RECT 1600.640 2794.310 1601.450 2794.610 ;
        RECT 1587.065 2794.295 1587.395 2794.300 ;
        RECT 1593.965 2794.295 1594.295 2794.310 ;
        RECT 1594.630 2794.300 1595.010 2794.310 ;
        RECT 1600.865 2794.300 1601.450 2794.310 ;
        RECT 1628.465 2794.610 1628.795 2794.625 ;
        RECT 1631.430 2794.610 1631.810 2794.620 ;
        RECT 1628.465 2794.310 1631.810 2794.610 ;
        RECT 1600.865 2794.295 1601.195 2794.300 ;
        RECT 1628.465 2794.295 1628.795 2794.310 ;
        RECT 1631.430 2794.300 1631.810 2794.310 ;
        RECT 1635.365 2794.610 1635.695 2794.625 ;
        RECT 1637.870 2794.610 1638.250 2794.620 ;
        RECT 1635.365 2794.310 1638.250 2794.610 ;
        RECT 1635.365 2794.295 1635.695 2794.310 ;
        RECT 1637.870 2794.300 1638.250 2794.310 ;
        RECT 1646.405 2794.610 1646.735 2794.625 ;
        RECT 1647.990 2794.610 1648.370 2794.620 ;
        RECT 1646.405 2794.310 1648.370 2794.610 ;
        RECT 1646.405 2794.295 1646.735 2794.310 ;
        RECT 1647.990 2794.300 1648.370 2794.310 ;
        RECT 1649.625 2794.610 1649.955 2794.625 ;
        RECT 1658.825 2794.620 1659.155 2794.625 ;
        RECT 1655.350 2794.610 1655.730 2794.620 ;
        RECT 1649.625 2794.310 1655.730 2794.610 ;
        RECT 1649.625 2794.295 1649.955 2794.310 ;
        RECT 1655.350 2794.300 1655.730 2794.310 ;
        RECT 1658.825 2794.610 1659.410 2794.620 ;
        RECT 1662.965 2794.610 1663.295 2794.625 ;
        RECT 1666.390 2794.610 1666.770 2794.620 ;
        RECT 1658.825 2794.310 1659.610 2794.610 ;
        RECT 1662.965 2794.310 1666.770 2794.610 ;
        RECT 1658.825 2794.300 1659.410 2794.310 ;
        RECT 1658.825 2794.295 1659.155 2794.300 ;
        RECT 1662.965 2794.295 1663.295 2794.310 ;
        RECT 1666.390 2794.300 1666.770 2794.310 ;
        RECT 1669.865 2794.610 1670.195 2794.625 ;
        RECT 1672.830 2794.610 1673.210 2794.620 ;
        RECT 1669.865 2794.310 1673.210 2794.610 ;
        RECT 1669.865 2794.295 1670.195 2794.310 ;
        RECT 1672.830 2794.300 1673.210 2794.310 ;
        RECT 1676.765 2794.610 1677.095 2794.625 ;
        RECT 1683.665 2794.620 1683.995 2794.625 ;
        RECT 1679.270 2794.610 1679.650 2794.620 ;
        RECT 1683.665 2794.610 1684.250 2794.620 ;
        RECT 1676.765 2794.310 1679.650 2794.610 ;
        RECT 1683.440 2794.310 1684.250 2794.610 ;
        RECT 1676.765 2794.295 1677.095 2794.310 ;
        RECT 1679.270 2794.300 1679.650 2794.310 ;
        RECT 1683.665 2794.300 1684.250 2794.310 ;
        RECT 1687.805 2794.610 1688.135 2794.625 ;
        RECT 1688.470 2794.610 1688.850 2794.620 ;
        RECT 1687.805 2794.310 1688.850 2794.610 ;
        RECT 1683.665 2794.295 1683.995 2794.300 ;
        RECT 1687.805 2794.295 1688.135 2794.310 ;
        RECT 1688.470 2794.300 1688.850 2794.310 ;
        RECT 1690.565 2794.610 1690.895 2794.625 ;
        RECT 1695.830 2794.610 1696.210 2794.620 ;
        RECT 1690.565 2794.310 1696.210 2794.610 ;
        RECT 1690.565 2794.295 1690.895 2794.310 ;
        RECT 1695.830 2794.300 1696.210 2794.310 ;
        RECT 1697.465 2794.610 1697.795 2794.625 ;
        RECT 1702.270 2794.610 1702.650 2794.620 ;
        RECT 1697.465 2794.310 1702.650 2794.610 ;
        RECT 1697.465 2794.295 1697.795 2794.310 ;
        RECT 1702.270 2794.300 1702.650 2794.310 ;
        RECT 1704.365 2794.610 1704.695 2794.625 ;
        RECT 1708.710 2794.610 1709.090 2794.620 ;
        RECT 1704.365 2794.310 1709.090 2794.610 ;
        RECT 1704.365 2794.295 1704.695 2794.310 ;
        RECT 1708.710 2794.300 1709.090 2794.310 ;
        RECT 1711.265 2794.610 1711.595 2794.625 ;
        RECT 1713.310 2794.610 1713.690 2794.620 ;
        RECT 1711.265 2794.310 1713.690 2794.610 ;
        RECT 1711.265 2794.295 1711.595 2794.310 ;
        RECT 1713.310 2794.300 1713.690 2794.310 ;
        RECT 1718.625 2794.610 1718.955 2794.625 ;
        RECT 1721.385 2794.620 1721.715 2794.625 ;
        RECT 1719.750 2794.610 1720.130 2794.620 ;
        RECT 1718.625 2794.310 1720.130 2794.610 ;
        RECT 1718.625 2794.295 1718.955 2794.310 ;
        RECT 1719.750 2794.300 1720.130 2794.310 ;
        RECT 1721.385 2794.610 1721.970 2794.620 ;
        RECT 1725.065 2794.610 1725.395 2794.625 ;
        RECT 1730.790 2794.610 1731.170 2794.620 ;
        RECT 1721.385 2794.310 1722.170 2794.610 ;
        RECT 1725.065 2794.310 1731.170 2794.610 ;
        RECT 1721.385 2794.300 1721.970 2794.310 ;
        RECT 1721.385 2794.295 1721.715 2794.300 ;
        RECT 1725.065 2794.295 1725.395 2794.310 ;
        RECT 1730.790 2794.300 1731.170 2794.310 ;
        RECT 1731.965 2794.610 1732.295 2794.625 ;
        RECT 1737.230 2794.610 1737.610 2794.620 ;
        RECT 1731.965 2794.310 1737.610 2794.610 ;
        RECT 1731.965 2794.295 1732.295 2794.310 ;
        RECT 1737.230 2794.300 1737.610 2794.310 ;
        RECT 1738.865 2794.610 1739.195 2794.625 ;
        RECT 1743.670 2794.610 1744.050 2794.620 ;
        RECT 1738.865 2794.310 1744.050 2794.610 ;
        RECT 1738.865 2794.295 1739.195 2794.310 ;
        RECT 1743.670 2794.300 1744.050 2794.310 ;
        RECT 1745.765 2794.610 1746.095 2794.625 ;
        RECT 1748.270 2794.610 1748.650 2794.620 ;
        RECT 1745.765 2794.310 1748.650 2794.610 ;
        RECT 1745.765 2794.295 1746.095 2794.310 ;
        RECT 1748.270 2794.300 1748.650 2794.310 ;
        RECT 1760.025 2794.610 1760.355 2794.625 ;
        RECT 1780.265 2794.620 1780.595 2794.625 ;
        RECT 1762.070 2794.610 1762.450 2794.620 ;
        RECT 1780.265 2794.610 1780.850 2794.620 ;
        RECT 1760.025 2794.310 1762.450 2794.610 ;
        RECT 1780.040 2794.310 1780.850 2794.610 ;
        RECT 1760.025 2794.295 1760.355 2794.310 ;
        RECT 1762.070 2794.300 1762.450 2794.310 ;
        RECT 1780.265 2794.300 1780.850 2794.310 ;
        RECT 2228.765 2794.610 2229.095 2794.625 ;
        RECT 2231.270 2794.610 2231.650 2794.620 ;
        RECT 2228.765 2794.310 2231.650 2794.610 ;
        RECT 1780.265 2794.295 1780.595 2794.300 ;
        RECT 2228.765 2794.295 2229.095 2794.310 ;
        RECT 2231.270 2794.300 2231.650 2794.310 ;
        RECT 2256.365 2794.610 2256.695 2794.625 ;
        RECT 2257.030 2794.610 2257.410 2794.620 ;
        RECT 2256.365 2794.310 2257.410 2794.610 ;
        RECT 2256.365 2794.295 2256.695 2794.310 ;
        RECT 2257.030 2794.300 2257.410 2794.310 ;
        RECT 2263.265 2794.610 2263.595 2794.625 ;
        RECT 2268.325 2794.620 2268.655 2794.625 ;
        RECT 2264.390 2794.610 2264.770 2794.620 ;
        RECT 2268.070 2794.610 2268.655 2794.620 ;
        RECT 2263.265 2794.310 2264.770 2794.610 ;
        RECT 2267.870 2794.310 2268.655 2794.610 ;
        RECT 2263.265 2794.295 2263.595 2794.310 ;
        RECT 2264.390 2794.300 2264.770 2794.310 ;
        RECT 2268.070 2794.300 2268.655 2794.310 ;
        RECT 2268.325 2794.295 2268.655 2794.300 ;
        RECT 2270.165 2794.610 2270.495 2794.625 ;
        RECT 2276.350 2794.610 2276.730 2794.620 ;
        RECT 2270.165 2794.310 2276.730 2794.610 ;
        RECT 2270.165 2794.295 2270.495 2794.310 ;
        RECT 2276.350 2794.300 2276.730 2794.310 ;
        RECT 2277.065 2794.610 2277.395 2794.625 ;
        RECT 2282.790 2794.610 2283.170 2794.620 ;
        RECT 2277.065 2794.310 2283.170 2794.610 ;
        RECT 2277.065 2794.295 2277.395 2794.310 ;
        RECT 2282.790 2794.300 2283.170 2794.310 ;
        RECT 2283.965 2794.610 2284.295 2794.625 ;
        RECT 2287.390 2794.610 2287.770 2794.620 ;
        RECT 2283.965 2794.310 2287.770 2794.610 ;
        RECT 2283.965 2794.295 2284.295 2794.310 ;
        RECT 2287.390 2794.300 2287.770 2794.310 ;
        RECT 2290.865 2794.610 2291.195 2794.625 ;
        RECT 2293.830 2794.610 2294.210 2794.620 ;
        RECT 2290.865 2794.310 2294.210 2794.610 ;
        RECT 2290.865 2794.295 2291.195 2794.310 ;
        RECT 2293.830 2794.300 2294.210 2794.310 ;
        RECT 2297.765 2794.610 2298.095 2794.625 ;
        RECT 2305.125 2794.620 2305.455 2794.625 ;
        RECT 2300.270 2794.610 2300.650 2794.620 ;
        RECT 2297.765 2794.310 2300.650 2794.610 ;
        RECT 2297.765 2794.295 2298.095 2794.310 ;
        RECT 2300.270 2794.300 2300.650 2794.310 ;
        RECT 2304.870 2794.610 2305.455 2794.620 ;
        RECT 2308.345 2794.620 2308.675 2794.625 ;
        RECT 2308.345 2794.610 2308.930 2794.620 ;
        RECT 2311.565 2794.610 2311.895 2794.625 ;
        RECT 2316.830 2794.610 2317.210 2794.620 ;
        RECT 2304.870 2794.310 2305.680 2794.610 ;
        RECT 2308.345 2794.310 2309.130 2794.610 ;
        RECT 2311.565 2794.310 2317.210 2794.610 ;
        RECT 2304.870 2794.300 2305.455 2794.310 ;
        RECT 2305.125 2794.295 2305.455 2794.300 ;
        RECT 2308.345 2794.300 2308.930 2794.310 ;
        RECT 2308.345 2794.295 2308.675 2794.300 ;
        RECT 2311.565 2794.295 2311.895 2794.310 ;
        RECT 2316.830 2794.300 2317.210 2794.310 ;
        RECT 2318.465 2794.610 2318.795 2794.625 ;
        RECT 2322.350 2794.610 2322.730 2794.620 ;
        RECT 2318.465 2794.310 2322.730 2794.610 ;
        RECT 2318.465 2794.295 2318.795 2794.310 ;
        RECT 2322.350 2794.300 2322.730 2794.310 ;
        RECT 2325.365 2794.610 2325.695 2794.625 ;
        RECT 2328.790 2794.610 2329.170 2794.620 ;
        RECT 2325.365 2794.310 2329.170 2794.610 ;
        RECT 2325.365 2794.295 2325.695 2794.310 ;
        RECT 2328.790 2794.300 2329.170 2794.310 ;
        RECT 2332.265 2794.610 2332.595 2794.625 ;
        RECT 2334.310 2794.610 2334.690 2794.620 ;
        RECT 2332.265 2794.310 2334.690 2794.610 ;
        RECT 2332.265 2794.295 2332.595 2794.310 ;
        RECT 2334.310 2794.300 2334.690 2794.310 ;
        RECT 2339.165 2794.610 2339.495 2794.625 ;
        RECT 2343.765 2794.620 2344.095 2794.625 ;
        RECT 2339.830 2794.610 2340.210 2794.620 ;
        RECT 2343.510 2794.610 2344.095 2794.620 ;
        RECT 2339.165 2794.310 2340.210 2794.610 ;
        RECT 2343.310 2794.310 2344.095 2794.610 ;
        RECT 2339.165 2794.295 2339.495 2794.310 ;
        RECT 2339.830 2794.300 2340.210 2794.310 ;
        RECT 2343.510 2794.300 2344.095 2794.310 ;
        RECT 2343.765 2794.295 2344.095 2794.300 ;
        RECT 2346.065 2794.610 2346.395 2794.625 ;
        RECT 2351.790 2794.610 2352.170 2794.620 ;
        RECT 2346.065 2794.310 2352.170 2794.610 ;
        RECT 2346.065 2794.295 2346.395 2794.310 ;
        RECT 2351.790 2794.300 2352.170 2794.310 ;
        RECT 2352.965 2794.610 2353.295 2794.625 ;
        RECT 2357.310 2794.610 2357.690 2794.620 ;
        RECT 2352.965 2794.310 2357.690 2794.610 ;
        RECT 2352.965 2794.295 2353.295 2794.310 ;
        RECT 2357.310 2794.300 2357.690 2794.310 ;
        RECT 2359.865 2794.610 2360.195 2794.625 ;
        RECT 2363.750 2794.610 2364.130 2794.620 ;
        RECT 2359.865 2794.310 2364.130 2794.610 ;
        RECT 2359.865 2794.295 2360.195 2794.310 ;
        RECT 2363.750 2794.300 2364.130 2794.310 ;
        RECT 2366.765 2794.610 2367.095 2794.625 ;
        RECT 2370.190 2794.610 2370.570 2794.620 ;
        RECT 2366.765 2794.310 2370.570 2794.610 ;
        RECT 2366.765 2794.295 2367.095 2794.310 ;
        RECT 2370.190 2794.300 2370.570 2794.310 ;
        RECT 2373.665 2794.610 2373.995 2794.625 ;
        RECT 2377.345 2794.620 2377.675 2794.625 ;
        RECT 2374.790 2794.610 2375.170 2794.620 ;
        RECT 2373.665 2794.310 2375.170 2794.610 ;
        RECT 2373.665 2794.295 2373.995 2794.310 ;
        RECT 2374.790 2794.300 2375.170 2794.310 ;
        RECT 2377.345 2794.610 2377.930 2794.620 ;
        RECT 2380.565 2794.610 2380.895 2794.625 ;
        RECT 2382.865 2794.620 2383.195 2794.625 ;
        RECT 2381.230 2794.610 2381.610 2794.620 ;
        RECT 2377.345 2794.310 2378.130 2794.610 ;
        RECT 2380.565 2794.310 2381.610 2794.610 ;
        RECT 2377.345 2794.300 2377.930 2794.310 ;
        RECT 2377.345 2794.295 2377.675 2794.300 ;
        RECT 2380.565 2794.295 2380.895 2794.310 ;
        RECT 2381.230 2794.300 2381.610 2794.310 ;
        RECT 2382.865 2794.610 2383.450 2794.620 ;
        RECT 2387.925 2794.610 2388.255 2794.625 ;
        RECT 2394.825 2794.620 2395.155 2794.625 ;
        RECT 2389.510 2794.610 2389.890 2794.620 ;
        RECT 2382.865 2794.310 2383.650 2794.610 ;
        RECT 2387.925 2794.310 2389.890 2794.610 ;
        RECT 2382.865 2794.300 2383.450 2794.310 ;
        RECT 2382.865 2794.295 2383.195 2794.300 ;
        RECT 2387.925 2794.295 2388.255 2794.310 ;
        RECT 2389.510 2794.300 2389.890 2794.310 ;
        RECT 2394.825 2794.610 2395.410 2794.620 ;
        RECT 2401.725 2794.610 2402.055 2794.625 ;
        RECT 2402.390 2794.610 2402.770 2794.620 ;
        RECT 2394.825 2794.310 2395.610 2794.610 ;
        RECT 2401.725 2794.310 2402.770 2794.610 ;
        RECT 2394.825 2794.300 2395.410 2794.310 ;
        RECT 2394.825 2794.295 2395.155 2794.300 ;
        RECT 2401.725 2794.295 2402.055 2794.310 ;
        RECT 2402.390 2794.300 2402.770 2794.310 ;
        RECT 1087.965 2793.940 1088.295 2793.945 ;
        RECT 1087.710 2793.930 1088.295 2793.940 ;
        RECT 1087.510 2793.630 1088.295 2793.930 ;
        RECT 1087.710 2793.620 1088.295 2793.630 ;
        RECT 1087.965 2793.615 1088.295 2793.620 ;
        RECT 1117.865 2793.940 1118.195 2793.945 ;
        RECT 1117.865 2793.930 1118.450 2793.940 ;
        RECT 1128.190 2793.930 1128.570 2793.940 ;
        RECT 1131.205 2793.930 1131.535 2793.945 ;
        RECT 1159.265 2793.940 1159.595 2793.945 ;
        RECT 1159.265 2793.930 1159.850 2793.940 ;
        RECT 1117.865 2793.630 1118.650 2793.930 ;
        RECT 1128.190 2793.630 1131.535 2793.930 ;
        RECT 1159.040 2793.630 1159.850 2793.930 ;
        RECT 1117.865 2793.620 1118.450 2793.630 ;
        RECT 1128.190 2793.620 1128.570 2793.630 ;
        RECT 1117.865 2793.615 1118.195 2793.620 ;
        RECT 1131.205 2793.615 1131.535 2793.630 ;
        RECT 1159.265 2793.620 1159.850 2793.630 ;
        RECT 1163.150 2793.930 1163.530 2793.940 ;
        RECT 1165.705 2793.930 1166.035 2793.945 ;
        RECT 1173.065 2793.940 1173.395 2793.945 ;
        RECT 1173.065 2793.930 1173.650 2793.940 ;
        RECT 1163.150 2793.630 1166.035 2793.930 ;
        RECT 1172.840 2793.630 1173.650 2793.930 ;
        RECT 1163.150 2793.620 1163.530 2793.630 ;
        RECT 1159.265 2793.615 1159.595 2793.620 ;
        RECT 1165.705 2793.615 1166.035 2793.630 ;
        RECT 1173.065 2793.620 1173.650 2793.630 ;
        RECT 1179.965 2793.930 1180.295 2793.945 ;
        RECT 1186.865 2793.940 1187.195 2793.945 ;
        RECT 1180.630 2793.930 1181.010 2793.940 ;
        RECT 1186.865 2793.930 1187.450 2793.940 ;
        RECT 1179.965 2793.630 1181.010 2793.930 ;
        RECT 1186.640 2793.630 1187.450 2793.930 ;
        RECT 1173.065 2793.615 1173.395 2793.620 ;
        RECT 1179.965 2793.615 1180.295 2793.630 ;
        RECT 1180.630 2793.620 1181.010 2793.630 ;
        RECT 1186.865 2793.620 1187.450 2793.630 ;
        RECT 1601.325 2793.930 1601.655 2793.945 ;
        RECT 1604.750 2793.930 1605.130 2793.940 ;
        RECT 1601.325 2793.630 1605.130 2793.930 ;
        RECT 1186.865 2793.615 1187.195 2793.620 ;
        RECT 1601.325 2793.615 1601.655 2793.630 ;
        RECT 1604.750 2793.620 1605.130 2793.630 ;
        RECT 1610.985 2793.930 1611.315 2793.945 ;
        RECT 1613.030 2793.930 1613.410 2793.940 ;
        RECT 1610.985 2793.630 1613.410 2793.930 ;
        RECT 1610.985 2793.615 1611.315 2793.630 ;
        RECT 1613.030 2793.620 1613.410 2793.630 ;
        RECT 1630.510 2793.930 1630.890 2793.940 ;
        RECT 1631.685 2793.930 1632.015 2793.945 ;
        RECT 1630.510 2793.630 1632.015 2793.930 ;
        RECT 1630.510 2793.620 1630.890 2793.630 ;
        RECT 1631.685 2793.615 1632.015 2793.630 ;
        RECT 1642.265 2793.930 1642.595 2793.945 ;
        RECT 1652.385 2793.940 1652.715 2793.945 ;
        RECT 1665.725 2793.940 1666.055 2793.945 ;
        RECT 1670.325 2793.940 1670.655 2793.945 ;
        RECT 1644.310 2793.930 1644.690 2793.940 ;
        RECT 1642.265 2793.630 1644.690 2793.930 ;
        RECT 1642.265 2793.615 1642.595 2793.630 ;
        RECT 1644.310 2793.620 1644.690 2793.630 ;
        RECT 1652.385 2793.930 1652.970 2793.940 ;
        RECT 1665.470 2793.930 1666.055 2793.940 ;
        RECT 1670.070 2793.930 1670.655 2793.940 ;
        RECT 1652.385 2793.630 1653.170 2793.930 ;
        RECT 1665.270 2793.630 1666.055 2793.930 ;
        RECT 1669.870 2793.630 1670.655 2793.930 ;
        RECT 1652.385 2793.620 1652.970 2793.630 ;
        RECT 1665.470 2793.620 1666.055 2793.630 ;
        RECT 1670.070 2793.620 1670.655 2793.630 ;
        RECT 1652.385 2793.615 1652.715 2793.620 ;
        RECT 1665.725 2793.615 1666.055 2793.620 ;
        RECT 1670.325 2793.615 1670.655 2793.620 ;
        RECT 1677.225 2793.940 1677.555 2793.945 ;
        RECT 1683.205 2793.940 1683.535 2793.945 ;
        RECT 1677.225 2793.930 1677.810 2793.940 ;
        RECT 1682.950 2793.930 1683.535 2793.940 ;
        RECT 1677.225 2793.630 1678.010 2793.930 ;
        RECT 1682.750 2793.630 1683.535 2793.930 ;
        RECT 1677.225 2793.620 1677.810 2793.630 ;
        RECT 1682.950 2793.620 1683.535 2793.630 ;
        RECT 1677.225 2793.615 1677.555 2793.620 ;
        RECT 1683.205 2793.615 1683.535 2793.620 ;
        RECT 1684.125 2793.930 1684.455 2793.945 ;
        RECT 1695.165 2793.940 1695.495 2793.945 ;
        RECT 1689.390 2793.930 1689.770 2793.940 ;
        RECT 1694.910 2793.930 1695.495 2793.940 ;
        RECT 1684.125 2793.630 1689.770 2793.930 ;
        RECT 1694.710 2793.630 1695.495 2793.930 ;
        RECT 1684.125 2793.615 1684.455 2793.630 ;
        RECT 1689.390 2793.620 1689.770 2793.630 ;
        RECT 1694.910 2793.620 1695.495 2793.630 ;
        RECT 1695.165 2793.615 1695.495 2793.620 ;
        RECT 1699.305 2793.940 1699.635 2793.945 ;
        RECT 1706.205 2793.940 1706.535 2793.945 ;
        RECT 1712.645 2793.940 1712.975 2793.945 ;
        RECT 1718.165 2793.940 1718.495 2793.945 ;
        RECT 1730.125 2793.940 1730.455 2793.945 ;
        RECT 1699.305 2793.930 1699.890 2793.940 ;
        RECT 1705.950 2793.930 1706.535 2793.940 ;
        RECT 1712.390 2793.930 1712.975 2793.940 ;
        RECT 1717.910 2793.930 1718.495 2793.940 ;
        RECT 1729.870 2793.930 1730.455 2793.940 ;
        RECT 1699.305 2793.630 1700.090 2793.930 ;
        RECT 1705.750 2793.630 1706.535 2793.930 ;
        RECT 1712.190 2793.630 1712.975 2793.930 ;
        RECT 1717.710 2793.630 1718.495 2793.930 ;
        RECT 1729.670 2793.630 1730.455 2793.930 ;
        RECT 1699.305 2793.620 1699.890 2793.630 ;
        RECT 1705.950 2793.620 1706.535 2793.630 ;
        RECT 1712.390 2793.620 1712.975 2793.630 ;
        RECT 1717.910 2793.620 1718.495 2793.630 ;
        RECT 1729.870 2793.620 1730.455 2793.630 ;
        RECT 1734.470 2793.930 1734.850 2793.940 ;
        RECT 1738.405 2793.930 1738.735 2793.945 ;
        RECT 1741.165 2793.940 1741.495 2793.945 ;
        RECT 1740.910 2793.930 1741.495 2793.940 ;
        RECT 1734.470 2793.630 1738.735 2793.930 ;
        RECT 1740.710 2793.630 1741.495 2793.930 ;
        RECT 1734.470 2793.620 1734.850 2793.630 ;
        RECT 1699.305 2793.615 1699.635 2793.620 ;
        RECT 1706.205 2793.615 1706.535 2793.620 ;
        RECT 1712.645 2793.615 1712.975 2793.620 ;
        RECT 1718.165 2793.615 1718.495 2793.620 ;
        RECT 1730.125 2793.615 1730.455 2793.620 ;
        RECT 1738.405 2793.615 1738.735 2793.630 ;
        RECT 1740.910 2793.620 1741.495 2793.630 ;
        RECT 1747.350 2793.930 1747.730 2793.940 ;
        RECT 1748.525 2793.930 1748.855 2793.945 ;
        RECT 1747.350 2793.630 1748.855 2793.930 ;
        RECT 1747.350 2793.620 1747.730 2793.630 ;
        RECT 1741.165 2793.615 1741.495 2793.620 ;
        RECT 1748.525 2793.615 1748.855 2793.630 ;
        RECT 1766.465 2793.930 1766.795 2793.945 ;
        RECT 1767.590 2793.930 1767.970 2793.940 ;
        RECT 1766.465 2793.630 1767.970 2793.930 ;
        RECT 1766.465 2793.615 1766.795 2793.630 ;
        RECT 1767.590 2793.620 1767.970 2793.630 ;
        RECT 1773.365 2793.930 1773.695 2793.945 ;
        RECT 1774.030 2793.930 1774.410 2793.940 ;
        RECT 1773.365 2793.630 1774.410 2793.930 ;
        RECT 1773.365 2793.615 1773.695 2793.630 ;
        RECT 1774.030 2793.620 1774.410 2793.630 ;
        RECT 2263.725 2793.930 2264.055 2793.945 ;
        RECT 2273.845 2793.940 2274.175 2793.945 ;
        RECT 2280.285 2793.940 2280.615 2793.945 ;
        RECT 2268.990 2793.930 2269.370 2793.940 ;
        RECT 2273.590 2793.930 2274.175 2793.940 ;
        RECT 2263.725 2793.630 2269.370 2793.930 ;
        RECT 2273.390 2793.630 2274.175 2793.930 ;
        RECT 2263.725 2793.615 2264.055 2793.630 ;
        RECT 2268.990 2793.620 2269.370 2793.630 ;
        RECT 2273.590 2793.620 2274.175 2793.630 ;
        RECT 2280.030 2793.930 2280.615 2793.940 ;
        RECT 2286.470 2793.930 2286.850 2793.940 ;
        RECT 2287.185 2793.930 2287.515 2793.945 ;
        RECT 2280.030 2793.630 2280.840 2793.930 ;
        RECT 2286.470 2793.630 2287.515 2793.930 ;
        RECT 2280.030 2793.620 2280.615 2793.630 ;
        RECT 2286.470 2793.620 2286.850 2793.630 ;
        RECT 2273.845 2793.615 2274.175 2793.620 ;
        RECT 2280.285 2793.615 2280.615 2793.620 ;
        RECT 2287.185 2793.615 2287.515 2793.630 ;
        RECT 2291.990 2793.930 2292.370 2793.940 ;
        RECT 2294.085 2793.930 2294.415 2793.945 ;
        RECT 2291.990 2793.630 2294.415 2793.930 ;
        RECT 2291.990 2793.620 2292.370 2793.630 ;
        RECT 2294.085 2793.615 2294.415 2793.630 ;
        RECT 2304.665 2793.930 2304.995 2793.945 ;
        RECT 2315.245 2793.940 2315.575 2793.945 ;
        RECT 2310.390 2793.930 2310.770 2793.940 ;
        RECT 2314.990 2793.930 2315.575 2793.940 ;
        RECT 2304.665 2793.630 2310.770 2793.930 ;
        RECT 2314.790 2793.630 2315.575 2793.930 ;
        RECT 2304.665 2793.615 2304.995 2793.630 ;
        RECT 2310.390 2793.620 2310.770 2793.630 ;
        RECT 2314.990 2793.620 2315.575 2793.630 ;
        RECT 2315.245 2793.615 2315.575 2793.620 ;
        RECT 2321.225 2793.940 2321.555 2793.945 ;
        RECT 2326.285 2793.940 2326.615 2793.945 ;
        RECT 2332.725 2793.940 2333.055 2793.945 ;
        RECT 2321.225 2793.930 2321.810 2793.940 ;
        RECT 2326.030 2793.930 2326.615 2793.940 ;
        RECT 2332.470 2793.930 2333.055 2793.940 ;
        RECT 2321.225 2793.630 2322.010 2793.930 ;
        RECT 2325.830 2793.630 2326.615 2793.930 ;
        RECT 2332.270 2793.630 2333.055 2793.930 ;
        RECT 2321.225 2793.620 2321.810 2793.630 ;
        RECT 2326.030 2793.620 2326.615 2793.630 ;
        RECT 2332.470 2793.620 2333.055 2793.630 ;
        RECT 2321.225 2793.615 2321.555 2793.620 ;
        RECT 2326.285 2793.615 2326.615 2793.620 ;
        RECT 2332.725 2793.615 2333.055 2793.620 ;
        RECT 2339.625 2793.930 2339.955 2793.945 ;
        RECT 2356.645 2793.940 2356.975 2793.945 ;
        RECT 2345.350 2793.930 2345.730 2793.940 ;
        RECT 2356.390 2793.930 2356.975 2793.940 ;
        RECT 2339.625 2793.630 2345.730 2793.930 ;
        RECT 2356.190 2793.630 2356.975 2793.930 ;
        RECT 2339.625 2793.615 2339.955 2793.630 ;
        RECT 2345.350 2793.620 2345.730 2793.630 ;
        RECT 2356.390 2793.620 2356.975 2793.630 ;
        RECT 2356.645 2793.615 2356.975 2793.620 ;
        RECT 2360.785 2793.940 2361.115 2793.945 ;
        RECT 2367.225 2793.940 2367.555 2793.945 ;
        RECT 2374.125 2793.940 2374.455 2793.945 ;
        RECT 2360.785 2793.930 2361.370 2793.940 ;
        RECT 2367.225 2793.930 2367.810 2793.940 ;
        RECT 2373.870 2793.930 2374.455 2793.940 ;
        RECT 2360.785 2793.630 2361.570 2793.930 ;
        RECT 2367.225 2793.630 2368.010 2793.930 ;
        RECT 2373.670 2793.630 2374.455 2793.930 ;
        RECT 2360.785 2793.620 2361.370 2793.630 ;
        RECT 2367.225 2793.620 2367.810 2793.630 ;
        RECT 2373.870 2793.620 2374.455 2793.630 ;
        RECT 2360.785 2793.615 2361.115 2793.620 ;
        RECT 2367.225 2793.615 2367.555 2793.620 ;
        RECT 2374.125 2793.615 2374.455 2793.620 ;
        RECT 2421.965 2793.930 2422.295 2793.945 ;
        RECT 2423.550 2793.930 2423.930 2793.940 ;
        RECT 2421.965 2793.630 2423.930 2793.930 ;
        RECT 2421.965 2793.615 2422.295 2793.630 ;
        RECT 2423.550 2793.620 2423.930 2793.630 ;
        RECT 348.950 2793.250 349.330 2793.260 ;
        RECT 351.045 2793.250 351.375 2793.265 ;
        RECT 379.565 2793.260 379.895 2793.265 ;
        RECT 392.445 2793.260 392.775 2793.265 ;
        RECT 397.045 2793.260 397.375 2793.265 ;
        RECT 379.310 2793.250 379.895 2793.260 ;
        RECT 392.190 2793.250 392.775 2793.260 ;
        RECT 396.790 2793.250 397.375 2793.260 ;
        RECT 348.950 2792.950 351.375 2793.250 ;
        RECT 379.110 2792.950 379.895 2793.250 ;
        RECT 391.990 2792.950 392.775 2793.250 ;
        RECT 396.590 2792.950 397.375 2793.250 ;
        RECT 348.950 2792.940 349.330 2792.950 ;
        RECT 351.045 2792.935 351.375 2792.950 ;
        RECT 379.310 2792.940 379.895 2792.950 ;
        RECT 392.190 2792.940 392.775 2792.950 ;
        RECT 396.790 2792.940 397.375 2792.950 ;
        RECT 379.565 2792.935 379.895 2792.940 ;
        RECT 392.445 2792.935 392.775 2792.940 ;
        RECT 397.045 2792.935 397.375 2792.940 ;
        RECT 426.945 2793.260 427.275 2793.265 ;
        RECT 426.945 2793.250 427.530 2793.260 ;
        RECT 430.830 2793.250 431.210 2793.260 ;
        RECT 434.305 2793.250 434.635 2793.265 ;
        RECT 426.945 2792.950 427.730 2793.250 ;
        RECT 430.830 2792.950 434.635 2793.250 ;
        RECT 426.945 2792.940 427.530 2792.950 ;
        RECT 430.830 2792.940 431.210 2792.950 ;
        RECT 426.945 2792.935 427.275 2792.940 ;
        RECT 434.305 2792.935 434.635 2792.950 ;
        RECT 455.465 2793.260 455.795 2793.265 ;
        RECT 455.465 2793.250 456.050 2793.260 ;
        RECT 465.790 2793.250 466.170 2793.260 ;
        RECT 468.345 2793.250 468.675 2793.265 ;
        RECT 455.465 2792.950 456.250 2793.250 ;
        RECT 465.790 2792.950 468.675 2793.250 ;
        RECT 455.465 2792.940 456.050 2792.950 ;
        RECT 465.790 2792.940 466.170 2792.950 ;
        RECT 455.465 2792.935 455.795 2792.940 ;
        RECT 468.345 2792.935 468.675 2792.950 ;
        RECT 473.865 2793.260 474.195 2793.265 ;
        RECT 531.365 2793.260 531.695 2793.265 ;
        RECT 473.865 2793.250 474.450 2793.260 ;
        RECT 531.110 2793.250 531.695 2793.260 ;
        RECT 1010.685 2793.250 1011.015 2793.265 ;
        RECT 1024.485 2793.260 1024.815 2793.265 ;
        RECT 1012.270 2793.250 1012.650 2793.260 ;
        RECT 1024.230 2793.250 1024.815 2793.260 ;
        RECT 473.865 2792.950 474.650 2793.250 ;
        RECT 531.110 2792.950 531.920 2793.250 ;
        RECT 1010.685 2792.950 1012.650 2793.250 ;
        RECT 1024.030 2792.950 1024.815 2793.250 ;
        RECT 473.865 2792.940 474.450 2792.950 ;
        RECT 531.110 2792.940 531.695 2792.950 ;
        RECT 473.865 2792.935 474.195 2792.940 ;
        RECT 531.365 2792.935 531.695 2792.940 ;
        RECT 1010.685 2792.935 1011.015 2792.950 ;
        RECT 1012.270 2792.940 1012.650 2792.950 ;
        RECT 1024.230 2792.940 1024.815 2792.950 ;
        RECT 1024.485 2792.935 1024.815 2792.940 ;
        RECT 1045.185 2793.250 1045.515 2793.265 ;
        RECT 1617.885 2793.260 1618.215 2793.265 ;
        RECT 1048.150 2793.250 1048.530 2793.260 ;
        RECT 1045.185 2792.950 1048.530 2793.250 ;
        RECT 1045.185 2792.935 1045.515 2792.950 ;
        RECT 1048.150 2792.940 1048.530 2792.950 ;
        RECT 1617.630 2793.250 1618.215 2793.260 ;
        RECT 1624.070 2793.250 1624.450 2793.260 ;
        RECT 1624.785 2793.250 1625.115 2793.265 ;
        RECT 1617.630 2792.950 1618.440 2793.250 ;
        RECT 1624.070 2792.950 1625.115 2793.250 ;
        RECT 1617.630 2792.940 1618.215 2792.950 ;
        RECT 1624.070 2792.940 1624.450 2792.950 ;
        RECT 1617.885 2792.935 1618.215 2792.940 ;
        RECT 1624.785 2792.935 1625.115 2792.950 ;
        RECT 1635.110 2793.250 1635.490 2793.260 ;
        RECT 1638.585 2793.250 1638.915 2793.265 ;
        RECT 1635.110 2792.950 1638.915 2793.250 ;
        RECT 1635.110 2792.940 1635.490 2792.950 ;
        RECT 1638.585 2792.935 1638.915 2792.950 ;
        RECT 1642.470 2793.250 1642.850 2793.260 ;
        RECT 1645.485 2793.250 1645.815 2793.265 ;
        RECT 1642.470 2792.950 1645.815 2793.250 ;
        RECT 1642.470 2792.940 1642.850 2792.950 ;
        RECT 1645.485 2792.935 1645.815 2792.950 ;
        RECT 2263.470 2793.250 2263.850 2793.260 ;
        RECT 2266.485 2793.250 2266.815 2793.265 ;
        RECT 2263.470 2792.950 2266.815 2793.250 ;
        RECT 2263.470 2792.940 2263.850 2792.950 ;
        RECT 2266.485 2792.935 2266.815 2792.950 ;
        RECT 2297.510 2793.250 2297.890 2793.260 ;
        RECT 2301.905 2793.250 2302.235 2793.265 ;
        RECT 2297.510 2792.950 2302.235 2793.250 ;
        RECT 2297.510 2792.940 2297.890 2792.950 ;
        RECT 2301.905 2792.935 2302.235 2792.950 ;
        RECT 2338.910 2793.250 2339.290 2793.260 ;
        RECT 2340.085 2793.250 2340.415 2793.265 ;
        RECT 2350.205 2793.260 2350.535 2793.265 ;
        RECT 2349.950 2793.250 2350.535 2793.260 ;
        RECT 2338.910 2792.950 2340.415 2793.250 ;
        RECT 2349.750 2792.950 2350.535 2793.250 ;
        RECT 2338.910 2792.940 2339.290 2792.950 ;
        RECT 2340.085 2792.935 2340.415 2792.950 ;
        RECT 2349.950 2792.940 2350.535 2792.950 ;
        RECT 2350.205 2792.935 2350.535 2792.940 ;
        RECT 2381.025 2793.250 2381.355 2793.265 ;
        RECT 2408.165 2793.260 2408.495 2793.265 ;
        RECT 2386.750 2793.250 2387.130 2793.260 ;
        RECT 2381.025 2792.950 2387.130 2793.250 ;
        RECT 2381.025 2792.935 2381.355 2792.950 ;
        RECT 2386.750 2792.940 2387.130 2792.950 ;
        RECT 2407.910 2793.250 2408.495 2793.260 ;
        RECT 2407.910 2792.950 2408.720 2793.250 ;
        RECT 2407.910 2792.940 2408.495 2792.950 ;
        RECT 2408.165 2792.935 2408.495 2792.940 ;
        RECT 497.325 2792.570 497.655 2792.585 ;
        RECT 497.990 2792.570 498.370 2792.580 ;
        RECT 501.925 2792.570 502.255 2792.585 ;
        RECT 497.325 2792.270 502.255 2792.570 ;
        RECT 497.325 2792.255 497.655 2792.270 ;
        RECT 497.990 2792.260 498.370 2792.270 ;
        RECT 501.925 2792.255 502.255 2792.270 ;
        RECT 542.405 2792.570 542.735 2792.585 ;
        RECT 543.070 2792.570 543.450 2792.580 ;
        RECT 542.405 2792.270 543.450 2792.570 ;
        RECT 542.405 2792.255 542.735 2792.270 ;
        RECT 543.070 2792.260 543.450 2792.270 ;
        RECT 544.910 2792.570 545.290 2792.580 ;
        RECT 551.605 2792.570 551.935 2792.585 ;
        RECT 544.910 2792.270 551.935 2792.570 ;
        RECT 544.910 2792.260 545.290 2792.270 ;
        RECT 551.605 2792.255 551.935 2792.270 ;
        RECT 1159.265 2792.570 1159.595 2792.585 ;
        RECT 1752.665 2792.580 1752.995 2792.585 ;
        RECT 1164.070 2792.570 1164.450 2792.580 ;
        RECT 1159.265 2792.270 1164.450 2792.570 ;
        RECT 1159.265 2792.255 1159.595 2792.270 ;
        RECT 1164.070 2792.260 1164.450 2792.270 ;
        RECT 1752.665 2792.570 1753.250 2792.580 ;
        RECT 1787.165 2792.570 1787.495 2792.585 ;
        RECT 1787.830 2792.570 1788.210 2792.580 ;
        RECT 1752.665 2792.270 1753.450 2792.570 ;
        RECT 1787.165 2792.270 1788.210 2792.570 ;
        RECT 1752.665 2792.260 1753.250 2792.270 ;
        RECT 1752.665 2792.255 1752.995 2792.260 ;
        RECT 1787.165 2792.255 1787.495 2792.270 ;
        RECT 1787.830 2792.260 1788.210 2792.270 ;
        RECT 2394.365 2792.570 2394.695 2792.585 ;
        RECT 2398.710 2792.570 2399.090 2792.580 ;
        RECT 2394.365 2792.270 2399.090 2792.570 ;
        RECT 2394.365 2792.255 2394.695 2792.270 ;
        RECT 2398.710 2792.260 2399.090 2792.270 ;
        RECT 2408.165 2792.570 2408.495 2792.585 ;
        RECT 2415.065 2792.580 2415.395 2792.585 ;
        RECT 2410.670 2792.570 2411.050 2792.580 ;
        RECT 2415.065 2792.570 2415.650 2792.580 ;
        RECT 2408.165 2792.270 2411.050 2792.570 ;
        RECT 2414.840 2792.270 2415.650 2792.570 ;
        RECT 2408.165 2792.255 2408.495 2792.270 ;
        RECT 2410.670 2792.260 2411.050 2792.270 ;
        RECT 2415.065 2792.260 2415.650 2792.270 ;
        RECT 2428.865 2792.570 2429.195 2792.585 ;
        RECT 2429.990 2792.570 2430.370 2792.580 ;
        RECT 2428.865 2792.270 2430.370 2792.570 ;
        RECT 2415.065 2792.255 2415.395 2792.260 ;
        RECT 2428.865 2792.255 2429.195 2792.270 ;
        RECT 2429.990 2792.260 2430.370 2792.270 ;
        RECT 2435.765 2792.570 2436.095 2792.585 ;
        RECT 2436.430 2792.570 2436.810 2792.580 ;
        RECT 2435.765 2792.270 2436.810 2792.570 ;
        RECT 2435.765 2792.255 2436.095 2792.270 ;
        RECT 2436.430 2792.260 2436.810 2792.270 ;
        RECT 310.105 2791.890 310.435 2791.905 ;
        RECT 986.510 2791.890 986.890 2791.900 ;
        RECT 310.105 2791.590 986.890 2791.890 ;
        RECT 310.105 2791.575 310.435 2791.590 ;
        RECT 986.510 2791.580 986.890 2791.590 ;
        RECT 1152.365 2791.890 1152.695 2791.905 ;
        RECT 1193.765 2791.900 1194.095 2791.905 ;
        RECT 1153.030 2791.890 1153.410 2791.900 ;
        RECT 1152.365 2791.590 1153.410 2791.890 ;
        RECT 1152.365 2791.575 1152.695 2791.590 ;
        RECT 1153.030 2791.580 1153.410 2791.590 ;
        RECT 1193.510 2791.890 1194.095 2791.900 ;
        RECT 1411.550 2791.890 1411.930 2791.900 ;
        RECT 2236.790 2791.890 2237.170 2791.900 ;
        RECT 1193.510 2791.590 1194.320 2791.890 ;
        RECT 1411.550 2791.590 2237.170 2791.890 ;
        RECT 1193.510 2791.580 1194.095 2791.590 ;
        RECT 1411.550 2791.580 1411.930 2791.590 ;
        RECT 2236.790 2791.580 2237.170 2791.590 ;
        RECT 2387.465 2791.890 2387.795 2791.905 ;
        RECT 2392.270 2791.890 2392.650 2791.900 ;
        RECT 2387.465 2791.590 2392.650 2791.890 ;
        RECT 1193.765 2791.575 1194.095 2791.580 ;
        RECT 2387.465 2791.575 2387.795 2791.590 ;
        RECT 2392.270 2791.580 2392.650 2791.590 ;
        RECT 2401.725 2791.890 2402.055 2791.905 ;
        RECT 2442.665 2791.900 2442.995 2791.905 ;
        RECT 2404.230 2791.890 2404.610 2791.900 ;
        RECT 2442.665 2791.890 2443.250 2791.900 ;
        RECT 2401.725 2791.590 2404.610 2791.890 ;
        RECT 2442.440 2791.590 2443.250 2791.890 ;
        RECT 2401.725 2791.575 2402.055 2791.590 ;
        RECT 2404.230 2791.580 2404.610 2791.590 ;
        RECT 2442.665 2791.580 2443.250 2791.590 ;
        RECT 2442.665 2791.575 2442.995 2791.580 ;
        RECT 317.005 2791.210 317.335 2791.225 ;
        RECT 993.870 2791.210 994.250 2791.220 ;
        RECT 317.005 2790.910 994.250 2791.210 ;
        RECT 317.005 2790.895 317.335 2790.910 ;
        RECT 993.870 2790.900 994.250 2790.910 ;
        RECT 1417.070 2791.210 1417.450 2791.220 ;
        RECT 2242.310 2791.210 2242.690 2791.220 ;
        RECT 1417.070 2790.910 2242.690 2791.210 ;
        RECT 1417.070 2790.900 1417.450 2790.910 ;
        RECT 2242.310 2790.900 2242.690 2790.910 ;
        RECT 2415.065 2791.210 2415.395 2791.225 ;
        RECT 2420.790 2791.210 2421.170 2791.220 ;
        RECT 2415.065 2790.910 2421.170 2791.210 ;
        RECT 2415.065 2790.895 2415.395 2790.910 ;
        RECT 2420.790 2790.900 2421.170 2790.910 ;
        RECT 1191.670 2790.530 1192.050 2790.540 ;
        RECT 1193.305 2790.530 1193.635 2790.545 ;
        RECT 1191.670 2790.230 1193.635 2790.530 ;
        RECT 1191.670 2790.220 1192.050 2790.230 ;
        RECT 1193.305 2790.215 1193.635 2790.230 ;
        RECT 1607.765 2790.530 1608.095 2790.545 ;
        RECT 1613.950 2790.530 1614.330 2790.540 ;
        RECT 1607.765 2790.230 1614.330 2790.530 ;
        RECT 1607.765 2790.215 1608.095 2790.230 ;
        RECT 1613.950 2790.220 1614.330 2790.230 ;
        RECT 1614.665 2790.530 1614.995 2790.545 ;
        RECT 1620.390 2790.530 1620.770 2790.540 ;
        RECT 1614.665 2790.230 1620.770 2790.530 ;
        RECT 1614.665 2790.215 1614.995 2790.230 ;
        RECT 1620.390 2790.220 1620.770 2790.230 ;
        RECT 2421.965 2790.530 2422.295 2790.545 ;
        RECT 2428.150 2790.530 2428.530 2790.540 ;
        RECT 2421.965 2790.230 2428.530 2790.530 ;
        RECT 2421.965 2790.215 2422.295 2790.230 ;
        RECT 2428.150 2790.220 2428.530 2790.230 ;
        RECT 413.605 2789.860 413.935 2789.865 ;
        RECT 413.350 2789.850 413.935 2789.860 ;
        RECT 538.470 2789.850 538.850 2789.860 ;
        RECT 541.485 2789.850 541.815 2789.865 ;
        RECT 1649.165 2789.860 1649.495 2789.865 ;
        RECT 413.350 2789.550 414.160 2789.850 ;
        RECT 538.470 2789.550 541.815 2789.850 ;
        RECT 413.350 2789.540 413.935 2789.550 ;
        RECT 538.470 2789.540 538.850 2789.550 ;
        RECT 413.605 2789.535 413.935 2789.540 ;
        RECT 541.485 2789.535 541.815 2789.550 ;
        RECT 1648.910 2789.850 1649.495 2789.860 ;
        RECT 2415.065 2789.850 2415.395 2789.865 ;
        RECT 2417.110 2789.850 2417.490 2789.860 ;
        RECT 1648.910 2789.550 1649.720 2789.850 ;
        RECT 2415.065 2789.550 2417.490 2789.850 ;
        RECT 1648.910 2789.540 1649.495 2789.550 ;
        RECT 1649.165 2789.535 1649.495 2789.540 ;
        RECT 2415.065 2789.535 2415.395 2789.550 ;
        RECT 2417.110 2789.540 2417.490 2789.550 ;
        RECT 2428.865 2789.850 2429.195 2789.865 ;
        RECT 2434.590 2789.850 2434.970 2789.860 ;
        RECT 2428.865 2789.550 2434.970 2789.850 ;
        RECT 2428.865 2789.535 2429.195 2789.550 ;
        RECT 2434.590 2789.540 2434.970 2789.550 ;
        RECT 504.225 2789.170 504.555 2789.185 ;
        RECT 506.985 2789.170 507.315 2789.185 ;
        RECT 1581.545 2789.180 1581.875 2789.185 ;
        RECT 508.110 2789.170 508.490 2789.180 ;
        RECT 1581.545 2789.170 1582.130 2789.180 ;
        RECT 504.225 2788.870 508.490 2789.170 ;
        RECT 1581.320 2788.870 1582.130 2789.170 ;
        RECT 504.225 2788.855 504.555 2788.870 ;
        RECT 506.985 2788.855 507.315 2788.870 ;
        RECT 508.110 2788.860 508.490 2788.870 ;
        RECT 1581.545 2788.860 1582.130 2788.870 ;
        RECT 1656.065 2789.170 1656.395 2789.185 ;
        RECT 2249.465 2789.180 2249.795 2789.185 ;
        RECT 1661.790 2789.170 1662.170 2789.180 ;
        RECT 2249.465 2789.170 2250.050 2789.180 ;
        RECT 1656.065 2788.870 1662.170 2789.170 ;
        RECT 2249.240 2788.870 2250.050 2789.170 ;
        RECT 1581.545 2788.855 1581.875 2788.860 ;
        RECT 1656.065 2788.855 1656.395 2788.870 ;
        RECT 1661.790 2788.860 1662.170 2788.870 ;
        RECT 2249.465 2788.860 2250.050 2788.870 ;
        RECT 2415.065 2789.170 2415.395 2789.185 ;
        RECT 2418.030 2789.170 2418.410 2789.180 ;
        RECT 2415.065 2788.870 2418.410 2789.170 ;
        RECT 2249.465 2788.855 2249.795 2788.860 ;
        RECT 2415.065 2788.855 2415.395 2788.870 ;
        RECT 2418.030 2788.860 2418.410 2788.870 ;
        RECT 2435.765 2789.170 2436.095 2789.185 ;
        RECT 2439.190 2789.170 2439.570 2789.180 ;
        RECT 2435.765 2788.870 2439.570 2789.170 ;
        RECT 2435.765 2788.855 2436.095 2788.870 ;
        RECT 2439.190 2788.860 2439.570 2788.870 ;
        RECT 500.085 2788.490 500.415 2788.505 ;
        RECT 500.750 2788.490 501.130 2788.500 ;
        RECT 500.085 2788.190 501.130 2788.490 ;
        RECT 500.085 2788.175 500.415 2788.190 ;
        RECT 500.750 2788.180 501.130 2788.190 ;
        RECT 531.110 2788.490 531.490 2788.500 ;
        RECT 534.585 2788.490 534.915 2788.505 ;
        RECT 1007.465 2788.500 1007.795 2788.505 ;
        RECT 1007.465 2788.490 1008.050 2788.500 ;
        RECT 531.110 2788.190 534.915 2788.490 ;
        RECT 1007.240 2788.190 1008.050 2788.490 ;
        RECT 531.110 2788.180 531.490 2788.190 ;
        RECT 534.585 2788.175 534.915 2788.190 ;
        RECT 1007.465 2788.180 1008.050 2788.190 ;
        RECT 1035.270 2788.490 1035.650 2788.500 ;
        RECT 1038.285 2788.490 1038.615 2788.505 ;
        RECT 1035.270 2788.190 1038.615 2788.490 ;
        RECT 1035.270 2788.180 1035.650 2788.190 ;
        RECT 1007.465 2788.175 1007.795 2788.180 ;
        RECT 1038.285 2788.175 1038.615 2788.190 ;
        RECT 1051.830 2788.490 1052.210 2788.500 ;
        RECT 1055.305 2788.490 1055.635 2788.505 ;
        RECT 1051.830 2788.190 1055.635 2788.490 ;
        RECT 1051.830 2788.180 1052.210 2788.190 ;
        RECT 1055.305 2788.175 1055.635 2788.190 ;
        RECT 1086.790 2788.490 1087.170 2788.500 ;
        RECT 1089.805 2788.490 1090.135 2788.505 ;
        RECT 1086.790 2788.190 1090.135 2788.490 ;
        RECT 1086.790 2788.180 1087.170 2788.190 ;
        RECT 1089.805 2788.175 1090.135 2788.190 ;
        RECT 1621.565 2788.490 1621.895 2788.505 ;
        RECT 1626.830 2788.490 1627.210 2788.500 ;
        RECT 1621.565 2788.190 1627.210 2788.490 ;
        RECT 1621.565 2788.175 1621.895 2788.190 ;
        RECT 1626.830 2788.180 1627.210 2788.190 ;
        RECT 1718.165 2788.490 1718.495 2788.505 ;
        RECT 1724.350 2788.490 1724.730 2788.500 ;
        RECT 1718.165 2788.190 1724.730 2788.490 ;
        RECT 1718.165 2788.175 1718.495 2788.190 ;
        RECT 1724.350 2788.180 1724.730 2788.190 ;
        RECT 1760.485 2788.490 1760.815 2788.505 ;
        RECT 2304.205 2788.500 2304.535 2788.505 ;
        RECT 1765.750 2788.490 1766.130 2788.500 ;
        RECT 2303.950 2788.490 2304.535 2788.500 ;
        RECT 1760.485 2788.190 1766.130 2788.490 ;
        RECT 2303.750 2788.190 2304.535 2788.490 ;
        RECT 1760.485 2788.175 1760.815 2788.190 ;
        RECT 1765.750 2788.180 1766.130 2788.190 ;
        RECT 2303.950 2788.180 2304.535 2788.190 ;
        RECT 2304.205 2788.175 2304.535 2788.180 ;
        RECT 2442.665 2788.490 2442.995 2788.505 ;
        RECT 2445.630 2788.490 2446.010 2788.500 ;
        RECT 2442.665 2788.190 2446.010 2788.490 ;
        RECT 2442.665 2788.175 2442.995 2788.190 ;
        RECT 2445.630 2788.180 2446.010 2788.190 ;
        RECT 507.190 2787.810 507.570 2787.820 ;
        RECT 510.205 2787.810 510.535 2787.825 ;
        RECT 513.885 2787.820 514.215 2787.825 ;
        RECT 513.630 2787.810 514.215 2787.820 ;
        RECT 507.190 2787.510 510.535 2787.810 ;
        RECT 513.430 2787.510 514.215 2787.810 ;
        RECT 507.190 2787.500 507.570 2787.510 ;
        RECT 510.205 2787.495 510.535 2787.510 ;
        RECT 513.630 2787.500 514.215 2787.510 ;
        RECT 516.390 2787.810 516.770 2787.820 ;
        RECT 517.105 2787.810 517.435 2787.825 ;
        RECT 516.390 2787.510 517.435 2787.810 ;
        RECT 516.390 2787.500 516.770 2787.510 ;
        RECT 513.885 2787.495 514.215 2787.500 ;
        RECT 517.105 2787.495 517.435 2787.510 ;
        RECT 520.070 2787.810 520.450 2787.820 ;
        RECT 520.785 2787.810 521.115 2787.825 ;
        RECT 520.070 2787.510 521.115 2787.810 ;
        RECT 520.070 2787.500 520.450 2787.510 ;
        RECT 520.785 2787.495 521.115 2787.510 ;
        RECT 526.510 2787.810 526.890 2787.820 ;
        RECT 527.685 2787.810 528.015 2787.825 ;
        RECT 526.510 2787.510 528.015 2787.810 ;
        RECT 526.510 2787.500 526.890 2787.510 ;
        RECT 527.685 2787.495 528.015 2787.510 ;
        RECT 530.190 2787.810 530.570 2787.820 ;
        RECT 530.905 2787.810 531.235 2787.825 ;
        RECT 1034.605 2787.820 1034.935 2787.825 ;
        RECT 530.190 2787.510 531.235 2787.810 ;
        RECT 530.190 2787.500 530.570 2787.510 ;
        RECT 530.905 2787.495 531.235 2787.510 ;
        RECT 1034.350 2787.810 1034.935 2787.820 ;
        RECT 1039.870 2787.810 1040.250 2787.820 ;
        RECT 1041.505 2787.810 1041.835 2787.825 ;
        RECT 1034.350 2787.510 1035.160 2787.810 ;
        RECT 1039.870 2787.510 1041.835 2787.810 ;
        RECT 1034.350 2787.500 1034.935 2787.510 ;
        RECT 1039.870 2787.500 1040.250 2787.510 ;
        RECT 1034.605 2787.495 1034.935 2787.500 ;
        RECT 1041.505 2787.495 1041.835 2787.510 ;
        RECT 1046.310 2787.810 1046.690 2787.820 ;
        RECT 1048.405 2787.810 1048.735 2787.825 ;
        RECT 1062.205 2787.820 1062.535 2787.825 ;
        RECT 1046.310 2787.510 1048.735 2787.810 ;
        RECT 1046.310 2787.500 1046.690 2787.510 ;
        RECT 1048.405 2787.495 1048.735 2787.510 ;
        RECT 1061.950 2787.810 1062.535 2787.820 ;
        RECT 1067.470 2787.810 1067.850 2787.820 ;
        RECT 1069.105 2787.810 1069.435 2787.825 ;
        RECT 1061.950 2787.510 1062.760 2787.810 ;
        RECT 1067.470 2787.510 1069.435 2787.810 ;
        RECT 1061.950 2787.500 1062.535 2787.510 ;
        RECT 1067.470 2787.500 1067.850 2787.510 ;
        RECT 1062.205 2787.495 1062.535 2787.500 ;
        RECT 1069.105 2787.495 1069.435 2787.510 ;
        RECT 1073.910 2787.810 1074.290 2787.820 ;
        RECT 1076.005 2787.810 1076.335 2787.825 ;
        RECT 1073.910 2787.510 1076.335 2787.810 ;
        RECT 1073.910 2787.500 1074.290 2787.510 ;
        RECT 1076.005 2787.495 1076.335 2787.510 ;
        RECT 1081.270 2787.810 1081.650 2787.820 ;
        RECT 1082.905 2787.810 1083.235 2787.825 ;
        RECT 1089.345 2787.820 1089.675 2787.825 ;
        RECT 1089.345 2787.810 1089.930 2787.820 ;
        RECT 1081.270 2787.510 1083.235 2787.810 ;
        RECT 1089.120 2787.510 1089.930 2787.810 ;
        RECT 1081.270 2787.500 1081.650 2787.510 ;
        RECT 1082.905 2787.495 1083.235 2787.510 ;
        RECT 1089.345 2787.500 1089.930 2787.510 ;
        RECT 1095.990 2787.810 1096.370 2787.820 ;
        RECT 1096.705 2787.810 1097.035 2787.825 ;
        RECT 1103.605 2787.820 1103.935 2787.825 ;
        RECT 1095.990 2787.510 1097.035 2787.810 ;
        RECT 1095.990 2787.500 1096.370 2787.510 ;
        RECT 1089.345 2787.495 1089.675 2787.500 ;
        RECT 1096.705 2787.495 1097.035 2787.510 ;
        RECT 1103.350 2787.810 1103.935 2787.820 ;
        RECT 1109.790 2787.810 1110.170 2787.820 ;
        RECT 1110.505 2787.810 1110.835 2787.825 ;
        RECT 1103.350 2787.510 1104.160 2787.810 ;
        RECT 1109.790 2787.510 1110.835 2787.810 ;
        RECT 1103.350 2787.500 1103.935 2787.510 ;
        RECT 1109.790 2787.500 1110.170 2787.510 ;
        RECT 1103.605 2787.495 1103.935 2787.500 ;
        RECT 1110.505 2787.495 1110.835 2787.510 ;
        RECT 1116.230 2787.810 1116.610 2787.820 ;
        RECT 1117.405 2787.810 1117.735 2787.825 ;
        RECT 1116.230 2787.510 1117.735 2787.810 ;
        RECT 1116.230 2787.500 1116.610 2787.510 ;
        RECT 1117.405 2787.495 1117.735 2787.510 ;
        RECT 1121.750 2787.810 1122.130 2787.820 ;
        RECT 1124.305 2787.810 1124.635 2787.825 ;
        RECT 1121.750 2787.510 1124.635 2787.810 ;
        RECT 1121.750 2787.500 1122.130 2787.510 ;
        RECT 1124.305 2787.495 1124.635 2787.510 ;
        RECT 1753.125 2787.810 1753.455 2787.825 ;
        RECT 1754.710 2787.810 1755.090 2787.820 ;
        RECT 1753.125 2787.510 1755.090 2787.810 ;
        RECT 1753.125 2787.495 1753.455 2787.510 ;
        RECT 1754.710 2787.500 1755.090 2787.510 ;
        RECT 1766.465 2787.810 1766.795 2787.825 ;
        RECT 1772.190 2787.810 1772.570 2787.820 ;
        RECT 1766.465 2787.510 1772.570 2787.810 ;
        RECT 1766.465 2787.495 1766.795 2787.510 ;
        RECT 1772.190 2787.500 1772.570 2787.510 ;
        RECT 1773.365 2787.810 1773.695 2787.825 ;
        RECT 1778.630 2787.810 1779.010 2787.820 ;
        RECT 1773.365 2787.510 1779.010 2787.810 ;
        RECT 1773.365 2787.495 1773.695 2787.510 ;
        RECT 1778.630 2787.500 1779.010 2787.510 ;
        RECT 1780.725 2787.810 1781.055 2787.825 ;
        RECT 1783.230 2787.810 1783.610 2787.820 ;
        RECT 1780.725 2787.510 1783.610 2787.810 ;
        RECT 1780.725 2787.495 1781.055 2787.510 ;
        RECT 1783.230 2787.500 1783.610 2787.510 ;
        RECT 1787.625 2787.810 1787.955 2787.825 ;
        RECT 1789.670 2787.810 1790.050 2787.820 ;
        RECT 1787.625 2787.510 1790.050 2787.810 ;
        RECT 1787.625 2787.495 1787.955 2787.510 ;
        RECT 1789.670 2787.500 1790.050 2787.510 ;
        RECT 1760.025 2777.610 1760.355 2777.625 ;
        RECT 1761.150 2777.610 1761.530 2777.620 ;
        RECT 1760.025 2777.310 1761.530 2777.610 ;
        RECT 1760.025 2777.295 1760.355 2777.310 ;
        RECT 1761.150 2777.300 1761.530 2777.310 ;
        RECT 1794.525 2777.610 1794.855 2777.625 ;
        RECT 1796.110 2777.610 1796.490 2777.620 ;
        RECT 1794.525 2777.310 1796.490 2777.610 ;
        RECT 1794.525 2777.295 1794.855 2777.310 ;
        RECT 1796.110 2777.300 1796.490 2777.310 ;
        RECT 700.185 2718.450 700.515 2718.465 ;
        RECT 1000.105 2718.450 1000.435 2718.465 ;
        RECT 700.185 2718.150 1000.435 2718.450 ;
        RECT 700.185 2718.135 700.515 2718.150 ;
        RECT 1000.105 2718.135 1000.435 2718.150 ;
        RECT 741.585 2717.770 741.915 2717.785 ;
        RECT 1052.085 2717.770 1052.415 2717.785 ;
        RECT 741.585 2717.470 1052.415 2717.770 ;
        RECT 741.585 2717.455 741.915 2717.470 ;
        RECT 1052.085 2717.455 1052.415 2717.470 ;
        RECT 707.085 2717.090 707.415 2717.105 ;
        RECT 1041.505 2717.090 1041.835 2717.105 ;
        RECT 707.085 2716.790 1041.835 2717.090 ;
        RECT 707.085 2716.775 707.415 2716.790 ;
        RECT 1041.505 2716.775 1041.835 2716.790 ;
        RECT 481.225 2716.410 481.555 2716.425 ;
        RECT 941.685 2716.410 942.015 2716.425 ;
        RECT 481.225 2716.110 942.015 2716.410 ;
        RECT 481.225 2716.095 481.555 2716.110 ;
        RECT 941.685 2716.095 942.015 2716.110 ;
        RECT 517.105 2715.730 517.435 2715.745 ;
        RECT 1010.225 2715.730 1010.555 2715.745 ;
        RECT 517.105 2715.430 1010.555 2715.730 ;
        RECT 517.105 2715.415 517.435 2715.430 ;
        RECT 1010.225 2715.415 1010.555 2715.430 ;
        RECT 387.845 2715.050 388.175 2715.065 ;
        RECT 944.905 2715.050 945.235 2715.065 ;
        RECT 387.845 2714.750 945.235 2715.050 ;
        RECT 387.845 2714.735 388.175 2714.750 ;
        RECT 944.905 2714.735 945.235 2714.750 ;
        RECT 1396.000 2697.370 1400.000 2697.480 ;
        RECT 1411.345 2697.370 1411.675 2697.385 ;
      LAYER met3 ;
        RECT 300.065 2696.480 1395.600 2697.340 ;
      LAYER met3 ;
        RECT 1396.000 2697.070 1411.675 2697.370 ;
        RECT 1396.000 2696.880 1400.000 2697.070 ;
        RECT 1411.345 2697.055 1411.675 2697.070 ;
      LAYER met3 ;
        RECT 300.065 2695.840 1396.000 2696.480 ;
      LAYER met3 ;
        RECT 300.000 2694.840 304.000 2695.440 ;
      LAYER met3 ;
        RECT 304.400 2694.440 1396.000 2695.840 ;
        RECT 300.065 2693.120 1396.000 2694.440 ;
        RECT 300.065 2691.720 1395.600 2693.120 ;
      LAYER met3 ;
        RECT 1396.000 2692.610 1400.000 2692.720 ;
        RECT 1414.105 2692.610 1414.435 2692.625 ;
        RECT 1396.000 2692.310 1414.435 2692.610 ;
        RECT 1396.000 2692.120 1400.000 2692.310 ;
        RECT 1414.105 2692.295 1414.435 2692.310 ;
      LAYER met3 ;
        RECT 300.065 2687.680 1396.000 2691.720 ;
        RECT 300.065 2686.320 1395.600 2687.680 ;
      LAYER met3 ;
        RECT 1396.000 2687.170 1400.000 2687.280 ;
        RECT 1414.105 2687.170 1414.435 2687.185 ;
        RECT 1396.000 2686.870 1414.435 2687.170 ;
        RECT 1396.000 2686.680 1400.000 2686.870 ;
        RECT 1414.105 2686.855 1414.435 2686.870 ;
      LAYER met3 ;
        RECT 304.400 2686.280 1395.600 2686.320 ;
      LAYER met3 ;
        RECT 300.000 2685.320 304.000 2685.920 ;
      LAYER met3 ;
        RECT 304.400 2684.920 1396.000 2686.280 ;
        RECT 300.065 2682.920 1396.000 2684.920 ;
        RECT 300.065 2681.520 1395.600 2682.920 ;
      LAYER met3 ;
        RECT 1396.000 2682.410 1400.000 2682.520 ;
        RECT 1414.105 2682.410 1414.435 2682.425 ;
        RECT 1396.000 2682.110 1414.435 2682.410 ;
        RECT 1396.000 2681.920 1400.000 2682.110 ;
        RECT 1414.105 2682.095 1414.435 2682.110 ;
      LAYER met3 ;
        RECT 300.065 2677.480 1396.000 2681.520 ;
        RECT 300.065 2676.800 1395.600 2677.480 ;
      LAYER met3 ;
        RECT 300.000 2675.800 304.000 2676.400 ;
      LAYER met3 ;
        RECT 304.400 2676.080 1395.600 2676.800 ;
      LAYER met3 ;
        RECT 1396.000 2676.970 1400.000 2677.080 ;
        RECT 1408.585 2676.970 1408.915 2676.985 ;
        RECT 1396.000 2676.670 1408.915 2676.970 ;
        RECT 1396.000 2676.480 1400.000 2676.670 ;
        RECT 1408.585 2676.655 1408.915 2676.670 ;
      LAYER met3 ;
        RECT 304.400 2675.400 1396.000 2676.080 ;
        RECT 300.065 2672.720 1396.000 2675.400 ;
        RECT 300.065 2671.320 1395.600 2672.720 ;
      LAYER met3 ;
        RECT 1396.000 2672.210 1400.000 2672.320 ;
        RECT 1410.425 2672.210 1410.755 2672.225 ;
        RECT 1396.000 2671.910 1410.755 2672.210 ;
        RECT 1396.000 2671.720 1400.000 2671.910 ;
        RECT 1410.425 2671.895 1410.755 2671.910 ;
      LAYER met3 ;
        RECT 300.065 2667.960 1396.000 2671.320 ;
        RECT 300.065 2667.280 1395.600 2667.960 ;
      LAYER met3 ;
        RECT 300.000 2666.280 304.000 2666.880 ;
      LAYER met3 ;
        RECT 304.400 2666.560 1395.600 2667.280 ;
      LAYER met3 ;
        RECT 1396.000 2667.450 1400.000 2667.560 ;
        RECT 1410.425 2667.450 1410.755 2667.465 ;
        RECT 1396.000 2667.150 1410.755 2667.450 ;
        RECT 1396.000 2666.960 1400.000 2667.150 ;
        RECT 1410.425 2667.135 1410.755 2667.150 ;
      LAYER met3 ;
        RECT 304.400 2665.880 1396.000 2666.560 ;
        RECT 300.065 2662.520 1396.000 2665.880 ;
        RECT 300.065 2661.120 1395.600 2662.520 ;
      LAYER met3 ;
        RECT 1396.000 2662.010 1400.000 2662.120 ;
        RECT 1411.345 2662.010 1411.675 2662.025 ;
        RECT 1396.000 2661.710 1411.675 2662.010 ;
        RECT 1396.000 2661.520 1400.000 2661.710 ;
        RECT 1411.345 2661.695 1411.675 2661.710 ;
      LAYER met3 ;
        RECT 300.065 2657.760 1396.000 2661.120 ;
      LAYER met3 ;
        RECT 300.000 2656.760 304.000 2657.360 ;
      LAYER met3 ;
        RECT 304.400 2656.360 1395.600 2657.760 ;
      LAYER met3 ;
        RECT 1396.000 2657.250 1400.000 2657.360 ;
        RECT 1414.105 2657.250 1414.435 2657.265 ;
        RECT 1396.000 2656.950 1414.435 2657.250 ;
        RECT 1396.000 2656.760 1400.000 2656.950 ;
        RECT 1414.105 2656.935 1414.435 2656.950 ;
      LAYER met3 ;
        RECT 300.065 2652.320 1396.000 2656.360 ;
        RECT 300.065 2650.920 1395.600 2652.320 ;
      LAYER met3 ;
        RECT 1396.000 2651.810 1400.000 2651.920 ;
        RECT 1414.105 2651.810 1414.435 2651.825 ;
        RECT 1396.000 2651.510 1414.435 2651.810 ;
        RECT 1396.000 2651.320 1400.000 2651.510 ;
        RECT 1414.105 2651.495 1414.435 2651.510 ;
      LAYER met3 ;
        RECT 300.065 2647.560 1396.000 2650.920 ;
      LAYER met3 ;
        RECT 300.000 2646.560 304.000 2647.160 ;
      LAYER met3 ;
        RECT 304.400 2646.160 1395.600 2647.560 ;
      LAYER met3 ;
        RECT 1396.000 2647.050 1400.000 2647.160 ;
        RECT 1414.105 2647.050 1414.435 2647.065 ;
        RECT 1396.000 2646.750 1414.435 2647.050 ;
        RECT 1396.000 2646.560 1400.000 2646.750 ;
        RECT 1414.105 2646.735 1414.435 2646.750 ;
      LAYER met3 ;
        RECT 300.065 2642.120 1396.000 2646.160 ;
        RECT 300.065 2640.720 1395.600 2642.120 ;
      LAYER met3 ;
        RECT 1396.000 2641.610 1400.000 2641.720 ;
        RECT 1411.345 2641.610 1411.675 2641.625 ;
        RECT 1396.000 2641.310 1411.675 2641.610 ;
        RECT 1396.000 2641.120 1400.000 2641.310 ;
        RECT 1411.345 2641.295 1411.675 2641.310 ;
      LAYER met3 ;
        RECT 300.065 2638.040 1396.000 2640.720 ;
      LAYER met3 ;
        RECT 300.000 2637.040 304.000 2637.640 ;
      LAYER met3 ;
        RECT 304.400 2637.360 1396.000 2638.040 ;
        RECT 304.400 2636.640 1395.600 2637.360 ;
        RECT 300.065 2635.960 1395.600 2636.640 ;
      LAYER met3 ;
        RECT 1396.000 2636.850 1400.000 2636.960 ;
        RECT 1414.105 2636.850 1414.435 2636.865 ;
        RECT 1396.000 2636.550 1414.435 2636.850 ;
        RECT 1396.000 2636.360 1400.000 2636.550 ;
        RECT 1414.105 2636.535 1414.435 2636.550 ;
      LAYER met3 ;
        RECT 300.065 2632.600 1396.000 2635.960 ;
        RECT 300.065 2631.200 1395.600 2632.600 ;
      LAYER met3 ;
        RECT 1396.000 2632.090 1400.000 2632.200 ;
        RECT 1409.505 2632.090 1409.835 2632.105 ;
        RECT 1396.000 2631.790 1409.835 2632.090 ;
        RECT 1396.000 2631.600 1400.000 2631.790 ;
        RECT 1409.505 2631.775 1409.835 2631.790 ;
      LAYER met3 ;
        RECT 300.065 2628.520 1396.000 2631.200 ;
      LAYER met3 ;
        RECT 300.000 2627.520 304.000 2628.120 ;
      LAYER met3 ;
        RECT 304.400 2627.160 1396.000 2628.520 ;
        RECT 304.400 2627.120 1395.600 2627.160 ;
        RECT 300.065 2625.760 1395.600 2627.120 ;
      LAYER met3 ;
        RECT 1396.000 2626.650 1400.000 2626.760 ;
        RECT 1414.105 2626.650 1414.435 2626.665 ;
        RECT 1396.000 2626.350 1414.435 2626.650 ;
        RECT 1396.000 2626.160 1400.000 2626.350 ;
        RECT 1414.105 2626.335 1414.435 2626.350 ;
      LAYER met3 ;
        RECT 300.065 2622.400 1396.000 2625.760 ;
        RECT 300.065 2621.000 1395.600 2622.400 ;
      LAYER met3 ;
        RECT 1396.000 2621.890 1400.000 2622.000 ;
        RECT 1411.805 2621.890 1412.135 2621.905 ;
        RECT 1396.000 2621.590 1412.135 2621.890 ;
        RECT 1396.000 2621.400 1400.000 2621.590 ;
        RECT 1411.805 2621.575 1412.135 2621.590 ;
      LAYER met3 ;
        RECT 300.065 2619.000 1396.000 2621.000 ;
      LAYER met3 ;
        RECT 300.000 2618.000 304.000 2618.600 ;
      LAYER met3 ;
        RECT 304.400 2617.600 1396.000 2619.000 ;
        RECT 300.065 2616.960 1396.000 2617.600 ;
        RECT 300.065 2615.560 1395.600 2616.960 ;
      LAYER met3 ;
        RECT 1396.000 2616.450 1400.000 2616.560 ;
        RECT 1414.105 2616.450 1414.435 2616.465 ;
        RECT 1396.000 2616.150 1414.435 2616.450 ;
        RECT 1396.000 2615.960 1400.000 2616.150 ;
        RECT 1414.105 2616.135 1414.435 2616.150 ;
      LAYER met3 ;
        RECT 300.065 2612.200 1396.000 2615.560 ;
        RECT 300.065 2610.800 1395.600 2612.200 ;
      LAYER met3 ;
        RECT 1396.000 2611.690 1400.000 2611.800 ;
        RECT 1414.105 2611.690 1414.435 2611.705 ;
        RECT 1396.000 2611.390 1414.435 2611.690 ;
        RECT 1396.000 2611.200 1400.000 2611.390 ;
        RECT 1414.105 2611.375 1414.435 2611.390 ;
      LAYER met3 ;
        RECT 300.065 2609.480 1396.000 2610.800 ;
      LAYER met3 ;
        RECT 300.000 2608.480 304.000 2609.080 ;
      LAYER met3 ;
        RECT 304.400 2608.080 1396.000 2609.480 ;
        RECT 300.065 2606.760 1396.000 2608.080 ;
        RECT 300.065 2605.360 1395.600 2606.760 ;
      LAYER met3 ;
        RECT 1396.000 2606.250 1400.000 2606.360 ;
        RECT 1417.785 2606.250 1418.115 2606.265 ;
        RECT 1396.000 2605.950 1418.115 2606.250 ;
        RECT 1396.000 2605.760 1400.000 2605.950 ;
        RECT 1417.785 2605.935 1418.115 2605.950 ;
      LAYER met3 ;
        RECT 300.065 2602.000 1396.000 2605.360 ;
        RECT 300.065 2600.600 1395.600 2602.000 ;
      LAYER met3 ;
        RECT 1396.000 2601.490 1400.000 2601.600 ;
        RECT 1414.105 2601.490 1414.435 2601.505 ;
        RECT 1396.000 2601.190 1414.435 2601.490 ;
        RECT 1396.000 2601.000 1400.000 2601.190 ;
        RECT 1414.105 2601.175 1414.435 2601.190 ;
      LAYER met3 ;
        RECT 300.065 2599.280 1396.000 2600.600 ;
      LAYER met3 ;
        RECT 300.000 2598.280 304.000 2598.880 ;
      LAYER met3 ;
        RECT 304.400 2597.880 1396.000 2599.280 ;
        RECT 300.065 2597.240 1396.000 2597.880 ;
        RECT 300.065 2595.840 1395.600 2597.240 ;
      LAYER met3 ;
        RECT 1396.000 2596.730 1400.000 2596.840 ;
        RECT 1408.585 2596.730 1408.915 2596.745 ;
        RECT 1396.000 2596.430 1408.915 2596.730 ;
        RECT 1396.000 2596.240 1400.000 2596.430 ;
        RECT 1408.585 2596.415 1408.915 2596.430 ;
      LAYER met3 ;
        RECT 300.065 2591.800 1396.000 2595.840 ;
        RECT 300.065 2590.400 1395.600 2591.800 ;
      LAYER met3 ;
        RECT 1396.000 2591.290 1400.000 2591.400 ;
        RECT 1410.425 2591.290 1410.755 2591.305 ;
        RECT 1396.000 2590.990 1410.755 2591.290 ;
        RECT 1396.000 2590.800 1400.000 2590.990 ;
        RECT 1410.425 2590.975 1410.755 2590.990 ;
      LAYER met3 ;
        RECT 300.065 2589.760 1396.000 2590.400 ;
      LAYER met3 ;
        RECT 300.000 2588.760 304.000 2589.360 ;
      LAYER met3 ;
        RECT 304.400 2588.360 1396.000 2589.760 ;
        RECT 300.065 2587.040 1396.000 2588.360 ;
        RECT 300.065 2585.640 1395.600 2587.040 ;
      LAYER met3 ;
        RECT 1396.000 2586.530 1400.000 2586.640 ;
        RECT 1411.345 2586.530 1411.675 2586.545 ;
        RECT 1396.000 2586.230 1411.675 2586.530 ;
        RECT 1396.000 2586.040 1400.000 2586.230 ;
        RECT 1411.345 2586.215 1411.675 2586.230 ;
      LAYER met3 ;
        RECT 300.065 2581.600 1396.000 2585.640 ;
        RECT 300.065 2580.240 1395.600 2581.600 ;
      LAYER met3 ;
        RECT 1396.000 2581.090 1400.000 2581.200 ;
        RECT 1414.105 2581.090 1414.435 2581.105 ;
        RECT 1396.000 2580.790 1414.435 2581.090 ;
        RECT 1396.000 2580.600 1400.000 2580.790 ;
        RECT 1414.105 2580.775 1414.435 2580.790 ;
      LAYER met3 ;
        RECT 304.400 2580.200 1395.600 2580.240 ;
      LAYER met3 ;
        RECT 300.000 2579.240 304.000 2579.840 ;
      LAYER met3 ;
        RECT 304.400 2578.840 1396.000 2580.200 ;
        RECT 300.065 2576.840 1396.000 2578.840 ;
        RECT 300.065 2575.440 1395.600 2576.840 ;
      LAYER met3 ;
        RECT 1396.000 2576.330 1400.000 2576.440 ;
        RECT 1414.105 2576.330 1414.435 2576.345 ;
        RECT 1396.000 2576.030 1414.435 2576.330 ;
        RECT 1396.000 2575.840 1400.000 2576.030 ;
        RECT 1414.105 2576.015 1414.435 2576.030 ;
      LAYER met3 ;
        RECT 300.065 2572.080 1396.000 2575.440 ;
        RECT 300.065 2570.720 1395.600 2572.080 ;
      LAYER met3 ;
        RECT 1396.000 2571.570 1400.000 2571.680 ;
        RECT 1411.345 2571.570 1411.675 2571.585 ;
        RECT 1396.000 2571.270 1411.675 2571.570 ;
        RECT 1396.000 2571.080 1400.000 2571.270 ;
        RECT 1411.345 2571.255 1411.675 2571.270 ;
      LAYER met3 ;
        RECT 304.400 2570.680 1395.600 2570.720 ;
      LAYER met3 ;
        RECT 300.000 2569.720 304.000 2570.320 ;
      LAYER met3 ;
        RECT 304.400 2569.320 1396.000 2570.680 ;
        RECT 300.065 2566.640 1396.000 2569.320 ;
        RECT 300.065 2565.240 1395.600 2566.640 ;
      LAYER met3 ;
        RECT 1396.000 2566.130 1400.000 2566.240 ;
        RECT 1413.645 2566.130 1413.975 2566.145 ;
        RECT 1396.000 2565.830 1413.975 2566.130 ;
        RECT 1396.000 2565.640 1400.000 2565.830 ;
        RECT 1413.645 2565.815 1413.975 2565.830 ;
      LAYER met3 ;
        RECT 300.065 2561.880 1396.000 2565.240 ;
        RECT 300.065 2561.200 1395.600 2561.880 ;
      LAYER met3 ;
        RECT 300.000 2560.200 304.000 2560.800 ;
      LAYER met3 ;
        RECT 304.400 2560.480 1395.600 2561.200 ;
      LAYER met3 ;
        RECT 1396.000 2561.370 1400.000 2561.480 ;
        RECT 1414.105 2561.370 1414.435 2561.385 ;
        RECT 1396.000 2561.070 1414.435 2561.370 ;
        RECT 1396.000 2560.880 1400.000 2561.070 ;
        RECT 1414.105 2561.055 1414.435 2561.070 ;
      LAYER met3 ;
        RECT 304.400 2559.800 1396.000 2560.480 ;
        RECT 300.065 2556.440 1396.000 2559.800 ;
        RECT 300.065 2555.040 1395.600 2556.440 ;
      LAYER met3 ;
        RECT 1396.000 2555.930 1400.000 2556.040 ;
        RECT 1408.585 2555.930 1408.915 2555.945 ;
        RECT 1396.000 2555.630 1408.915 2555.930 ;
        RECT 1396.000 2555.440 1400.000 2555.630 ;
        RECT 1408.585 2555.615 1408.915 2555.630 ;
      LAYER met3 ;
        RECT 300.065 2551.680 1396.000 2555.040 ;
        RECT 300.065 2551.000 1395.600 2551.680 ;
      LAYER met3 ;
        RECT 300.000 2550.000 304.000 2550.600 ;
      LAYER met3 ;
        RECT 304.400 2550.280 1395.600 2551.000 ;
      LAYER met3 ;
        RECT 1396.000 2551.170 1400.000 2551.280 ;
        RECT 1411.345 2551.170 1411.675 2551.185 ;
        RECT 1396.000 2550.870 1411.675 2551.170 ;
        RECT 1396.000 2550.680 1400.000 2550.870 ;
        RECT 1411.345 2550.855 1411.675 2550.870 ;
      LAYER met3 ;
        RECT 304.400 2549.600 1396.000 2550.280 ;
        RECT 300.065 2546.240 1396.000 2549.600 ;
        RECT 300.065 2544.840 1395.600 2546.240 ;
      LAYER met3 ;
        RECT 1396.000 2545.730 1400.000 2545.840 ;
        RECT 1412.725 2545.730 1413.055 2545.745 ;
        RECT 1396.000 2545.430 1413.055 2545.730 ;
        RECT 1396.000 2545.240 1400.000 2545.430 ;
        RECT 1412.725 2545.415 1413.055 2545.430 ;
      LAYER met3 ;
        RECT 300.065 2541.480 1396.000 2544.840 ;
      LAYER met3 ;
        RECT 300.000 2540.480 304.000 2541.080 ;
      LAYER met3 ;
        RECT 304.400 2540.080 1395.600 2541.480 ;
      LAYER met3 ;
        RECT 1396.000 2540.970 1400.000 2541.080 ;
        RECT 1414.105 2540.970 1414.435 2540.985 ;
        RECT 1396.000 2540.670 1414.435 2540.970 ;
        RECT 1396.000 2540.480 1400.000 2540.670 ;
        RECT 1414.105 2540.655 1414.435 2540.670 ;
      LAYER met3 ;
        RECT 300.065 2536.720 1396.000 2540.080 ;
        RECT 300.065 2535.320 1395.600 2536.720 ;
      LAYER met3 ;
        RECT 1396.000 2536.210 1400.000 2536.320 ;
        RECT 1410.425 2536.210 1410.755 2536.225 ;
        RECT 1396.000 2535.910 1410.755 2536.210 ;
        RECT 1396.000 2535.720 1400.000 2535.910 ;
        RECT 1410.425 2535.895 1410.755 2535.910 ;
      LAYER met3 ;
        RECT 300.065 2531.960 1396.000 2535.320 ;
      LAYER met3 ;
        RECT 300.000 2530.960 304.000 2531.560 ;
      LAYER met3 ;
        RECT 304.400 2531.280 1396.000 2531.960 ;
        RECT 304.400 2530.560 1395.600 2531.280 ;
        RECT 300.065 2529.880 1395.600 2530.560 ;
      LAYER met3 ;
        RECT 1396.000 2530.770 1400.000 2530.880 ;
        RECT 1413.645 2530.770 1413.975 2530.785 ;
        RECT 1396.000 2530.470 1413.975 2530.770 ;
        RECT 1396.000 2530.280 1400.000 2530.470 ;
        RECT 1413.645 2530.455 1413.975 2530.470 ;
      LAYER met3 ;
        RECT 300.065 2526.520 1396.000 2529.880 ;
        RECT 300.065 2525.120 1395.600 2526.520 ;
      LAYER met3 ;
        RECT 1396.000 2526.010 1400.000 2526.120 ;
        RECT 1414.105 2526.010 1414.435 2526.025 ;
        RECT 1396.000 2525.710 1414.435 2526.010 ;
        RECT 1396.000 2525.520 1400.000 2525.710 ;
        RECT 1414.105 2525.695 1414.435 2525.710 ;
      LAYER met3 ;
        RECT 300.065 2522.440 1396.000 2525.120 ;
      LAYER met3 ;
        RECT 300.000 2521.440 304.000 2522.040 ;
      LAYER met3 ;
        RECT 304.400 2521.080 1396.000 2522.440 ;
        RECT 304.400 2521.040 1395.600 2521.080 ;
        RECT 300.065 2519.680 1395.600 2521.040 ;
      LAYER met3 ;
        RECT 1396.000 2520.570 1400.000 2520.680 ;
        RECT 1414.105 2520.570 1414.435 2520.585 ;
        RECT 1396.000 2520.270 1414.435 2520.570 ;
        RECT 1396.000 2520.080 1400.000 2520.270 ;
        RECT 1414.105 2520.255 1414.435 2520.270 ;
      LAYER met3 ;
        RECT 300.065 2516.320 1396.000 2519.680 ;
        RECT 300.065 2514.920 1395.600 2516.320 ;
      LAYER met3 ;
        RECT 1396.000 2515.810 1400.000 2515.920 ;
        RECT 1414.105 2515.810 1414.435 2515.825 ;
        RECT 1396.000 2515.510 1414.435 2515.810 ;
        RECT 1396.000 2515.320 1400.000 2515.510 ;
        RECT 1414.105 2515.495 1414.435 2515.510 ;
      LAYER met3 ;
        RECT 300.065 2512.920 1396.000 2514.920 ;
      LAYER met3 ;
        RECT 300.000 2511.920 304.000 2512.520 ;
      LAYER met3 ;
        RECT 304.400 2511.520 1396.000 2512.920 ;
        RECT 300.065 2510.880 1396.000 2511.520 ;
        RECT 300.065 2509.480 1395.600 2510.880 ;
      LAYER met3 ;
        RECT 1396.000 2510.370 1400.000 2510.480 ;
        RECT 1411.345 2510.370 1411.675 2510.385 ;
        RECT 1396.000 2510.070 1411.675 2510.370 ;
        RECT 1396.000 2509.880 1400.000 2510.070 ;
        RECT 1411.345 2510.055 1411.675 2510.070 ;
      LAYER met3 ;
        RECT 300.065 2506.120 1396.000 2509.480 ;
        RECT 300.065 2504.720 1395.600 2506.120 ;
      LAYER met3 ;
        RECT 1396.000 2505.610 1400.000 2505.720 ;
        RECT 1414.105 2505.610 1414.435 2505.625 ;
        RECT 1396.000 2505.310 1414.435 2505.610 ;
        RECT 1396.000 2505.120 1400.000 2505.310 ;
        RECT 1414.105 2505.295 1414.435 2505.310 ;
      LAYER met3 ;
        RECT 300.065 2502.720 1396.000 2504.720 ;
      LAYER met3 ;
        RECT 300.000 2501.720 304.000 2502.320 ;
      LAYER met3 ;
        RECT 304.400 2501.360 1396.000 2502.720 ;
        RECT 304.400 2501.320 1395.600 2501.360 ;
        RECT 300.065 2499.960 1395.600 2501.320 ;
      LAYER met3 ;
        RECT 1396.000 2500.360 1400.000 2500.960 ;
      LAYER met3 ;
        RECT 300.065 2495.920 1396.000 2499.960 ;
        RECT 300.065 2494.520 1395.600 2495.920 ;
      LAYER met3 ;
        RECT 1396.000 2495.410 1400.000 2495.520 ;
        RECT 1414.105 2495.410 1414.435 2495.425 ;
        RECT 1396.000 2495.110 1414.435 2495.410 ;
        RECT 1396.000 2494.920 1400.000 2495.110 ;
        RECT 1414.105 2495.095 1414.435 2495.110 ;
      LAYER met3 ;
        RECT 300.065 2493.200 1396.000 2494.520 ;
      LAYER met3 ;
        RECT 300.000 2492.200 304.000 2492.800 ;
      LAYER met3 ;
        RECT 304.400 2491.800 1396.000 2493.200 ;
        RECT 300.065 2491.160 1396.000 2491.800 ;
        RECT 300.065 2489.760 1395.600 2491.160 ;
      LAYER met3 ;
        RECT 1396.000 2490.160 1400.000 2490.760 ;
      LAYER met3 ;
        RECT 300.065 2485.720 1396.000 2489.760 ;
        RECT 300.065 2484.320 1395.600 2485.720 ;
      LAYER met3 ;
        RECT 1396.000 2485.210 1400.000 2485.320 ;
        RECT 1414.105 2485.210 1414.435 2485.225 ;
        RECT 1396.000 2484.910 1414.435 2485.210 ;
        RECT 1396.000 2484.720 1400.000 2484.910 ;
        RECT 1414.105 2484.895 1414.435 2484.910 ;
      LAYER met3 ;
        RECT 300.065 2483.680 1396.000 2484.320 ;
      LAYER met3 ;
        RECT 300.000 2482.680 304.000 2483.280 ;
      LAYER met3 ;
        RECT 304.400 2482.280 1396.000 2483.680 ;
        RECT 300.065 2480.960 1396.000 2482.280 ;
        RECT 300.065 2479.560 1395.600 2480.960 ;
      LAYER met3 ;
        RECT 1396.000 2480.450 1400.000 2480.560 ;
        RECT 1409.505 2480.450 1409.835 2480.465 ;
        RECT 1396.000 2480.150 1409.835 2480.450 ;
        RECT 1396.000 2479.960 1400.000 2480.150 ;
        RECT 1409.505 2480.135 1409.835 2480.150 ;
      LAYER met3 ;
        RECT 300.065 2476.200 1396.000 2479.560 ;
        RECT 300.065 2474.800 1395.600 2476.200 ;
      LAYER met3 ;
        RECT 1396.000 2475.690 1400.000 2475.800 ;
        RECT 1414.105 2475.690 1414.435 2475.705 ;
        RECT 1396.000 2475.390 1414.435 2475.690 ;
        RECT 1396.000 2475.200 1400.000 2475.390 ;
        RECT 1414.105 2475.375 1414.435 2475.390 ;
      LAYER met3 ;
        RECT 300.065 2474.160 1396.000 2474.800 ;
      LAYER met3 ;
        RECT 300.000 2473.160 304.000 2473.760 ;
      LAYER met3 ;
        RECT 304.400 2472.760 1396.000 2474.160 ;
        RECT 300.065 2470.760 1396.000 2472.760 ;
        RECT 300.065 2469.360 1395.600 2470.760 ;
      LAYER met3 ;
        RECT 1396.000 2470.250 1400.000 2470.360 ;
        RECT 1411.805 2470.250 1412.135 2470.265 ;
        RECT 1396.000 2469.950 1412.135 2470.250 ;
        RECT 1396.000 2469.760 1400.000 2469.950 ;
        RECT 1411.805 2469.935 1412.135 2469.950 ;
      LAYER met3 ;
        RECT 300.065 2466.000 1396.000 2469.360 ;
        RECT 300.065 2464.640 1395.600 2466.000 ;
      LAYER met3 ;
        RECT 1396.000 2465.490 1400.000 2465.600 ;
        RECT 1414.105 2465.490 1414.435 2465.505 ;
        RECT 1396.000 2465.190 1414.435 2465.490 ;
        RECT 1396.000 2465.000 1400.000 2465.190 ;
        RECT 1414.105 2465.175 1414.435 2465.190 ;
      LAYER met3 ;
        RECT 304.400 2464.600 1395.600 2464.640 ;
      LAYER met3 ;
        RECT 300.000 2463.640 304.000 2464.240 ;
      LAYER met3 ;
        RECT 304.400 2463.240 1396.000 2464.600 ;
        RECT 300.065 2460.560 1396.000 2463.240 ;
        RECT 300.065 2459.160 1395.600 2460.560 ;
      LAYER met3 ;
        RECT 1396.000 2460.050 1400.000 2460.160 ;
        RECT 1414.105 2460.050 1414.435 2460.065 ;
        RECT 1396.000 2459.750 1414.435 2460.050 ;
        RECT 1396.000 2459.560 1400.000 2459.750 ;
        RECT 1414.105 2459.735 1414.435 2459.750 ;
      LAYER met3 ;
        RECT 300.065 2455.800 1396.000 2459.160 ;
        RECT 300.065 2454.440 1395.600 2455.800 ;
      LAYER met3 ;
        RECT 1396.000 2455.290 1400.000 2455.400 ;
        RECT 1411.345 2455.290 1411.675 2455.305 ;
        RECT 1396.000 2454.990 1411.675 2455.290 ;
        RECT 1396.000 2454.800 1400.000 2454.990 ;
        RECT 1411.345 2454.975 1411.675 2454.990 ;
      LAYER met3 ;
        RECT 304.400 2454.400 1395.600 2454.440 ;
      LAYER met3 ;
        RECT 300.000 2453.440 304.000 2454.040 ;
      LAYER met3 ;
        RECT 304.400 2453.040 1396.000 2454.400 ;
        RECT 300.065 2450.360 1396.000 2453.040 ;
        RECT 300.065 2448.960 1395.600 2450.360 ;
      LAYER met3 ;
        RECT 1396.000 2449.850 1400.000 2449.960 ;
        RECT 1414.105 2449.850 1414.435 2449.865 ;
        RECT 1396.000 2449.550 1414.435 2449.850 ;
        RECT 1396.000 2449.360 1400.000 2449.550 ;
        RECT 1414.105 2449.535 1414.435 2449.550 ;
      LAYER met3 ;
        RECT 300.065 2445.600 1396.000 2448.960 ;
        RECT 300.065 2444.920 1395.600 2445.600 ;
      LAYER met3 ;
        RECT 300.000 2443.920 304.000 2444.520 ;
      LAYER met3 ;
        RECT 304.400 2444.200 1395.600 2444.920 ;
      LAYER met3 ;
        RECT 1396.000 2445.090 1400.000 2445.200 ;
        RECT 1411.345 2445.090 1411.675 2445.105 ;
        RECT 1396.000 2444.790 1411.675 2445.090 ;
        RECT 1396.000 2444.600 1400.000 2444.790 ;
        RECT 1411.345 2444.775 1411.675 2444.790 ;
      LAYER met3 ;
        RECT 304.400 2443.520 1396.000 2444.200 ;
        RECT 300.065 2440.840 1396.000 2443.520 ;
        RECT 300.065 2439.440 1395.600 2440.840 ;
      LAYER met3 ;
        RECT 1396.000 2440.330 1400.000 2440.440 ;
        RECT 1414.105 2440.330 1414.435 2440.345 ;
        RECT 1396.000 2440.030 1414.435 2440.330 ;
        RECT 1396.000 2439.840 1400.000 2440.030 ;
        RECT 1414.105 2440.015 1414.435 2440.030 ;
      LAYER met3 ;
        RECT 300.065 2435.400 1396.000 2439.440 ;
      LAYER met3 ;
        RECT 300.000 2434.400 304.000 2435.000 ;
      LAYER met3 ;
        RECT 304.400 2434.000 1395.600 2435.400 ;
      LAYER met3 ;
        RECT 1396.000 2434.890 1400.000 2435.000 ;
        RECT 1411.345 2434.890 1411.675 2434.905 ;
        RECT 1396.000 2434.590 1411.675 2434.890 ;
        RECT 1396.000 2434.400 1400.000 2434.590 ;
        RECT 1411.345 2434.575 1411.675 2434.590 ;
      LAYER met3 ;
        RECT 300.065 2430.640 1396.000 2434.000 ;
        RECT 300.065 2429.240 1395.600 2430.640 ;
      LAYER met3 ;
        RECT 1396.000 2430.130 1400.000 2430.240 ;
        RECT 1414.105 2430.130 1414.435 2430.145 ;
        RECT 1396.000 2429.830 1414.435 2430.130 ;
        RECT 1396.000 2429.640 1400.000 2429.830 ;
        RECT 1414.105 2429.815 1414.435 2429.830 ;
      LAYER met3 ;
        RECT 300.065 2425.880 1396.000 2429.240 ;
      LAYER met3 ;
        RECT 300.000 2424.880 304.000 2425.480 ;
      LAYER met3 ;
        RECT 304.400 2425.200 1396.000 2425.880 ;
        RECT 304.400 2424.480 1395.600 2425.200 ;
        RECT 300.065 2423.800 1395.600 2424.480 ;
      LAYER met3 ;
        RECT 1396.000 2424.690 1400.000 2424.800 ;
        RECT 1408.585 2424.690 1408.915 2424.705 ;
        RECT 1396.000 2424.390 1408.915 2424.690 ;
        RECT 1396.000 2424.200 1400.000 2424.390 ;
        RECT 1408.585 2424.375 1408.915 2424.390 ;
      LAYER met3 ;
        RECT 300.065 2420.440 1396.000 2423.800 ;
        RECT 300.065 2419.040 1395.600 2420.440 ;
      LAYER met3 ;
        RECT 1396.000 2419.930 1400.000 2420.040 ;
        RECT 1411.345 2419.930 1411.675 2419.945 ;
        RECT 1396.000 2419.630 1411.675 2419.930 ;
        RECT 1396.000 2419.440 1400.000 2419.630 ;
        RECT 1411.345 2419.615 1411.675 2419.630 ;
      LAYER met3 ;
        RECT 300.065 2416.360 1396.000 2419.040 ;
      LAYER met3 ;
        RECT 300.000 2415.360 304.000 2415.960 ;
      LAYER met3 ;
        RECT 304.400 2415.000 1396.000 2416.360 ;
        RECT 304.400 2414.960 1395.600 2415.000 ;
        RECT 300.065 2413.600 1395.600 2414.960 ;
      LAYER met3 ;
        RECT 1396.000 2414.490 1400.000 2414.600 ;
        RECT 1412.725 2414.490 1413.055 2414.505 ;
        RECT 1396.000 2414.190 1413.055 2414.490 ;
        RECT 1396.000 2414.000 1400.000 2414.190 ;
        RECT 1412.725 2414.175 1413.055 2414.190 ;
      LAYER met3 ;
        RECT 300.065 2410.240 1396.000 2413.600 ;
        RECT 300.065 2408.840 1395.600 2410.240 ;
      LAYER met3 ;
        RECT 1396.000 2409.730 1400.000 2409.840 ;
        RECT 1414.105 2409.730 1414.435 2409.745 ;
        RECT 1396.000 2409.430 1414.435 2409.730 ;
        RECT 1396.000 2409.240 1400.000 2409.430 ;
        RECT 1414.105 2409.415 1414.435 2409.430 ;
      LAYER met3 ;
        RECT 300.065 2406.840 1396.000 2408.840 ;
      LAYER met3 ;
        RECT 300.000 2405.840 304.000 2406.440 ;
      LAYER met3 ;
        RECT 304.400 2405.480 1396.000 2406.840 ;
        RECT 304.400 2405.440 1395.600 2405.480 ;
        RECT 300.065 2404.080 1395.600 2405.440 ;
      LAYER met3 ;
        RECT 1396.000 2404.970 1400.000 2405.080 ;
        RECT 1410.425 2404.970 1410.755 2404.985 ;
        RECT 1396.000 2404.670 1410.755 2404.970 ;
        RECT 1396.000 2404.480 1400.000 2404.670 ;
        RECT 1410.425 2404.655 1410.755 2404.670 ;
      LAYER met3 ;
        RECT 300.065 2400.040 1396.000 2404.080 ;
        RECT 300.065 2398.640 1395.600 2400.040 ;
      LAYER met3 ;
        RECT 1396.000 2399.530 1400.000 2399.640 ;
        RECT 1413.645 2399.530 1413.975 2399.545 ;
        RECT 1396.000 2399.230 1413.975 2399.530 ;
        RECT 1396.000 2399.040 1400.000 2399.230 ;
        RECT 1413.645 2399.215 1413.975 2399.230 ;
      LAYER met3 ;
        RECT 300.065 2396.640 1396.000 2398.640 ;
      LAYER met3 ;
        RECT 300.000 2395.640 304.000 2396.240 ;
      LAYER met3 ;
        RECT 304.400 2395.280 1396.000 2396.640 ;
        RECT 304.400 2395.240 1395.600 2395.280 ;
        RECT 300.065 2393.880 1395.600 2395.240 ;
      LAYER met3 ;
        RECT 1396.000 2394.770 1400.000 2394.880 ;
        RECT 1414.105 2394.770 1414.435 2394.785 ;
        RECT 1396.000 2394.470 1414.435 2394.770 ;
        RECT 1396.000 2394.280 1400.000 2394.470 ;
        RECT 1414.105 2394.455 1414.435 2394.470 ;
      LAYER met3 ;
        RECT 300.065 2389.840 1396.000 2393.880 ;
        RECT 300.065 2388.440 1395.600 2389.840 ;
      LAYER met3 ;
        RECT 1396.000 2389.330 1400.000 2389.440 ;
        RECT 1414.105 2389.330 1414.435 2389.345 ;
        RECT 1396.000 2389.030 1414.435 2389.330 ;
        RECT 1396.000 2388.840 1400.000 2389.030 ;
        RECT 1414.105 2389.015 1414.435 2389.030 ;
      LAYER met3 ;
        RECT 300.065 2387.120 1396.000 2388.440 ;
      LAYER met3 ;
        RECT 300.000 2386.120 304.000 2386.720 ;
      LAYER met3 ;
        RECT 304.400 2385.720 1396.000 2387.120 ;
        RECT 300.065 2385.080 1396.000 2385.720 ;
        RECT 300.065 2383.680 1395.600 2385.080 ;
      LAYER met3 ;
        RECT 1396.000 2384.570 1400.000 2384.680 ;
        RECT 1410.425 2384.570 1410.755 2384.585 ;
        RECT 1396.000 2384.270 1410.755 2384.570 ;
        RECT 1396.000 2384.080 1400.000 2384.270 ;
        RECT 1410.425 2384.255 1410.755 2384.270 ;
      LAYER met3 ;
        RECT 300.065 2379.640 1396.000 2383.680 ;
        RECT 300.065 2378.240 1395.600 2379.640 ;
      LAYER met3 ;
        RECT 1396.000 2379.130 1400.000 2379.240 ;
        RECT 1411.345 2379.130 1411.675 2379.145 ;
        RECT 1396.000 2378.830 1411.675 2379.130 ;
        RECT 1396.000 2378.640 1400.000 2378.830 ;
        RECT 1411.345 2378.815 1411.675 2378.830 ;
      LAYER met3 ;
        RECT 300.065 2377.600 1396.000 2378.240 ;
      LAYER met3 ;
        RECT 300.000 2376.600 304.000 2377.200 ;
      LAYER met3 ;
        RECT 304.400 2376.200 1396.000 2377.600 ;
        RECT 300.065 2374.880 1396.000 2376.200 ;
        RECT 300.065 2373.480 1395.600 2374.880 ;
      LAYER met3 ;
        RECT 1396.000 2374.370 1400.000 2374.480 ;
        RECT 1414.105 2374.370 1414.435 2374.385 ;
        RECT 1396.000 2374.070 1414.435 2374.370 ;
        RECT 1396.000 2373.880 1400.000 2374.070 ;
        RECT 1414.105 2374.055 1414.435 2374.070 ;
      LAYER met3 ;
        RECT 300.065 2370.120 1396.000 2373.480 ;
        RECT 300.065 2368.720 1395.600 2370.120 ;
      LAYER met3 ;
        RECT 1396.000 2369.610 1400.000 2369.720 ;
        RECT 1408.585 2369.610 1408.915 2369.625 ;
        RECT 1396.000 2369.310 1408.915 2369.610 ;
        RECT 1396.000 2369.120 1400.000 2369.310 ;
        RECT 1408.585 2369.295 1408.915 2369.310 ;
      LAYER met3 ;
        RECT 300.065 2368.080 1396.000 2368.720 ;
      LAYER met3 ;
        RECT 300.000 2367.080 304.000 2367.680 ;
      LAYER met3 ;
        RECT 304.400 2366.680 1396.000 2368.080 ;
        RECT 300.065 2364.680 1396.000 2366.680 ;
        RECT 300.065 2363.280 1395.600 2364.680 ;
      LAYER met3 ;
        RECT 1396.000 2364.170 1400.000 2364.280 ;
        RECT 1410.425 2364.170 1410.755 2364.185 ;
        RECT 1396.000 2363.870 1410.755 2364.170 ;
        RECT 1396.000 2363.680 1400.000 2363.870 ;
        RECT 1410.425 2363.855 1410.755 2363.870 ;
      LAYER met3 ;
        RECT 300.065 2359.920 1396.000 2363.280 ;
        RECT 300.065 2358.560 1395.600 2359.920 ;
      LAYER met3 ;
        RECT 1396.000 2359.410 1400.000 2359.520 ;
        RECT 1413.645 2359.410 1413.975 2359.425 ;
        RECT 1396.000 2359.110 1413.975 2359.410 ;
        RECT 1396.000 2358.920 1400.000 2359.110 ;
        RECT 1413.645 2359.095 1413.975 2359.110 ;
      LAYER met3 ;
        RECT 304.400 2358.520 1395.600 2358.560 ;
      LAYER met3 ;
        RECT 300.000 2357.560 304.000 2358.160 ;
      LAYER met3 ;
        RECT 304.400 2357.160 1396.000 2358.520 ;
        RECT 300.065 2354.480 1396.000 2357.160 ;
        RECT 300.065 2353.080 1395.600 2354.480 ;
      LAYER met3 ;
        RECT 1396.000 2353.970 1400.000 2354.080 ;
        RECT 1414.105 2353.970 1414.435 2353.985 ;
        RECT 1396.000 2353.670 1414.435 2353.970 ;
        RECT 1396.000 2353.480 1400.000 2353.670 ;
        RECT 1414.105 2353.655 1414.435 2353.670 ;
      LAYER met3 ;
        RECT 300.065 2349.720 1396.000 2353.080 ;
        RECT 300.065 2348.360 1395.600 2349.720 ;
      LAYER met3 ;
        RECT 1396.000 2349.210 1400.000 2349.320 ;
        RECT 1409.505 2349.210 1409.835 2349.225 ;
        RECT 1396.000 2348.910 1409.835 2349.210 ;
        RECT 1396.000 2348.720 1400.000 2348.910 ;
        RECT 1409.505 2348.895 1409.835 2348.910 ;
      LAYER met3 ;
        RECT 304.400 2348.320 1395.600 2348.360 ;
      LAYER met3 ;
        RECT 300.000 2347.360 304.000 2347.960 ;
      LAYER met3 ;
        RECT 304.400 2346.960 1396.000 2348.320 ;
        RECT 300.065 2344.960 1396.000 2346.960 ;
        RECT 300.065 2343.560 1395.600 2344.960 ;
      LAYER met3 ;
        RECT 1396.000 2344.450 1400.000 2344.560 ;
        RECT 1414.105 2344.450 1414.435 2344.465 ;
        RECT 1396.000 2344.150 1414.435 2344.450 ;
        RECT 1396.000 2343.960 1400.000 2344.150 ;
        RECT 1414.105 2344.135 1414.435 2344.150 ;
      LAYER met3 ;
        RECT 300.065 2339.520 1396.000 2343.560 ;
        RECT 300.065 2338.840 1395.600 2339.520 ;
      LAYER met3 ;
        RECT 300.000 2337.840 304.000 2338.440 ;
      LAYER met3 ;
        RECT 304.400 2338.120 1395.600 2338.840 ;
      LAYER met3 ;
        RECT 1396.000 2339.010 1400.000 2339.120 ;
        RECT 1413.645 2339.010 1413.975 2339.025 ;
        RECT 1396.000 2338.710 1413.975 2339.010 ;
        RECT 1396.000 2338.520 1400.000 2338.710 ;
        RECT 1413.645 2338.695 1413.975 2338.710 ;
      LAYER met3 ;
        RECT 304.400 2337.440 1396.000 2338.120 ;
        RECT 300.065 2334.760 1396.000 2337.440 ;
        RECT 300.065 2333.360 1395.600 2334.760 ;
      LAYER met3 ;
        RECT 1396.000 2334.250 1400.000 2334.360 ;
        RECT 1414.105 2334.250 1414.435 2334.265 ;
        RECT 1396.000 2333.950 1414.435 2334.250 ;
        RECT 1396.000 2333.760 1400.000 2333.950 ;
        RECT 1414.105 2333.935 1414.435 2333.950 ;
      LAYER met3 ;
        RECT 300.065 2329.320 1396.000 2333.360 ;
      LAYER met3 ;
        RECT 300.000 2328.320 304.000 2328.920 ;
      LAYER met3 ;
        RECT 304.400 2327.920 1395.600 2329.320 ;
      LAYER met3 ;
        RECT 1396.000 2328.810 1400.000 2328.920 ;
        RECT 1414.105 2328.810 1414.435 2328.825 ;
        RECT 1396.000 2328.510 1414.435 2328.810 ;
        RECT 1396.000 2328.320 1400.000 2328.510 ;
        RECT 1414.105 2328.495 1414.435 2328.510 ;
      LAYER met3 ;
        RECT 300.065 2324.560 1396.000 2327.920 ;
        RECT 300.065 2323.160 1395.600 2324.560 ;
      LAYER met3 ;
        RECT 1396.000 2324.050 1400.000 2324.160 ;
        RECT 1413.645 2324.050 1413.975 2324.065 ;
        RECT 1396.000 2323.750 1413.975 2324.050 ;
        RECT 1396.000 2323.560 1400.000 2323.750 ;
        RECT 1413.645 2323.735 1413.975 2323.750 ;
      LAYER met3 ;
        RECT 300.065 2319.800 1396.000 2323.160 ;
      LAYER met3 ;
        RECT 300.000 2318.800 304.000 2319.400 ;
      LAYER met3 ;
        RECT 304.400 2319.120 1396.000 2319.800 ;
        RECT 304.400 2318.400 1395.600 2319.120 ;
        RECT 300.065 2317.720 1395.600 2318.400 ;
      LAYER met3 ;
        RECT 1396.000 2318.610 1400.000 2318.720 ;
        RECT 1414.105 2318.610 1414.435 2318.625 ;
        RECT 1396.000 2318.310 1414.435 2318.610 ;
        RECT 1396.000 2318.120 1400.000 2318.310 ;
        RECT 1414.105 2318.295 1414.435 2318.310 ;
      LAYER met3 ;
        RECT 300.065 2314.360 1396.000 2317.720 ;
        RECT 300.065 2312.960 1395.600 2314.360 ;
      LAYER met3 ;
        RECT 1396.000 2313.850 1400.000 2313.960 ;
        RECT 1414.105 2313.850 1414.435 2313.865 ;
        RECT 1396.000 2313.550 1414.435 2313.850 ;
        RECT 1396.000 2313.360 1400.000 2313.550 ;
        RECT 1414.105 2313.535 1414.435 2313.550 ;
      LAYER met3 ;
        RECT 300.065 2310.280 1396.000 2312.960 ;
      LAYER met3 ;
        RECT 300.000 2309.280 304.000 2309.880 ;
      LAYER met3 ;
        RECT 304.400 2309.600 1396.000 2310.280 ;
        RECT 304.400 2308.880 1395.600 2309.600 ;
        RECT 300.065 2308.200 1395.600 2308.880 ;
      LAYER met3 ;
        RECT 1396.000 2309.090 1400.000 2309.200 ;
        RECT 1414.105 2309.090 1414.435 2309.105 ;
        RECT 1396.000 2308.790 1414.435 2309.090 ;
        RECT 1396.000 2308.600 1400.000 2308.790 ;
        RECT 1414.105 2308.775 1414.435 2308.790 ;
      LAYER met3 ;
        RECT 300.065 2304.160 1396.000 2308.200 ;
        RECT 300.065 2302.760 1395.600 2304.160 ;
      LAYER met3 ;
        RECT 1396.000 2303.650 1400.000 2303.760 ;
        RECT 1414.105 2303.650 1414.435 2303.665 ;
        RECT 1396.000 2303.350 1414.435 2303.650 ;
        RECT 1396.000 2303.160 1400.000 2303.350 ;
        RECT 1414.105 2303.335 1414.435 2303.350 ;
      LAYER met3 ;
        RECT 300.065 2300.080 1396.000 2302.760 ;
      LAYER met3 ;
        RECT 300.000 2299.080 304.000 2299.680 ;
      LAYER met3 ;
        RECT 304.400 2299.400 1396.000 2300.080 ;
        RECT 304.400 2298.680 1395.600 2299.400 ;
        RECT 300.065 2298.000 1395.600 2298.680 ;
      LAYER met3 ;
        RECT 1396.000 2298.890 1400.000 2299.000 ;
        RECT 1413.645 2298.890 1413.975 2298.905 ;
        RECT 1396.000 2298.590 1413.975 2298.890 ;
        RECT 1396.000 2298.400 1400.000 2298.590 ;
        RECT 1413.645 2298.575 1413.975 2298.590 ;
      LAYER met3 ;
        RECT 300.065 2293.960 1396.000 2298.000 ;
        RECT 300.065 2292.560 1395.600 2293.960 ;
      LAYER met3 ;
        RECT 1396.000 2293.450 1400.000 2293.560 ;
        RECT 1408.585 2293.450 1408.915 2293.465 ;
        RECT 1396.000 2293.150 1408.915 2293.450 ;
        RECT 1396.000 2292.960 1400.000 2293.150 ;
        RECT 1408.585 2293.135 1408.915 2293.150 ;
      LAYER met3 ;
        RECT 300.065 2290.560 1396.000 2292.560 ;
      LAYER met3 ;
        RECT 300.000 2289.560 304.000 2290.160 ;
      LAYER met3 ;
        RECT 304.400 2289.200 1396.000 2290.560 ;
        RECT 304.400 2289.160 1395.600 2289.200 ;
        RECT 300.065 2287.800 1395.600 2289.160 ;
      LAYER met3 ;
        RECT 1396.000 2288.690 1400.000 2288.800 ;
        RECT 1410.425 2288.690 1410.755 2288.705 ;
        RECT 1396.000 2288.390 1410.755 2288.690 ;
        RECT 1396.000 2288.200 1400.000 2288.390 ;
        RECT 1410.425 2288.375 1410.755 2288.390 ;
      LAYER met3 ;
        RECT 300.065 2283.760 1396.000 2287.800 ;
        RECT 300.065 2282.360 1395.600 2283.760 ;
      LAYER met3 ;
        RECT 1396.000 2283.250 1400.000 2283.360 ;
        RECT 1408.125 2283.250 1408.455 2283.265 ;
        RECT 1396.000 2282.950 1408.455 2283.250 ;
        RECT 1396.000 2282.760 1400.000 2282.950 ;
        RECT 1408.125 2282.935 1408.455 2282.950 ;
      LAYER met3 ;
        RECT 300.065 2281.040 1396.000 2282.360 ;
      LAYER met3 ;
        RECT 300.000 2280.040 304.000 2280.640 ;
      LAYER met3 ;
        RECT 304.400 2279.640 1396.000 2281.040 ;
        RECT 300.065 2279.000 1396.000 2279.640 ;
        RECT 300.065 2277.600 1395.600 2279.000 ;
      LAYER met3 ;
        RECT 1396.000 2278.490 1400.000 2278.600 ;
        RECT 1414.105 2278.490 1414.435 2278.505 ;
        RECT 1396.000 2278.190 1414.435 2278.490 ;
        RECT 1396.000 2278.000 1400.000 2278.190 ;
        RECT 1414.105 2278.175 1414.435 2278.190 ;
      LAYER met3 ;
        RECT 300.065 2274.240 1396.000 2277.600 ;
        RECT 300.065 2272.840 1395.600 2274.240 ;
      LAYER met3 ;
        RECT 1396.000 2273.730 1400.000 2273.840 ;
        RECT 1408.125 2273.730 1408.455 2273.745 ;
        RECT 1396.000 2273.430 1408.455 2273.730 ;
        RECT 1396.000 2273.240 1400.000 2273.430 ;
        RECT 1408.125 2273.415 1408.455 2273.430 ;
      LAYER met3 ;
        RECT 300.065 2271.520 1396.000 2272.840 ;
      LAYER met3 ;
        RECT 300.000 2270.520 304.000 2271.120 ;
      LAYER met3 ;
        RECT 304.400 2270.120 1396.000 2271.520 ;
        RECT 300.065 2268.800 1396.000 2270.120 ;
        RECT 300.065 2267.400 1395.600 2268.800 ;
      LAYER met3 ;
        RECT 1396.000 2268.290 1400.000 2268.400 ;
        RECT 1412.265 2268.290 1412.595 2268.305 ;
        RECT 1396.000 2267.990 1412.595 2268.290 ;
        RECT 1396.000 2267.800 1400.000 2267.990 ;
        RECT 1412.265 2267.975 1412.595 2267.990 ;
      LAYER met3 ;
        RECT 300.065 2264.040 1396.000 2267.400 ;
        RECT 300.065 2262.640 1395.600 2264.040 ;
      LAYER met3 ;
        RECT 1396.000 2263.530 1400.000 2263.640 ;
        RECT 1411.345 2263.530 1411.675 2263.545 ;
        RECT 1396.000 2263.230 1411.675 2263.530 ;
        RECT 1396.000 2263.040 1400.000 2263.230 ;
        RECT 1411.345 2263.215 1411.675 2263.230 ;
      LAYER met3 ;
        RECT 300.065 2262.000 1396.000 2262.640 ;
      LAYER met3 ;
        RECT 300.000 2261.000 304.000 2261.600 ;
      LAYER met3 ;
        RECT 304.400 2260.600 1396.000 2262.000 ;
        RECT 300.065 2258.600 1396.000 2260.600 ;
        RECT 300.065 2257.200 1395.600 2258.600 ;
      LAYER met3 ;
        RECT 1396.000 2258.090 1400.000 2258.200 ;
        RECT 1411.805 2258.090 1412.135 2258.105 ;
        RECT 1396.000 2257.790 1412.135 2258.090 ;
        RECT 1396.000 2257.600 1400.000 2257.790 ;
        RECT 1411.805 2257.775 1412.135 2257.790 ;
      LAYER met3 ;
        RECT 300.065 2253.840 1396.000 2257.200 ;
        RECT 300.065 2252.440 1395.600 2253.840 ;
      LAYER met3 ;
        RECT 1396.000 2253.330 1400.000 2253.440 ;
        RECT 1412.725 2253.330 1413.055 2253.345 ;
        RECT 1396.000 2253.030 1413.055 2253.330 ;
        RECT 1396.000 2252.840 1400.000 2253.030 ;
        RECT 1412.725 2253.015 1413.055 2253.030 ;
      LAYER met3 ;
        RECT 300.065 2251.800 1396.000 2252.440 ;
      LAYER met3 ;
        RECT 300.000 2250.800 304.000 2251.400 ;
      LAYER met3 ;
        RECT 304.400 2250.400 1396.000 2251.800 ;
        RECT 300.065 2249.080 1396.000 2250.400 ;
        RECT 300.065 2247.680 1395.600 2249.080 ;
      LAYER met3 ;
        RECT 1396.000 2248.570 1400.000 2248.680 ;
        RECT 1414.105 2248.570 1414.435 2248.585 ;
        RECT 1396.000 2248.270 1414.435 2248.570 ;
        RECT 1396.000 2248.080 1400.000 2248.270 ;
        RECT 1414.105 2248.255 1414.435 2248.270 ;
      LAYER met3 ;
        RECT 300.065 2243.640 1396.000 2247.680 ;
        RECT 300.065 2242.280 1395.600 2243.640 ;
      LAYER met3 ;
        RECT 1396.000 2243.130 1400.000 2243.240 ;
        RECT 1413.185 2243.130 1413.515 2243.145 ;
        RECT 1396.000 2242.830 1413.515 2243.130 ;
        RECT 1396.000 2242.640 1400.000 2242.830 ;
        RECT 1413.185 2242.815 1413.515 2242.830 ;
      LAYER met3 ;
        RECT 304.400 2242.240 1395.600 2242.280 ;
      LAYER met3 ;
        RECT 300.000 2241.280 304.000 2241.880 ;
      LAYER met3 ;
        RECT 304.400 2240.880 1396.000 2242.240 ;
        RECT 300.065 2238.880 1396.000 2240.880 ;
        RECT 300.065 2237.480 1395.600 2238.880 ;
      LAYER met3 ;
        RECT 1396.000 2238.370 1400.000 2238.480 ;
        RECT 1413.645 2238.370 1413.975 2238.385 ;
        RECT 1396.000 2238.070 1413.975 2238.370 ;
        RECT 1396.000 2237.880 1400.000 2238.070 ;
        RECT 1413.645 2238.055 1413.975 2238.070 ;
      LAYER met3 ;
        RECT 300.065 2233.440 1396.000 2237.480 ;
        RECT 300.065 2232.760 1395.600 2233.440 ;
      LAYER met3 ;
        RECT 300.000 2231.760 304.000 2232.360 ;
      LAYER met3 ;
        RECT 304.400 2232.040 1395.600 2232.760 ;
      LAYER met3 ;
        RECT 1396.000 2232.930 1400.000 2233.040 ;
        RECT 1410.425 2232.930 1410.755 2232.945 ;
        RECT 1396.000 2232.630 1410.755 2232.930 ;
        RECT 1396.000 2232.440 1400.000 2232.630 ;
        RECT 1410.425 2232.615 1410.755 2232.630 ;
      LAYER met3 ;
        RECT 304.400 2231.360 1396.000 2232.040 ;
        RECT 300.065 2228.680 1396.000 2231.360 ;
        RECT 300.065 2227.280 1395.600 2228.680 ;
      LAYER met3 ;
        RECT 1396.000 2228.170 1400.000 2228.280 ;
        RECT 1409.045 2228.170 1409.375 2228.185 ;
        RECT 1396.000 2227.870 1409.375 2228.170 ;
        RECT 1396.000 2227.680 1400.000 2227.870 ;
        RECT 1409.045 2227.855 1409.375 2227.870 ;
      LAYER met3 ;
        RECT 300.065 2223.240 1396.000 2227.280 ;
      LAYER met3 ;
        RECT 300.000 2222.240 304.000 2222.840 ;
      LAYER met3 ;
        RECT 304.400 2221.840 1395.600 2223.240 ;
      LAYER met3 ;
        RECT 1396.000 2222.730 1400.000 2222.840 ;
        RECT 1409.965 2222.730 1410.295 2222.745 ;
        RECT 1396.000 2222.430 1410.295 2222.730 ;
        RECT 1396.000 2222.240 1400.000 2222.430 ;
        RECT 1409.965 2222.415 1410.295 2222.430 ;
      LAYER met3 ;
        RECT 300.065 2218.480 1396.000 2221.840 ;
        RECT 300.065 2217.080 1395.600 2218.480 ;
      LAYER met3 ;
        RECT 1396.000 2217.970 1400.000 2218.080 ;
        RECT 1409.505 2217.970 1409.835 2217.985 ;
        RECT 1396.000 2217.670 1409.835 2217.970 ;
        RECT 1396.000 2217.480 1400.000 2217.670 ;
        RECT 1409.505 2217.655 1409.835 2217.670 ;
      LAYER met3 ;
        RECT 300.065 2213.720 1396.000 2217.080 ;
      LAYER met3 ;
        RECT 300.000 2212.720 304.000 2213.320 ;
      LAYER met3 ;
        RECT 304.400 2212.320 1395.600 2213.720 ;
      LAYER met3 ;
        RECT 1396.000 2213.210 1400.000 2213.320 ;
        RECT 1408.585 2213.210 1408.915 2213.225 ;
        RECT 1396.000 2212.910 1408.915 2213.210 ;
        RECT 1396.000 2212.720 1400.000 2212.910 ;
        RECT 1408.585 2212.895 1408.915 2212.910 ;
      LAYER met3 ;
        RECT 300.065 2208.280 1396.000 2212.320 ;
        RECT 300.065 2206.880 1395.600 2208.280 ;
      LAYER met3 ;
        RECT 1396.000 2207.280 1400.000 2207.880 ;
      LAYER met3 ;
        RECT 300.065 2203.520 1396.000 2206.880 ;
      LAYER met3 ;
        RECT 1399.630 2205.050 1399.930 2207.280 ;
        RECT 1407.205 2205.050 1407.535 2205.065 ;
        RECT 1399.630 2204.750 1407.535 2205.050 ;
        RECT 1407.205 2204.735 1407.535 2204.750 ;
        RECT 300.000 2202.520 304.000 2203.120 ;
      LAYER met3 ;
        RECT 304.400 2202.120 1395.600 2203.520 ;
      LAYER met3 ;
        RECT 1396.000 2203.010 1400.000 2203.120 ;
        RECT 1410.885 2203.010 1411.215 2203.025 ;
        RECT 1396.000 2202.710 1411.215 2203.010 ;
        RECT 1396.000 2202.520 1400.000 2202.710 ;
        RECT 1410.885 2202.695 1411.215 2202.710 ;
      LAYER met3 ;
        RECT 300.065 2198.080 1396.000 2202.120 ;
        RECT 300.065 2196.680 1395.600 2198.080 ;
      LAYER met3 ;
        RECT 1396.000 2197.570 1400.000 2197.680 ;
        RECT 1410.885 2197.570 1411.215 2197.585 ;
        RECT 1396.000 2197.270 1411.215 2197.570 ;
        RECT 1396.000 2197.080 1400.000 2197.270 ;
        RECT 1410.885 2197.255 1411.215 2197.270 ;
      LAYER met3 ;
        RECT 300.065 2194.000 1396.000 2196.680 ;
      LAYER met3 ;
        RECT 300.000 2193.000 304.000 2193.600 ;
      LAYER met3 ;
        RECT 304.400 2193.320 1396.000 2194.000 ;
        RECT 304.400 2192.600 1395.600 2193.320 ;
        RECT 300.065 2191.920 1395.600 2192.600 ;
      LAYER met3 ;
        RECT 1396.000 2192.810 1400.000 2192.920 ;
        RECT 1417.325 2192.810 1417.655 2192.825 ;
        RECT 1396.000 2192.510 1417.655 2192.810 ;
        RECT 1396.000 2192.320 1400.000 2192.510 ;
        RECT 1417.325 2192.495 1417.655 2192.510 ;
      LAYER met3 ;
        RECT 300.065 2187.880 1396.000 2191.920 ;
        RECT 300.065 2186.480 1395.600 2187.880 ;
      LAYER met3 ;
        RECT 1396.000 2187.370 1400.000 2187.480 ;
        RECT 1410.885 2187.370 1411.215 2187.385 ;
        RECT 1396.000 2187.070 1411.215 2187.370 ;
        RECT 1396.000 2186.880 1400.000 2187.070 ;
        RECT 1410.885 2187.055 1411.215 2187.070 ;
      LAYER met3 ;
        RECT 300.065 2184.480 1396.000 2186.480 ;
      LAYER met3 ;
        RECT 300.000 2183.480 304.000 2184.080 ;
      LAYER met3 ;
        RECT 304.400 2183.120 1396.000 2184.480 ;
        RECT 304.400 2183.080 1395.600 2183.120 ;
        RECT 300.065 2181.720 1395.600 2183.080 ;
      LAYER met3 ;
        RECT 1396.000 2182.610 1400.000 2182.720 ;
        RECT 1410.885 2182.610 1411.215 2182.625 ;
        RECT 1396.000 2182.310 1411.215 2182.610 ;
        RECT 1396.000 2182.120 1400.000 2182.310 ;
        RECT 1410.885 2182.295 1411.215 2182.310 ;
      LAYER met3 ;
        RECT 300.065 2178.360 1396.000 2181.720 ;
        RECT 300.065 2176.960 1395.600 2178.360 ;
      LAYER met3 ;
        RECT 1396.000 2177.850 1400.000 2177.960 ;
        RECT 1410.885 2177.850 1411.215 2177.865 ;
        RECT 1396.000 2177.550 1411.215 2177.850 ;
        RECT 1396.000 2177.360 1400.000 2177.550 ;
        RECT 1410.885 2177.535 1411.215 2177.550 ;
      LAYER met3 ;
        RECT 300.065 2174.960 1396.000 2176.960 ;
      LAYER met3 ;
        RECT 300.000 2173.960 304.000 2174.560 ;
      LAYER met3 ;
        RECT 304.400 2173.560 1396.000 2174.960 ;
        RECT 300.065 2172.920 1396.000 2173.560 ;
        RECT 300.065 2171.520 1395.600 2172.920 ;
      LAYER met3 ;
        RECT 1396.000 2172.410 1400.000 2172.520 ;
        RECT 1410.885 2172.410 1411.215 2172.425 ;
        RECT 1396.000 2172.110 1411.215 2172.410 ;
        RECT 1396.000 2171.920 1400.000 2172.110 ;
        RECT 1410.885 2172.095 1411.215 2172.110 ;
      LAYER met3 ;
        RECT 300.065 2168.160 1396.000 2171.520 ;
        RECT 300.065 2166.760 1395.600 2168.160 ;
      LAYER met3 ;
        RECT 1396.000 2167.650 1400.000 2167.760 ;
        RECT 1416.865 2167.650 1417.195 2167.665 ;
        RECT 1396.000 2167.350 1417.195 2167.650 ;
        RECT 1396.000 2167.160 1400.000 2167.350 ;
        RECT 1416.865 2167.335 1417.195 2167.350 ;
      LAYER met3 ;
        RECT 300.065 2165.440 1396.000 2166.760 ;
      LAYER met3 ;
        RECT 300.000 2164.440 304.000 2165.040 ;
      LAYER met3 ;
        RECT 304.400 2164.040 1396.000 2165.440 ;
        RECT 300.065 2162.720 1396.000 2164.040 ;
        RECT 300.065 2161.320 1395.600 2162.720 ;
      LAYER met3 ;
        RECT 1396.000 2162.210 1400.000 2162.320 ;
        RECT 1410.885 2162.210 1411.215 2162.225 ;
        RECT 1396.000 2161.910 1411.215 2162.210 ;
        RECT 1396.000 2161.720 1400.000 2161.910 ;
        RECT 1410.885 2161.895 1411.215 2161.910 ;
      LAYER met3 ;
        RECT 300.065 2157.960 1396.000 2161.320 ;
        RECT 300.065 2156.560 1395.600 2157.960 ;
      LAYER met3 ;
        RECT 1396.000 2157.450 1400.000 2157.560 ;
        RECT 1411.345 2157.450 1411.675 2157.465 ;
        RECT 1396.000 2157.150 1411.675 2157.450 ;
        RECT 1396.000 2156.960 1400.000 2157.150 ;
        RECT 1411.345 2157.135 1411.675 2157.150 ;
      LAYER met3 ;
        RECT 300.065 2155.920 1396.000 2156.560 ;
      LAYER met3 ;
        RECT 300.000 2154.920 304.000 2155.520 ;
      LAYER met3 ;
        RECT 304.400 2154.520 1396.000 2155.920 ;
        RECT 300.065 2153.200 1396.000 2154.520 ;
        RECT 300.065 2151.800 1395.600 2153.200 ;
      LAYER met3 ;
        RECT 1396.000 2152.200 1400.000 2152.800 ;
      LAYER met3 ;
        RECT 300.065 2147.760 1396.000 2151.800 ;
      LAYER met3 ;
        RECT 1399.630 2149.970 1399.930 2152.200 ;
        RECT 1407.205 2149.970 1407.535 2149.985 ;
        RECT 1399.630 2149.670 1407.535 2149.970 ;
        RECT 1407.205 2149.655 1407.535 2149.670 ;
      LAYER met3 ;
        RECT 300.065 2146.360 1395.600 2147.760 ;
      LAYER met3 ;
        RECT 1396.000 2147.250 1400.000 2147.360 ;
        RECT 1411.345 2147.250 1411.675 2147.265 ;
        RECT 1396.000 2146.950 1411.675 2147.250 ;
        RECT 1396.000 2146.760 1400.000 2146.950 ;
        RECT 1411.345 2146.935 1411.675 2146.950 ;
      LAYER met3 ;
        RECT 300.065 2145.720 1396.000 2146.360 ;
      LAYER met3 ;
        RECT 300.000 2144.720 304.000 2145.320 ;
      LAYER met3 ;
        RECT 304.400 2144.320 1396.000 2145.720 ;
        RECT 300.065 2143.000 1396.000 2144.320 ;
        RECT 300.065 2141.600 1395.600 2143.000 ;
      LAYER met3 ;
        RECT 1396.000 2142.490 1400.000 2142.600 ;
        RECT 1411.345 2142.490 1411.675 2142.505 ;
        RECT 1396.000 2142.190 1411.675 2142.490 ;
        RECT 1396.000 2142.000 1400.000 2142.190 ;
        RECT 1411.345 2142.175 1411.675 2142.190 ;
      LAYER met3 ;
        RECT 300.065 2137.560 1396.000 2141.600 ;
        RECT 300.065 2136.200 1395.600 2137.560 ;
      LAYER met3 ;
        RECT 1396.000 2137.050 1400.000 2137.160 ;
        RECT 1411.345 2137.050 1411.675 2137.065 ;
        RECT 1396.000 2136.750 1411.675 2137.050 ;
        RECT 1396.000 2136.560 1400.000 2136.750 ;
        RECT 1411.345 2136.735 1411.675 2136.750 ;
      LAYER met3 ;
        RECT 304.400 2136.160 1395.600 2136.200 ;
      LAYER met3 ;
        RECT 300.000 2135.200 304.000 2135.800 ;
      LAYER met3 ;
        RECT 304.400 2134.800 1396.000 2136.160 ;
      LAYER met3 ;
        RECT 1411.345 2135.010 1411.675 2135.025 ;
      LAYER met3 ;
        RECT 300.065 2132.800 1396.000 2134.800 ;
      LAYER met3 ;
        RECT 1399.630 2134.710 1411.675 2135.010 ;
      LAYER met3 ;
        RECT 300.065 2131.400 1395.600 2132.800 ;
      LAYER met3 ;
        RECT 1399.630 2132.400 1399.930 2134.710 ;
        RECT 1411.345 2134.695 1411.675 2134.710 ;
        RECT 1396.000 2131.800 1400.000 2132.400 ;
      LAYER met3 ;
        RECT 300.065 2127.360 1396.000 2131.400 ;
        RECT 300.065 2126.680 1395.600 2127.360 ;
      LAYER met3 ;
        RECT 300.000 2125.680 304.000 2126.280 ;
      LAYER met3 ;
        RECT 304.400 2125.960 1395.600 2126.680 ;
      LAYER met3 ;
        RECT 1396.000 2126.850 1400.000 2126.960 ;
        RECT 1411.345 2126.850 1411.675 2126.865 ;
        RECT 1396.000 2126.550 1411.675 2126.850 ;
        RECT 1396.000 2126.360 1400.000 2126.550 ;
        RECT 1411.345 2126.535 1411.675 2126.550 ;
      LAYER met3 ;
        RECT 304.400 2125.280 1396.000 2125.960 ;
        RECT 300.065 2122.600 1396.000 2125.280 ;
        RECT 300.065 2121.200 1395.600 2122.600 ;
      LAYER met3 ;
        RECT 1396.000 2122.090 1400.000 2122.200 ;
        RECT 1411.345 2122.090 1411.675 2122.105 ;
        RECT 1396.000 2121.790 1411.675 2122.090 ;
        RECT 1396.000 2121.600 1400.000 2121.790 ;
        RECT 1411.345 2121.775 1411.675 2121.790 ;
      LAYER met3 ;
        RECT 300.065 2117.840 1396.000 2121.200 ;
        RECT 300.065 2117.160 1395.600 2117.840 ;
      LAYER met3 ;
        RECT 300.000 2116.160 304.000 2116.760 ;
      LAYER met3 ;
        RECT 304.400 2116.440 1395.600 2117.160 ;
      LAYER met3 ;
        RECT 1396.000 2117.330 1400.000 2117.440 ;
        RECT 1411.345 2117.330 1411.675 2117.345 ;
        RECT 1396.000 2117.030 1411.675 2117.330 ;
        RECT 1396.000 2116.840 1400.000 2117.030 ;
        RECT 1411.345 2117.015 1411.675 2117.030 ;
      LAYER met3 ;
        RECT 304.400 2115.760 1396.000 2116.440 ;
        RECT 300.065 2112.400 1396.000 2115.760 ;
        RECT 300.065 2111.000 1395.600 2112.400 ;
      LAYER met3 ;
        RECT 1396.000 2111.890 1400.000 2112.000 ;
        RECT 1411.345 2111.890 1411.675 2111.905 ;
        RECT 1396.000 2111.590 1411.675 2111.890 ;
        RECT 1396.000 2111.400 1400.000 2111.590 ;
        RECT 1411.345 2111.575 1411.675 2111.590 ;
      LAYER met3 ;
        RECT 300.065 2107.640 1396.000 2111.000 ;
      LAYER met3 ;
        RECT 300.000 2106.640 304.000 2107.240 ;
      LAYER met3 ;
        RECT 304.400 2106.240 1395.600 2107.640 ;
      LAYER met3 ;
        RECT 1396.000 2107.130 1400.000 2107.240 ;
        RECT 1411.345 2107.130 1411.675 2107.145 ;
        RECT 1396.000 2106.830 1411.675 2107.130 ;
        RECT 1396.000 2106.640 1400.000 2106.830 ;
        RECT 1411.345 2106.815 1411.675 2106.830 ;
      LAYER met3 ;
        RECT 300.065 2102.200 1396.000 2106.240 ;
        RECT 300.065 2100.800 1395.600 2102.200 ;
      LAYER met3 ;
        RECT 1396.000 2101.690 1400.000 2101.800 ;
        RECT 1414.105 2101.690 1414.435 2101.705 ;
        RECT 1396.000 2101.390 1414.435 2101.690 ;
        RECT 1396.000 2101.200 1400.000 2101.390 ;
        RECT 1414.105 2101.375 1414.435 2101.390 ;
      LAYER met3 ;
        RECT 300.065 2097.440 1396.000 2100.800 ;
      LAYER met3 ;
        RECT 300.000 2096.440 304.000 2097.040 ;
      LAYER met3 ;
        RECT 304.400 2096.040 1395.600 2097.440 ;
      LAYER met3 ;
        RECT 1396.000 2096.930 1400.000 2097.040 ;
        RECT 1414.105 2096.930 1414.435 2096.945 ;
        RECT 1396.000 2096.630 1414.435 2096.930 ;
        RECT 1396.000 2096.440 1400.000 2096.630 ;
        RECT 1414.105 2096.615 1414.435 2096.630 ;
      LAYER met3 ;
        RECT 300.065 2092.000 1396.000 2096.040 ;
        RECT 300.065 2090.600 1395.600 2092.000 ;
      LAYER met3 ;
        RECT 1396.000 2091.490 1400.000 2091.600 ;
        RECT 1412.725 2091.490 1413.055 2091.505 ;
        RECT 1396.000 2091.190 1413.055 2091.490 ;
        RECT 1396.000 2091.000 1400.000 2091.190 ;
        RECT 1412.725 2091.175 1413.055 2091.190 ;
      LAYER met3 ;
        RECT 300.065 2087.920 1396.000 2090.600 ;
      LAYER met3 ;
        RECT 300.000 2086.920 304.000 2087.520 ;
      LAYER met3 ;
        RECT 304.400 2087.240 1396.000 2087.920 ;
        RECT 304.400 2086.520 1395.600 2087.240 ;
        RECT 300.065 2085.840 1395.600 2086.520 ;
      LAYER met3 ;
        RECT 1396.000 2086.730 1400.000 2086.840 ;
        RECT 1414.105 2086.730 1414.435 2086.745 ;
        RECT 1396.000 2086.430 1414.435 2086.730 ;
        RECT 1396.000 2086.240 1400.000 2086.430 ;
        RECT 1414.105 2086.415 1414.435 2086.430 ;
      LAYER met3 ;
        RECT 300.065 2082.480 1396.000 2085.840 ;
        RECT 300.065 2081.080 1395.600 2082.480 ;
      LAYER met3 ;
        RECT 1396.000 2081.970 1400.000 2082.080 ;
        RECT 1414.105 2081.970 1414.435 2081.985 ;
        RECT 1396.000 2081.670 1414.435 2081.970 ;
        RECT 1396.000 2081.480 1400.000 2081.670 ;
        RECT 1414.105 2081.655 1414.435 2081.670 ;
      LAYER met3 ;
        RECT 300.065 2078.400 1396.000 2081.080 ;
      LAYER met3 ;
        RECT 300.000 2077.400 304.000 2078.000 ;
      LAYER met3 ;
        RECT 304.400 2077.040 1396.000 2078.400 ;
        RECT 304.400 2077.000 1395.600 2077.040 ;
        RECT 300.065 2075.640 1395.600 2077.000 ;
      LAYER met3 ;
        RECT 1396.000 2076.530 1400.000 2076.640 ;
        RECT 1414.105 2076.530 1414.435 2076.545 ;
        RECT 1396.000 2076.230 1414.435 2076.530 ;
        RECT 1396.000 2076.040 1400.000 2076.230 ;
        RECT 1414.105 2076.215 1414.435 2076.230 ;
      LAYER met3 ;
        RECT 300.065 2072.280 1396.000 2075.640 ;
        RECT 300.065 2070.880 1395.600 2072.280 ;
      LAYER met3 ;
        RECT 1396.000 2071.770 1400.000 2071.880 ;
        RECT 1411.345 2071.770 1411.675 2071.785 ;
        RECT 1396.000 2071.470 1411.675 2071.770 ;
        RECT 1396.000 2071.280 1400.000 2071.470 ;
        RECT 1411.345 2071.455 1411.675 2071.470 ;
      LAYER met3 ;
        RECT 300.065 2068.880 1396.000 2070.880 ;
      LAYER met3 ;
        RECT 1859.385 2070.410 1859.715 2070.425 ;
        RECT 1859.385 2070.110 1866.370 2070.410 ;
        RECT 1859.385 2070.095 1859.715 2070.110 ;
        RECT 1835.465 2069.730 1835.795 2069.745 ;
        RECT 1841.190 2069.730 1841.570 2069.740 ;
        RECT 1835.465 2069.430 1841.570 2069.730 ;
        RECT 1835.465 2069.415 1835.795 2069.430 ;
        RECT 1841.190 2069.420 1841.570 2069.430 ;
        RECT 1842.825 2069.730 1843.155 2069.745 ;
        RECT 1844.870 2069.730 1845.250 2069.740 ;
        RECT 1842.825 2069.430 1845.250 2069.730 ;
        RECT 1842.825 2069.415 1843.155 2069.430 ;
        RECT 1844.870 2069.420 1845.250 2069.430 ;
        RECT 1849.725 2069.730 1850.055 2069.745 ;
        RECT 1851.310 2069.730 1851.690 2069.740 ;
        RECT 1849.725 2069.430 1851.690 2069.730 ;
        RECT 1849.725 2069.415 1850.055 2069.430 ;
        RECT 1851.310 2069.420 1851.690 2069.430 ;
        RECT 1856.165 2069.730 1856.495 2069.745 ;
        RECT 1859.590 2069.730 1859.970 2069.740 ;
        RECT 1856.165 2069.430 1859.970 2069.730 ;
        RECT 1856.165 2069.415 1856.495 2069.430 ;
        RECT 1859.590 2069.420 1859.970 2069.430 ;
        RECT 1863.065 2069.730 1863.395 2069.745 ;
        RECT 1865.110 2069.730 1865.490 2069.740 ;
        RECT 1863.065 2069.430 1865.490 2069.730 ;
        RECT 1866.070 2069.730 1866.370 2070.110 ;
        RECT 1897.350 2070.110 1902.250 2070.410 ;
        RECT 1897.350 2069.730 1897.650 2070.110 ;
        RECT 1866.070 2069.430 1897.650 2069.730 ;
        RECT 1898.025 2069.730 1898.355 2069.745 ;
        RECT 1900.990 2069.730 1901.370 2069.740 ;
        RECT 1898.025 2069.430 1901.370 2069.730 ;
        RECT 1901.950 2069.730 1902.250 2070.110 ;
        RECT 1923.070 2069.730 1923.450 2069.740 ;
        RECT 1901.950 2069.430 1904.090 2069.730 ;
        RECT 1863.065 2069.415 1863.395 2069.430 ;
        RECT 1865.110 2069.420 1865.490 2069.430 ;
        RECT 1898.025 2069.415 1898.355 2069.430 ;
        RECT 1900.990 2069.420 1901.370 2069.430 ;
        RECT 300.000 2067.880 304.000 2068.480 ;
      LAYER met3 ;
        RECT 304.400 2067.480 1396.000 2068.880 ;
      LAYER met3 ;
        RECT 1770.605 2069.050 1770.935 2069.065 ;
        RECT 1903.085 2069.050 1903.415 2069.065 ;
        RECT 1770.605 2068.750 1903.415 2069.050 ;
        RECT 1903.790 2069.050 1904.090 2069.430 ;
        RECT 1907.470 2069.430 1923.450 2069.730 ;
        RECT 1907.470 2069.050 1907.770 2069.430 ;
        RECT 1923.070 2069.420 1923.450 2069.430 ;
        RECT 1939.425 2069.730 1939.755 2069.745 ;
        RECT 1953.225 2069.740 1953.555 2069.745 ;
        RECT 1941.470 2069.730 1941.850 2069.740 ;
        RECT 1953.225 2069.730 1953.810 2069.740 ;
        RECT 1939.425 2069.430 1941.850 2069.730 ;
        RECT 1953.000 2069.430 1953.810 2069.730 ;
        RECT 1939.425 2069.415 1939.755 2069.430 ;
        RECT 1941.470 2069.420 1941.850 2069.430 ;
        RECT 1953.225 2069.420 1953.810 2069.430 ;
        RECT 1960.125 2069.730 1960.455 2069.745 ;
        RECT 2014.865 2069.740 2015.195 2069.745 ;
        RECT 2038.785 2069.740 2039.115 2069.745 ;
        RECT 2052.585 2069.740 2052.915 2069.745 ;
        RECT 1964.470 2069.730 1964.850 2069.740 ;
        RECT 1989.310 2069.730 1989.690 2069.740 ;
        RECT 1960.125 2069.430 1964.850 2069.730 ;
        RECT 1953.225 2069.415 1953.555 2069.420 ;
        RECT 1960.125 2069.415 1960.455 2069.430 ;
        RECT 1964.470 2069.420 1964.850 2069.430 ;
        RECT 1965.430 2069.430 1989.690 2069.730 ;
        RECT 1903.790 2068.750 1907.770 2069.050 ;
        RECT 1921.485 2069.050 1921.815 2069.065 ;
        RECT 1959.665 2069.050 1959.995 2069.065 ;
        RECT 1960.790 2069.050 1961.170 2069.060 ;
        RECT 1921.485 2068.750 1948.250 2069.050 ;
        RECT 1770.605 2068.735 1770.935 2068.750 ;
        RECT 1903.085 2068.735 1903.415 2068.750 ;
        RECT 1921.485 2068.735 1921.815 2068.750 ;
        RECT 1417.785 2068.370 1418.115 2068.385 ;
        RECT 1946.990 2068.370 1947.370 2068.380 ;
        RECT 1417.785 2068.070 1947.370 2068.370 ;
        RECT 1947.950 2068.370 1948.250 2068.750 ;
        RECT 1959.665 2068.750 1961.170 2069.050 ;
        RECT 1959.665 2068.735 1959.995 2068.750 ;
        RECT 1960.790 2068.740 1961.170 2068.750 ;
        RECT 1965.430 2068.370 1965.730 2069.430 ;
        RECT 1989.310 2069.420 1989.690 2069.430 ;
        RECT 2014.865 2069.730 2015.450 2069.740 ;
        RECT 2038.785 2069.730 2039.370 2069.740 ;
        RECT 2014.865 2069.430 2015.650 2069.730 ;
        RECT 2038.560 2069.430 2039.370 2069.730 ;
        RECT 2014.865 2069.420 2015.450 2069.430 ;
        RECT 2038.785 2069.420 2039.370 2069.430 ;
        RECT 2052.585 2069.730 2053.170 2069.740 ;
        RECT 2353.425 2069.730 2353.755 2069.745 ;
        RECT 2374.125 2069.740 2374.455 2069.745 ;
        RECT 2354.550 2069.730 2354.930 2069.740 ;
        RECT 2373.870 2069.730 2374.455 2069.740 ;
        RECT 2052.585 2069.430 2053.370 2069.730 ;
        RECT 2353.425 2069.430 2354.930 2069.730 ;
        RECT 2373.670 2069.430 2374.455 2069.730 ;
        RECT 2052.585 2069.420 2053.170 2069.430 ;
        RECT 2014.865 2069.415 2015.195 2069.420 ;
        RECT 2038.785 2069.415 2039.115 2069.420 ;
        RECT 2052.585 2069.415 2052.915 2069.420 ;
        RECT 2353.425 2069.415 2353.755 2069.430 ;
        RECT 2354.550 2069.420 2354.930 2069.430 ;
        RECT 2373.870 2069.420 2374.455 2069.430 ;
        RECT 2374.125 2069.415 2374.455 2069.420 ;
        RECT 2387.925 2069.730 2388.255 2069.745 ;
        RECT 2391.350 2069.730 2391.730 2069.740 ;
        RECT 2387.925 2069.430 2391.730 2069.730 ;
        RECT 2387.925 2069.415 2388.255 2069.430 ;
        RECT 2391.350 2069.420 2391.730 2069.430 ;
        RECT 1980.365 2069.060 1980.695 2069.065 ;
        RECT 1980.110 2069.050 1980.695 2069.060 ;
        RECT 2380.565 2069.050 2380.895 2069.065 ;
        RECT 2387.465 2069.060 2387.795 2069.065 ;
        RECT 2381.230 2069.050 2381.610 2069.060 ;
        RECT 2387.465 2069.050 2388.050 2069.060 ;
        RECT 1980.110 2068.750 1980.920 2069.050 ;
        RECT 2380.565 2068.750 2381.610 2069.050 ;
        RECT 2387.240 2068.750 2388.050 2069.050 ;
        RECT 1980.110 2068.740 1980.695 2068.750 ;
        RECT 1980.365 2068.735 1980.695 2068.740 ;
        RECT 2380.565 2068.735 2380.895 2068.750 ;
        RECT 2381.230 2068.740 2381.610 2068.750 ;
        RECT 2387.465 2068.740 2388.050 2068.750 ;
        RECT 2525.465 2069.050 2525.795 2069.065 ;
        RECT 2528.430 2069.050 2528.810 2069.060 ;
        RECT 2525.465 2068.750 2528.810 2069.050 ;
        RECT 2387.465 2068.735 2387.795 2068.740 ;
        RECT 2525.465 2068.735 2525.795 2068.750 ;
        RECT 2528.430 2068.740 2528.810 2068.750 ;
        RECT 1947.950 2068.070 1965.730 2068.370 ;
        RECT 2394.365 2068.370 2394.695 2068.385 ;
        RECT 2396.870 2068.370 2397.250 2068.380 ;
        RECT 2394.365 2068.070 2397.250 2068.370 ;
        RECT 1417.785 2068.055 1418.115 2068.070 ;
        RECT 1946.990 2068.060 1947.370 2068.070 ;
        RECT 2394.365 2068.055 2394.695 2068.070 ;
        RECT 2396.870 2068.060 2397.250 2068.070 ;
        RECT 2532.365 2068.370 2532.695 2068.385 ;
        RECT 2534.870 2068.370 2535.250 2068.380 ;
        RECT 2532.365 2068.070 2535.250 2068.370 ;
        RECT 2532.365 2068.055 2532.695 2068.070 ;
        RECT 2534.870 2068.060 2535.250 2068.070 ;
      LAYER met3 ;
        RECT 300.065 2066.840 1396.000 2067.480 ;
      LAYER met3 ;
        RECT 1418.705 2067.690 1419.035 2067.705 ;
        RECT 1926.545 2067.690 1926.875 2067.705 ;
        RECT 1932.065 2067.700 1932.395 2067.705 ;
        RECT 1945.865 2067.700 1946.195 2067.705 ;
        RECT 1932.065 2067.690 1932.650 2067.700 ;
        RECT 1945.865 2067.690 1946.450 2067.700 ;
        RECT 1418.705 2067.390 1926.875 2067.690 ;
        RECT 1931.840 2067.390 1932.650 2067.690 ;
        RECT 1945.640 2067.390 1946.450 2067.690 ;
        RECT 1418.705 2067.375 1419.035 2067.390 ;
        RECT 1926.545 2067.375 1926.875 2067.390 ;
        RECT 1932.065 2067.380 1932.650 2067.390 ;
        RECT 1945.865 2067.380 1946.450 2067.390 ;
        RECT 1946.785 2067.690 1947.115 2067.705 ;
        RECT 1973.465 2067.700 1973.795 2067.705 ;
        RECT 2021.765 2067.700 2022.095 2067.705 ;
        RECT 1973.465 2067.690 1974.050 2067.700 ;
        RECT 2007.710 2067.690 2008.090 2067.700 ;
        RECT 1946.785 2067.390 1965.730 2067.690 ;
        RECT 1973.240 2067.390 1974.050 2067.690 ;
        RECT 1932.065 2067.375 1932.395 2067.380 ;
        RECT 1945.865 2067.375 1946.195 2067.380 ;
        RECT 1946.785 2067.375 1947.115 2067.390 ;
        RECT 1416.865 2067.010 1417.195 2067.025 ;
        RECT 1435.265 2067.010 1435.595 2067.025 ;
      LAYER met3 ;
        RECT 300.065 2065.440 1395.600 2066.840 ;
      LAYER met3 ;
        RECT 1416.865 2066.710 1435.595 2067.010 ;
        RECT 1416.865 2066.695 1417.195 2066.710 ;
        RECT 1435.265 2066.695 1435.595 2066.710 ;
        RECT 1483.105 2067.010 1483.435 2067.025 ;
        RECT 1531.865 2067.010 1532.195 2067.025 ;
        RECT 1483.105 2066.710 1532.195 2067.010 ;
        RECT 1483.105 2066.695 1483.435 2066.710 ;
        RECT 1531.865 2066.695 1532.195 2066.710 ;
        RECT 1579.705 2067.010 1580.035 2067.025 ;
        RECT 1676.305 2067.010 1676.635 2067.025 ;
        RECT 1772.905 2067.010 1773.235 2067.025 ;
        RECT 1821.665 2067.010 1821.995 2067.025 ;
        RECT 1579.705 2066.710 1605.090 2067.010 ;
        RECT 1579.705 2066.695 1580.035 2066.710 ;
        RECT 1396.000 2066.330 1400.000 2066.440 ;
        RECT 1414.105 2066.330 1414.435 2066.345 ;
        RECT 1396.000 2066.030 1414.435 2066.330 ;
        RECT 1396.000 2065.840 1400.000 2066.030 ;
        RECT 1414.105 2066.015 1414.435 2066.030 ;
        RECT 1419.625 2066.330 1419.955 2066.345 ;
        RECT 1435.725 2066.330 1436.055 2066.345 ;
        RECT 1419.625 2066.030 1436.055 2066.330 ;
        RECT 1419.625 2066.015 1419.955 2066.030 ;
        RECT 1435.725 2066.015 1436.055 2066.030 ;
        RECT 1482.645 2066.330 1482.975 2066.345 ;
        RECT 1532.325 2066.330 1532.655 2066.345 ;
        RECT 1482.645 2066.030 1532.655 2066.330 ;
        RECT 1482.645 2066.015 1482.975 2066.030 ;
        RECT 1532.325 2066.015 1532.655 2066.030 ;
        RECT 1579.245 2066.330 1579.575 2066.345 ;
        RECT 1579.245 2066.030 1603.250 2066.330 ;
        RECT 1579.245 2066.015 1579.575 2066.030 ;
        RECT 1435.265 2065.650 1435.595 2065.665 ;
        RECT 1483.105 2065.650 1483.435 2065.665 ;
      LAYER met3 ;
        RECT 300.065 2062.080 1396.000 2065.440 ;
      LAYER met3 ;
        RECT 1435.265 2065.350 1483.435 2065.650 ;
        RECT 1435.265 2065.335 1435.595 2065.350 ;
        RECT 1483.105 2065.335 1483.435 2065.350 ;
        RECT 1531.865 2065.650 1532.195 2065.665 ;
        RECT 1579.705 2065.650 1580.035 2065.665 ;
        RECT 1531.865 2065.350 1580.035 2065.650 ;
        RECT 1531.865 2065.335 1532.195 2065.350 ;
        RECT 1579.705 2065.335 1580.035 2065.350 ;
        RECT 1435.265 2064.970 1435.595 2064.985 ;
        RECT 1483.105 2064.970 1483.435 2064.985 ;
        RECT 1435.265 2064.670 1483.435 2064.970 ;
        RECT 1435.265 2064.655 1435.595 2064.670 ;
        RECT 1483.105 2064.655 1483.435 2064.670 ;
        RECT 1531.865 2064.970 1532.195 2064.985 ;
        RECT 1579.705 2064.970 1580.035 2064.985 ;
        RECT 1531.865 2064.670 1580.035 2064.970 ;
        RECT 1531.865 2064.655 1532.195 2064.670 ;
        RECT 1579.705 2064.655 1580.035 2064.670 ;
        RECT 1435.725 2064.290 1436.055 2064.305 ;
        RECT 1482.645 2064.290 1482.975 2064.305 ;
        RECT 1435.725 2063.990 1482.975 2064.290 ;
        RECT 1435.725 2063.975 1436.055 2063.990 ;
        RECT 1482.645 2063.975 1482.975 2063.990 ;
        RECT 1532.325 2064.290 1532.655 2064.305 ;
        RECT 1579.245 2064.290 1579.575 2064.305 ;
        RECT 1532.325 2063.990 1579.575 2064.290 ;
        RECT 1602.950 2064.290 1603.250 2066.030 ;
        RECT 1604.790 2065.650 1605.090 2066.710 ;
        RECT 1676.305 2066.710 1702.610 2067.010 ;
        RECT 1676.305 2066.695 1676.635 2066.710 ;
        RECT 1675.845 2066.330 1676.175 2066.345 ;
        RECT 1675.845 2066.030 1700.770 2066.330 ;
        RECT 1675.845 2066.015 1676.175 2066.030 ;
        RECT 1676.305 2065.650 1676.635 2065.665 ;
        RECT 1604.790 2065.350 1676.635 2065.650 ;
        RECT 1676.305 2065.335 1676.635 2065.350 ;
        RECT 1655.605 2064.970 1655.935 2064.985 ;
        RECT 1676.305 2064.970 1676.635 2064.985 ;
        RECT 1655.605 2064.670 1676.635 2064.970 ;
        RECT 1700.470 2064.970 1700.770 2066.030 ;
        RECT 1702.310 2065.650 1702.610 2066.710 ;
        RECT 1772.905 2066.710 1821.995 2067.010 ;
        RECT 1772.905 2066.695 1773.235 2066.710 ;
        RECT 1821.665 2066.695 1821.995 2066.710 ;
        RECT 1869.505 2067.010 1869.835 2067.025 ;
        RECT 1898.945 2067.010 1899.275 2067.025 ;
        RECT 1869.505 2066.710 1899.275 2067.010 ;
        RECT 1869.505 2066.695 1869.835 2066.710 ;
        RECT 1898.945 2066.695 1899.275 2066.710 ;
        RECT 1904.925 2067.010 1905.255 2067.025 ;
        RECT 1907.430 2067.010 1907.810 2067.020 ;
        RECT 1904.925 2066.710 1907.810 2067.010 ;
        RECT 1904.925 2066.695 1905.255 2066.710 ;
        RECT 1907.430 2066.700 1907.810 2066.710 ;
        RECT 1911.365 2067.010 1911.695 2067.025 ;
        RECT 1912.030 2067.010 1912.410 2067.020 ;
        RECT 1911.365 2066.710 1912.410 2067.010 ;
        RECT 1911.365 2066.695 1911.695 2066.710 ;
        RECT 1912.030 2066.700 1912.410 2066.710 ;
        RECT 1772.445 2066.330 1772.775 2066.345 ;
        RECT 1869.965 2066.330 1870.295 2066.345 ;
        RECT 1876.865 2066.340 1877.195 2066.345 ;
        RECT 1871.550 2066.330 1871.930 2066.340 ;
        RECT 1876.865 2066.330 1877.450 2066.340 ;
        RECT 1772.445 2066.030 1823.130 2066.330 ;
        RECT 1772.445 2066.015 1772.775 2066.030 ;
        RECT 1772.905 2065.650 1773.235 2065.665 ;
        RECT 1702.310 2065.350 1773.235 2065.650 ;
        RECT 1772.905 2065.335 1773.235 2065.350 ;
        RECT 1821.665 2065.650 1821.995 2065.665 ;
        RECT 1822.830 2065.650 1823.130 2066.030 ;
        RECT 1869.965 2066.030 1871.930 2066.330 ;
        RECT 1876.640 2066.030 1877.450 2066.330 ;
        RECT 1869.965 2066.015 1870.295 2066.030 ;
        RECT 1871.550 2066.020 1871.930 2066.030 ;
        RECT 1876.865 2066.020 1877.450 2066.030 ;
        RECT 1877.785 2066.330 1878.115 2066.345 ;
        RECT 1879.830 2066.330 1880.210 2066.340 ;
        RECT 1877.785 2066.030 1880.210 2066.330 ;
        RECT 1876.865 2066.015 1877.195 2066.020 ;
        RECT 1877.785 2066.015 1878.115 2066.030 ;
        RECT 1879.830 2066.020 1880.210 2066.030 ;
        RECT 1883.765 2066.330 1884.095 2066.345 ;
        RECT 1889.030 2066.330 1889.410 2066.340 ;
        RECT 1883.765 2066.030 1889.410 2066.330 ;
        RECT 1883.765 2066.015 1884.095 2066.030 ;
        RECT 1889.030 2066.020 1889.410 2066.030 ;
        RECT 1891.125 2066.330 1891.455 2066.345 ;
        RECT 1894.550 2066.330 1894.930 2066.340 ;
        RECT 1891.125 2066.030 1894.930 2066.330 ;
        RECT 1891.125 2066.015 1891.455 2066.030 ;
        RECT 1894.550 2066.020 1894.930 2066.030 ;
        RECT 1903.085 2066.330 1903.415 2066.345 ;
        RECT 1935.950 2066.330 1936.330 2066.340 ;
        RECT 1903.085 2066.030 1936.330 2066.330 ;
        RECT 1965.430 2066.330 1965.730 2067.390 ;
        RECT 1973.465 2067.380 1974.050 2067.390 ;
        RECT 1985.670 2067.390 2008.090 2067.690 ;
        RECT 1973.465 2067.375 1973.795 2067.380 ;
        RECT 1966.105 2067.010 1966.435 2067.025 ;
        RECT 1985.670 2067.010 1985.970 2067.390 ;
        RECT 2007.710 2067.380 2008.090 2067.390 ;
        RECT 2021.510 2067.690 2022.095 2067.700 ;
        RECT 2402.185 2067.690 2402.515 2067.705 ;
        RECT 2428.865 2067.700 2429.195 2067.705 ;
        RECT 2403.310 2067.690 2403.690 2067.700 ;
        RECT 2428.865 2067.690 2429.450 2067.700 ;
        RECT 2021.510 2067.390 2022.320 2067.690 ;
        RECT 2402.185 2067.390 2403.690 2067.690 ;
        RECT 2428.640 2067.390 2429.450 2067.690 ;
        RECT 2021.510 2067.380 2022.095 2067.390 ;
        RECT 2021.765 2067.375 2022.095 2067.380 ;
        RECT 2402.185 2067.375 2402.515 2067.390 ;
        RECT 2403.310 2067.380 2403.690 2067.390 ;
        RECT 2428.865 2067.380 2429.450 2067.390 ;
        RECT 2428.865 2067.375 2429.195 2067.380 ;
        RECT 1987.265 2067.020 1987.595 2067.025 ;
        RECT 1987.265 2067.010 1987.850 2067.020 ;
        RECT 1966.105 2066.710 1985.970 2067.010 ;
        RECT 1987.040 2066.710 1987.850 2067.010 ;
        RECT 1966.105 2066.695 1966.435 2066.710 ;
        RECT 1987.265 2066.700 1987.850 2066.710 ;
        RECT 2007.965 2067.010 2008.295 2067.025 ;
        RECT 2011.390 2067.010 2011.770 2067.020 ;
        RECT 2007.965 2066.710 2011.770 2067.010 ;
        RECT 1987.265 2066.695 1987.595 2066.700 ;
        RECT 2007.965 2066.695 2008.295 2066.710 ;
        RECT 2011.390 2066.700 2011.770 2066.710 ;
        RECT 2408.165 2067.010 2408.495 2067.025 ;
        RECT 2409.750 2067.010 2410.130 2067.020 ;
        RECT 2408.165 2066.710 2410.130 2067.010 ;
        RECT 2408.165 2066.695 2408.495 2066.710 ;
        RECT 2409.750 2066.700 2410.130 2066.710 ;
        RECT 2415.065 2067.010 2415.395 2067.025 ;
        RECT 2417.110 2067.010 2417.490 2067.020 ;
        RECT 2415.065 2066.710 2417.490 2067.010 ;
        RECT 2415.065 2066.695 2415.395 2066.710 ;
        RECT 2417.110 2066.700 2417.490 2066.710 ;
        RECT 2023.350 2066.330 2023.730 2066.340 ;
        RECT 1965.430 2066.030 2023.730 2066.330 ;
        RECT 1903.085 2066.015 1903.415 2066.030 ;
        RECT 1935.950 2066.020 1936.330 2066.030 ;
        RECT 2023.350 2066.020 2023.730 2066.030 ;
        RECT 2421.965 2066.330 2422.295 2066.345 ;
        RECT 2442.665 2066.340 2442.995 2066.345 ;
        RECT 2422.630 2066.330 2423.010 2066.340 ;
        RECT 2442.665 2066.330 2443.250 2066.340 ;
        RECT 2421.965 2066.030 2423.010 2066.330 ;
        RECT 2442.440 2066.030 2443.250 2066.330 ;
        RECT 2421.965 2066.015 2422.295 2066.030 ;
        RECT 2422.630 2066.020 2423.010 2066.030 ;
        RECT 2442.665 2066.020 2443.250 2066.030 ;
        RECT 2442.665 2066.015 2442.995 2066.020 ;
        RECT 1841.445 2065.650 1841.775 2065.665 ;
        RECT 1821.665 2065.335 1822.210 2065.650 ;
        RECT 1822.830 2065.350 1841.775 2065.650 ;
        RECT 1841.445 2065.335 1841.775 2065.350 ;
        RECT 1842.365 2065.650 1842.695 2065.665 ;
        RECT 1847.630 2065.650 1848.010 2065.660 ;
        RECT 1842.365 2065.350 1848.010 2065.650 ;
        RECT 1842.365 2065.335 1842.695 2065.350 ;
        RECT 1847.630 2065.340 1848.010 2065.350 ;
        RECT 1849.265 2065.650 1849.595 2065.665 ;
        RECT 1854.070 2065.650 1854.450 2065.660 ;
        RECT 1849.265 2065.350 1854.450 2065.650 ;
        RECT 1849.265 2065.335 1849.595 2065.350 ;
        RECT 1854.070 2065.340 1854.450 2065.350 ;
        RECT 1854.785 2065.650 1855.115 2065.665 ;
        RECT 1877.325 2065.650 1877.655 2065.665 ;
        RECT 1910.905 2065.660 1911.235 2065.665 ;
        RECT 1882.590 2065.650 1882.970 2065.660 ;
        RECT 1910.905 2065.650 1911.490 2065.660 ;
        RECT 1854.785 2065.350 1876.490 2065.650 ;
        RECT 1854.785 2065.335 1855.115 2065.350 ;
        RECT 1752.205 2064.970 1752.535 2064.985 ;
        RECT 1772.905 2064.970 1773.235 2064.985 ;
        RECT 1700.470 2064.670 1728.370 2064.970 ;
        RECT 1655.605 2064.655 1655.935 2064.670 ;
        RECT 1676.305 2064.655 1676.635 2064.670 ;
        RECT 1675.845 2064.290 1676.175 2064.305 ;
        RECT 1602.950 2063.990 1676.175 2064.290 ;
        RECT 1728.070 2064.290 1728.370 2064.670 ;
        RECT 1752.205 2064.670 1773.235 2064.970 ;
        RECT 1821.910 2064.970 1822.210 2065.335 ;
        RECT 1869.505 2064.970 1869.835 2064.985 ;
        RECT 1821.910 2064.670 1869.835 2064.970 ;
        RECT 1876.190 2064.970 1876.490 2065.350 ;
        RECT 1877.325 2065.350 1882.970 2065.650 ;
        RECT 1910.680 2065.350 1911.490 2065.650 ;
        RECT 1877.325 2065.335 1877.655 2065.350 ;
        RECT 1882.590 2065.340 1882.970 2065.350 ;
        RECT 1910.905 2065.340 1911.490 2065.350 ;
        RECT 1911.825 2065.650 1912.155 2065.665 ;
        RECT 1913.870 2065.650 1914.250 2065.660 ;
        RECT 1911.825 2065.350 1914.250 2065.650 ;
        RECT 1910.905 2065.335 1911.235 2065.340 ;
        RECT 1911.825 2065.335 1912.155 2065.350 ;
        RECT 1913.870 2065.340 1914.250 2065.350 ;
        RECT 1925.165 2065.650 1925.495 2065.665 ;
        RECT 1925.830 2065.650 1926.210 2065.660 ;
        RECT 1925.165 2065.350 1926.210 2065.650 ;
        RECT 1925.165 2065.335 1925.495 2065.350 ;
        RECT 1925.830 2065.340 1926.210 2065.350 ;
        RECT 1926.545 2065.650 1926.875 2065.665 ;
        RECT 1958.950 2065.650 1959.330 2065.660 ;
        RECT 1926.545 2065.350 1959.330 2065.650 ;
        RECT 1926.545 2065.335 1926.875 2065.350 ;
        RECT 1958.950 2065.340 1959.330 2065.350 ;
        RECT 1987.725 2065.650 1988.055 2065.665 ;
        RECT 1990.230 2065.650 1990.610 2065.660 ;
        RECT 1987.725 2065.350 1990.610 2065.650 ;
        RECT 1987.725 2065.335 1988.055 2065.350 ;
        RECT 1990.230 2065.340 1990.610 2065.350 ;
        RECT 1994.165 2065.650 1994.495 2065.665 ;
        RECT 1999.430 2065.650 1999.810 2065.660 ;
        RECT 1994.165 2065.350 1999.810 2065.650 ;
        RECT 1994.165 2065.335 1994.495 2065.350 ;
        RECT 1999.430 2065.340 1999.810 2065.350 ;
        RECT 2435.765 2065.650 2436.095 2065.665 ;
        RECT 2436.430 2065.650 2436.810 2065.660 ;
        RECT 2435.765 2065.350 2436.810 2065.650 ;
        RECT 2435.765 2065.335 2436.095 2065.350 ;
        RECT 2436.430 2065.340 2436.810 2065.350 ;
        RECT 1945.405 2064.970 1945.735 2064.985 ;
        RECT 1876.190 2064.670 1945.735 2064.970 ;
        RECT 1752.205 2064.655 1752.535 2064.670 ;
        RECT 1772.905 2064.655 1773.235 2064.670 ;
        RECT 1869.505 2064.655 1869.835 2064.670 ;
        RECT 1945.405 2064.655 1945.735 2064.670 ;
        RECT 1946.325 2064.970 1946.655 2064.985 ;
        RECT 1948.830 2064.970 1949.210 2064.980 ;
        RECT 1946.325 2064.670 1949.210 2064.970 ;
        RECT 1946.325 2064.655 1946.655 2064.670 ;
        RECT 1948.830 2064.660 1949.210 2064.670 ;
        RECT 1952.765 2064.970 1953.095 2064.985 ;
        RECT 1955.270 2064.970 1955.650 2064.980 ;
        RECT 1952.765 2064.670 1955.650 2064.970 ;
        RECT 1952.765 2064.655 1953.095 2064.670 ;
        RECT 1955.270 2064.660 1955.650 2064.670 ;
        RECT 1966.565 2064.970 1966.895 2064.985 ;
        RECT 1967.230 2064.970 1967.610 2064.980 ;
        RECT 1966.565 2064.670 1967.610 2064.970 ;
        RECT 1966.565 2064.655 1966.895 2064.670 ;
        RECT 1967.230 2064.660 1967.610 2064.670 ;
        RECT 1980.365 2064.970 1980.695 2064.985 ;
        RECT 1981.950 2064.970 1982.330 2064.980 ;
        RECT 1980.365 2064.670 1982.330 2064.970 ;
        RECT 1980.365 2064.655 1980.695 2064.670 ;
        RECT 1981.950 2064.660 1982.330 2064.670 ;
        RECT 1987.265 2064.970 1987.595 2064.985 ;
        RECT 1992.990 2064.970 1993.370 2064.980 ;
        RECT 1987.265 2064.670 1993.370 2064.970 ;
        RECT 1987.265 2064.655 1987.595 2064.670 ;
        RECT 1992.990 2064.660 1993.370 2064.670 ;
        RECT 2449.565 2064.970 2449.895 2064.985 ;
        RECT 2456.465 2064.980 2456.795 2064.985 ;
        RECT 2450.230 2064.970 2450.610 2064.980 ;
        RECT 2456.465 2064.970 2457.050 2064.980 ;
        RECT 2449.565 2064.670 2450.610 2064.970 ;
        RECT 2456.240 2064.670 2457.050 2064.970 ;
        RECT 2449.565 2064.655 2449.895 2064.670 ;
        RECT 2450.230 2064.660 2450.610 2064.670 ;
        RECT 2456.465 2064.660 2457.050 2064.670 ;
        RECT 2456.465 2064.655 2456.795 2064.660 ;
        RECT 1772.445 2064.290 1772.775 2064.305 ;
        RECT 1728.070 2063.990 1772.775 2064.290 ;
        RECT 1532.325 2063.975 1532.655 2063.990 ;
        RECT 1579.245 2063.975 1579.575 2063.990 ;
        RECT 1675.845 2063.975 1676.175 2063.990 ;
        RECT 1772.445 2063.975 1772.775 2063.990 ;
        RECT 1821.665 2064.290 1821.995 2064.305 ;
        RECT 1856.625 2064.290 1856.955 2064.305 ;
        RECT 1869.965 2064.300 1870.295 2064.305 ;
        RECT 1821.665 2063.990 1856.955 2064.290 ;
        RECT 1821.665 2063.975 1821.995 2063.990 ;
        RECT 1856.625 2063.975 1856.955 2063.990 ;
        RECT 1869.710 2064.290 1870.295 2064.300 ;
        RECT 1883.765 2064.290 1884.095 2064.305 ;
        RECT 1890.665 2064.300 1890.995 2064.305 ;
        RECT 1898.025 2064.300 1898.355 2064.305 ;
        RECT 1886.270 2064.290 1886.650 2064.300 ;
        RECT 1890.665 2064.290 1891.250 2064.300 ;
        RECT 1898.025 2064.290 1898.610 2064.300 ;
        RECT 1869.710 2063.990 1870.520 2064.290 ;
        RECT 1883.765 2063.990 1886.650 2064.290 ;
        RECT 1890.440 2063.990 1891.250 2064.290 ;
        RECT 1897.800 2063.990 1898.610 2064.290 ;
        RECT 1869.710 2063.980 1870.295 2063.990 ;
        RECT 1869.965 2063.975 1870.295 2063.980 ;
        RECT 1883.765 2063.975 1884.095 2063.990 ;
        RECT 1886.270 2063.980 1886.650 2063.990 ;
        RECT 1890.665 2063.980 1891.250 2063.990 ;
        RECT 1898.025 2063.980 1898.610 2063.990 ;
        RECT 1898.945 2064.290 1899.275 2064.305 ;
        RECT 1966.105 2064.290 1966.435 2064.305 ;
        RECT 1898.945 2063.990 1966.435 2064.290 ;
        RECT 1890.665 2063.975 1890.995 2063.980 ;
        RECT 1898.025 2063.975 1898.355 2063.980 ;
        RECT 1898.945 2063.975 1899.275 2063.990 ;
        RECT 1966.105 2063.975 1966.435 2063.990 ;
        RECT 1973.465 2064.290 1973.795 2064.305 ;
        RECT 1976.430 2064.290 1976.810 2064.300 ;
        RECT 1973.465 2063.990 1976.810 2064.290 ;
        RECT 1973.465 2063.975 1973.795 2063.990 ;
        RECT 1976.430 2063.980 1976.810 2063.990 ;
        RECT 2001.065 2064.290 2001.395 2064.305 ;
        RECT 2002.190 2064.290 2002.570 2064.300 ;
        RECT 2001.065 2063.990 2002.570 2064.290 ;
        RECT 2001.065 2063.975 2001.395 2063.990 ;
        RECT 2002.190 2063.980 2002.570 2063.990 ;
        RECT 2015.785 2064.290 2016.115 2064.305 ;
        RECT 2016.910 2064.290 2017.290 2064.300 ;
        RECT 2015.785 2063.990 2017.290 2064.290 ;
        RECT 2015.785 2063.975 2016.115 2063.990 ;
        RECT 2016.910 2063.980 2017.290 2063.990 ;
        RECT 1835.465 2063.610 1835.795 2063.625 ;
        RECT 1838.430 2063.610 1838.810 2063.620 ;
        RECT 1835.465 2063.310 1838.810 2063.610 ;
        RECT 1835.465 2063.295 1835.795 2063.310 ;
        RECT 1838.430 2063.300 1838.810 2063.310 ;
        RECT 1841.445 2063.610 1841.775 2063.625 ;
        RECT 1854.785 2063.610 1855.115 2063.625 ;
        RECT 1841.445 2063.310 1855.115 2063.610 ;
        RECT 1841.445 2063.295 1841.775 2063.310 ;
        RECT 1854.785 2063.295 1855.115 2063.310 ;
        RECT 1856.165 2063.610 1856.495 2063.625 ;
        RECT 1863.065 2063.620 1863.395 2063.625 ;
        RECT 1856.830 2063.610 1857.210 2063.620 ;
        RECT 1863.065 2063.610 1863.650 2063.620 ;
        RECT 1856.165 2063.310 1857.210 2063.610 ;
        RECT 1862.840 2063.310 1863.650 2063.610 ;
        RECT 1856.165 2063.295 1856.495 2063.310 ;
        RECT 1856.830 2063.300 1857.210 2063.310 ;
        RECT 1863.065 2063.300 1863.650 2063.310 ;
        RECT 1870.885 2063.610 1871.215 2063.625 ;
        RECT 1904.465 2063.620 1904.795 2063.625 ;
        RECT 1873.390 2063.610 1873.770 2063.620 ;
        RECT 1904.465 2063.610 1905.050 2063.620 ;
        RECT 1870.885 2063.310 1873.770 2063.610 ;
        RECT 1904.240 2063.310 1905.050 2063.610 ;
        RECT 1863.065 2063.295 1863.395 2063.300 ;
        RECT 1870.885 2063.295 1871.215 2063.310 ;
        RECT 1873.390 2063.300 1873.770 2063.310 ;
        RECT 1904.465 2063.300 1905.050 2063.310 ;
        RECT 1911.365 2063.610 1911.695 2063.625 ;
        RECT 1917.550 2063.610 1917.930 2063.620 ;
        RECT 1911.365 2063.310 1917.930 2063.610 ;
        RECT 1904.465 2063.295 1904.795 2063.300 ;
        RECT 1911.365 2063.295 1911.695 2063.310 ;
        RECT 1917.550 2063.300 1917.930 2063.310 ;
        RECT 1918.265 2063.610 1918.595 2063.625 ;
        RECT 1920.310 2063.610 1920.690 2063.620 ;
        RECT 1918.265 2063.310 1920.690 2063.610 ;
        RECT 1918.265 2063.295 1918.595 2063.310 ;
        RECT 1920.310 2063.300 1920.690 2063.310 ;
        RECT 1925.165 2063.610 1925.495 2063.625 ;
        RECT 1929.510 2063.610 1929.890 2063.620 ;
        RECT 1925.165 2063.310 1929.890 2063.610 ;
        RECT 1925.165 2063.295 1925.495 2063.310 ;
        RECT 1929.510 2063.300 1929.890 2063.310 ;
        RECT 1935.285 2063.610 1935.615 2063.625 ;
        RECT 1938.965 2063.610 1939.295 2063.625 ;
        RECT 1940.550 2063.610 1940.930 2063.620 ;
        RECT 1970.910 2063.610 1971.290 2063.620 ;
        RECT 1935.285 2063.310 1938.130 2063.610 ;
        RECT 1935.285 2063.295 1935.615 2063.310 ;
        RECT 1937.830 2062.930 1938.130 2063.310 ;
        RECT 1938.965 2063.310 1940.930 2063.610 ;
        RECT 1938.965 2063.295 1939.295 2063.310 ;
        RECT 1940.550 2063.300 1940.930 2063.310 ;
        RECT 1941.510 2063.310 1971.290 2063.610 ;
        RECT 1941.510 2062.930 1941.810 2063.310 ;
        RECT 1970.910 2063.300 1971.290 2063.310 ;
        RECT 1994.165 2063.610 1994.495 2063.625 ;
        RECT 1995.750 2063.610 1996.130 2063.620 ;
        RECT 1994.165 2063.310 1996.130 2063.610 ;
        RECT 1994.165 2063.295 1994.495 2063.310 ;
        RECT 1995.750 2063.300 1996.130 2063.310 ;
        RECT 2001.065 2063.610 2001.395 2063.625 ;
        RECT 2340.545 2063.620 2340.875 2063.625 ;
        RECT 2346.985 2063.620 2347.315 2063.625 ;
        RECT 2359.865 2063.620 2360.195 2063.625 ;
        RECT 2005.870 2063.610 2006.250 2063.620 ;
        RECT 2001.065 2063.310 2006.250 2063.610 ;
        RECT 2001.065 2063.295 2001.395 2063.310 ;
        RECT 2005.870 2063.300 2006.250 2063.310 ;
        RECT 2340.545 2063.610 2341.130 2063.620 ;
        RECT 2346.985 2063.610 2347.570 2063.620 ;
        RECT 2359.865 2063.610 2360.450 2063.620 ;
        RECT 2456.925 2063.610 2457.255 2063.625 ;
        RECT 2459.430 2063.610 2459.810 2063.620 ;
        RECT 2340.545 2063.310 2341.330 2063.610 ;
        RECT 2346.985 2063.310 2347.770 2063.610 ;
        RECT 2359.865 2063.310 2360.650 2063.610 ;
        RECT 2456.925 2063.310 2459.810 2063.610 ;
        RECT 2340.545 2063.300 2341.130 2063.310 ;
        RECT 2346.985 2063.300 2347.570 2063.310 ;
        RECT 2359.865 2063.300 2360.450 2063.310 ;
        RECT 2340.545 2063.295 2340.875 2063.300 ;
        RECT 2346.985 2063.295 2347.315 2063.300 ;
        RECT 2359.865 2063.295 2360.195 2063.300 ;
        RECT 2456.925 2063.295 2457.255 2063.310 ;
        RECT 2459.430 2063.300 2459.810 2063.310 ;
        RECT 2463.365 2063.610 2463.695 2063.625 ;
        RECT 2465.870 2063.610 2466.250 2063.620 ;
        RECT 2463.365 2063.310 2466.250 2063.610 ;
        RECT 2463.365 2063.295 2463.695 2063.310 ;
        RECT 2465.870 2063.300 2466.250 2063.310 ;
        RECT 2470.265 2063.610 2470.595 2063.625 ;
        RECT 2478.545 2063.620 2478.875 2063.625 ;
        RECT 2484.065 2063.620 2484.395 2063.625 ;
        RECT 2491.425 2063.620 2491.755 2063.625 ;
        RECT 2497.865 2063.620 2498.195 2063.625 ;
        RECT 2505.225 2063.620 2505.555 2063.625 ;
        RECT 2472.310 2063.610 2472.690 2063.620 ;
        RECT 2470.265 2063.310 2472.690 2063.610 ;
        RECT 2470.265 2063.295 2470.595 2063.310 ;
        RECT 2472.310 2063.300 2472.690 2063.310 ;
        RECT 2478.545 2063.610 2479.130 2063.620 ;
        RECT 2484.065 2063.610 2484.650 2063.620 ;
        RECT 2491.425 2063.610 2492.010 2063.620 ;
        RECT 2497.865 2063.610 2498.450 2063.620 ;
        RECT 2505.225 2063.610 2505.810 2063.620 ;
        RECT 2512.585 2063.610 2512.915 2063.625 ;
        RECT 2518.565 2063.620 2518.895 2063.625 ;
        RECT 2513.710 2063.610 2514.090 2063.620 ;
        RECT 2518.310 2063.610 2518.895 2063.620 ;
        RECT 2478.545 2063.310 2479.330 2063.610 ;
        RECT 2484.065 2063.310 2484.850 2063.610 ;
        RECT 2491.425 2063.310 2492.210 2063.610 ;
        RECT 2497.865 2063.310 2498.650 2063.610 ;
        RECT 2505.225 2063.310 2506.010 2063.610 ;
        RECT 2512.585 2063.310 2514.090 2063.610 ;
        RECT 2518.110 2063.310 2518.895 2063.610 ;
        RECT 2478.545 2063.300 2479.130 2063.310 ;
        RECT 2484.065 2063.300 2484.650 2063.310 ;
        RECT 2491.425 2063.300 2492.010 2063.310 ;
        RECT 2497.865 2063.300 2498.450 2063.310 ;
        RECT 2505.225 2063.300 2505.810 2063.310 ;
        RECT 2478.545 2063.295 2478.875 2063.300 ;
        RECT 2484.065 2063.295 2484.395 2063.300 ;
        RECT 2491.425 2063.295 2491.755 2063.300 ;
        RECT 2497.865 2063.295 2498.195 2063.300 ;
        RECT 2505.225 2063.295 2505.555 2063.300 ;
        RECT 2512.585 2063.295 2512.915 2063.310 ;
        RECT 2513.710 2063.300 2514.090 2063.310 ;
        RECT 2518.310 2063.300 2518.895 2063.310 ;
        RECT 2518.565 2063.295 2518.895 2063.300 ;
        RECT 2519.945 2063.610 2520.275 2063.625 ;
        RECT 2521.990 2063.610 2522.370 2063.620 ;
        RECT 2519.945 2063.310 2522.370 2063.610 ;
        RECT 2519.945 2063.295 2520.275 2063.310 ;
        RECT 2521.990 2063.300 2522.370 2063.310 ;
        RECT 2587.565 2063.610 2587.895 2063.625 ;
        RECT 2590.070 2063.610 2590.450 2063.620 ;
        RECT 2587.565 2063.310 2590.450 2063.610 ;
        RECT 2587.565 2063.295 2587.895 2063.310 ;
        RECT 2590.070 2063.300 2590.450 2063.310 ;
        RECT 1937.830 2062.630 1941.810 2062.930 ;
      LAYER met3 ;
        RECT 300.065 2060.680 1395.600 2062.080 ;
      LAYER met3 ;
        RECT 1396.000 2061.570 1400.000 2061.680 ;
        RECT 1414.105 2061.570 1414.435 2061.585 ;
        RECT 1396.000 2061.270 1414.435 2061.570 ;
        RECT 1396.000 2061.080 1400.000 2061.270 ;
        RECT 1414.105 2061.255 1414.435 2061.270 ;
      LAYER met3 ;
        RECT 300.065 2059.360 1396.000 2060.680 ;
      LAYER met3 ;
        RECT 300.000 2058.360 304.000 2058.960 ;
      LAYER met3 ;
        RECT 304.400 2057.960 1396.000 2059.360 ;
        RECT 300.065 2056.640 1396.000 2057.960 ;
      LAYER met3 ;
        RECT 2028.665 2057.500 2028.995 2057.505 ;
        RECT 2028.665 2057.490 2029.150 2057.500 ;
        RECT 2028.665 2057.190 2029.450 2057.490 ;
        RECT 2028.665 2057.180 2029.150 2057.190 ;
        RECT 2028.665 2057.175 2028.995 2057.180 ;
      LAYER met3 ;
        RECT 300.065 2055.240 1395.600 2056.640 ;
      LAYER met3 ;
        RECT 1396.000 2056.130 1400.000 2056.240 ;
        RECT 1414.105 2056.130 1414.435 2056.145 ;
        RECT 1396.000 2055.830 1414.435 2056.130 ;
        RECT 1396.000 2055.640 1400.000 2055.830 ;
        RECT 1414.105 2055.815 1414.435 2055.830 ;
      LAYER met3 ;
        RECT 300.065 2051.880 1396.000 2055.240 ;
      LAYER met3 ;
        RECT 2367.225 2052.060 2367.555 2052.065 ;
        RECT 2367.200 2052.050 2367.580 2052.060 ;
      LAYER met3 ;
        RECT 300.065 2050.480 1395.600 2051.880 ;
      LAYER met3 ;
        RECT 2366.770 2051.750 2367.580 2052.050 ;
        RECT 2367.200 2051.740 2367.580 2051.750 ;
        RECT 2367.225 2051.735 2367.555 2051.740 ;
        RECT 1396.000 2051.370 1400.000 2051.480 ;
        RECT 1413.645 2051.370 1413.975 2051.385 ;
        RECT 1396.000 2051.070 1413.975 2051.370 ;
        RECT 2609.280 2051.235 2611.020 2052.140 ;
        RECT 1396.000 2050.880 1400.000 2051.070 ;
        RECT 1413.645 2051.055 1413.975 2051.070 ;
      LAYER met3 ;
        RECT 300.065 2049.160 1396.000 2050.480 ;
      LAYER met3 ;
        RECT 300.000 2048.160 304.000 2048.760 ;
      LAYER met3 ;
        RECT 304.400 2047.760 1396.000 2049.160 ;
        RECT 300.065 2047.120 1396.000 2047.760 ;
        RECT 300.065 2045.720 1395.600 2047.120 ;
      LAYER met3 ;
        RECT 1396.000 2046.610 1400.000 2046.720 ;
        RECT 1408.585 2046.610 1408.915 2046.625 ;
        RECT 1396.000 2046.310 1408.915 2046.610 ;
        RECT 1396.000 2046.120 1400.000 2046.310 ;
        RECT 1408.585 2046.295 1408.915 2046.310 ;
      LAYER met3 ;
        RECT 300.065 2041.680 1396.000 2045.720 ;
        RECT 300.065 2040.280 1395.600 2041.680 ;
      LAYER met3 ;
        RECT 1396.000 2041.170 1400.000 2041.280 ;
        RECT 1408.585 2041.170 1408.915 2041.185 ;
        RECT 1396.000 2040.870 1408.915 2041.170 ;
        RECT 1396.000 2040.680 1400.000 2040.870 ;
        RECT 1408.585 2040.855 1408.915 2040.870 ;
      LAYER met3 ;
        RECT 300.065 2039.640 1396.000 2040.280 ;
      LAYER met3 ;
        RECT 300.000 2038.640 304.000 2039.240 ;
      LAYER met3 ;
        RECT 304.400 2038.240 1396.000 2039.640 ;
        RECT 300.065 2036.920 1396.000 2038.240 ;
        RECT 300.065 2035.520 1395.600 2036.920 ;
      LAYER met3 ;
        RECT 1396.000 2036.410 1400.000 2036.520 ;
        RECT 1414.105 2036.410 1414.435 2036.425 ;
        RECT 1396.000 2036.110 1414.435 2036.410 ;
        RECT 1396.000 2035.920 1400.000 2036.110 ;
        RECT 1414.105 2036.095 1414.435 2036.110 ;
      LAYER met3 ;
        RECT 300.065 2031.480 1396.000 2035.520 ;
        RECT 300.065 2030.120 1395.600 2031.480 ;
      LAYER met3 ;
        RECT 1396.000 2030.970 1400.000 2031.080 ;
        RECT 1411.805 2030.970 1412.135 2030.985 ;
        RECT 1396.000 2030.670 1412.135 2030.970 ;
        RECT 1396.000 2030.480 1400.000 2030.670 ;
        RECT 1411.805 2030.655 1412.135 2030.670 ;
      LAYER met3 ;
        RECT 304.400 2030.080 1395.600 2030.120 ;
      LAYER met3 ;
        RECT 300.000 2029.120 304.000 2029.720 ;
      LAYER met3 ;
        RECT 304.400 2028.720 1396.000 2030.080 ;
        RECT 300.065 2026.720 1396.000 2028.720 ;
        RECT 300.065 2025.320 1395.600 2026.720 ;
      LAYER met3 ;
        RECT 1396.000 2026.210 1400.000 2026.320 ;
        RECT 1414.105 2026.210 1414.435 2026.225 ;
        RECT 1396.000 2025.910 1414.435 2026.210 ;
        RECT 1396.000 2025.720 1400.000 2025.910 ;
        RECT 1414.105 2025.895 1414.435 2025.910 ;
      LAYER met3 ;
        RECT 300.065 2021.960 1396.000 2025.320 ;
        RECT 300.065 2020.600 1395.600 2021.960 ;
      LAYER met3 ;
        RECT 1396.000 2021.450 1400.000 2021.560 ;
        RECT 1414.105 2021.450 1414.435 2021.465 ;
        RECT 1396.000 2021.150 1414.435 2021.450 ;
        RECT 1396.000 2020.960 1400.000 2021.150 ;
        RECT 1414.105 2021.135 1414.435 2021.150 ;
      LAYER met3 ;
        RECT 304.400 2020.560 1395.600 2020.600 ;
      LAYER met3 ;
        RECT 300.000 2019.600 304.000 2020.200 ;
      LAYER met3 ;
        RECT 304.400 2019.200 1396.000 2020.560 ;
        RECT 300.065 2016.520 1396.000 2019.200 ;
        RECT 300.065 2015.120 1395.600 2016.520 ;
      LAYER met3 ;
        RECT 1396.000 2016.010 1400.000 2016.120 ;
        RECT 1408.125 2016.010 1408.455 2016.025 ;
        RECT 1396.000 2015.710 1408.455 2016.010 ;
        RECT 1396.000 2015.520 1400.000 2015.710 ;
        RECT 1408.125 2015.695 1408.455 2015.710 ;
      LAYER met3 ;
        RECT 300.065 2011.760 1396.000 2015.120 ;
        RECT 300.065 2011.080 1395.600 2011.760 ;
      LAYER met3 ;
        RECT 300.000 2010.080 304.000 2010.680 ;
      LAYER met3 ;
        RECT 304.400 2010.360 1395.600 2011.080 ;
      LAYER met3 ;
        RECT 1396.000 2011.250 1400.000 2011.360 ;
        RECT 1414.105 2011.250 1414.435 2011.265 ;
        RECT 1396.000 2010.950 1414.435 2011.250 ;
        RECT 1396.000 2010.760 1400.000 2010.950 ;
        RECT 1414.105 2010.935 1414.435 2010.950 ;
      LAYER met3 ;
        RECT 304.400 2009.680 1396.000 2010.360 ;
        RECT 300.065 2006.320 1396.000 2009.680 ;
        RECT 300.065 2004.920 1395.600 2006.320 ;
      LAYER met3 ;
        RECT 1396.000 2005.810 1400.000 2005.920 ;
        RECT 1414.105 2005.810 1414.435 2005.825 ;
        RECT 1396.000 2005.510 1414.435 2005.810 ;
        RECT 1396.000 2005.320 1400.000 2005.510 ;
        RECT 1414.105 2005.495 1414.435 2005.510 ;
      LAYER met3 ;
        RECT 300.065 2001.560 1396.000 2004.920 ;
        RECT 300.065 2000.880 1395.600 2001.560 ;
      LAYER met3 ;
        RECT 300.000 1999.880 304.000 2000.480 ;
      LAYER met3 ;
        RECT 304.400 2000.160 1395.600 2000.880 ;
      LAYER met3 ;
        RECT 1396.000 2001.050 1400.000 2001.160 ;
        RECT 1414.105 2001.050 1414.435 2001.065 ;
        RECT 1396.000 2000.750 1414.435 2001.050 ;
        RECT 1396.000 2000.560 1400.000 2000.750 ;
        RECT 1414.105 2000.735 1414.435 2000.750 ;
      LAYER met3 ;
        RECT 304.400 1999.480 1396.000 2000.160 ;
        RECT 300.065 1996.120 1396.000 1999.480 ;
        RECT 300.065 1994.720 1395.600 1996.120 ;
      LAYER met3 ;
        RECT 1396.000 1995.610 1400.000 1995.720 ;
        RECT 1411.345 1995.610 1411.675 1995.625 ;
        RECT 1396.000 1995.310 1411.675 1995.610 ;
        RECT 1396.000 1995.120 1400.000 1995.310 ;
        RECT 1411.345 1995.295 1411.675 1995.310 ;
      LAYER met3 ;
        RECT 300.065 1991.360 1396.000 1994.720 ;
      LAYER met3 ;
        RECT 300.000 1990.360 304.000 1990.960 ;
      LAYER met3 ;
        RECT 304.400 1989.960 1395.600 1991.360 ;
      LAYER met3 ;
        RECT 1396.000 1990.850 1400.000 1990.960 ;
        RECT 1408.125 1990.850 1408.455 1990.865 ;
        RECT 1396.000 1990.550 1408.455 1990.850 ;
        RECT 1396.000 1990.360 1400.000 1990.550 ;
        RECT 1408.125 1990.535 1408.455 1990.550 ;
      LAYER met3 ;
        RECT 300.065 1986.600 1396.000 1989.960 ;
        RECT 300.065 1985.200 1395.600 1986.600 ;
      LAYER met3 ;
        RECT 1396.000 1986.090 1400.000 1986.200 ;
        RECT 1408.125 1986.090 1408.455 1986.105 ;
        RECT 1396.000 1985.790 1408.455 1986.090 ;
        RECT 1396.000 1985.600 1400.000 1985.790 ;
        RECT 1408.125 1985.775 1408.455 1985.790 ;
      LAYER met3 ;
        RECT 300.065 1981.840 1396.000 1985.200 ;
      LAYER met3 ;
        RECT 300.000 1980.840 304.000 1981.440 ;
      LAYER met3 ;
        RECT 304.400 1981.160 1396.000 1981.840 ;
        RECT 304.400 1980.440 1395.600 1981.160 ;
        RECT 300.065 1979.760 1395.600 1980.440 ;
      LAYER met3 ;
        RECT 1396.000 1980.650 1400.000 1980.760 ;
        RECT 1408.125 1980.650 1408.455 1980.665 ;
        RECT 1396.000 1980.350 1408.455 1980.650 ;
        RECT 1396.000 1980.160 1400.000 1980.350 ;
        RECT 1408.125 1980.335 1408.455 1980.350 ;
      LAYER met3 ;
        RECT 300.065 1976.400 1396.000 1979.760 ;
        RECT 300.065 1975.000 1395.600 1976.400 ;
      LAYER met3 ;
        RECT 1396.000 1975.890 1400.000 1976.000 ;
        RECT 1408.125 1975.890 1408.455 1975.905 ;
        RECT 1396.000 1975.590 1408.455 1975.890 ;
        RECT 1396.000 1975.400 1400.000 1975.590 ;
        RECT 1408.125 1975.575 1408.455 1975.590 ;
      LAYER met3 ;
        RECT 300.065 1972.320 1396.000 1975.000 ;
      LAYER met3 ;
        RECT 300.000 1971.320 304.000 1971.920 ;
      LAYER met3 ;
        RECT 304.400 1970.960 1396.000 1972.320 ;
        RECT 304.400 1970.920 1395.600 1970.960 ;
        RECT 300.065 1969.560 1395.600 1970.920 ;
      LAYER met3 ;
        RECT 1396.000 1970.450 1400.000 1970.560 ;
        RECT 1408.125 1970.450 1408.455 1970.465 ;
        RECT 1396.000 1970.150 1408.455 1970.450 ;
        RECT 1396.000 1969.960 1400.000 1970.150 ;
        RECT 1408.125 1970.135 1408.455 1970.150 ;
      LAYER met3 ;
        RECT 300.065 1966.200 1396.000 1969.560 ;
        RECT 300.065 1964.800 1395.600 1966.200 ;
      LAYER met3 ;
        RECT 1396.000 1965.690 1400.000 1965.800 ;
        RECT 1408.125 1965.690 1408.455 1965.705 ;
        RECT 1396.000 1965.390 1408.455 1965.690 ;
        RECT 1396.000 1965.200 1400.000 1965.390 ;
        RECT 1408.125 1965.375 1408.455 1965.390 ;
      LAYER met3 ;
        RECT 300.065 1962.800 1396.000 1964.800 ;
      LAYER met3 ;
        RECT 300.000 1961.800 304.000 1962.400 ;
      LAYER met3 ;
        RECT 304.400 1961.400 1396.000 1962.800 ;
        RECT 300.065 1960.760 1396.000 1961.400 ;
        RECT 300.065 1959.360 1395.600 1960.760 ;
      LAYER met3 ;
        RECT 1396.000 1960.250 1400.000 1960.360 ;
        RECT 1408.125 1960.250 1408.455 1960.265 ;
        RECT 1396.000 1959.950 1408.455 1960.250 ;
        RECT 1396.000 1959.760 1400.000 1959.950 ;
        RECT 1408.125 1959.935 1408.455 1959.950 ;
      LAYER met3 ;
        RECT 300.065 1956.000 1396.000 1959.360 ;
        RECT 300.065 1954.600 1395.600 1956.000 ;
      LAYER met3 ;
        RECT 1396.000 1955.490 1400.000 1955.600 ;
        RECT 1408.125 1955.490 1408.455 1955.505 ;
        RECT 1396.000 1955.190 1408.455 1955.490 ;
        RECT 1396.000 1955.000 1400.000 1955.190 ;
        RECT 1408.125 1955.175 1408.455 1955.190 ;
      LAYER met3 ;
        RECT 300.065 1952.600 1396.000 1954.600 ;
      LAYER met3 ;
        RECT 300.000 1951.600 304.000 1952.200 ;
      LAYER met3 ;
        RECT 304.400 1951.240 1396.000 1952.600 ;
      LAYER met3 ;
        RECT 1700.000 1951.445 1704.600 1951.745 ;
      LAYER met3 ;
        RECT 304.400 1951.200 1395.600 1951.240 ;
        RECT 300.065 1949.840 1395.600 1951.200 ;
      LAYER met3 ;
        RECT 1396.000 1950.730 1400.000 1950.840 ;
        RECT 1408.125 1950.730 1408.455 1950.745 ;
        RECT 1396.000 1950.430 1408.455 1950.730 ;
        RECT 1396.000 1950.240 1400.000 1950.430 ;
        RECT 1408.125 1950.415 1408.455 1950.430 ;
      LAYER met3 ;
        RECT 300.065 1945.800 1396.000 1949.840 ;
      LAYER met3 ;
        RECT 1700.000 1945.805 1704.600 1946.105 ;
      LAYER met3 ;
        RECT 300.065 1944.400 1395.600 1945.800 ;
      LAYER met3 ;
        RECT 1396.000 1945.290 1400.000 1945.400 ;
        RECT 1408.125 1945.290 1408.455 1945.305 ;
        RECT 1396.000 1944.990 1408.455 1945.290 ;
        RECT 1396.000 1944.800 1400.000 1944.990 ;
        RECT 1408.125 1944.975 1408.455 1944.990 ;
      LAYER met3 ;
        RECT 300.065 1943.080 1396.000 1944.400 ;
      LAYER met3 ;
        RECT 300.000 1942.080 304.000 1942.680 ;
      LAYER met3 ;
        RECT 304.400 1941.680 1396.000 1943.080 ;
        RECT 300.065 1941.040 1396.000 1941.680 ;
        RECT 300.065 1939.640 1395.600 1941.040 ;
      LAYER met3 ;
        RECT 1396.000 1940.530 1400.000 1940.640 ;
        RECT 1408.125 1940.530 1408.455 1940.545 ;
        RECT 1396.000 1940.230 1408.455 1940.530 ;
        RECT 1396.000 1940.040 1400.000 1940.230 ;
        RECT 1408.125 1940.215 1408.455 1940.230 ;
      LAYER met3 ;
        RECT 300.065 1935.600 1396.000 1939.640 ;
      LAYER met3 ;
        RECT 1700.000 1937.305 1704.600 1937.605 ;
      LAYER met3 ;
        RECT 300.065 1934.200 1395.600 1935.600 ;
      LAYER met3 ;
        RECT 1396.000 1935.090 1400.000 1935.200 ;
        RECT 1408.125 1935.090 1408.455 1935.105 ;
        RECT 1396.000 1934.790 1408.455 1935.090 ;
        RECT 1396.000 1934.600 1400.000 1934.790 ;
        RECT 1408.125 1934.775 1408.455 1934.790 ;
      LAYER met3 ;
        RECT 300.065 1933.560 1396.000 1934.200 ;
      LAYER met3 ;
        RECT 300.000 1932.560 304.000 1933.160 ;
      LAYER met3 ;
        RECT 304.400 1932.160 1396.000 1933.560 ;
        RECT 300.065 1930.840 1396.000 1932.160 ;
      LAYER met3 ;
        RECT 1700.000 1931.665 1704.600 1931.965 ;
      LAYER met3 ;
        RECT 300.065 1929.440 1395.600 1930.840 ;
      LAYER met3 ;
        RECT 1396.000 1930.330 1400.000 1930.440 ;
        RECT 1408.125 1930.330 1408.455 1930.345 ;
        RECT 1396.000 1930.030 1408.455 1930.330 ;
        RECT 1396.000 1929.840 1400.000 1930.030 ;
        RECT 1408.125 1930.015 1408.455 1930.030 ;
      LAYER met3 ;
        RECT 300.065 1926.080 1396.000 1929.440 ;
        RECT 300.065 1924.680 1395.600 1926.080 ;
      LAYER met3 ;
        RECT 1396.000 1925.570 1400.000 1925.680 ;
        RECT 1408.125 1925.570 1408.455 1925.585 ;
        RECT 1396.000 1925.270 1408.455 1925.570 ;
        RECT 1396.000 1925.080 1400.000 1925.270 ;
        RECT 1408.125 1925.255 1408.455 1925.270 ;
      LAYER met3 ;
        RECT 300.065 1924.040 1396.000 1924.680 ;
      LAYER met3 ;
        RECT 300.000 1923.040 304.000 1923.640 ;
      LAYER met3 ;
        RECT 304.400 1922.640 1396.000 1924.040 ;
      LAYER met3 ;
        RECT 1700.000 1923.165 1704.600 1923.465 ;
      LAYER met3 ;
        RECT 300.065 1920.640 1396.000 1922.640 ;
        RECT 300.065 1919.240 1395.600 1920.640 ;
      LAYER met3 ;
        RECT 1396.000 1920.130 1400.000 1920.240 ;
        RECT 1408.125 1920.130 1408.455 1920.145 ;
        RECT 1396.000 1919.830 1408.455 1920.130 ;
        RECT 1396.000 1919.640 1400.000 1919.830 ;
        RECT 1408.125 1919.815 1408.455 1919.830 ;
      LAYER met3 ;
        RECT 300.065 1915.880 1396.000 1919.240 ;
      LAYER met3 ;
        RECT 1700.000 1917.525 1704.600 1917.825 ;
      LAYER met3 ;
        RECT 300.065 1914.520 1395.600 1915.880 ;
      LAYER met3 ;
        RECT 1396.000 1915.370 1400.000 1915.480 ;
        RECT 1408.125 1915.370 1408.455 1915.385 ;
        RECT 1396.000 1915.070 1408.455 1915.370 ;
        RECT 1396.000 1914.880 1400.000 1915.070 ;
        RECT 1408.125 1915.055 1408.455 1915.070 ;
      LAYER met3 ;
        RECT 304.400 1914.480 1395.600 1914.520 ;
      LAYER met3 ;
        RECT 300.000 1913.520 304.000 1914.120 ;
      LAYER met3 ;
        RECT 304.400 1913.120 1396.000 1914.480 ;
        RECT 300.065 1910.440 1396.000 1913.120 ;
        RECT 300.065 1909.040 1395.600 1910.440 ;
      LAYER met3 ;
        RECT 1396.000 1909.930 1400.000 1910.040 ;
        RECT 1408.125 1909.930 1408.455 1909.945 ;
        RECT 1396.000 1909.630 1408.455 1909.930 ;
        RECT 1396.000 1909.440 1400.000 1909.630 ;
        RECT 1408.125 1909.615 1408.455 1909.630 ;
      LAYER met3 ;
        RECT 300.065 1905.680 1396.000 1909.040 ;
      LAYER met3 ;
        RECT 1700.000 1909.025 1704.600 1909.325 ;
      LAYER met3 ;
        RECT 300.065 1904.320 1395.600 1905.680 ;
      LAYER met3 ;
        RECT 1396.000 1905.170 1400.000 1905.280 ;
        RECT 1409.045 1905.170 1409.375 1905.185 ;
        RECT 1396.000 1904.870 1409.375 1905.170 ;
        RECT 1396.000 1904.680 1400.000 1904.870 ;
        RECT 1409.045 1904.855 1409.375 1904.870 ;
      LAYER met3 ;
        RECT 304.400 1904.280 1395.600 1904.320 ;
      LAYER met3 ;
        RECT 300.000 1903.320 304.000 1903.920 ;
      LAYER met3 ;
        RECT 304.400 1902.920 1396.000 1904.280 ;
        RECT 300.065 1900.240 1396.000 1902.920 ;
        RECT 300.065 1898.840 1395.600 1900.240 ;
      LAYER met3 ;
        RECT 1396.000 1899.730 1400.000 1899.840 ;
        RECT 1408.125 1899.730 1408.455 1899.745 ;
        RECT 1396.000 1899.430 1408.455 1899.730 ;
        RECT 1396.000 1899.240 1400.000 1899.430 ;
        RECT 1408.125 1899.415 1408.455 1899.430 ;
      LAYER met3 ;
        RECT 300.065 1895.480 1396.000 1898.840 ;
        RECT 300.065 1894.800 1395.600 1895.480 ;
      LAYER met3 ;
        RECT 300.000 1893.800 304.000 1894.400 ;
      LAYER met3 ;
        RECT 304.400 1894.080 1395.600 1894.800 ;
      LAYER met3 ;
        RECT 1396.000 1894.970 1400.000 1895.080 ;
        RECT 1408.125 1894.970 1408.455 1894.985 ;
        RECT 1396.000 1894.670 1408.455 1894.970 ;
        RECT 1396.000 1894.480 1400.000 1894.670 ;
        RECT 1408.125 1894.655 1408.455 1894.670 ;
      LAYER met3 ;
        RECT 304.400 1893.400 1396.000 1894.080 ;
        RECT 300.065 1890.720 1396.000 1893.400 ;
        RECT 300.065 1889.320 1395.600 1890.720 ;
      LAYER met3 ;
        RECT 1396.000 1890.210 1400.000 1890.320 ;
        RECT 1408.125 1890.210 1408.455 1890.225 ;
        RECT 1396.000 1889.910 1408.455 1890.210 ;
        RECT 1396.000 1889.720 1400.000 1889.910 ;
        RECT 1408.125 1889.895 1408.455 1889.910 ;
      LAYER met3 ;
        RECT 300.065 1885.280 1396.000 1889.320 ;
      LAYER met3 ;
        RECT 300.000 1884.280 304.000 1884.880 ;
      LAYER met3 ;
        RECT 304.400 1883.880 1395.600 1885.280 ;
      LAYER met3 ;
        RECT 1396.000 1884.770 1400.000 1884.880 ;
        RECT 1409.045 1884.770 1409.375 1884.785 ;
        RECT 1396.000 1884.470 1409.375 1884.770 ;
        RECT 1396.000 1884.280 1400.000 1884.470 ;
        RECT 1409.045 1884.455 1409.375 1884.470 ;
      LAYER met3 ;
        RECT 300.065 1880.520 1396.000 1883.880 ;
        RECT 300.065 1879.120 1395.600 1880.520 ;
      LAYER met3 ;
        RECT 1396.000 1880.010 1400.000 1880.120 ;
        RECT 1408.125 1880.010 1408.455 1880.025 ;
        RECT 1396.000 1879.710 1408.455 1880.010 ;
        RECT 1396.000 1879.520 1400.000 1879.710 ;
        RECT 1408.125 1879.695 1408.455 1879.710 ;
      LAYER met3 ;
        RECT 300.065 1875.760 1396.000 1879.120 ;
      LAYER met3 ;
        RECT 300.000 1874.760 304.000 1875.360 ;
      LAYER met3 ;
        RECT 304.400 1875.080 1396.000 1875.760 ;
        RECT 304.400 1874.360 1395.600 1875.080 ;
        RECT 300.065 1873.680 1395.600 1874.360 ;
      LAYER met3 ;
        RECT 1396.000 1874.570 1400.000 1874.680 ;
        RECT 1408.125 1874.570 1408.455 1874.585 ;
        RECT 1396.000 1874.270 1408.455 1874.570 ;
        RECT 1396.000 1874.080 1400.000 1874.270 ;
        RECT 1408.125 1874.255 1408.455 1874.270 ;
      LAYER met3 ;
        RECT 300.065 1870.320 1396.000 1873.680 ;
        RECT 300.065 1868.920 1395.600 1870.320 ;
      LAYER met3 ;
        RECT 1396.000 1869.810 1400.000 1869.920 ;
        RECT 1408.125 1869.810 1408.455 1869.825 ;
        RECT 1396.000 1869.510 1408.455 1869.810 ;
        RECT 1396.000 1869.320 1400.000 1869.510 ;
        RECT 1408.125 1869.495 1408.455 1869.510 ;
      LAYER met3 ;
        RECT 300.065 1866.240 1396.000 1868.920 ;
      LAYER met3 ;
        RECT 300.000 1865.240 304.000 1865.840 ;
      LAYER met3 ;
        RECT 304.400 1864.880 1396.000 1866.240 ;
        RECT 304.400 1864.840 1395.600 1864.880 ;
        RECT 300.065 1863.480 1395.600 1864.840 ;
      LAYER met3 ;
        RECT 1396.000 1864.370 1400.000 1864.480 ;
        RECT 1409.045 1864.370 1409.375 1864.385 ;
        RECT 1396.000 1864.070 1409.375 1864.370 ;
        RECT 1396.000 1863.880 1400.000 1864.070 ;
        RECT 1409.045 1864.055 1409.375 1864.070 ;
      LAYER met3 ;
        RECT 300.065 1860.120 1396.000 1863.480 ;
        RECT 300.065 1858.720 1395.600 1860.120 ;
      LAYER met3 ;
        RECT 1396.000 1859.610 1400.000 1859.720 ;
        RECT 1408.125 1859.610 1408.455 1859.625 ;
        RECT 1396.000 1859.310 1408.455 1859.610 ;
        RECT 1396.000 1859.120 1400.000 1859.310 ;
        RECT 1408.125 1859.295 1408.455 1859.310 ;
      LAYER met3 ;
        RECT 300.065 1856.720 1396.000 1858.720 ;
      LAYER met3 ;
        RECT 300.000 1855.720 304.000 1856.320 ;
      LAYER met3 ;
        RECT 304.400 1855.360 1396.000 1856.720 ;
        RECT 304.400 1855.320 1395.600 1855.360 ;
        RECT 300.065 1853.960 1395.600 1855.320 ;
      LAYER met3 ;
        RECT 1396.000 1854.850 1400.000 1854.960 ;
        RECT 1408.125 1854.850 1408.455 1854.865 ;
        RECT 1396.000 1854.550 1408.455 1854.850 ;
        RECT 1396.000 1854.360 1400.000 1854.550 ;
        RECT 1408.125 1854.535 1408.455 1854.550 ;
      LAYER met3 ;
        RECT 300.065 1849.920 1396.000 1853.960 ;
        RECT 300.065 1848.520 1395.600 1849.920 ;
      LAYER met3 ;
        RECT 1396.000 1849.410 1400.000 1849.520 ;
        RECT 1409.045 1849.410 1409.375 1849.425 ;
        RECT 1396.000 1849.110 1409.375 1849.410 ;
        RECT 1396.000 1848.920 1400.000 1849.110 ;
        RECT 1409.045 1849.095 1409.375 1849.110 ;
      LAYER met3 ;
        RECT 300.065 1846.520 1396.000 1848.520 ;
      LAYER met3 ;
        RECT 300.000 1845.520 304.000 1846.120 ;
      LAYER met3 ;
        RECT 304.400 1845.160 1396.000 1846.520 ;
        RECT 304.400 1845.120 1395.600 1845.160 ;
        RECT 300.065 1843.760 1395.600 1845.120 ;
      LAYER met3 ;
        RECT 1396.000 1844.650 1400.000 1844.760 ;
        RECT 1408.125 1844.650 1408.455 1844.665 ;
        RECT 1396.000 1844.350 1408.455 1844.650 ;
        RECT 1396.000 1844.160 1400.000 1844.350 ;
        RECT 1408.125 1844.335 1408.455 1844.350 ;
      LAYER met3 ;
        RECT 300.065 1839.720 1396.000 1843.760 ;
        RECT 300.065 1838.320 1395.600 1839.720 ;
      LAYER met3 ;
        RECT 1396.000 1839.210 1400.000 1839.320 ;
        RECT 1408.125 1839.210 1408.455 1839.225 ;
        RECT 1396.000 1838.910 1408.455 1839.210 ;
        RECT 1396.000 1838.720 1400.000 1838.910 ;
        RECT 1408.125 1838.895 1408.455 1838.910 ;
      LAYER met3 ;
        RECT 300.065 1837.000 1396.000 1838.320 ;
      LAYER met3 ;
        RECT 300.000 1836.000 304.000 1836.600 ;
      LAYER met3 ;
        RECT 304.400 1835.600 1396.000 1837.000 ;
        RECT 300.065 1834.960 1396.000 1835.600 ;
        RECT 300.065 1833.560 1395.600 1834.960 ;
      LAYER met3 ;
        RECT 1396.000 1834.450 1400.000 1834.560 ;
        RECT 1422.385 1834.450 1422.715 1834.465 ;
        RECT 1396.000 1834.150 1422.715 1834.450 ;
        RECT 1396.000 1833.960 1400.000 1834.150 ;
        RECT 1422.385 1834.135 1422.715 1834.150 ;
      LAYER met3 ;
        RECT 300.065 1829.520 1396.000 1833.560 ;
        RECT 300.065 1828.120 1395.600 1829.520 ;
      LAYER met3 ;
        RECT 1396.000 1829.010 1400.000 1829.120 ;
        RECT 1425.605 1829.010 1425.935 1829.025 ;
        RECT 1396.000 1828.710 1425.935 1829.010 ;
        RECT 1396.000 1828.520 1400.000 1828.710 ;
        RECT 1425.605 1828.695 1425.935 1828.710 ;
      LAYER met3 ;
        RECT 300.065 1827.480 1396.000 1828.120 ;
      LAYER met3 ;
        RECT 300.000 1826.480 304.000 1827.080 ;
      LAYER met3 ;
        RECT 304.400 1826.080 1396.000 1827.480 ;
        RECT 300.065 1824.760 1396.000 1826.080 ;
        RECT 300.065 1823.360 1395.600 1824.760 ;
      LAYER met3 ;
        RECT 1396.000 1824.250 1400.000 1824.360 ;
        RECT 1408.125 1824.250 1408.455 1824.265 ;
        RECT 1396.000 1823.950 1408.455 1824.250 ;
        RECT 1396.000 1823.760 1400.000 1823.950 ;
        RECT 1408.125 1823.935 1408.455 1823.950 ;
      LAYER met3 ;
        RECT 300.065 1820.000 1396.000 1823.360 ;
        RECT 300.065 1818.600 1395.600 1820.000 ;
      LAYER met3 ;
        RECT 1396.000 1819.490 1400.000 1819.600 ;
        RECT 1408.125 1819.490 1408.455 1819.505 ;
        RECT 1396.000 1819.190 1408.455 1819.490 ;
        RECT 1396.000 1819.000 1400.000 1819.190 ;
        RECT 1408.125 1819.175 1408.455 1819.190 ;
      LAYER met3 ;
        RECT 300.065 1817.960 1396.000 1818.600 ;
      LAYER met3 ;
        RECT 300.000 1816.960 304.000 1817.560 ;
      LAYER met3 ;
        RECT 304.400 1816.560 1396.000 1817.960 ;
        RECT 300.065 1814.560 1396.000 1816.560 ;
        RECT 300.065 1813.160 1395.600 1814.560 ;
      LAYER met3 ;
        RECT 1396.000 1814.050 1400.000 1814.160 ;
        RECT 1408.125 1814.050 1408.455 1814.065 ;
        RECT 1396.000 1813.750 1408.455 1814.050 ;
        RECT 1396.000 1813.560 1400.000 1813.750 ;
        RECT 1408.125 1813.735 1408.455 1813.750 ;
      LAYER met3 ;
        RECT 300.065 1809.800 1396.000 1813.160 ;
        RECT 300.065 1808.440 1395.600 1809.800 ;
      LAYER met3 ;
        RECT 1396.000 1809.290 1400.000 1809.400 ;
        RECT 1409.045 1809.290 1409.375 1809.305 ;
        RECT 1396.000 1808.990 1409.375 1809.290 ;
        RECT 1396.000 1808.800 1400.000 1808.990 ;
        RECT 1409.045 1808.975 1409.375 1808.990 ;
      LAYER met3 ;
        RECT 304.400 1808.400 1395.600 1808.440 ;
      LAYER met3 ;
        RECT 300.000 1807.440 304.000 1808.040 ;
      LAYER met3 ;
        RECT 304.400 1807.040 1396.000 1808.400 ;
        RECT 300.065 1804.360 1396.000 1807.040 ;
        RECT 300.065 1802.960 1395.600 1804.360 ;
      LAYER met3 ;
        RECT 1396.000 1803.850 1400.000 1803.960 ;
        RECT 1408.125 1803.850 1408.455 1803.865 ;
        RECT 1396.000 1803.550 1408.455 1803.850 ;
        RECT 1396.000 1803.360 1400.000 1803.550 ;
        RECT 1408.125 1803.535 1408.455 1803.550 ;
      LAYER met3 ;
        RECT 300.065 1799.600 1396.000 1802.960 ;
        RECT 300.065 1798.240 1395.600 1799.600 ;
      LAYER met3 ;
        RECT 1396.000 1799.090 1400.000 1799.200 ;
        RECT 1408.125 1799.090 1408.455 1799.105 ;
        RECT 1396.000 1798.790 1408.455 1799.090 ;
        RECT 1396.000 1798.600 1400.000 1798.790 ;
        RECT 1408.125 1798.775 1408.455 1798.790 ;
      LAYER met3 ;
        RECT 304.400 1798.200 1395.600 1798.240 ;
      LAYER met3 ;
        RECT 300.000 1797.240 304.000 1797.840 ;
      LAYER met3 ;
        RECT 304.400 1796.840 1396.000 1798.200 ;
        RECT 300.065 1794.840 1396.000 1796.840 ;
        RECT 300.065 1793.440 1395.600 1794.840 ;
      LAYER met3 ;
        RECT 1396.000 1794.330 1400.000 1794.440 ;
        RECT 1409.045 1794.330 1409.375 1794.345 ;
        RECT 1396.000 1794.030 1409.375 1794.330 ;
        RECT 1396.000 1793.840 1400.000 1794.030 ;
        RECT 1409.045 1794.015 1409.375 1794.030 ;
      LAYER met3 ;
        RECT 300.065 1789.400 1396.000 1793.440 ;
        RECT 300.065 1788.720 1395.600 1789.400 ;
      LAYER met3 ;
        RECT 300.000 1787.720 304.000 1788.320 ;
      LAYER met3 ;
        RECT 304.400 1788.000 1395.600 1788.720 ;
      LAYER met3 ;
        RECT 1396.000 1788.890 1400.000 1789.000 ;
        RECT 1408.125 1788.890 1408.455 1788.905 ;
        RECT 1396.000 1788.590 1408.455 1788.890 ;
        RECT 1396.000 1788.400 1400.000 1788.590 ;
        RECT 1408.125 1788.575 1408.455 1788.590 ;
      LAYER met3 ;
        RECT 304.400 1787.320 1396.000 1788.000 ;
        RECT 300.065 1784.640 1396.000 1787.320 ;
        RECT 300.065 1783.240 1395.600 1784.640 ;
      LAYER met3 ;
        RECT 1396.000 1784.130 1400.000 1784.240 ;
        RECT 1413.185 1784.130 1413.515 1784.145 ;
        RECT 1396.000 1783.830 1413.515 1784.130 ;
        RECT 1396.000 1783.640 1400.000 1783.830 ;
        RECT 1413.185 1783.815 1413.515 1783.830 ;
      LAYER met3 ;
        RECT 300.065 1779.200 1396.000 1783.240 ;
      LAYER met3 ;
        RECT 300.000 1778.200 304.000 1778.800 ;
      LAYER met3 ;
        RECT 304.400 1777.800 1395.600 1779.200 ;
      LAYER met3 ;
        RECT 1396.000 1778.690 1400.000 1778.800 ;
        RECT 1412.725 1778.690 1413.055 1778.705 ;
        RECT 1396.000 1778.390 1413.055 1778.690 ;
        RECT 1396.000 1778.200 1400.000 1778.390 ;
        RECT 1412.725 1778.375 1413.055 1778.390 ;
      LAYER met3 ;
        RECT 300.065 1774.440 1396.000 1777.800 ;
        RECT 300.065 1773.040 1395.600 1774.440 ;
      LAYER met3 ;
        RECT 1396.000 1773.930 1400.000 1774.040 ;
        RECT 1411.345 1773.930 1411.675 1773.945 ;
        RECT 1396.000 1773.630 1411.675 1773.930 ;
        RECT 1396.000 1773.440 1400.000 1773.630 ;
        RECT 1411.345 1773.615 1411.675 1773.630 ;
      LAYER met3 ;
        RECT 300.065 1769.680 1396.000 1773.040 ;
      LAYER met3 ;
        RECT 300.000 1768.680 304.000 1769.280 ;
      LAYER met3 ;
        RECT 304.400 1769.000 1396.000 1769.680 ;
        RECT 304.400 1768.280 1395.600 1769.000 ;
        RECT 300.065 1767.600 1395.600 1768.280 ;
      LAYER met3 ;
        RECT 1396.000 1768.490 1400.000 1768.600 ;
        RECT 1412.265 1768.490 1412.595 1768.505 ;
        RECT 1396.000 1768.190 1412.595 1768.490 ;
        RECT 1396.000 1768.000 1400.000 1768.190 ;
        RECT 1412.265 1768.175 1412.595 1768.190 ;
      LAYER met3 ;
        RECT 300.065 1764.240 1396.000 1767.600 ;
        RECT 300.065 1762.840 1395.600 1764.240 ;
      LAYER met3 ;
        RECT 1396.000 1763.730 1400.000 1763.840 ;
        RECT 1411.805 1763.730 1412.135 1763.745 ;
        RECT 1396.000 1763.430 1412.135 1763.730 ;
        RECT 1396.000 1763.240 1400.000 1763.430 ;
        RECT 1411.805 1763.415 1412.135 1763.430 ;
      LAYER met3 ;
        RECT 300.065 1760.160 1396.000 1762.840 ;
      LAYER met3 ;
        RECT 300.000 1759.160 304.000 1759.760 ;
      LAYER met3 ;
        RECT 304.400 1759.480 1396.000 1760.160 ;
        RECT 304.400 1758.760 1395.600 1759.480 ;
        RECT 300.065 1758.080 1395.600 1758.760 ;
      LAYER met3 ;
        RECT 1396.000 1758.970 1400.000 1759.080 ;
        RECT 1408.125 1758.970 1408.455 1758.985 ;
        RECT 1396.000 1758.670 1408.455 1758.970 ;
        RECT 1396.000 1758.480 1400.000 1758.670 ;
        RECT 1408.125 1758.655 1408.455 1758.670 ;
      LAYER met3 ;
        RECT 300.065 1754.040 1396.000 1758.080 ;
        RECT 300.065 1752.640 1395.600 1754.040 ;
      LAYER met3 ;
        RECT 1396.000 1753.530 1400.000 1753.640 ;
        RECT 1408.125 1753.530 1408.455 1753.545 ;
        RECT 1396.000 1753.230 1408.455 1753.530 ;
        RECT 1396.000 1753.040 1400.000 1753.230 ;
        RECT 1408.125 1753.215 1408.455 1753.230 ;
      LAYER met3 ;
        RECT 300.065 1749.960 1396.000 1752.640 ;
      LAYER met3 ;
        RECT 300.000 1748.960 304.000 1749.560 ;
      LAYER met3 ;
        RECT 304.400 1749.280 1396.000 1749.960 ;
        RECT 304.400 1748.560 1395.600 1749.280 ;
        RECT 300.065 1747.880 1395.600 1748.560 ;
      LAYER met3 ;
        RECT 1396.000 1748.770 1400.000 1748.880 ;
        RECT 1408.125 1748.770 1408.455 1748.785 ;
        RECT 1396.000 1748.470 1408.455 1748.770 ;
        RECT 1396.000 1748.280 1400.000 1748.470 ;
        RECT 1408.125 1748.455 1408.455 1748.470 ;
      LAYER met3 ;
        RECT 300.065 1743.840 1396.000 1747.880 ;
        RECT 300.065 1742.440 1395.600 1743.840 ;
      LAYER met3 ;
        RECT 1396.000 1743.330 1400.000 1743.440 ;
        RECT 1408.125 1743.330 1408.455 1743.345 ;
        RECT 1396.000 1743.030 1408.455 1743.330 ;
        RECT 1396.000 1742.840 1400.000 1743.030 ;
        RECT 1408.125 1743.015 1408.455 1743.030 ;
      LAYER met3 ;
        RECT 300.065 1740.440 1396.000 1742.440 ;
      LAYER met3 ;
        RECT 300.000 1739.440 304.000 1740.040 ;
      LAYER met3 ;
        RECT 304.400 1739.080 1396.000 1740.440 ;
        RECT 304.400 1739.040 1395.600 1739.080 ;
        RECT 300.065 1737.680 1395.600 1739.040 ;
      LAYER met3 ;
        RECT 1396.000 1738.570 1400.000 1738.680 ;
        RECT 1408.125 1738.570 1408.455 1738.585 ;
        RECT 1396.000 1738.270 1408.455 1738.570 ;
        RECT 1396.000 1738.080 1400.000 1738.270 ;
        RECT 1408.125 1738.255 1408.455 1738.270 ;
      LAYER met3 ;
        RECT 300.065 1733.640 1396.000 1737.680 ;
        RECT 300.065 1732.240 1395.600 1733.640 ;
      LAYER met3 ;
        RECT 1396.000 1733.130 1400.000 1733.240 ;
        RECT 1408.125 1733.130 1408.455 1733.145 ;
        RECT 1396.000 1732.830 1408.455 1733.130 ;
        RECT 1396.000 1732.640 1400.000 1732.830 ;
        RECT 1408.125 1732.815 1408.455 1732.830 ;
      LAYER met3 ;
        RECT 300.065 1730.920 1396.000 1732.240 ;
      LAYER met3 ;
        RECT 300.000 1729.920 304.000 1730.520 ;
      LAYER met3 ;
        RECT 304.400 1729.520 1396.000 1730.920 ;
        RECT 300.065 1728.880 1396.000 1729.520 ;
        RECT 300.065 1727.480 1395.600 1728.880 ;
      LAYER met3 ;
        RECT 1396.000 1728.370 1400.000 1728.480 ;
        RECT 1408.125 1728.370 1408.455 1728.385 ;
        RECT 1396.000 1728.070 1408.455 1728.370 ;
        RECT 1396.000 1727.880 1400.000 1728.070 ;
        RECT 1408.125 1728.055 1408.455 1728.070 ;
      LAYER met3 ;
        RECT 300.065 1724.120 1396.000 1727.480 ;
        RECT 300.065 1722.720 1395.600 1724.120 ;
      LAYER met3 ;
        RECT 1396.000 1723.610 1400.000 1723.720 ;
        RECT 1408.125 1723.610 1408.455 1723.625 ;
        RECT 1396.000 1723.310 1408.455 1723.610 ;
        RECT 1396.000 1723.120 1400.000 1723.310 ;
        RECT 1408.125 1723.295 1408.455 1723.310 ;
      LAYER met3 ;
        RECT 300.065 1721.400 1396.000 1722.720 ;
      LAYER met3 ;
        RECT 300.000 1720.400 304.000 1721.000 ;
      LAYER met3 ;
        RECT 304.400 1720.000 1396.000 1721.400 ;
        RECT 300.065 1718.680 1396.000 1720.000 ;
        RECT 300.065 1717.280 1395.600 1718.680 ;
      LAYER met3 ;
        RECT 1396.000 1718.170 1400.000 1718.280 ;
        RECT 1408.125 1718.170 1408.455 1718.185 ;
        RECT 1396.000 1717.870 1408.455 1718.170 ;
        RECT 1396.000 1717.680 1400.000 1717.870 ;
        RECT 1408.125 1717.855 1408.455 1717.870 ;
      LAYER met3 ;
        RECT 300.065 1713.920 1396.000 1717.280 ;
        RECT 300.065 1712.520 1395.600 1713.920 ;
      LAYER met3 ;
        RECT 1396.000 1713.410 1400.000 1713.520 ;
        RECT 1409.045 1713.410 1409.375 1713.425 ;
        RECT 1396.000 1713.110 1409.375 1713.410 ;
        RECT 1396.000 1712.920 1400.000 1713.110 ;
        RECT 1409.045 1713.095 1409.375 1713.110 ;
      LAYER met3 ;
        RECT 300.065 1711.880 1396.000 1712.520 ;
      LAYER met3 ;
        RECT 300.000 1710.880 304.000 1711.480 ;
      LAYER met3 ;
        RECT 304.400 1710.480 1396.000 1711.880 ;
        RECT 300.065 1708.480 1396.000 1710.480 ;
        RECT 300.065 1707.080 1395.600 1708.480 ;
      LAYER met3 ;
        RECT 1396.000 1707.970 1400.000 1708.080 ;
        RECT 1408.125 1707.970 1408.455 1707.985 ;
        RECT 1396.000 1707.670 1408.455 1707.970 ;
        RECT 1396.000 1707.480 1400.000 1707.670 ;
        RECT 1408.125 1707.655 1408.455 1707.670 ;
      LAYER met3 ;
        RECT 300.065 1703.720 1396.000 1707.080 ;
        RECT 300.065 1702.320 1395.600 1703.720 ;
      LAYER met3 ;
        RECT 1396.000 1703.210 1400.000 1703.320 ;
        RECT 1408.125 1703.210 1408.455 1703.225 ;
        RECT 1396.000 1702.910 1408.455 1703.210 ;
        RECT 1396.000 1702.720 1400.000 1702.910 ;
        RECT 1408.125 1702.895 1408.455 1702.910 ;
      LAYER met3 ;
        RECT 300.065 1701.680 1396.000 1702.320 ;
      LAYER met3 ;
        RECT 300.000 1700.680 304.000 1701.280 ;
      LAYER met3 ;
        RECT 304.400 1700.280 1396.000 1701.680 ;
        RECT 300.065 1698.960 1396.000 1700.280 ;
        RECT 300.065 1697.560 1395.600 1698.960 ;
      LAYER met3 ;
        RECT 1396.000 1698.450 1400.000 1698.560 ;
        RECT 1408.585 1698.450 1408.915 1698.465 ;
        RECT 1396.000 1698.150 1408.915 1698.450 ;
        RECT 1396.000 1697.960 1400.000 1698.150 ;
        RECT 1408.585 1698.135 1408.915 1698.150 ;
      LAYER met3 ;
        RECT 300.065 1693.520 1396.000 1697.560 ;
        RECT 300.065 1692.160 1395.600 1693.520 ;
      LAYER met3 ;
        RECT 1396.000 1693.010 1400.000 1693.120 ;
        RECT 1408.125 1693.010 1408.455 1693.025 ;
        RECT 1396.000 1692.710 1408.455 1693.010 ;
        RECT 1396.000 1692.520 1400.000 1692.710 ;
        RECT 1408.125 1692.695 1408.455 1692.710 ;
      LAYER met3 ;
        RECT 304.400 1692.120 1395.600 1692.160 ;
      LAYER met3 ;
        RECT 300.000 1691.160 304.000 1691.760 ;
      LAYER met3 ;
        RECT 304.400 1690.760 1396.000 1692.120 ;
        RECT 300.065 1688.760 1396.000 1690.760 ;
        RECT 300.065 1687.360 1395.600 1688.760 ;
      LAYER met3 ;
        RECT 1396.000 1688.250 1400.000 1688.360 ;
        RECT 1408.125 1688.250 1408.455 1688.265 ;
        RECT 1396.000 1687.950 1408.455 1688.250 ;
        RECT 1396.000 1687.760 1400.000 1687.950 ;
        RECT 1408.125 1687.935 1408.455 1687.950 ;
      LAYER met3 ;
        RECT 300.065 1683.320 1396.000 1687.360 ;
        RECT 300.065 1682.640 1395.600 1683.320 ;
      LAYER met3 ;
        RECT 300.000 1681.640 304.000 1682.240 ;
      LAYER met3 ;
        RECT 304.400 1681.920 1395.600 1682.640 ;
      LAYER met3 ;
        RECT 1396.000 1682.810 1400.000 1682.920 ;
        RECT 1408.125 1682.810 1408.455 1682.825 ;
        RECT 1396.000 1682.510 1408.455 1682.810 ;
        RECT 1396.000 1682.320 1400.000 1682.510 ;
        RECT 1408.125 1682.495 1408.455 1682.510 ;
      LAYER met3 ;
        RECT 304.400 1681.240 1396.000 1681.920 ;
        RECT 300.065 1678.560 1396.000 1681.240 ;
        RECT 300.065 1677.160 1395.600 1678.560 ;
      LAYER met3 ;
        RECT 1396.000 1678.050 1400.000 1678.160 ;
        RECT 1408.585 1678.050 1408.915 1678.065 ;
        RECT 1396.000 1677.750 1408.915 1678.050 ;
        RECT 1396.000 1677.560 1400.000 1677.750 ;
        RECT 1408.585 1677.735 1408.915 1677.750 ;
      LAYER met3 ;
        RECT 300.065 1673.120 1396.000 1677.160 ;
      LAYER met3 ;
        RECT 300.000 1672.120 304.000 1672.720 ;
      LAYER met3 ;
        RECT 304.400 1671.720 1395.600 1673.120 ;
      LAYER met3 ;
        RECT 1396.000 1672.610 1400.000 1672.720 ;
        RECT 1408.125 1672.610 1408.455 1672.625 ;
        RECT 1396.000 1672.310 1408.455 1672.610 ;
        RECT 1396.000 1672.120 1400.000 1672.310 ;
        RECT 1408.125 1672.295 1408.455 1672.310 ;
      LAYER met3 ;
        RECT 300.065 1668.360 1396.000 1671.720 ;
        RECT 300.065 1666.960 1395.600 1668.360 ;
      LAYER met3 ;
        RECT 1396.000 1667.850 1400.000 1667.960 ;
        RECT 1408.125 1667.850 1408.455 1667.865 ;
        RECT 1396.000 1667.550 1408.455 1667.850 ;
        RECT 1396.000 1667.360 1400.000 1667.550 ;
        RECT 1408.125 1667.535 1408.455 1667.550 ;
      LAYER met3 ;
        RECT 300.065 1663.600 1396.000 1666.960 ;
      LAYER met3 ;
        RECT 300.000 1662.600 304.000 1663.200 ;
      LAYER met3 ;
        RECT 304.400 1662.200 1395.600 1663.600 ;
      LAYER met3 ;
        RECT 1396.000 1663.090 1400.000 1663.200 ;
        RECT 1408.585 1663.090 1408.915 1663.105 ;
        RECT 1396.000 1662.790 1408.915 1663.090 ;
        RECT 1396.000 1662.600 1400.000 1662.790 ;
        RECT 1408.585 1662.775 1408.915 1662.790 ;
      LAYER met3 ;
        RECT 300.065 1658.160 1396.000 1662.200 ;
        RECT 300.065 1656.760 1395.600 1658.160 ;
      LAYER met3 ;
        RECT 1396.000 1657.650 1400.000 1657.760 ;
        RECT 1409.505 1657.650 1409.835 1657.665 ;
        RECT 1396.000 1657.350 1409.835 1657.650 ;
        RECT 1396.000 1657.160 1400.000 1657.350 ;
        RECT 1409.505 1657.335 1409.835 1657.350 ;
      LAYER met3 ;
        RECT 300.065 1653.400 1396.000 1656.760 ;
      LAYER met3 ;
        RECT 300.000 1652.400 304.000 1653.000 ;
      LAYER met3 ;
        RECT 304.400 1652.000 1395.600 1653.400 ;
      LAYER met3 ;
        RECT 1396.000 1652.890 1400.000 1653.000 ;
        RECT 1408.125 1652.890 1408.455 1652.905 ;
        RECT 1396.000 1652.590 1408.455 1652.890 ;
        RECT 1396.000 1652.400 1400.000 1652.590 ;
        RECT 1408.125 1652.575 1408.455 1652.590 ;
      LAYER met3 ;
        RECT 300.065 1647.960 1396.000 1652.000 ;
        RECT 300.065 1646.560 1395.600 1647.960 ;
      LAYER met3 ;
        RECT 1396.000 1647.450 1400.000 1647.560 ;
        RECT 1407.665 1647.450 1407.995 1647.465 ;
        RECT 1396.000 1647.150 1407.995 1647.450 ;
        RECT 1396.000 1646.960 1400.000 1647.150 ;
        RECT 1407.665 1647.135 1407.995 1647.150 ;
      LAYER met3 ;
        RECT 300.065 1643.880 1396.000 1646.560 ;
      LAYER met3 ;
        RECT 300.000 1642.880 304.000 1643.480 ;
      LAYER met3 ;
        RECT 304.400 1643.200 1396.000 1643.880 ;
        RECT 304.400 1642.480 1395.600 1643.200 ;
        RECT 300.065 1641.800 1395.600 1642.480 ;
      LAYER met3 ;
        RECT 1396.000 1642.690 1400.000 1642.800 ;
        RECT 1408.125 1642.690 1408.455 1642.705 ;
        RECT 1396.000 1642.390 1408.455 1642.690 ;
        RECT 1396.000 1642.200 1400.000 1642.390 ;
        RECT 1408.125 1642.375 1408.455 1642.390 ;
      LAYER met3 ;
        RECT 300.065 1637.760 1396.000 1641.800 ;
        RECT 300.065 1636.360 1395.600 1637.760 ;
      LAYER met3 ;
        RECT 1396.000 1637.250 1400.000 1637.360 ;
        RECT 1407.665 1637.250 1407.995 1637.265 ;
        RECT 1396.000 1636.950 1407.995 1637.250 ;
        RECT 1396.000 1636.760 1400.000 1636.950 ;
        RECT 1407.665 1636.935 1407.995 1636.950 ;
      LAYER met3 ;
        RECT 300.065 1634.360 1396.000 1636.360 ;
      LAYER met3 ;
        RECT 300.000 1633.360 304.000 1633.960 ;
      LAYER met3 ;
        RECT 304.400 1633.000 1396.000 1634.360 ;
        RECT 304.400 1632.960 1395.600 1633.000 ;
        RECT 300.065 1631.600 1395.600 1632.960 ;
      LAYER met3 ;
        RECT 1396.000 1632.490 1400.000 1632.600 ;
        RECT 1411.805 1632.490 1412.135 1632.505 ;
        RECT 1396.000 1632.190 1412.135 1632.490 ;
        RECT 1396.000 1632.000 1400.000 1632.190 ;
        RECT 1411.805 1632.175 1412.135 1632.190 ;
      LAYER met3 ;
        RECT 300.065 1628.240 1396.000 1631.600 ;
        RECT 300.065 1626.840 1395.600 1628.240 ;
      LAYER met3 ;
        RECT 1396.000 1627.730 1400.000 1627.840 ;
        RECT 1407.665 1627.730 1407.995 1627.745 ;
        RECT 1396.000 1627.430 1407.995 1627.730 ;
        RECT 1396.000 1627.240 1400.000 1627.430 ;
        RECT 1407.665 1627.415 1407.995 1627.430 ;
      LAYER met3 ;
        RECT 300.065 1624.840 1396.000 1626.840 ;
      LAYER met3 ;
        RECT 300.000 1623.840 304.000 1624.440 ;
      LAYER met3 ;
        RECT 304.400 1623.440 1396.000 1624.840 ;
        RECT 300.065 1622.800 1396.000 1623.440 ;
        RECT 300.065 1621.400 1395.600 1622.800 ;
      LAYER met3 ;
        RECT 1396.000 1622.290 1400.000 1622.400 ;
        RECT 1417.070 1622.290 1417.450 1622.300 ;
        RECT 1396.000 1621.990 1417.450 1622.290 ;
        RECT 1396.000 1621.800 1400.000 1621.990 ;
        RECT 1417.070 1621.980 1417.450 1621.990 ;
      LAYER met3 ;
        RECT 300.065 1618.040 1396.000 1621.400 ;
        RECT 300.065 1616.640 1395.600 1618.040 ;
      LAYER met3 ;
        RECT 1396.000 1617.530 1400.000 1617.640 ;
        RECT 1411.550 1617.530 1411.930 1617.540 ;
        RECT 1396.000 1617.230 1411.930 1617.530 ;
        RECT 1396.000 1617.040 1400.000 1617.230 ;
        RECT 1411.550 1617.220 1411.930 1617.230 ;
      LAYER met3 ;
        RECT 300.065 1615.320 1396.000 1616.640 ;
      LAYER met3 ;
        RECT 300.000 1614.320 304.000 1614.920 ;
      LAYER met3 ;
        RECT 304.400 1613.920 1396.000 1615.320 ;
        RECT 300.065 1612.600 1396.000 1613.920 ;
        RECT 300.065 1611.200 1395.600 1612.600 ;
      LAYER met3 ;
        RECT 1396.000 1612.090 1400.000 1612.200 ;
        RECT 1408.585 1612.090 1408.915 1612.105 ;
        RECT 1396.000 1611.790 1408.915 1612.090 ;
        RECT 1396.000 1611.600 1400.000 1611.790 ;
        RECT 1408.585 1611.775 1408.915 1611.790 ;
      LAYER met3 ;
        RECT 300.065 1607.840 1396.000 1611.200 ;
        RECT 300.065 1606.440 1395.600 1607.840 ;
      LAYER met3 ;
        RECT 1700.000 1607.670 1704.600 1607.970 ;
        RECT 1396.000 1607.330 1400.000 1607.440 ;
        RECT 1414.105 1607.330 1414.435 1607.345 ;
        RECT 1396.000 1607.030 1414.435 1607.330 ;
        RECT 1396.000 1606.840 1400.000 1607.030 ;
        RECT 1414.105 1607.015 1414.435 1607.030 ;
      LAYER met3 ;
        RECT 300.065 1605.800 1396.000 1606.440 ;
      LAYER met3 ;
        RECT 300.000 1604.800 304.000 1605.400 ;
      LAYER met3 ;
        RECT 304.400 1604.400 1396.000 1605.800 ;
        RECT 1705.000 1605.000 2081.480 2051.235 ;
      LAYER met3 ;
        RECT 2250.000 2032.785 2254.600 2033.085 ;
        RECT 2250.000 2027.145 2254.600 2027.445 ;
        RECT 2250.000 2018.645 2254.600 2018.945 ;
        RECT 2250.000 2013.005 2254.600 2013.305 ;
        RECT 2250.000 2004.505 2254.600 2004.805 ;
        RECT 2250.000 1998.865 2254.600 1999.165 ;
        RECT 2250.000 1990.365 2254.600 1990.665 ;
        RECT 2083.865 1965.010 2084.195 1965.025 ;
        RECT 2083.865 1964.695 2084.410 1965.010 ;
        RECT 2084.110 1963.610 2084.410 1964.695 ;
        RECT 2081.880 1963.310 2086.480 1963.610 ;
        RECT 2082.025 1956.850 2082.355 1956.865 ;
        RECT 2082.025 1956.535 2082.570 1956.850 ;
        RECT 2082.270 1955.110 2082.570 1956.535 ;
        RECT 2081.880 1954.810 2086.480 1955.110 ;
        RECT 2100.425 1746.050 2100.755 1746.065 ;
        RECT 2103.390 1746.050 2103.770 1746.060 ;
        RECT 2100.425 1745.750 2103.770 1746.050 ;
        RECT 2100.425 1745.735 2100.755 1745.750 ;
        RECT 2103.390 1745.740 2103.770 1745.750 ;
        RECT 2099.505 1733.140 2099.835 1733.145 ;
        RECT 2099.505 1733.130 2100.090 1733.140 ;
        RECT 2099.505 1732.830 2100.290 1733.130 ;
        RECT 2099.505 1732.820 2100.090 1732.830 ;
        RECT 2099.505 1732.815 2099.835 1732.820 ;
        RECT 2099.965 1732.450 2100.295 1732.465 ;
        RECT 2103.390 1732.450 2103.770 1732.460 ;
        RECT 2099.965 1732.150 2103.770 1732.450 ;
        RECT 2099.965 1732.135 2100.295 1732.150 ;
        RECT 2103.390 1732.140 2103.770 1732.150 ;
        RECT 2114.430 1732.450 2114.810 1732.460 ;
        RECT 2139.270 1732.450 2139.650 1732.460 ;
        RECT 2114.430 1732.150 2139.650 1732.450 ;
        RECT 2114.430 1732.140 2114.810 1732.150 ;
        RECT 2139.270 1732.140 2139.650 1732.150 ;
        RECT 2234.030 1732.450 2234.410 1732.460 ;
        RECT 2238.630 1732.450 2239.010 1732.460 ;
        RECT 2234.030 1732.150 2239.010 1732.450 ;
        RECT 2234.030 1732.140 2234.410 1732.150 ;
        RECT 2238.630 1732.140 2239.010 1732.150 ;
        RECT 2189.870 1729.050 2190.250 1729.060 ;
        RECT 2235.870 1729.050 2236.250 1729.060 ;
        RECT 2189.870 1728.750 2236.250 1729.050 ;
        RECT 2189.870 1728.740 2190.250 1728.750 ;
        RECT 2235.870 1728.740 2236.250 1728.750 ;
        RECT 2099.045 1722.250 2099.375 1722.265 ;
        RECT 2188.950 1722.250 2189.330 1722.260 ;
        RECT 2099.045 1721.950 2189.330 1722.250 ;
        RECT 2099.045 1721.935 2099.375 1721.950 ;
        RECT 2188.950 1721.940 2189.330 1721.950 ;
        RECT 2098.585 1718.850 2098.915 1718.865 ;
        RECT 2103.390 1718.850 2103.770 1718.860 ;
        RECT 2098.585 1718.550 2103.770 1718.850 ;
        RECT 2098.585 1718.535 2098.915 1718.550 ;
        RECT 2103.390 1718.540 2103.770 1718.550 ;
        RECT 2188.030 1715.450 2188.410 1715.460 ;
        RECT 2240.470 1715.450 2240.850 1715.460 ;
        RECT 2188.030 1715.150 2240.850 1715.450 ;
        RECT 2188.030 1715.140 2188.410 1715.150 ;
        RECT 2240.470 1715.140 2240.850 1715.150 ;
        RECT 2247.830 1715.450 2248.210 1715.460 ;
        RECT 2253.350 1715.450 2253.730 1715.460 ;
        RECT 2247.830 1715.150 2253.730 1715.450 ;
        RECT 2247.830 1715.140 2248.210 1715.150 ;
        RECT 2253.350 1715.140 2253.730 1715.150 ;
        RECT 2098.125 1708.650 2098.455 1708.665 ;
        RECT 2102.470 1708.650 2102.850 1708.660 ;
        RECT 2098.125 1708.350 2102.850 1708.650 ;
        RECT 2098.125 1708.335 2098.455 1708.350 ;
        RECT 2102.470 1708.340 2102.850 1708.350 ;
        RECT 2139.270 1705.930 2139.650 1705.940 ;
        RECT 2197.230 1705.930 2197.610 1705.940 ;
        RECT 2139.270 1705.630 2197.610 1705.930 ;
        RECT 2139.270 1705.620 2139.650 1705.630 ;
        RECT 2197.230 1705.620 2197.610 1705.630 ;
        RECT 2097.665 1705.250 2097.995 1705.265 ;
        RECT 2102.470 1705.250 2102.850 1705.260 ;
        RECT 2097.665 1704.950 2102.850 1705.250 ;
        RECT 2097.665 1704.935 2097.995 1704.950 ;
        RECT 2102.470 1704.940 2102.850 1704.950 ;
        RECT 2222.070 1701.850 2222.450 1701.860 ;
        RECT 2227.590 1701.850 2227.970 1701.860 ;
        RECT 2222.070 1701.550 2227.970 1701.850 ;
        RECT 2222.070 1701.540 2222.450 1701.550 ;
        RECT 2227.590 1701.540 2227.970 1701.550 ;
        RECT 2250.000 1701.125 2254.600 1701.425 ;
        RECT 2250.000 1692.625 2254.600 1692.925 ;
        RECT 2100.425 1668.530 2100.755 1668.545 ;
        RECT 2085.950 1668.230 2100.755 1668.530 ;
        RECT 2085.950 1665.870 2086.250 1668.230 ;
        RECT 2100.425 1668.215 2100.755 1668.230 ;
        RECT 2081.880 1665.570 2086.480 1665.870 ;
        RECT 2099.965 1660.370 2100.295 1660.385 ;
        RECT 2085.950 1660.070 2100.295 1660.370 ;
        RECT 2085.950 1657.370 2086.250 1660.070 ;
        RECT 2099.965 1660.055 2100.295 1660.070 ;
        RECT 2081.880 1657.070 2086.480 1657.370 ;
        RECT 2099.505 1654.930 2099.835 1654.945 ;
        RECT 2085.950 1654.630 2099.835 1654.930 ;
        RECT 2085.950 1651.730 2086.250 1654.630 ;
        RECT 2099.505 1654.615 2099.835 1654.630 ;
        RECT 2081.880 1651.430 2086.480 1651.730 ;
        RECT 2099.045 1646.090 2099.375 1646.105 ;
        RECT 2085.950 1645.790 2099.375 1646.090 ;
        RECT 2085.950 1643.230 2086.250 1645.790 ;
        RECT 2099.045 1645.775 2099.375 1645.790 ;
        RECT 2081.880 1642.930 2086.480 1643.230 ;
        RECT 2098.585 1640.650 2098.915 1640.665 ;
        RECT 2085.950 1640.350 2098.915 1640.650 ;
        RECT 2085.950 1637.590 2086.250 1640.350 ;
        RECT 2098.585 1640.335 2098.915 1640.350 ;
        RECT 2081.880 1637.290 2086.480 1637.590 ;
        RECT 2098.125 1629.090 2098.455 1629.105 ;
        RECT 2081.880 1628.790 2098.455 1629.090 ;
        RECT 2098.125 1628.775 2098.455 1628.790 ;
        RECT 2097.665 1625.690 2097.995 1625.705 ;
        RECT 2085.950 1625.390 2097.995 1625.690 ;
        RECT 2085.950 1623.450 2086.250 1625.390 ;
        RECT 2097.665 1625.375 2097.995 1625.390 ;
        RECT 2081.880 1623.150 2086.480 1623.450 ;
      LAYER met3 ;
        RECT 2255.000 1605.000 2631.480 2051.235 ;
      LAYER met3 ;
        RECT 2632.185 2050.010 2632.515 2050.025 ;
        RECT 2632.185 2049.695 2632.730 2050.010 ;
        RECT 2632.430 2048.565 2632.730 2049.695 ;
        RECT 2631.880 2048.265 2636.480 2048.565 ;
        RECT 2631.880 1746.910 2636.480 1747.210 ;
        RECT 2636.110 1746.050 2636.410 1746.910 ;
        RECT 2637.910 1746.050 2638.290 1746.060 ;
        RECT 2636.110 1745.750 2638.290 1746.050 ;
        RECT 2637.910 1745.740 2638.290 1745.750 ;
        RECT 2631.880 1738.410 2636.480 1738.710 ;
        RECT 2636.110 1735.850 2636.410 1738.410 ;
        RECT 2639.750 1735.850 2640.130 1735.860 ;
        RECT 2636.110 1735.550 2640.130 1735.850 ;
        RECT 2639.750 1735.540 2640.130 1735.550 ;
        RECT 2631.880 1732.770 2636.480 1733.070 ;
        RECT 2636.110 1732.450 2636.410 1732.770 ;
        RECT 2637.910 1732.450 2638.290 1732.460 ;
        RECT 2636.110 1732.150 2638.290 1732.450 ;
        RECT 2637.910 1732.140 2638.290 1732.150 ;
        RECT 2637.910 1724.570 2638.290 1724.580 ;
        RECT 2631.880 1724.270 2638.290 1724.570 ;
        RECT 2637.910 1724.260 2638.290 1724.270 ;
        RECT 2631.880 1718.630 2636.480 1718.930 ;
        RECT 2636.110 1716.130 2636.410 1718.630 ;
        RECT 2639.750 1716.130 2640.130 1716.140 ;
        RECT 2636.110 1715.830 2640.130 1716.130 ;
        RECT 2639.750 1715.820 2640.130 1715.830 ;
        RECT 2631.880 1710.130 2636.480 1710.430 ;
        RECT 2636.110 1708.650 2636.410 1710.130 ;
        RECT 2637.910 1710.010 2638.290 1710.020 ;
        RECT 2637.910 1709.710 2639.170 1710.010 ;
        RECT 2637.910 1709.700 2638.290 1709.710 ;
        RECT 2637.910 1708.650 2638.290 1708.660 ;
        RECT 2636.110 1708.350 2638.290 1708.650 ;
        RECT 2637.910 1708.340 2638.290 1708.350 ;
        RECT 2638.870 1707.970 2639.170 1709.710 ;
        RECT 2636.110 1707.670 2639.170 1707.970 ;
        RECT 2636.110 1704.790 2636.410 1707.670 ;
        RECT 2631.880 1704.490 2636.480 1704.790 ;
      LAYER met3 ;
        RECT 300.065 1603.080 1396.000 1604.400 ;
      LAYER met3 ;
        RECT 1396.625 1604.610 1396.955 1604.625 ;
        RECT 1396.625 1604.295 1397.170 1604.610 ;
      LAYER met3 ;
        RECT 300.065 1602.215 1395.600 1603.080 ;
      LAYER met3 ;
        RECT 1396.870 1602.680 1397.170 1604.295 ;
        RECT 1725.460 1604.095 1727.200 1605.000 ;
        RECT 1396.000 1602.080 1400.000 1602.680 ;
      LAYER met3 ;
        RECT 1550.065 1496.480 2645.600 1497.340 ;
      LAYER met3 ;
        RECT 2646.000 1496.880 2650.000 1497.480 ;
      LAYER met3 ;
        RECT 1550.065 1495.840 2646.000 1496.480 ;
      LAYER met3 ;
        RECT 1550.000 1494.840 1554.000 1495.440 ;
      LAYER met3 ;
        RECT 1554.400 1494.440 2646.000 1495.840 ;
        RECT 1550.065 1493.120 2646.000 1494.440 ;
        RECT 1550.065 1491.720 2645.600 1493.120 ;
      LAYER met3 ;
        RECT 2646.000 1492.120 2650.000 1492.720 ;
      LAYER met3 ;
        RECT 1550.065 1487.680 2646.000 1491.720 ;
        RECT 1550.065 1486.320 2645.600 1487.680 ;
      LAYER met3 ;
        RECT 2646.000 1486.680 2650.000 1487.280 ;
      LAYER met3 ;
        RECT 1554.400 1486.280 2645.600 1486.320 ;
      LAYER met3 ;
        RECT 1550.000 1485.320 1554.000 1485.920 ;
      LAYER met3 ;
        RECT 1554.400 1484.920 2646.000 1486.280 ;
        RECT 1550.065 1482.920 2646.000 1484.920 ;
        RECT 1550.065 1481.520 2645.600 1482.920 ;
      LAYER met3 ;
        RECT 2646.000 1481.920 2650.000 1482.520 ;
      LAYER met3 ;
        RECT 1550.065 1477.480 2646.000 1481.520 ;
        RECT 1550.065 1476.800 2645.600 1477.480 ;
      LAYER met3 ;
        RECT 1550.000 1475.800 1554.000 1476.400 ;
      LAYER met3 ;
        RECT 1554.400 1476.080 2645.600 1476.800 ;
      LAYER met3 ;
        RECT 2646.000 1476.480 2650.000 1477.080 ;
      LAYER met3 ;
        RECT 1554.400 1475.400 2646.000 1476.080 ;
        RECT 1550.065 1472.720 2646.000 1475.400 ;
        RECT 1550.065 1471.320 2645.600 1472.720 ;
      LAYER met3 ;
        RECT 2646.000 1471.720 2650.000 1472.320 ;
      LAYER met3 ;
        RECT 1550.065 1467.960 2646.000 1471.320 ;
        RECT 1550.065 1467.280 2645.600 1467.960 ;
      LAYER met3 ;
        RECT 1550.000 1466.280 1554.000 1466.880 ;
      LAYER met3 ;
        RECT 1554.400 1466.560 2645.600 1467.280 ;
      LAYER met3 ;
        RECT 2646.000 1466.960 2650.000 1467.560 ;
      LAYER met3 ;
        RECT 1554.400 1465.880 2646.000 1466.560 ;
        RECT 1550.065 1462.520 2646.000 1465.880 ;
        RECT 1550.065 1461.120 2645.600 1462.520 ;
      LAYER met3 ;
        RECT 2646.000 1461.520 2650.000 1462.120 ;
      LAYER met3 ;
        RECT 1550.065 1457.760 2646.000 1461.120 ;
      LAYER met3 ;
        RECT 1550.000 1456.760 1554.000 1457.360 ;
      LAYER met3 ;
        RECT 1554.400 1456.360 2645.600 1457.760 ;
      LAYER met3 ;
        RECT 2646.000 1456.760 2650.000 1457.360 ;
      LAYER met3 ;
        RECT 1550.065 1452.320 2646.000 1456.360 ;
        RECT 1550.065 1450.920 2645.600 1452.320 ;
      LAYER met3 ;
        RECT 2646.000 1451.320 2650.000 1451.920 ;
      LAYER met3 ;
        RECT 1550.065 1447.560 2646.000 1450.920 ;
      LAYER met3 ;
        RECT 1550.000 1446.560 1554.000 1447.160 ;
      LAYER met3 ;
        RECT 1554.400 1446.160 2645.600 1447.560 ;
      LAYER met3 ;
        RECT 2646.000 1446.560 2650.000 1447.160 ;
      LAYER met3 ;
        RECT 1550.065 1442.120 2646.000 1446.160 ;
        RECT 1550.065 1440.720 2645.600 1442.120 ;
      LAYER met3 ;
        RECT 2646.000 1441.120 2650.000 1441.720 ;
      LAYER met3 ;
        RECT 1550.065 1438.040 2646.000 1440.720 ;
      LAYER met3 ;
        RECT 1550.000 1437.040 1554.000 1437.640 ;
      LAYER met3 ;
        RECT 1554.400 1437.360 2646.000 1438.040 ;
        RECT 1554.400 1436.640 2645.600 1437.360 ;
        RECT 1550.065 1435.960 2645.600 1436.640 ;
      LAYER met3 ;
        RECT 2646.000 1436.360 2650.000 1436.960 ;
      LAYER met3 ;
        RECT 1550.065 1432.600 2646.000 1435.960 ;
        RECT 1550.065 1431.200 2645.600 1432.600 ;
      LAYER met3 ;
        RECT 2646.000 1431.600 2650.000 1432.200 ;
      LAYER met3 ;
        RECT 1550.065 1428.520 2646.000 1431.200 ;
      LAYER met3 ;
        RECT 1550.000 1427.520 1554.000 1428.120 ;
      LAYER met3 ;
        RECT 1554.400 1427.160 2646.000 1428.520 ;
        RECT 1554.400 1427.120 2645.600 1427.160 ;
        RECT 1550.065 1425.760 2645.600 1427.120 ;
      LAYER met3 ;
        RECT 2646.000 1426.160 2650.000 1426.760 ;
      LAYER met3 ;
        RECT 1550.065 1422.400 2646.000 1425.760 ;
        RECT 1550.065 1421.000 2645.600 1422.400 ;
      LAYER met3 ;
        RECT 2646.000 1421.400 2650.000 1422.000 ;
      LAYER met3 ;
        RECT 1550.065 1419.000 2646.000 1421.000 ;
      LAYER met3 ;
        RECT 1550.000 1418.000 1554.000 1418.600 ;
      LAYER met3 ;
        RECT 1554.400 1417.600 2646.000 1419.000 ;
        RECT 1550.065 1416.960 2646.000 1417.600 ;
        RECT 1550.065 1415.560 2645.600 1416.960 ;
      LAYER met3 ;
        RECT 2646.000 1415.960 2650.000 1416.560 ;
      LAYER met3 ;
        RECT 1550.065 1412.200 2646.000 1415.560 ;
        RECT 1550.065 1410.800 2645.600 1412.200 ;
      LAYER met3 ;
        RECT 2646.000 1411.200 2650.000 1411.800 ;
      LAYER met3 ;
        RECT 1550.065 1409.480 2646.000 1410.800 ;
      LAYER met3 ;
        RECT 1550.000 1408.480 1554.000 1409.080 ;
      LAYER met3 ;
        RECT 1554.400 1408.080 2646.000 1409.480 ;
        RECT 1550.065 1406.760 2646.000 1408.080 ;
        RECT 1550.065 1405.360 2645.600 1406.760 ;
      LAYER met3 ;
        RECT 2646.000 1405.760 2650.000 1406.360 ;
      LAYER met3 ;
        RECT 1550.065 1402.000 2646.000 1405.360 ;
        RECT 1550.065 1400.600 2645.600 1402.000 ;
      LAYER met3 ;
        RECT 2646.000 1401.000 2650.000 1401.600 ;
      LAYER met3 ;
        RECT 1550.065 1399.280 2646.000 1400.600 ;
      LAYER met3 ;
        RECT 1550.000 1398.280 1554.000 1398.880 ;
      LAYER met3 ;
        RECT 1554.400 1397.880 2646.000 1399.280 ;
        RECT 1550.065 1397.240 2646.000 1397.880 ;
        RECT 1550.065 1395.840 2645.600 1397.240 ;
      LAYER met3 ;
        RECT 2646.000 1396.240 2650.000 1396.840 ;
      LAYER met3 ;
        RECT 1550.065 1391.800 2646.000 1395.840 ;
        RECT 1550.065 1390.400 2645.600 1391.800 ;
      LAYER met3 ;
        RECT 2646.000 1390.800 2650.000 1391.400 ;
      LAYER met3 ;
        RECT 1550.065 1389.760 2646.000 1390.400 ;
      LAYER met3 ;
        RECT 1550.000 1388.760 1554.000 1389.360 ;
      LAYER met3 ;
        RECT 1554.400 1388.360 2646.000 1389.760 ;
        RECT 1550.065 1387.040 2646.000 1388.360 ;
        RECT 1550.065 1385.640 2645.600 1387.040 ;
      LAYER met3 ;
        RECT 2646.000 1386.040 2650.000 1386.640 ;
      LAYER met3 ;
        RECT 1550.065 1381.600 2646.000 1385.640 ;
        RECT 1550.065 1380.240 2645.600 1381.600 ;
      LAYER met3 ;
        RECT 2646.000 1380.600 2650.000 1381.200 ;
      LAYER met3 ;
        RECT 1554.400 1380.200 2645.600 1380.240 ;
      LAYER met3 ;
        RECT 1550.000 1379.240 1554.000 1379.840 ;
      LAYER met3 ;
        RECT 1554.400 1378.840 2646.000 1380.200 ;
        RECT 1550.065 1376.840 2646.000 1378.840 ;
        RECT 1550.065 1375.440 2645.600 1376.840 ;
      LAYER met3 ;
        RECT 2646.000 1375.840 2650.000 1376.440 ;
      LAYER met3 ;
        RECT 1550.065 1372.080 2646.000 1375.440 ;
        RECT 1550.065 1370.720 2645.600 1372.080 ;
      LAYER met3 ;
        RECT 2646.000 1371.080 2650.000 1371.680 ;
      LAYER met3 ;
        RECT 1554.400 1370.680 2645.600 1370.720 ;
      LAYER met3 ;
        RECT 1550.000 1369.720 1554.000 1370.320 ;
      LAYER met3 ;
        RECT 1554.400 1369.320 2646.000 1370.680 ;
        RECT 1550.065 1366.640 2646.000 1369.320 ;
        RECT 1550.065 1365.240 2645.600 1366.640 ;
      LAYER met3 ;
        RECT 2646.000 1365.640 2650.000 1366.240 ;
      LAYER met3 ;
        RECT 1550.065 1361.880 2646.000 1365.240 ;
        RECT 1550.065 1361.200 2645.600 1361.880 ;
      LAYER met3 ;
        RECT 1550.000 1360.200 1554.000 1360.800 ;
      LAYER met3 ;
        RECT 1554.400 1360.480 2645.600 1361.200 ;
      LAYER met3 ;
        RECT 2646.000 1360.880 2650.000 1361.480 ;
      LAYER met3 ;
        RECT 1554.400 1359.800 2646.000 1360.480 ;
        RECT 1550.065 1356.440 2646.000 1359.800 ;
        RECT 1550.065 1355.040 2645.600 1356.440 ;
      LAYER met3 ;
        RECT 2646.000 1355.440 2650.000 1356.040 ;
      LAYER met3 ;
        RECT 1550.065 1351.680 2646.000 1355.040 ;
        RECT 1550.065 1351.000 2645.600 1351.680 ;
      LAYER met3 ;
        RECT 1550.000 1350.000 1554.000 1350.600 ;
      LAYER met3 ;
        RECT 1554.400 1350.280 2645.600 1351.000 ;
      LAYER met3 ;
        RECT 2646.000 1350.680 2650.000 1351.280 ;
      LAYER met3 ;
        RECT 1554.400 1349.600 2646.000 1350.280 ;
        RECT 1550.065 1346.240 2646.000 1349.600 ;
        RECT 1550.065 1344.840 2645.600 1346.240 ;
      LAYER met3 ;
        RECT 2646.000 1345.240 2650.000 1345.840 ;
      LAYER met3 ;
        RECT 1550.065 1341.480 2646.000 1344.840 ;
      LAYER met3 ;
        RECT 1550.000 1340.480 1554.000 1341.080 ;
      LAYER met3 ;
        RECT 1554.400 1340.080 2645.600 1341.480 ;
      LAYER met3 ;
        RECT 2646.000 1340.480 2650.000 1341.080 ;
      LAYER met3 ;
        RECT 1550.065 1336.720 2646.000 1340.080 ;
        RECT 1550.065 1335.320 2645.600 1336.720 ;
      LAYER met3 ;
        RECT 2646.000 1335.720 2650.000 1336.320 ;
      LAYER met3 ;
        RECT 1550.065 1331.960 2646.000 1335.320 ;
      LAYER met3 ;
        RECT 1550.000 1330.960 1554.000 1331.560 ;
      LAYER met3 ;
        RECT 1554.400 1331.280 2646.000 1331.960 ;
        RECT 1554.400 1330.560 2645.600 1331.280 ;
        RECT 1550.065 1329.880 2645.600 1330.560 ;
      LAYER met3 ;
        RECT 2646.000 1330.280 2650.000 1330.880 ;
      LAYER met3 ;
        RECT 1550.065 1326.520 2646.000 1329.880 ;
        RECT 1550.065 1325.120 2645.600 1326.520 ;
      LAYER met3 ;
        RECT 2646.000 1325.520 2650.000 1326.120 ;
      LAYER met3 ;
        RECT 1550.065 1322.440 2646.000 1325.120 ;
      LAYER met3 ;
        RECT 1550.000 1321.440 1554.000 1322.040 ;
      LAYER met3 ;
        RECT 1554.400 1321.080 2646.000 1322.440 ;
        RECT 1554.400 1321.040 2645.600 1321.080 ;
        RECT 1550.065 1319.680 2645.600 1321.040 ;
      LAYER met3 ;
        RECT 2646.000 1320.080 2650.000 1320.680 ;
      LAYER met3 ;
        RECT 1550.065 1316.320 2646.000 1319.680 ;
        RECT 1550.065 1314.920 2645.600 1316.320 ;
      LAYER met3 ;
        RECT 2646.000 1315.320 2650.000 1315.920 ;
      LAYER met3 ;
        RECT 1550.065 1312.920 2646.000 1314.920 ;
      LAYER met3 ;
        RECT 1550.000 1311.920 1554.000 1312.520 ;
      LAYER met3 ;
        RECT 1554.400 1311.520 2646.000 1312.920 ;
        RECT 1550.065 1310.880 2646.000 1311.520 ;
        RECT 1550.065 1309.480 2645.600 1310.880 ;
      LAYER met3 ;
        RECT 2646.000 1309.880 2650.000 1310.480 ;
      LAYER met3 ;
        RECT 1550.065 1306.120 2646.000 1309.480 ;
        RECT 1550.065 1304.720 2645.600 1306.120 ;
      LAYER met3 ;
        RECT 2646.000 1305.120 2650.000 1305.720 ;
      LAYER met3 ;
        RECT 1550.065 1302.720 2646.000 1304.720 ;
      LAYER met3 ;
        RECT 1550.000 1301.720 1554.000 1302.320 ;
      LAYER met3 ;
        RECT 1554.400 1301.360 2646.000 1302.720 ;
        RECT 1554.400 1301.320 2645.600 1301.360 ;
        RECT 1550.065 1299.960 2645.600 1301.320 ;
      LAYER met3 ;
        RECT 2646.000 1300.360 2650.000 1300.960 ;
      LAYER met3 ;
        RECT 1550.065 1295.920 2646.000 1299.960 ;
        RECT 1550.065 1294.520 2645.600 1295.920 ;
      LAYER met3 ;
        RECT 2646.000 1294.920 2650.000 1295.520 ;
      LAYER met3 ;
        RECT 1550.065 1293.200 2646.000 1294.520 ;
      LAYER met3 ;
        RECT 1550.000 1292.200 1554.000 1292.800 ;
      LAYER met3 ;
        RECT 1554.400 1291.800 2646.000 1293.200 ;
        RECT 1550.065 1291.160 2646.000 1291.800 ;
        RECT 1550.065 1289.760 2645.600 1291.160 ;
      LAYER met3 ;
        RECT 2646.000 1290.160 2650.000 1290.760 ;
      LAYER met3 ;
        RECT 1550.065 1285.720 2646.000 1289.760 ;
        RECT 1550.065 1284.320 2645.600 1285.720 ;
      LAYER met3 ;
        RECT 2646.000 1284.720 2650.000 1285.320 ;
      LAYER met3 ;
        RECT 1550.065 1283.680 2646.000 1284.320 ;
      LAYER met3 ;
        RECT 1550.000 1282.680 1554.000 1283.280 ;
      LAYER met3 ;
        RECT 1554.400 1282.280 2646.000 1283.680 ;
        RECT 1550.065 1280.960 2646.000 1282.280 ;
        RECT 1550.065 1279.560 2645.600 1280.960 ;
      LAYER met3 ;
        RECT 2646.000 1279.960 2650.000 1280.560 ;
      LAYER met3 ;
        RECT 1550.065 1276.200 2646.000 1279.560 ;
        RECT 1550.065 1274.800 2645.600 1276.200 ;
      LAYER met3 ;
        RECT 2646.000 1275.200 2650.000 1275.800 ;
      LAYER met3 ;
        RECT 1550.065 1274.160 2646.000 1274.800 ;
      LAYER met3 ;
        RECT 1550.000 1273.160 1554.000 1273.760 ;
      LAYER met3 ;
        RECT 1554.400 1272.760 2646.000 1274.160 ;
        RECT 1550.065 1270.760 2646.000 1272.760 ;
        RECT 1550.065 1269.360 2645.600 1270.760 ;
      LAYER met3 ;
        RECT 2646.000 1269.760 2650.000 1270.360 ;
      LAYER met3 ;
        RECT 1550.065 1266.000 2646.000 1269.360 ;
        RECT 1550.065 1264.640 2645.600 1266.000 ;
      LAYER met3 ;
        RECT 2646.000 1265.000 2650.000 1265.600 ;
      LAYER met3 ;
        RECT 1554.400 1264.600 2645.600 1264.640 ;
      LAYER met3 ;
        RECT 1550.000 1263.640 1554.000 1264.240 ;
      LAYER met3 ;
        RECT 1554.400 1263.240 2646.000 1264.600 ;
        RECT 1550.065 1260.560 2646.000 1263.240 ;
        RECT 1550.065 1259.160 2645.600 1260.560 ;
      LAYER met3 ;
        RECT 2646.000 1259.560 2650.000 1260.160 ;
      LAYER met3 ;
        RECT 1550.065 1255.800 2646.000 1259.160 ;
        RECT 1550.065 1254.440 2645.600 1255.800 ;
      LAYER met3 ;
        RECT 2646.000 1254.800 2650.000 1255.400 ;
      LAYER met3 ;
        RECT 1554.400 1254.400 2645.600 1254.440 ;
      LAYER met3 ;
        RECT 1550.000 1253.440 1554.000 1254.040 ;
      LAYER met3 ;
        RECT 1554.400 1253.040 2646.000 1254.400 ;
        RECT 1550.065 1250.360 2646.000 1253.040 ;
        RECT 1550.065 1248.960 2645.600 1250.360 ;
      LAYER met3 ;
        RECT 2646.000 1249.360 2650.000 1249.960 ;
      LAYER met3 ;
        RECT 1550.065 1245.600 2646.000 1248.960 ;
        RECT 1550.065 1244.920 2645.600 1245.600 ;
      LAYER met3 ;
        RECT 1550.000 1243.920 1554.000 1244.520 ;
      LAYER met3 ;
        RECT 1554.400 1244.200 2645.600 1244.920 ;
      LAYER met3 ;
        RECT 2646.000 1244.600 2650.000 1245.200 ;
      LAYER met3 ;
        RECT 1554.400 1243.520 2646.000 1244.200 ;
        RECT 1550.065 1240.840 2646.000 1243.520 ;
        RECT 1550.065 1239.440 2645.600 1240.840 ;
      LAYER met3 ;
        RECT 2646.000 1239.840 2650.000 1240.440 ;
      LAYER met3 ;
        RECT 1550.065 1235.400 2646.000 1239.440 ;
      LAYER met3 ;
        RECT 1550.000 1234.400 1554.000 1235.000 ;
      LAYER met3 ;
        RECT 1554.400 1234.000 2645.600 1235.400 ;
      LAYER met3 ;
        RECT 2646.000 1234.400 2650.000 1235.000 ;
      LAYER met3 ;
        RECT 1550.065 1230.640 2646.000 1234.000 ;
        RECT 1550.065 1229.240 2645.600 1230.640 ;
      LAYER met3 ;
        RECT 2646.000 1229.640 2650.000 1230.240 ;
      LAYER met3 ;
        RECT 1550.065 1225.880 2646.000 1229.240 ;
      LAYER met3 ;
        RECT 1550.000 1224.880 1554.000 1225.480 ;
      LAYER met3 ;
        RECT 1554.400 1225.200 2646.000 1225.880 ;
        RECT 1554.400 1224.480 2645.600 1225.200 ;
        RECT 1550.065 1223.800 2645.600 1224.480 ;
      LAYER met3 ;
        RECT 2646.000 1224.200 2650.000 1224.800 ;
      LAYER met3 ;
        RECT 1550.065 1220.440 2646.000 1223.800 ;
        RECT 1550.065 1219.040 2645.600 1220.440 ;
      LAYER met3 ;
        RECT 2646.000 1219.440 2650.000 1220.040 ;
      LAYER met3 ;
        RECT 1550.065 1216.360 2646.000 1219.040 ;
      LAYER met3 ;
        RECT 1550.000 1215.360 1554.000 1215.960 ;
      LAYER met3 ;
        RECT 1554.400 1215.000 2646.000 1216.360 ;
        RECT 1554.400 1214.960 2645.600 1215.000 ;
        RECT 1550.065 1213.600 2645.600 1214.960 ;
      LAYER met3 ;
        RECT 2646.000 1214.000 2650.000 1214.600 ;
      LAYER met3 ;
        RECT 1550.065 1210.240 2646.000 1213.600 ;
        RECT 1550.065 1208.840 2645.600 1210.240 ;
      LAYER met3 ;
        RECT 2646.000 1209.240 2650.000 1209.840 ;
      LAYER met3 ;
        RECT 1550.065 1206.840 2646.000 1208.840 ;
      LAYER met3 ;
        RECT 1550.000 1205.840 1554.000 1206.440 ;
      LAYER met3 ;
        RECT 1554.400 1205.480 2646.000 1206.840 ;
        RECT 1554.400 1205.440 2645.600 1205.480 ;
        RECT 1550.065 1204.080 2645.600 1205.440 ;
      LAYER met3 ;
        RECT 2646.000 1204.480 2650.000 1205.080 ;
      LAYER met3 ;
        RECT 1550.065 1200.040 2646.000 1204.080 ;
        RECT 1550.065 1198.640 2645.600 1200.040 ;
      LAYER met3 ;
        RECT 2646.000 1199.040 2650.000 1199.640 ;
      LAYER met3 ;
        RECT 1550.065 1196.640 2646.000 1198.640 ;
      LAYER met3 ;
        RECT 1550.000 1195.640 1554.000 1196.240 ;
      LAYER met3 ;
        RECT 1554.400 1195.280 2646.000 1196.640 ;
        RECT 1554.400 1195.240 2645.600 1195.280 ;
        RECT 1550.065 1193.880 2645.600 1195.240 ;
      LAYER met3 ;
        RECT 2646.000 1194.280 2650.000 1194.880 ;
      LAYER met3 ;
        RECT 1550.065 1189.840 2646.000 1193.880 ;
        RECT 1550.065 1188.440 2645.600 1189.840 ;
      LAYER met3 ;
        RECT 2646.000 1188.840 2650.000 1189.440 ;
      LAYER met3 ;
        RECT 1550.065 1187.120 2646.000 1188.440 ;
      LAYER met3 ;
        RECT 1550.000 1186.120 1554.000 1186.720 ;
      LAYER met3 ;
        RECT 1554.400 1185.720 2646.000 1187.120 ;
        RECT 1550.065 1185.080 2646.000 1185.720 ;
        RECT 1550.065 1183.680 2645.600 1185.080 ;
      LAYER met3 ;
        RECT 2646.000 1184.080 2650.000 1184.680 ;
      LAYER met3 ;
        RECT 1550.065 1179.640 2646.000 1183.680 ;
        RECT 1550.065 1178.240 2645.600 1179.640 ;
      LAYER met3 ;
        RECT 2646.000 1178.640 2650.000 1179.240 ;
      LAYER met3 ;
        RECT 1550.065 1177.600 2646.000 1178.240 ;
      LAYER met3 ;
        RECT 1550.000 1176.600 1554.000 1177.200 ;
      LAYER met3 ;
        RECT 1554.400 1176.200 2646.000 1177.600 ;
        RECT 1550.065 1174.880 2646.000 1176.200 ;
        RECT 1550.065 1173.480 2645.600 1174.880 ;
      LAYER met3 ;
        RECT 2646.000 1173.880 2650.000 1174.480 ;
      LAYER met3 ;
        RECT 1550.065 1170.120 2646.000 1173.480 ;
        RECT 1550.065 1168.720 2645.600 1170.120 ;
      LAYER met3 ;
        RECT 2646.000 1169.120 2650.000 1169.720 ;
      LAYER met3 ;
        RECT 1550.065 1168.080 2646.000 1168.720 ;
      LAYER met3 ;
        RECT 1550.000 1167.080 1554.000 1167.680 ;
      LAYER met3 ;
        RECT 1554.400 1166.680 2646.000 1168.080 ;
        RECT 1550.065 1164.680 2646.000 1166.680 ;
        RECT 1550.065 1163.280 2645.600 1164.680 ;
      LAYER met3 ;
        RECT 2646.000 1163.680 2650.000 1164.280 ;
      LAYER met3 ;
        RECT 1550.065 1159.920 2646.000 1163.280 ;
        RECT 1550.065 1158.560 2645.600 1159.920 ;
      LAYER met3 ;
        RECT 2646.000 1158.920 2650.000 1159.520 ;
      LAYER met3 ;
        RECT 1554.400 1158.520 2645.600 1158.560 ;
      LAYER met3 ;
        RECT 1550.000 1157.560 1554.000 1158.160 ;
      LAYER met3 ;
        RECT 1554.400 1157.160 2646.000 1158.520 ;
        RECT 1550.065 1154.480 2646.000 1157.160 ;
        RECT 1550.065 1153.080 2645.600 1154.480 ;
      LAYER met3 ;
        RECT 2646.000 1153.480 2650.000 1154.080 ;
      LAYER met3 ;
        RECT 1550.065 1149.720 2646.000 1153.080 ;
        RECT 1550.065 1148.360 2645.600 1149.720 ;
      LAYER met3 ;
        RECT 2646.000 1148.720 2650.000 1149.320 ;
      LAYER met3 ;
        RECT 1554.400 1148.320 2645.600 1148.360 ;
      LAYER met3 ;
        RECT 1550.000 1147.360 1554.000 1147.960 ;
      LAYER met3 ;
        RECT 1554.400 1146.960 2646.000 1148.320 ;
        RECT 1550.065 1144.960 2646.000 1146.960 ;
        RECT 1550.065 1143.560 2645.600 1144.960 ;
      LAYER met3 ;
        RECT 2646.000 1143.960 2650.000 1144.560 ;
      LAYER met3 ;
        RECT 1550.065 1139.520 2646.000 1143.560 ;
        RECT 1550.065 1138.840 2645.600 1139.520 ;
      LAYER met3 ;
        RECT 1550.000 1137.840 1554.000 1138.440 ;
      LAYER met3 ;
        RECT 1554.400 1138.120 2645.600 1138.840 ;
      LAYER met3 ;
        RECT 2646.000 1138.520 2650.000 1139.120 ;
      LAYER met3 ;
        RECT 1554.400 1137.440 2646.000 1138.120 ;
        RECT 1550.065 1134.760 2646.000 1137.440 ;
        RECT 1550.065 1133.360 2645.600 1134.760 ;
      LAYER met3 ;
        RECT 2646.000 1133.760 2650.000 1134.360 ;
      LAYER met3 ;
        RECT 1550.065 1129.320 2646.000 1133.360 ;
      LAYER met3 ;
        RECT 1550.000 1128.320 1554.000 1128.920 ;
      LAYER met3 ;
        RECT 1554.400 1127.920 2645.600 1129.320 ;
      LAYER met3 ;
        RECT 2646.000 1128.320 2650.000 1128.920 ;
      LAYER met3 ;
        RECT 1550.065 1124.560 2646.000 1127.920 ;
        RECT 1550.065 1123.160 2645.600 1124.560 ;
      LAYER met3 ;
        RECT 2646.000 1123.560 2650.000 1124.160 ;
      LAYER met3 ;
        RECT 1550.065 1119.800 2646.000 1123.160 ;
      LAYER met3 ;
        RECT 1550.000 1118.800 1554.000 1119.400 ;
      LAYER met3 ;
        RECT 1554.400 1119.120 2646.000 1119.800 ;
        RECT 1554.400 1118.400 2645.600 1119.120 ;
        RECT 1550.065 1117.720 2645.600 1118.400 ;
      LAYER met3 ;
        RECT 2646.000 1118.120 2650.000 1118.720 ;
      LAYER met3 ;
        RECT 1550.065 1114.360 2646.000 1117.720 ;
        RECT 1550.065 1112.960 2645.600 1114.360 ;
      LAYER met3 ;
        RECT 2646.000 1113.360 2650.000 1113.960 ;
      LAYER met3 ;
        RECT 1550.065 1110.280 2646.000 1112.960 ;
      LAYER met3 ;
        RECT 1550.000 1109.280 1554.000 1109.880 ;
      LAYER met3 ;
        RECT 1554.400 1109.600 2646.000 1110.280 ;
        RECT 1554.400 1108.880 2645.600 1109.600 ;
        RECT 1550.065 1108.200 2645.600 1108.880 ;
      LAYER met3 ;
        RECT 2646.000 1108.600 2650.000 1109.200 ;
      LAYER met3 ;
        RECT 1550.065 1104.160 2646.000 1108.200 ;
        RECT 1550.065 1102.760 2645.600 1104.160 ;
      LAYER met3 ;
        RECT 2646.000 1103.160 2650.000 1103.760 ;
      LAYER met3 ;
        RECT 1550.065 1100.080 2646.000 1102.760 ;
      LAYER met3 ;
        RECT 1550.000 1099.080 1554.000 1099.680 ;
      LAYER met3 ;
        RECT 1554.400 1099.400 2646.000 1100.080 ;
        RECT 1554.400 1098.680 2645.600 1099.400 ;
        RECT 1550.065 1098.000 2645.600 1098.680 ;
      LAYER met3 ;
        RECT 2646.000 1098.400 2650.000 1099.000 ;
      LAYER met3 ;
        RECT 1550.065 1093.960 2646.000 1098.000 ;
        RECT 1550.065 1092.560 2645.600 1093.960 ;
      LAYER met3 ;
        RECT 2646.000 1092.960 2650.000 1093.560 ;
      LAYER met3 ;
        RECT 1550.065 1090.560 2646.000 1092.560 ;
      LAYER met3 ;
        RECT 1550.000 1089.560 1554.000 1090.160 ;
      LAYER met3 ;
        RECT 1554.400 1089.200 2646.000 1090.560 ;
        RECT 1554.400 1089.160 2645.600 1089.200 ;
        RECT 1550.065 1087.800 2645.600 1089.160 ;
      LAYER met3 ;
        RECT 2646.000 1088.200 2650.000 1088.800 ;
      LAYER met3 ;
        RECT 1550.065 1083.760 2646.000 1087.800 ;
        RECT 1550.065 1082.360 2645.600 1083.760 ;
      LAYER met3 ;
        RECT 2646.000 1082.760 2650.000 1083.360 ;
      LAYER met3 ;
        RECT 1550.065 1081.040 2646.000 1082.360 ;
      LAYER met3 ;
        RECT 1550.000 1080.040 1554.000 1080.640 ;
      LAYER met3 ;
        RECT 1554.400 1079.640 2646.000 1081.040 ;
        RECT 1550.065 1079.000 2646.000 1079.640 ;
        RECT 1550.065 1077.600 2645.600 1079.000 ;
      LAYER met3 ;
        RECT 2646.000 1078.000 2650.000 1078.600 ;
      LAYER met3 ;
        RECT 1550.065 1074.240 2646.000 1077.600 ;
        RECT 1550.065 1072.840 2645.600 1074.240 ;
      LAYER met3 ;
        RECT 2646.000 1073.240 2650.000 1073.840 ;
      LAYER met3 ;
        RECT 1550.065 1071.520 2646.000 1072.840 ;
      LAYER met3 ;
        RECT 1550.000 1070.520 1554.000 1071.120 ;
      LAYER met3 ;
        RECT 1554.400 1070.120 2646.000 1071.520 ;
        RECT 1550.065 1068.800 2646.000 1070.120 ;
        RECT 1550.065 1067.400 2645.600 1068.800 ;
      LAYER met3 ;
        RECT 2646.000 1067.800 2650.000 1068.400 ;
      LAYER met3 ;
        RECT 1550.065 1064.040 2646.000 1067.400 ;
        RECT 1550.065 1062.640 2645.600 1064.040 ;
      LAYER met3 ;
        RECT 2646.000 1063.040 2650.000 1063.640 ;
      LAYER met3 ;
        RECT 1550.065 1062.000 2646.000 1062.640 ;
      LAYER met3 ;
        RECT 1550.000 1061.000 1554.000 1061.600 ;
      LAYER met3 ;
        RECT 1554.400 1060.600 2646.000 1062.000 ;
        RECT 1550.065 1058.600 2646.000 1060.600 ;
        RECT 1550.065 1057.200 2645.600 1058.600 ;
      LAYER met3 ;
        RECT 2646.000 1057.600 2650.000 1058.200 ;
      LAYER met3 ;
        RECT 1550.065 1053.840 2646.000 1057.200 ;
        RECT 1550.065 1052.440 2645.600 1053.840 ;
      LAYER met3 ;
        RECT 2646.000 1052.840 2650.000 1053.440 ;
      LAYER met3 ;
        RECT 1550.065 1051.800 2646.000 1052.440 ;
      LAYER met3 ;
        RECT 1550.000 1050.800 1554.000 1051.400 ;
      LAYER met3 ;
        RECT 1554.400 1050.400 2646.000 1051.800 ;
        RECT 1550.065 1049.080 2646.000 1050.400 ;
        RECT 1550.065 1047.680 2645.600 1049.080 ;
      LAYER met3 ;
        RECT 2646.000 1048.080 2650.000 1048.680 ;
      LAYER met3 ;
        RECT 1550.065 1043.640 2646.000 1047.680 ;
        RECT 1550.065 1042.280 2645.600 1043.640 ;
      LAYER met3 ;
        RECT 2646.000 1042.640 2650.000 1043.240 ;
      LAYER met3 ;
        RECT 1554.400 1042.240 2645.600 1042.280 ;
      LAYER met3 ;
        RECT 1550.000 1041.280 1554.000 1041.880 ;
      LAYER met3 ;
        RECT 1554.400 1040.880 2646.000 1042.240 ;
        RECT 1550.065 1038.880 2646.000 1040.880 ;
        RECT 1550.065 1037.480 2645.600 1038.880 ;
      LAYER met3 ;
        RECT 2646.000 1037.880 2650.000 1038.480 ;
      LAYER met3 ;
        RECT 1550.065 1033.440 2646.000 1037.480 ;
        RECT 1550.065 1032.760 2645.600 1033.440 ;
      LAYER met3 ;
        RECT 1550.000 1031.760 1554.000 1032.360 ;
      LAYER met3 ;
        RECT 1554.400 1032.040 2645.600 1032.760 ;
      LAYER met3 ;
        RECT 2646.000 1032.440 2650.000 1033.040 ;
      LAYER met3 ;
        RECT 1554.400 1031.360 2646.000 1032.040 ;
        RECT 1550.065 1028.680 2646.000 1031.360 ;
        RECT 1550.065 1027.280 2645.600 1028.680 ;
      LAYER met3 ;
        RECT 2646.000 1027.680 2650.000 1028.280 ;
      LAYER met3 ;
        RECT 1550.065 1023.240 2646.000 1027.280 ;
      LAYER met3 ;
        RECT 1550.000 1022.240 1554.000 1022.840 ;
      LAYER met3 ;
        RECT 1554.400 1021.840 2645.600 1023.240 ;
      LAYER met3 ;
        RECT 2646.000 1022.240 2650.000 1022.840 ;
      LAYER met3 ;
        RECT 1550.065 1018.480 2646.000 1021.840 ;
        RECT 1550.065 1017.080 2645.600 1018.480 ;
      LAYER met3 ;
        RECT 2646.000 1017.480 2650.000 1018.080 ;
      LAYER met3 ;
        RECT 1550.065 1013.720 2646.000 1017.080 ;
      LAYER met3 ;
        RECT 1550.000 1012.720 1554.000 1013.320 ;
      LAYER met3 ;
        RECT 1554.400 1012.320 2645.600 1013.720 ;
      LAYER met3 ;
        RECT 2646.000 1012.720 2650.000 1013.320 ;
      LAYER met3 ;
        RECT 1550.065 1008.280 2646.000 1012.320 ;
        RECT 1550.065 1006.880 2645.600 1008.280 ;
      LAYER met3 ;
        RECT 2646.000 1007.280 2650.000 1007.880 ;
      LAYER met3 ;
        RECT 1550.065 1003.520 2646.000 1006.880 ;
      LAYER met3 ;
        RECT 1550.000 1002.520 1554.000 1003.120 ;
      LAYER met3 ;
        RECT 1554.400 1002.120 2645.600 1003.520 ;
      LAYER met3 ;
        RECT 2646.000 1002.520 2650.000 1003.120 ;
      LAYER met3 ;
        RECT 1550.065 998.080 2646.000 1002.120 ;
        RECT 1550.065 996.680 2645.600 998.080 ;
      LAYER met3 ;
        RECT 2646.000 997.080 2650.000 997.680 ;
      LAYER met3 ;
        RECT 1550.065 994.000 2646.000 996.680 ;
      LAYER met3 ;
        RECT 1550.000 993.000 1554.000 993.600 ;
      LAYER met3 ;
        RECT 1554.400 993.320 2646.000 994.000 ;
        RECT 1554.400 992.600 2645.600 993.320 ;
        RECT 1550.065 991.920 2645.600 992.600 ;
      LAYER met3 ;
        RECT 2646.000 992.320 2650.000 992.920 ;
      LAYER met3 ;
        RECT 1550.065 987.880 2646.000 991.920 ;
        RECT 1550.065 986.480 2645.600 987.880 ;
      LAYER met3 ;
        RECT 2646.000 986.880 2650.000 987.480 ;
      LAYER met3 ;
        RECT 1550.065 984.480 2646.000 986.480 ;
      LAYER met3 ;
        RECT 1550.000 983.480 1554.000 984.080 ;
      LAYER met3 ;
        RECT 1554.400 983.120 2646.000 984.480 ;
        RECT 1554.400 983.080 2645.600 983.120 ;
        RECT 1550.065 981.720 2645.600 983.080 ;
      LAYER met3 ;
        RECT 2646.000 982.120 2650.000 982.720 ;
      LAYER met3 ;
        RECT 1550.065 978.360 2646.000 981.720 ;
        RECT 1550.065 976.960 2645.600 978.360 ;
      LAYER met3 ;
        RECT 2646.000 977.360 2650.000 977.960 ;
      LAYER met3 ;
        RECT 1550.065 974.960 2646.000 976.960 ;
      LAYER met3 ;
        RECT 1550.000 973.960 1554.000 974.560 ;
      LAYER met3 ;
        RECT 1554.400 973.560 2646.000 974.960 ;
        RECT 1550.065 972.920 2646.000 973.560 ;
        RECT 1550.065 971.520 2645.600 972.920 ;
      LAYER met3 ;
        RECT 2646.000 971.920 2650.000 972.520 ;
      LAYER met3 ;
        RECT 1550.065 968.160 2646.000 971.520 ;
        RECT 1550.065 966.760 2645.600 968.160 ;
      LAYER met3 ;
        RECT 2646.000 967.160 2650.000 967.760 ;
      LAYER met3 ;
        RECT 1550.065 965.440 2646.000 966.760 ;
      LAYER met3 ;
        RECT 1550.000 964.440 1554.000 965.040 ;
      LAYER met3 ;
        RECT 1554.400 964.040 2646.000 965.440 ;
        RECT 1550.065 962.720 2646.000 964.040 ;
        RECT 1550.065 961.320 2645.600 962.720 ;
      LAYER met3 ;
        RECT 2646.000 961.720 2650.000 962.320 ;
      LAYER met3 ;
        RECT 1550.065 957.960 2646.000 961.320 ;
        RECT 1550.065 956.560 2645.600 957.960 ;
      LAYER met3 ;
        RECT 2646.000 956.960 2650.000 957.560 ;
      LAYER met3 ;
        RECT 1550.065 955.920 2646.000 956.560 ;
      LAYER met3 ;
        RECT 1550.000 954.920 1554.000 955.520 ;
      LAYER met3 ;
        RECT 1554.400 954.520 2646.000 955.920 ;
        RECT 1550.065 953.200 2646.000 954.520 ;
        RECT 1550.065 951.800 2645.600 953.200 ;
      LAYER met3 ;
        RECT 2646.000 952.200 2650.000 952.800 ;
      LAYER met3 ;
        RECT 1550.065 947.760 2646.000 951.800 ;
        RECT 1550.065 946.360 2645.600 947.760 ;
      LAYER met3 ;
        RECT 2646.000 946.760 2650.000 947.360 ;
      LAYER met3 ;
        RECT 1550.065 945.720 2646.000 946.360 ;
      LAYER met3 ;
        RECT 1550.000 944.720 1554.000 945.320 ;
      LAYER met3 ;
        RECT 1554.400 944.320 2646.000 945.720 ;
        RECT 1550.065 943.000 2646.000 944.320 ;
        RECT 1550.065 941.600 2645.600 943.000 ;
      LAYER met3 ;
        RECT 2646.000 942.000 2650.000 942.600 ;
      LAYER met3 ;
        RECT 1550.065 937.560 2646.000 941.600 ;
        RECT 1550.065 936.200 2645.600 937.560 ;
      LAYER met3 ;
        RECT 2646.000 936.560 2650.000 937.160 ;
      LAYER met3 ;
        RECT 1554.400 936.160 2645.600 936.200 ;
      LAYER met3 ;
        RECT 1550.000 935.200 1554.000 935.800 ;
      LAYER met3 ;
        RECT 1554.400 934.800 2646.000 936.160 ;
        RECT 1550.065 932.800 2646.000 934.800 ;
        RECT 1550.065 931.400 2645.600 932.800 ;
      LAYER met3 ;
        RECT 2646.000 931.800 2650.000 932.400 ;
      LAYER met3 ;
        RECT 1550.065 927.360 2646.000 931.400 ;
        RECT 1550.065 926.680 2645.600 927.360 ;
      LAYER met3 ;
        RECT 1550.000 925.680 1554.000 926.280 ;
      LAYER met3 ;
        RECT 1554.400 925.960 2645.600 926.680 ;
      LAYER met3 ;
        RECT 2646.000 926.360 2650.000 926.960 ;
      LAYER met3 ;
        RECT 1554.400 925.280 2646.000 925.960 ;
        RECT 1550.065 922.600 2646.000 925.280 ;
        RECT 1550.065 921.200 2645.600 922.600 ;
      LAYER met3 ;
        RECT 2646.000 921.600 2650.000 922.200 ;
      LAYER met3 ;
        RECT 1550.065 917.840 2646.000 921.200 ;
        RECT 1550.065 917.160 2645.600 917.840 ;
      LAYER met3 ;
        RECT 1550.000 916.160 1554.000 916.760 ;
      LAYER met3 ;
        RECT 1554.400 916.440 2645.600 917.160 ;
      LAYER met3 ;
        RECT 2646.000 916.840 2650.000 917.440 ;
      LAYER met3 ;
        RECT 1554.400 915.760 2646.000 916.440 ;
        RECT 1550.065 912.400 2646.000 915.760 ;
        RECT 1550.065 911.000 2645.600 912.400 ;
      LAYER met3 ;
        RECT 2646.000 911.400 2650.000 912.000 ;
      LAYER met3 ;
        RECT 1550.065 907.640 2646.000 911.000 ;
      LAYER met3 ;
        RECT 1550.000 906.640 1554.000 907.240 ;
      LAYER met3 ;
        RECT 1554.400 906.240 2645.600 907.640 ;
      LAYER met3 ;
        RECT 2646.000 906.640 2650.000 907.240 ;
      LAYER met3 ;
        RECT 1550.065 902.200 2646.000 906.240 ;
        RECT 1550.065 900.800 2645.600 902.200 ;
      LAYER met3 ;
        RECT 2646.000 901.200 2650.000 901.800 ;
      LAYER met3 ;
        RECT 1550.065 897.440 2646.000 900.800 ;
      LAYER met3 ;
        RECT 1550.000 896.440 1554.000 897.040 ;
      LAYER met3 ;
        RECT 1554.400 896.040 2645.600 897.440 ;
      LAYER met3 ;
        RECT 2646.000 896.440 2650.000 897.040 ;
      LAYER met3 ;
        RECT 1550.065 892.000 2646.000 896.040 ;
        RECT 1550.065 890.600 2645.600 892.000 ;
      LAYER met3 ;
        RECT 2646.000 891.000 2650.000 891.600 ;
      LAYER met3 ;
        RECT 1550.065 887.920 2646.000 890.600 ;
      LAYER met3 ;
        RECT 1550.000 886.920 1554.000 887.520 ;
      LAYER met3 ;
        RECT 1554.400 887.240 2646.000 887.920 ;
        RECT 1554.400 886.520 2645.600 887.240 ;
        RECT 1550.065 885.840 2645.600 886.520 ;
      LAYER met3 ;
        RECT 2646.000 886.240 2650.000 886.840 ;
      LAYER met3 ;
        RECT 1550.065 882.480 2646.000 885.840 ;
        RECT 1550.065 881.080 2645.600 882.480 ;
      LAYER met3 ;
        RECT 2646.000 881.480 2650.000 882.080 ;
      LAYER met3 ;
        RECT 1550.065 878.400 2646.000 881.080 ;
      LAYER met3 ;
        RECT 1550.000 877.400 1554.000 878.000 ;
      LAYER met3 ;
        RECT 1554.400 877.040 2646.000 878.400 ;
        RECT 1554.400 877.000 2645.600 877.040 ;
        RECT 1550.065 875.640 2645.600 877.000 ;
      LAYER met3 ;
        RECT 2646.000 876.040 2650.000 876.640 ;
      LAYER met3 ;
        RECT 1550.065 872.280 2646.000 875.640 ;
        RECT 1550.065 870.880 2645.600 872.280 ;
      LAYER met3 ;
        RECT 2646.000 871.280 2650.000 871.880 ;
      LAYER met3 ;
        RECT 1550.065 868.880 2646.000 870.880 ;
      LAYER met3 ;
        RECT 1550.000 867.880 1554.000 868.480 ;
      LAYER met3 ;
        RECT 1554.400 867.480 2646.000 868.880 ;
        RECT 1550.065 866.840 2646.000 867.480 ;
        RECT 1550.065 865.440 2645.600 866.840 ;
      LAYER met3 ;
        RECT 2646.000 865.840 2650.000 866.440 ;
      LAYER met3 ;
        RECT 1550.065 862.080 2646.000 865.440 ;
        RECT 1550.065 860.680 2645.600 862.080 ;
      LAYER met3 ;
        RECT 2646.000 861.080 2650.000 861.680 ;
      LAYER met3 ;
        RECT 1550.065 859.360 2646.000 860.680 ;
      LAYER met3 ;
        RECT 1550.000 858.360 1554.000 858.960 ;
      LAYER met3 ;
        RECT 1554.400 857.960 2646.000 859.360 ;
        RECT 1550.065 856.640 2646.000 857.960 ;
        RECT 1550.065 855.240 2645.600 856.640 ;
      LAYER met3 ;
        RECT 2646.000 855.640 2650.000 856.240 ;
      LAYER met3 ;
        RECT 1550.065 851.880 2646.000 855.240 ;
        RECT 1550.065 850.480 2645.600 851.880 ;
      LAYER met3 ;
        RECT 2646.000 850.880 2650.000 851.480 ;
      LAYER met3 ;
        RECT 1550.065 849.160 2646.000 850.480 ;
      LAYER met3 ;
        RECT 1550.000 848.160 1554.000 848.760 ;
      LAYER met3 ;
        RECT 1554.400 847.760 2646.000 849.160 ;
        RECT 1550.065 847.120 2646.000 847.760 ;
        RECT 1550.065 845.720 2645.600 847.120 ;
      LAYER met3 ;
        RECT 2646.000 846.120 2650.000 846.720 ;
      LAYER met3 ;
        RECT 1550.065 841.680 2646.000 845.720 ;
        RECT 1550.065 840.280 2645.600 841.680 ;
      LAYER met3 ;
        RECT 2646.000 840.680 2650.000 841.280 ;
      LAYER met3 ;
        RECT 1550.065 839.640 2646.000 840.280 ;
      LAYER met3 ;
        RECT 1550.000 838.640 1554.000 839.240 ;
      LAYER met3 ;
        RECT 1554.400 838.240 2646.000 839.640 ;
        RECT 1550.065 836.920 2646.000 838.240 ;
        RECT 1550.065 835.520 2645.600 836.920 ;
      LAYER met3 ;
        RECT 2646.000 835.920 2650.000 836.520 ;
      LAYER met3 ;
        RECT 1550.065 831.480 2646.000 835.520 ;
        RECT 1550.065 830.120 2645.600 831.480 ;
      LAYER met3 ;
        RECT 2646.000 830.480 2650.000 831.080 ;
      LAYER met3 ;
        RECT 1554.400 830.080 2645.600 830.120 ;
      LAYER met3 ;
        RECT 1550.000 829.120 1554.000 829.720 ;
      LAYER met3 ;
        RECT 1554.400 828.720 2646.000 830.080 ;
        RECT 1550.065 826.720 2646.000 828.720 ;
        RECT 1550.065 825.320 2645.600 826.720 ;
      LAYER met3 ;
        RECT 2646.000 825.720 2650.000 826.320 ;
      LAYER met3 ;
        RECT 1550.065 821.960 2646.000 825.320 ;
        RECT 1550.065 820.600 2645.600 821.960 ;
      LAYER met3 ;
        RECT 2646.000 820.960 2650.000 821.560 ;
      LAYER met3 ;
        RECT 1554.400 820.560 2645.600 820.600 ;
      LAYER met3 ;
        RECT 1550.000 819.600 1554.000 820.200 ;
      LAYER met3 ;
        RECT 1554.400 819.200 2646.000 820.560 ;
        RECT 1550.065 816.520 2646.000 819.200 ;
        RECT 1550.065 815.120 2645.600 816.520 ;
      LAYER met3 ;
        RECT 2646.000 815.520 2650.000 816.120 ;
      LAYER met3 ;
        RECT 1550.065 811.760 2646.000 815.120 ;
        RECT 1550.065 811.080 2645.600 811.760 ;
      LAYER met3 ;
        RECT 1550.000 810.080 1554.000 810.680 ;
      LAYER met3 ;
        RECT 1554.400 810.360 2645.600 811.080 ;
      LAYER met3 ;
        RECT 2646.000 810.760 2650.000 811.360 ;
      LAYER met3 ;
        RECT 1554.400 809.680 2646.000 810.360 ;
        RECT 1550.065 806.320 2646.000 809.680 ;
        RECT 1550.065 804.920 2645.600 806.320 ;
      LAYER met3 ;
        RECT 2646.000 805.320 2650.000 805.920 ;
      LAYER met3 ;
        RECT 1550.065 801.560 2646.000 804.920 ;
        RECT 1550.065 800.880 2645.600 801.560 ;
      LAYER met3 ;
        RECT 1550.000 799.880 1554.000 800.480 ;
      LAYER met3 ;
        RECT 1554.400 800.160 2645.600 800.880 ;
      LAYER met3 ;
        RECT 2646.000 800.560 2650.000 801.160 ;
      LAYER met3 ;
        RECT 1554.400 799.480 2646.000 800.160 ;
        RECT 1550.065 796.120 2646.000 799.480 ;
        RECT 1550.065 794.720 2645.600 796.120 ;
      LAYER met3 ;
        RECT 2646.000 795.120 2650.000 795.720 ;
      LAYER met3 ;
        RECT 1550.065 791.360 2646.000 794.720 ;
      LAYER met3 ;
        RECT 1550.000 790.360 1554.000 790.960 ;
      LAYER met3 ;
        RECT 1554.400 789.960 2645.600 791.360 ;
      LAYER met3 ;
        RECT 2646.000 790.360 2650.000 790.960 ;
      LAYER met3 ;
        RECT 1550.065 786.600 2646.000 789.960 ;
        RECT 1550.065 785.200 2645.600 786.600 ;
      LAYER met3 ;
        RECT 2646.000 785.600 2650.000 786.200 ;
      LAYER met3 ;
        RECT 1550.065 781.840 2646.000 785.200 ;
      LAYER met3 ;
        RECT 1550.000 780.840 1554.000 781.440 ;
      LAYER met3 ;
        RECT 1554.400 781.160 2646.000 781.840 ;
        RECT 1554.400 780.440 2645.600 781.160 ;
        RECT 1550.065 779.760 2645.600 780.440 ;
      LAYER met3 ;
        RECT 2646.000 780.160 2650.000 780.760 ;
      LAYER met3 ;
        RECT 1550.065 776.400 2646.000 779.760 ;
        RECT 1550.065 775.000 2645.600 776.400 ;
      LAYER met3 ;
        RECT 2646.000 775.400 2650.000 776.000 ;
      LAYER met3 ;
        RECT 1550.065 772.320 2646.000 775.000 ;
      LAYER met3 ;
        RECT 1550.000 771.320 1554.000 771.920 ;
      LAYER met3 ;
        RECT 1554.400 770.960 2646.000 772.320 ;
        RECT 1554.400 770.920 2645.600 770.960 ;
        RECT 1550.065 769.560 2645.600 770.920 ;
      LAYER met3 ;
        RECT 2646.000 769.960 2650.000 770.560 ;
      LAYER met3 ;
        RECT 1550.065 766.200 2646.000 769.560 ;
        RECT 1550.065 764.800 2645.600 766.200 ;
      LAYER met3 ;
        RECT 2646.000 765.200 2650.000 765.800 ;
      LAYER met3 ;
        RECT 1550.065 762.800 2646.000 764.800 ;
      LAYER met3 ;
        RECT 1550.000 761.800 1554.000 762.400 ;
      LAYER met3 ;
        RECT 1554.400 761.400 2646.000 762.800 ;
        RECT 1550.065 760.760 2646.000 761.400 ;
        RECT 1550.065 759.360 2645.600 760.760 ;
      LAYER met3 ;
        RECT 2646.000 759.760 2650.000 760.360 ;
      LAYER met3 ;
        RECT 1550.065 756.000 2646.000 759.360 ;
        RECT 1550.065 754.600 2645.600 756.000 ;
      LAYER met3 ;
        RECT 2646.000 755.000 2650.000 755.600 ;
      LAYER met3 ;
        RECT 1550.065 752.600 2646.000 754.600 ;
      LAYER met3 ;
        RECT 1550.000 751.600 1554.000 752.200 ;
      LAYER met3 ;
        RECT 1554.400 751.240 2646.000 752.600 ;
        RECT 1554.400 751.200 2645.600 751.240 ;
        RECT 1550.065 749.840 2645.600 751.200 ;
      LAYER met3 ;
        RECT 2646.000 750.240 2650.000 750.840 ;
      LAYER met3 ;
        RECT 1550.065 745.800 2646.000 749.840 ;
        RECT 1550.065 744.400 2645.600 745.800 ;
      LAYER met3 ;
        RECT 2646.000 744.800 2650.000 745.400 ;
      LAYER met3 ;
        RECT 1550.065 743.080 2646.000 744.400 ;
      LAYER met3 ;
        RECT 1550.000 742.080 1554.000 742.680 ;
      LAYER met3 ;
        RECT 1554.400 741.680 2646.000 743.080 ;
        RECT 1550.065 741.040 2646.000 741.680 ;
        RECT 1550.065 739.640 2645.600 741.040 ;
      LAYER met3 ;
        RECT 2646.000 740.040 2650.000 740.640 ;
      LAYER met3 ;
        RECT 1550.065 735.600 2646.000 739.640 ;
        RECT 1550.065 734.200 2645.600 735.600 ;
      LAYER met3 ;
        RECT 2646.000 734.600 2650.000 735.200 ;
      LAYER met3 ;
        RECT 1550.065 733.560 2646.000 734.200 ;
      LAYER met3 ;
        RECT 1550.000 732.560 1554.000 733.160 ;
      LAYER met3 ;
        RECT 1554.400 732.160 2646.000 733.560 ;
        RECT 1550.065 730.840 2646.000 732.160 ;
        RECT 1550.065 729.440 2645.600 730.840 ;
      LAYER met3 ;
        RECT 2646.000 729.840 2650.000 730.440 ;
      LAYER met3 ;
        RECT 1550.065 726.080 2646.000 729.440 ;
        RECT 1550.065 724.680 2645.600 726.080 ;
      LAYER met3 ;
        RECT 2646.000 725.080 2650.000 725.680 ;
      LAYER met3 ;
        RECT 1550.065 724.040 2646.000 724.680 ;
      LAYER met3 ;
        RECT 1550.000 723.040 1554.000 723.640 ;
      LAYER met3 ;
        RECT 1554.400 722.640 2646.000 724.040 ;
        RECT 1550.065 720.640 2646.000 722.640 ;
        RECT 1550.065 719.240 2645.600 720.640 ;
      LAYER met3 ;
        RECT 2646.000 719.640 2650.000 720.240 ;
      LAYER met3 ;
        RECT 1550.065 715.880 2646.000 719.240 ;
        RECT 1550.065 714.520 2645.600 715.880 ;
      LAYER met3 ;
        RECT 2646.000 714.880 2650.000 715.480 ;
      LAYER met3 ;
        RECT 1554.400 714.480 2645.600 714.520 ;
      LAYER met3 ;
        RECT 1550.000 713.520 1554.000 714.120 ;
      LAYER met3 ;
        RECT 1554.400 713.120 2646.000 714.480 ;
        RECT 1550.065 710.440 2646.000 713.120 ;
        RECT 1550.065 709.040 2645.600 710.440 ;
      LAYER met3 ;
        RECT 2646.000 709.440 2650.000 710.040 ;
      LAYER met3 ;
        RECT 1550.065 705.680 2646.000 709.040 ;
        RECT 1550.065 704.320 2645.600 705.680 ;
      LAYER met3 ;
        RECT 2646.000 704.680 2650.000 705.280 ;
      LAYER met3 ;
        RECT 1554.400 704.280 2645.600 704.320 ;
      LAYER met3 ;
        RECT 1550.000 703.320 1554.000 703.920 ;
      LAYER met3 ;
        RECT 1554.400 702.920 2646.000 704.280 ;
        RECT 1550.065 700.240 2646.000 702.920 ;
        RECT 1550.065 698.840 2645.600 700.240 ;
      LAYER met3 ;
        RECT 2646.000 699.240 2650.000 699.840 ;
      LAYER met3 ;
        RECT 1550.065 695.480 2646.000 698.840 ;
        RECT 1550.065 694.800 2645.600 695.480 ;
      LAYER met3 ;
        RECT 1550.000 693.800 1554.000 694.400 ;
      LAYER met3 ;
        RECT 1554.400 694.080 2645.600 694.800 ;
      LAYER met3 ;
        RECT 2646.000 694.480 2650.000 695.080 ;
      LAYER met3 ;
        RECT 1554.400 693.400 2646.000 694.080 ;
        RECT 1550.065 690.720 2646.000 693.400 ;
        RECT 1550.065 689.320 2645.600 690.720 ;
      LAYER met3 ;
        RECT 2646.000 689.720 2650.000 690.320 ;
      LAYER met3 ;
        RECT 1550.065 685.280 2646.000 689.320 ;
      LAYER met3 ;
        RECT 1550.000 684.280 1554.000 684.880 ;
      LAYER met3 ;
        RECT 1554.400 683.880 2645.600 685.280 ;
      LAYER met3 ;
        RECT 2646.000 684.280 2650.000 684.880 ;
      LAYER met3 ;
        RECT 1550.065 680.520 2646.000 683.880 ;
        RECT 1550.065 679.120 2645.600 680.520 ;
      LAYER met3 ;
        RECT 2646.000 679.520 2650.000 680.120 ;
      LAYER met3 ;
        RECT 1550.065 675.760 2646.000 679.120 ;
      LAYER met3 ;
        RECT 1550.000 674.760 1554.000 675.360 ;
      LAYER met3 ;
        RECT 1554.400 675.080 2646.000 675.760 ;
        RECT 1554.400 674.360 2645.600 675.080 ;
        RECT 1550.065 673.680 2645.600 674.360 ;
      LAYER met3 ;
        RECT 2646.000 674.080 2650.000 674.680 ;
      LAYER met3 ;
        RECT 1550.065 670.320 2646.000 673.680 ;
        RECT 1550.065 668.920 2645.600 670.320 ;
      LAYER met3 ;
        RECT 2646.000 669.320 2650.000 669.920 ;
      LAYER met3 ;
        RECT 1550.065 666.240 2646.000 668.920 ;
      LAYER met3 ;
        RECT 1550.000 665.240 1554.000 665.840 ;
      LAYER met3 ;
        RECT 1554.400 664.880 2646.000 666.240 ;
        RECT 1554.400 664.840 2645.600 664.880 ;
        RECT 1550.065 663.480 2645.600 664.840 ;
      LAYER met3 ;
        RECT 2646.000 663.880 2650.000 664.480 ;
      LAYER met3 ;
        RECT 1550.065 660.120 2646.000 663.480 ;
        RECT 1550.065 658.720 2645.600 660.120 ;
      LAYER met3 ;
        RECT 2646.000 659.120 2650.000 659.720 ;
      LAYER met3 ;
        RECT 1550.065 656.720 2646.000 658.720 ;
      LAYER met3 ;
        RECT 1550.000 655.720 1554.000 656.320 ;
      LAYER met3 ;
        RECT 1554.400 655.360 2646.000 656.720 ;
        RECT 1554.400 655.320 2645.600 655.360 ;
        RECT 1550.065 653.960 2645.600 655.320 ;
      LAYER met3 ;
        RECT 2646.000 654.360 2650.000 654.960 ;
      LAYER met3 ;
        RECT 1550.065 649.920 2646.000 653.960 ;
        RECT 1550.065 648.520 2645.600 649.920 ;
      LAYER met3 ;
        RECT 2646.000 648.920 2650.000 649.520 ;
      LAYER met3 ;
        RECT 1550.065 646.520 2646.000 648.520 ;
      LAYER met3 ;
        RECT 1550.000 645.520 1554.000 646.120 ;
      LAYER met3 ;
        RECT 1554.400 645.160 2646.000 646.520 ;
        RECT 1554.400 645.120 2645.600 645.160 ;
        RECT 1550.065 643.760 2645.600 645.120 ;
      LAYER met3 ;
        RECT 2646.000 644.160 2650.000 644.760 ;
      LAYER met3 ;
        RECT 1550.065 639.720 2646.000 643.760 ;
        RECT 1550.065 638.320 2645.600 639.720 ;
      LAYER met3 ;
        RECT 2646.000 638.720 2650.000 639.320 ;
      LAYER met3 ;
        RECT 1550.065 637.000 2646.000 638.320 ;
      LAYER met3 ;
        RECT 1550.000 636.000 1554.000 636.600 ;
      LAYER met3 ;
        RECT 1554.400 635.600 2646.000 637.000 ;
        RECT 1550.065 634.960 2646.000 635.600 ;
        RECT 1550.065 633.560 2645.600 634.960 ;
      LAYER met3 ;
        RECT 2646.000 633.960 2650.000 634.560 ;
      LAYER met3 ;
        RECT 1550.065 629.520 2646.000 633.560 ;
        RECT 1550.065 628.120 2645.600 629.520 ;
      LAYER met3 ;
        RECT 2646.000 628.520 2650.000 629.120 ;
      LAYER met3 ;
        RECT 1550.065 627.480 2646.000 628.120 ;
      LAYER met3 ;
        RECT 1550.000 626.480 1554.000 627.080 ;
      LAYER met3 ;
        RECT 1554.400 626.080 2646.000 627.480 ;
        RECT 1550.065 624.760 2646.000 626.080 ;
        RECT 1550.065 623.360 2645.600 624.760 ;
      LAYER met3 ;
        RECT 2646.000 623.760 2650.000 624.360 ;
      LAYER met3 ;
        RECT 1550.065 620.000 2646.000 623.360 ;
        RECT 1550.065 618.600 2645.600 620.000 ;
      LAYER met3 ;
        RECT 2646.000 619.000 2650.000 619.600 ;
      LAYER met3 ;
        RECT 1550.065 617.960 2646.000 618.600 ;
      LAYER met3 ;
        RECT 1550.000 616.960 1554.000 617.560 ;
      LAYER met3 ;
        RECT 1554.400 616.560 2646.000 617.960 ;
        RECT 1550.065 614.560 2646.000 616.560 ;
        RECT 1550.065 613.160 2645.600 614.560 ;
      LAYER met3 ;
        RECT 2646.000 613.560 2650.000 614.160 ;
      LAYER met3 ;
        RECT 1550.065 609.800 2646.000 613.160 ;
        RECT 1550.065 608.440 2645.600 609.800 ;
      LAYER met3 ;
        RECT 2646.000 608.800 2650.000 609.400 ;
      LAYER met3 ;
        RECT 1554.400 608.400 2645.600 608.440 ;
      LAYER met3 ;
        RECT 1550.000 607.440 1554.000 608.040 ;
      LAYER met3 ;
        RECT 1554.400 607.040 2646.000 608.400 ;
        RECT 1550.065 604.360 2646.000 607.040 ;
        RECT 1550.065 602.960 2645.600 604.360 ;
      LAYER met3 ;
        RECT 2646.000 603.360 2650.000 603.960 ;
      LAYER met3 ;
        RECT 1550.065 599.600 2646.000 602.960 ;
        RECT 1550.065 598.240 2645.600 599.600 ;
      LAYER met3 ;
        RECT 2646.000 598.600 2650.000 599.200 ;
      LAYER met3 ;
        RECT 1554.400 598.200 2645.600 598.240 ;
      LAYER met3 ;
        RECT 1550.000 597.240 1554.000 597.840 ;
      LAYER met3 ;
        RECT 1554.400 596.840 2646.000 598.200 ;
        RECT 1550.065 594.840 2646.000 596.840 ;
        RECT 1550.065 593.440 2645.600 594.840 ;
      LAYER met3 ;
        RECT 2646.000 593.840 2650.000 594.440 ;
      LAYER met3 ;
        RECT 1550.065 589.400 2646.000 593.440 ;
        RECT 1550.065 588.720 2645.600 589.400 ;
      LAYER met3 ;
        RECT 1550.000 587.720 1554.000 588.320 ;
      LAYER met3 ;
        RECT 1554.400 588.000 2645.600 588.720 ;
      LAYER met3 ;
        RECT 2646.000 588.400 2650.000 589.000 ;
      LAYER met3 ;
        RECT 1554.400 587.320 2646.000 588.000 ;
        RECT 1550.065 584.640 2646.000 587.320 ;
        RECT 1550.065 583.240 2645.600 584.640 ;
      LAYER met3 ;
        RECT 2646.000 583.640 2650.000 584.240 ;
      LAYER met3 ;
        RECT 1550.065 579.200 2646.000 583.240 ;
      LAYER met3 ;
        RECT 1550.000 578.200 1554.000 578.800 ;
      LAYER met3 ;
        RECT 1554.400 577.800 2645.600 579.200 ;
      LAYER met3 ;
        RECT 2646.000 578.200 2650.000 578.800 ;
      LAYER met3 ;
        RECT 1550.065 574.440 2646.000 577.800 ;
        RECT 1550.065 573.040 2645.600 574.440 ;
      LAYER met3 ;
        RECT 2646.000 573.440 2650.000 574.040 ;
      LAYER met3 ;
        RECT 1550.065 569.680 2646.000 573.040 ;
      LAYER met3 ;
        RECT 1550.000 568.680 1554.000 569.280 ;
      LAYER met3 ;
        RECT 1554.400 569.000 2646.000 569.680 ;
        RECT 1554.400 568.280 2645.600 569.000 ;
        RECT 1550.065 567.600 2645.600 568.280 ;
      LAYER met3 ;
        RECT 2646.000 568.000 2650.000 568.600 ;
      LAYER met3 ;
        RECT 1550.065 564.240 2646.000 567.600 ;
        RECT 1550.065 562.840 2645.600 564.240 ;
      LAYER met3 ;
        RECT 2646.000 563.240 2650.000 563.840 ;
      LAYER met3 ;
        RECT 1550.065 560.160 2646.000 562.840 ;
      LAYER met3 ;
        RECT 1550.000 559.160 1554.000 559.760 ;
      LAYER met3 ;
        RECT 1554.400 559.480 2646.000 560.160 ;
        RECT 1554.400 558.760 2645.600 559.480 ;
        RECT 1550.065 558.080 2645.600 558.760 ;
      LAYER met3 ;
        RECT 2646.000 558.480 2650.000 559.080 ;
      LAYER met3 ;
        RECT 1550.065 554.040 2646.000 558.080 ;
        RECT 1550.065 552.640 2645.600 554.040 ;
      LAYER met3 ;
        RECT 2646.000 553.040 2650.000 553.640 ;
      LAYER met3 ;
        RECT 1550.065 549.960 2646.000 552.640 ;
      LAYER met3 ;
        RECT 1550.000 548.960 1554.000 549.560 ;
      LAYER met3 ;
        RECT 1554.400 549.280 2646.000 549.960 ;
        RECT 1554.400 548.560 2645.600 549.280 ;
        RECT 1550.065 547.880 2645.600 548.560 ;
      LAYER met3 ;
        RECT 2646.000 548.280 2650.000 548.880 ;
      LAYER met3 ;
        RECT 1550.065 543.840 2646.000 547.880 ;
        RECT 1550.065 542.440 2645.600 543.840 ;
      LAYER met3 ;
        RECT 2646.000 542.840 2650.000 543.440 ;
      LAYER met3 ;
        RECT 1550.065 540.440 2646.000 542.440 ;
      LAYER met3 ;
        RECT 1550.000 539.440 1554.000 540.040 ;
      LAYER met3 ;
        RECT 1554.400 539.080 2646.000 540.440 ;
        RECT 1554.400 539.040 2645.600 539.080 ;
        RECT 1550.065 537.680 2645.600 539.040 ;
      LAYER met3 ;
        RECT 2646.000 538.080 2650.000 538.680 ;
      LAYER met3 ;
        RECT 1550.065 533.640 2646.000 537.680 ;
        RECT 1550.065 532.240 2645.600 533.640 ;
      LAYER met3 ;
        RECT 2646.000 532.640 2650.000 533.240 ;
      LAYER met3 ;
        RECT 1550.065 530.920 2646.000 532.240 ;
      LAYER met3 ;
        RECT 1550.000 529.920 1554.000 530.520 ;
      LAYER met3 ;
        RECT 1554.400 529.520 2646.000 530.920 ;
        RECT 1550.065 528.880 2646.000 529.520 ;
        RECT 1550.065 527.480 2645.600 528.880 ;
      LAYER met3 ;
        RECT 2646.000 527.880 2650.000 528.480 ;
      LAYER met3 ;
        RECT 1550.065 524.120 2646.000 527.480 ;
        RECT 1550.065 522.720 2645.600 524.120 ;
      LAYER met3 ;
        RECT 2646.000 523.120 2650.000 523.720 ;
      LAYER met3 ;
        RECT 1550.065 521.400 2646.000 522.720 ;
      LAYER met3 ;
        RECT 1550.000 520.400 1554.000 521.000 ;
      LAYER met3 ;
        RECT 1554.400 520.000 2646.000 521.400 ;
        RECT 1550.065 518.680 2646.000 520.000 ;
        RECT 1550.065 517.280 2645.600 518.680 ;
      LAYER met3 ;
        RECT 2646.000 517.680 2650.000 518.280 ;
      LAYER met3 ;
        RECT 1550.065 513.920 2646.000 517.280 ;
        RECT 1550.065 512.520 2645.600 513.920 ;
      LAYER met3 ;
        RECT 2646.000 512.920 2650.000 513.520 ;
      LAYER met3 ;
        RECT 1550.065 511.880 2646.000 512.520 ;
      LAYER met3 ;
        RECT 1550.000 510.880 1554.000 511.480 ;
      LAYER met3 ;
        RECT 1554.400 510.480 2646.000 511.880 ;
        RECT 1550.065 508.480 2646.000 510.480 ;
        RECT 1550.065 507.080 2645.600 508.480 ;
      LAYER met3 ;
        RECT 2646.000 507.480 2650.000 508.080 ;
      LAYER met3 ;
        RECT 1550.065 503.720 2646.000 507.080 ;
        RECT 1550.065 502.320 2645.600 503.720 ;
      LAYER met3 ;
        RECT 2646.000 502.720 2650.000 503.320 ;
      LAYER met3 ;
        RECT 1550.065 501.680 2646.000 502.320 ;
      LAYER met3 ;
        RECT 1550.000 500.680 1554.000 501.280 ;
      LAYER met3 ;
        RECT 1554.400 500.280 2646.000 501.680 ;
        RECT 1550.065 498.960 2646.000 500.280 ;
        RECT 1550.065 497.560 2645.600 498.960 ;
      LAYER met3 ;
        RECT 2646.000 497.960 2650.000 498.560 ;
      LAYER met3 ;
        RECT 1550.065 493.520 2646.000 497.560 ;
        RECT 1550.065 492.160 2645.600 493.520 ;
      LAYER met3 ;
        RECT 2646.000 492.520 2650.000 493.120 ;
      LAYER met3 ;
        RECT 1554.400 492.120 2645.600 492.160 ;
      LAYER met3 ;
        RECT 1550.000 491.160 1554.000 491.760 ;
      LAYER met3 ;
        RECT 1554.400 490.760 2646.000 492.120 ;
        RECT 1550.065 488.760 2646.000 490.760 ;
        RECT 1550.065 487.360 2645.600 488.760 ;
      LAYER met3 ;
        RECT 2646.000 487.760 2650.000 488.360 ;
      LAYER met3 ;
        RECT 1550.065 483.320 2646.000 487.360 ;
        RECT 1550.065 482.640 2645.600 483.320 ;
      LAYER met3 ;
        RECT 1550.000 481.640 1554.000 482.240 ;
      LAYER met3 ;
        RECT 1554.400 481.920 2645.600 482.640 ;
      LAYER met3 ;
        RECT 2646.000 482.320 2650.000 482.920 ;
      LAYER met3 ;
        RECT 1554.400 481.240 2646.000 481.920 ;
        RECT 1550.065 478.560 2646.000 481.240 ;
        RECT 1550.065 477.160 2645.600 478.560 ;
      LAYER met3 ;
        RECT 2646.000 477.560 2650.000 478.160 ;
      LAYER met3 ;
        RECT 1550.065 473.120 2646.000 477.160 ;
      LAYER met3 ;
        RECT 1550.000 472.120 1554.000 472.720 ;
      LAYER met3 ;
        RECT 1554.400 471.720 2645.600 473.120 ;
      LAYER met3 ;
        RECT 2646.000 472.120 2650.000 472.720 ;
      LAYER met3 ;
        RECT 1550.065 468.360 2646.000 471.720 ;
        RECT 1550.065 466.960 2645.600 468.360 ;
      LAYER met3 ;
        RECT 2646.000 467.360 2650.000 467.960 ;
      LAYER met3 ;
        RECT 1550.065 463.600 2646.000 466.960 ;
      LAYER met3 ;
        RECT 1550.000 462.600 1554.000 463.200 ;
      LAYER met3 ;
        RECT 1554.400 462.200 2645.600 463.600 ;
      LAYER met3 ;
        RECT 2646.000 462.600 2650.000 463.200 ;
      LAYER met3 ;
        RECT 1550.065 458.160 2646.000 462.200 ;
        RECT 1550.065 456.760 2645.600 458.160 ;
      LAYER met3 ;
        RECT 2646.000 457.160 2650.000 457.760 ;
      LAYER met3 ;
        RECT 1550.065 453.400 2646.000 456.760 ;
      LAYER met3 ;
        RECT 1550.000 452.400 1554.000 453.000 ;
      LAYER met3 ;
        RECT 1554.400 452.000 2645.600 453.400 ;
      LAYER met3 ;
        RECT 2646.000 452.400 2650.000 453.000 ;
      LAYER met3 ;
        RECT 1550.065 447.960 2646.000 452.000 ;
        RECT 1550.065 446.560 2645.600 447.960 ;
      LAYER met3 ;
        RECT 2646.000 446.960 2650.000 447.560 ;
      LAYER met3 ;
        RECT 1550.065 443.880 2646.000 446.560 ;
      LAYER met3 ;
        RECT 1550.000 442.880 1554.000 443.480 ;
      LAYER met3 ;
        RECT 1554.400 443.200 2646.000 443.880 ;
        RECT 1554.400 442.480 2645.600 443.200 ;
        RECT 1550.065 441.800 2645.600 442.480 ;
      LAYER met3 ;
        RECT 2646.000 442.200 2650.000 442.800 ;
      LAYER met3 ;
        RECT 1550.065 437.760 2646.000 441.800 ;
        RECT 1550.065 436.360 2645.600 437.760 ;
      LAYER met3 ;
        RECT 2646.000 436.760 2650.000 437.360 ;
      LAYER met3 ;
        RECT 1550.065 434.360 2646.000 436.360 ;
      LAYER met3 ;
        RECT 1550.000 433.360 1554.000 433.960 ;
      LAYER met3 ;
        RECT 1554.400 433.000 2646.000 434.360 ;
        RECT 1554.400 432.960 2645.600 433.000 ;
        RECT 1550.065 431.600 2645.600 432.960 ;
      LAYER met3 ;
        RECT 2646.000 432.000 2650.000 432.600 ;
      LAYER met3 ;
        RECT 1550.065 428.240 2646.000 431.600 ;
        RECT 1550.065 426.840 2645.600 428.240 ;
      LAYER met3 ;
        RECT 2646.000 427.240 2650.000 427.840 ;
      LAYER met3 ;
        RECT 1550.065 424.840 2646.000 426.840 ;
      LAYER met3 ;
        RECT 1550.000 423.840 1554.000 424.440 ;
      LAYER met3 ;
        RECT 1554.400 423.440 2646.000 424.840 ;
        RECT 1550.065 422.800 2646.000 423.440 ;
        RECT 1550.065 421.400 2645.600 422.800 ;
      LAYER met3 ;
        RECT 2646.000 421.800 2650.000 422.400 ;
      LAYER met3 ;
        RECT 1550.065 418.040 2646.000 421.400 ;
        RECT 1550.065 416.640 2645.600 418.040 ;
      LAYER met3 ;
        RECT 2646.000 417.040 2650.000 417.640 ;
      LAYER met3 ;
        RECT 1550.065 415.320 2646.000 416.640 ;
      LAYER met3 ;
        RECT 1550.000 414.320 1554.000 414.920 ;
      LAYER met3 ;
        RECT 1554.400 413.920 2646.000 415.320 ;
        RECT 1550.065 412.600 2646.000 413.920 ;
        RECT 1550.065 411.200 2645.600 412.600 ;
      LAYER met3 ;
        RECT 2646.000 411.600 2650.000 412.200 ;
      LAYER met3 ;
        RECT 1550.065 407.840 2646.000 411.200 ;
        RECT 1550.065 406.440 2645.600 407.840 ;
      LAYER met3 ;
        RECT 2646.000 406.840 2650.000 407.440 ;
      LAYER met3 ;
        RECT 1550.065 405.800 2646.000 406.440 ;
      LAYER met3 ;
        RECT 1550.000 404.800 1554.000 405.400 ;
      LAYER met3 ;
        RECT 1554.400 404.400 2646.000 405.800 ;
        RECT 1550.065 403.080 2646.000 404.400 ;
        RECT 1550.065 402.215 2645.600 403.080 ;
      LAYER met3 ;
        RECT 2646.000 402.080 2650.000 402.680 ;
      LAYER via3 ;
        RECT 1890.900 3264.180 1891.220 3264.500 ;
        RECT 1917.580 3264.180 1917.900 3264.500 ;
        RECT 2542.260 3264.180 2542.580 3264.500 ;
        RECT 2567.100 3264.180 2567.420 3264.500 ;
        RECT 1292.880 3258.060 1293.200 3258.380 ;
        RECT 1317.855 3258.060 1318.175 3258.380 ;
        RECT 646.140 3255.340 646.460 3255.660 ;
        RECT 669.140 3255.340 669.460 3255.660 ;
        RECT 302.980 2894.940 303.300 2895.260 ;
        RECT 944.220 2894.940 944.540 2895.260 ;
        RECT 1351.780 2935.740 1352.100 2936.060 ;
        RECT 1412.500 2894.940 1412.820 2895.260 ;
        RECT 1551.420 2894.940 1551.740 2895.260 ;
        RECT 1937.820 2935.740 1938.140 2936.060 ;
        RECT 1946.100 2904.460 1946.420 2904.780 ;
        RECT 2187.140 2894.940 2187.460 2895.260 ;
        RECT 2594.700 2904.460 2595.020 2904.780 ;
        RECT 1055.540 2799.740 1055.860 2800.060 ;
        RECT 1759.340 2796.340 1759.660 2796.660 ;
        RECT 1794.300 2796.340 1794.620 2796.660 ;
        RECT 337.020 2794.300 337.340 2794.620 ;
        RECT 342.540 2794.300 342.860 2794.620 ;
        RECT 350.820 2794.300 351.140 2794.620 ;
        RECT 358.180 2794.300 358.500 2794.620 ;
        RECT 361.860 2794.300 362.180 2794.620 ;
        RECT 364.620 2794.300 364.940 2794.620 ;
        RECT 368.300 2794.300 368.620 2794.620 ;
        RECT 371.060 2794.300 371.380 2794.620 ;
        RECT 374.740 2794.300 375.060 2794.620 ;
        RECT 378.420 2794.300 378.740 2794.620 ;
        RECT 383.940 2794.300 384.260 2794.620 ;
        RECT 386.700 2794.300 387.020 2794.620 ;
        RECT 390.380 2794.300 390.700 2794.620 ;
        RECT 395.900 2794.300 396.220 2794.620 ;
        RECT 399.580 2794.300 399.900 2794.620 ;
        RECT 403.260 2794.300 403.580 2794.620 ;
        RECT 406.020 2794.300 406.340 2794.620 ;
        RECT 409.700 2794.300 410.020 2794.620 ;
        RECT 414.300 2794.300 414.620 2794.620 ;
        RECT 418.900 2794.300 419.220 2794.620 ;
        RECT 420.740 2794.300 421.060 2794.620 ;
        RECT 425.340 2794.300 425.660 2794.620 ;
        RECT 431.780 2794.300 432.100 2794.620 ;
        RECT 433.620 2794.300 433.940 2794.620 ;
        RECT 439.140 2794.300 439.460 2794.620 ;
        RECT 440.980 2794.300 441.300 2794.620 ;
        RECT 444.660 2794.300 444.980 2794.620 ;
        RECT 445.580 2794.300 445.900 2794.620 ;
        RECT 449.260 2794.300 449.580 2794.620 ;
        RECT 454.780 2794.300 455.100 2794.620 ;
        RECT 459.380 2794.300 459.700 2794.620 ;
        RECT 462.140 2794.300 462.460 2794.620 ;
        RECT 466.740 2794.300 467.060 2794.620 ;
        RECT 468.580 2794.300 468.900 2794.620 ;
        RECT 475.020 2794.300 475.340 2794.620 ;
        RECT 478.700 2794.300 479.020 2794.620 ;
        RECT 482.380 2794.300 482.700 2794.620 ;
        RECT 485.140 2794.300 485.460 2794.620 ;
        RECT 488.820 2794.300 489.140 2794.620 ;
        RECT 491.580 2794.300 491.900 2794.620 ;
        RECT 495.260 2794.300 495.580 2794.620 ;
        RECT 499.860 2794.300 500.180 2794.620 ;
        RECT 509.980 2794.300 510.300 2794.620 ;
        RECT 523.780 2794.300 524.100 2794.620 ;
        RECT 535.740 2794.300 536.060 2794.620 ;
        RECT 542.180 2794.300 542.500 2794.620 ;
        RECT 981.020 2794.300 981.340 2794.620 ;
        RECT 1001.260 2794.300 1001.580 2794.620 ;
        RECT 1013.220 2794.300 1013.540 2794.620 ;
        RECT 1018.740 2794.300 1019.060 2794.620 ;
        RECT 1019.660 2794.300 1019.980 2794.620 ;
        RECT 1027.020 2794.300 1027.340 2794.620 ;
        RECT 1030.700 2794.300 1031.020 2794.620 ;
        RECT 1041.740 2794.300 1042.060 2794.620 ;
        RECT 1052.780 2794.300 1053.100 2794.620 ;
        RECT 1059.220 2794.300 1059.540 2794.620 ;
        RECT 1065.660 2794.300 1065.980 2794.620 ;
        RECT 1070.260 2794.300 1070.580 2794.620 ;
        RECT 1076.700 2794.300 1077.020 2794.620 ;
        RECT 1083.140 2794.300 1083.460 2794.620 ;
        RECT 1094.180 2794.300 1094.500 2794.620 ;
        RECT 1100.620 2794.300 1100.940 2794.620 ;
        RECT 1105.220 2794.300 1105.540 2794.620 ;
        RECT 1111.660 2794.300 1111.980 2794.620 ;
        RECT 1122.700 2794.300 1123.020 2794.620 ;
        RECT 1129.140 2794.300 1129.460 2794.620 ;
        RECT 1130.980 2794.300 1131.300 2794.620 ;
        RECT 1135.580 2794.300 1135.900 2794.620 ;
        RECT 1137.420 2794.300 1137.740 2794.620 ;
        RECT 1140.180 2794.300 1140.500 2794.620 ;
        RECT 1143.860 2794.300 1144.180 2794.620 ;
        RECT 1147.540 2794.300 1147.860 2794.620 ;
        RECT 1151.220 2794.300 1151.540 2794.620 ;
        RECT 1153.980 2794.300 1154.300 2794.620 ;
        RECT 1165.020 2794.300 1165.340 2794.620 ;
        RECT 1167.780 2794.300 1168.100 2794.620 ;
        RECT 1172.380 2794.300 1172.700 2794.620 ;
        RECT 1178.820 2794.300 1179.140 2794.620 ;
        RECT 1186.180 2794.300 1186.500 2794.620 ;
        RECT 1198.140 2794.300 1198.460 2794.620 ;
        RECT 1587.300 2794.300 1587.620 2794.620 ;
        RECT 1594.660 2794.300 1594.980 2794.620 ;
        RECT 1601.100 2794.300 1601.420 2794.620 ;
        RECT 1631.460 2794.300 1631.780 2794.620 ;
        RECT 1637.900 2794.300 1638.220 2794.620 ;
        RECT 1648.020 2794.300 1648.340 2794.620 ;
        RECT 1655.380 2794.300 1655.700 2794.620 ;
        RECT 1659.060 2794.300 1659.380 2794.620 ;
        RECT 1666.420 2794.300 1666.740 2794.620 ;
        RECT 1672.860 2794.300 1673.180 2794.620 ;
        RECT 1679.300 2794.300 1679.620 2794.620 ;
        RECT 1683.900 2794.300 1684.220 2794.620 ;
        RECT 1688.500 2794.300 1688.820 2794.620 ;
        RECT 1695.860 2794.300 1696.180 2794.620 ;
        RECT 1702.300 2794.300 1702.620 2794.620 ;
        RECT 1708.740 2794.300 1709.060 2794.620 ;
        RECT 1713.340 2794.300 1713.660 2794.620 ;
        RECT 1719.780 2794.300 1720.100 2794.620 ;
        RECT 1721.620 2794.300 1721.940 2794.620 ;
        RECT 1730.820 2794.300 1731.140 2794.620 ;
        RECT 1737.260 2794.300 1737.580 2794.620 ;
        RECT 1743.700 2794.300 1744.020 2794.620 ;
        RECT 1748.300 2794.300 1748.620 2794.620 ;
        RECT 1762.100 2794.300 1762.420 2794.620 ;
        RECT 1780.500 2794.300 1780.820 2794.620 ;
        RECT 2231.300 2794.300 2231.620 2794.620 ;
        RECT 2257.060 2794.300 2257.380 2794.620 ;
        RECT 2264.420 2794.300 2264.740 2794.620 ;
        RECT 2268.100 2794.300 2268.420 2794.620 ;
        RECT 2276.380 2794.300 2276.700 2794.620 ;
        RECT 2282.820 2794.300 2283.140 2794.620 ;
        RECT 2287.420 2794.300 2287.740 2794.620 ;
        RECT 2293.860 2794.300 2294.180 2794.620 ;
        RECT 2300.300 2794.300 2300.620 2794.620 ;
        RECT 2304.900 2794.300 2305.220 2794.620 ;
        RECT 2308.580 2794.300 2308.900 2794.620 ;
        RECT 2316.860 2794.300 2317.180 2794.620 ;
        RECT 2322.380 2794.300 2322.700 2794.620 ;
        RECT 2328.820 2794.300 2329.140 2794.620 ;
        RECT 2334.340 2794.300 2334.660 2794.620 ;
        RECT 2339.860 2794.300 2340.180 2794.620 ;
        RECT 2343.540 2794.300 2343.860 2794.620 ;
        RECT 2351.820 2794.300 2352.140 2794.620 ;
        RECT 2357.340 2794.300 2357.660 2794.620 ;
        RECT 2363.780 2794.300 2364.100 2794.620 ;
        RECT 2370.220 2794.300 2370.540 2794.620 ;
        RECT 2374.820 2794.300 2375.140 2794.620 ;
        RECT 2377.580 2794.300 2377.900 2794.620 ;
        RECT 2381.260 2794.300 2381.580 2794.620 ;
        RECT 2383.100 2794.300 2383.420 2794.620 ;
        RECT 2389.540 2794.300 2389.860 2794.620 ;
        RECT 2395.060 2794.300 2395.380 2794.620 ;
        RECT 2402.420 2794.300 2402.740 2794.620 ;
        RECT 1087.740 2793.620 1088.060 2793.940 ;
        RECT 1118.100 2793.620 1118.420 2793.940 ;
        RECT 1128.220 2793.620 1128.540 2793.940 ;
        RECT 1159.500 2793.620 1159.820 2793.940 ;
        RECT 1163.180 2793.620 1163.500 2793.940 ;
        RECT 1173.300 2793.620 1173.620 2793.940 ;
        RECT 1180.660 2793.620 1180.980 2793.940 ;
        RECT 1187.100 2793.620 1187.420 2793.940 ;
        RECT 1604.780 2793.620 1605.100 2793.940 ;
        RECT 1613.060 2793.620 1613.380 2793.940 ;
        RECT 1630.540 2793.620 1630.860 2793.940 ;
        RECT 1644.340 2793.620 1644.660 2793.940 ;
        RECT 1652.620 2793.620 1652.940 2793.940 ;
        RECT 1665.500 2793.620 1665.820 2793.940 ;
        RECT 1670.100 2793.620 1670.420 2793.940 ;
        RECT 1677.460 2793.620 1677.780 2793.940 ;
        RECT 1682.980 2793.620 1683.300 2793.940 ;
        RECT 1689.420 2793.620 1689.740 2793.940 ;
        RECT 1694.940 2793.620 1695.260 2793.940 ;
        RECT 1699.540 2793.620 1699.860 2793.940 ;
        RECT 1705.980 2793.620 1706.300 2793.940 ;
        RECT 1712.420 2793.620 1712.740 2793.940 ;
        RECT 1717.940 2793.620 1718.260 2793.940 ;
        RECT 1729.900 2793.620 1730.220 2793.940 ;
        RECT 1734.500 2793.620 1734.820 2793.940 ;
        RECT 1740.940 2793.620 1741.260 2793.940 ;
        RECT 1747.380 2793.620 1747.700 2793.940 ;
        RECT 1767.620 2793.620 1767.940 2793.940 ;
        RECT 1774.060 2793.620 1774.380 2793.940 ;
        RECT 2269.020 2793.620 2269.340 2793.940 ;
        RECT 2273.620 2793.620 2273.940 2793.940 ;
        RECT 2280.060 2793.620 2280.380 2793.940 ;
        RECT 2286.500 2793.620 2286.820 2793.940 ;
        RECT 2292.020 2793.620 2292.340 2793.940 ;
        RECT 2310.420 2793.620 2310.740 2793.940 ;
        RECT 2315.020 2793.620 2315.340 2793.940 ;
        RECT 2321.460 2793.620 2321.780 2793.940 ;
        RECT 2326.060 2793.620 2326.380 2793.940 ;
        RECT 2332.500 2793.620 2332.820 2793.940 ;
        RECT 2345.380 2793.620 2345.700 2793.940 ;
        RECT 2356.420 2793.620 2356.740 2793.940 ;
        RECT 2361.020 2793.620 2361.340 2793.940 ;
        RECT 2367.460 2793.620 2367.780 2793.940 ;
        RECT 2373.900 2793.620 2374.220 2793.940 ;
        RECT 2423.580 2793.620 2423.900 2793.940 ;
        RECT 348.980 2792.940 349.300 2793.260 ;
        RECT 379.340 2792.940 379.660 2793.260 ;
        RECT 392.220 2792.940 392.540 2793.260 ;
        RECT 396.820 2792.940 397.140 2793.260 ;
        RECT 427.180 2792.940 427.500 2793.260 ;
        RECT 430.860 2792.940 431.180 2793.260 ;
        RECT 455.700 2792.940 456.020 2793.260 ;
        RECT 465.820 2792.940 466.140 2793.260 ;
        RECT 474.100 2792.940 474.420 2793.260 ;
        RECT 531.140 2792.940 531.460 2793.260 ;
        RECT 1012.300 2792.940 1012.620 2793.260 ;
        RECT 1024.260 2792.940 1024.580 2793.260 ;
        RECT 1048.180 2792.940 1048.500 2793.260 ;
        RECT 1617.660 2792.940 1617.980 2793.260 ;
        RECT 1624.100 2792.940 1624.420 2793.260 ;
        RECT 1635.140 2792.940 1635.460 2793.260 ;
        RECT 1642.500 2792.940 1642.820 2793.260 ;
        RECT 2263.500 2792.940 2263.820 2793.260 ;
        RECT 2297.540 2792.940 2297.860 2793.260 ;
        RECT 2338.940 2792.940 2339.260 2793.260 ;
        RECT 2349.980 2792.940 2350.300 2793.260 ;
        RECT 2386.780 2792.940 2387.100 2793.260 ;
        RECT 2407.940 2792.940 2408.260 2793.260 ;
        RECT 498.020 2792.260 498.340 2792.580 ;
        RECT 543.100 2792.260 543.420 2792.580 ;
        RECT 544.940 2792.260 545.260 2792.580 ;
        RECT 1164.100 2792.260 1164.420 2792.580 ;
        RECT 1752.900 2792.260 1753.220 2792.580 ;
        RECT 1787.860 2792.260 1788.180 2792.580 ;
        RECT 2398.740 2792.260 2399.060 2792.580 ;
        RECT 2410.700 2792.260 2411.020 2792.580 ;
        RECT 2415.300 2792.260 2415.620 2792.580 ;
        RECT 2430.020 2792.260 2430.340 2792.580 ;
        RECT 2436.460 2792.260 2436.780 2792.580 ;
        RECT 986.540 2791.580 986.860 2791.900 ;
        RECT 1153.060 2791.580 1153.380 2791.900 ;
        RECT 1193.540 2791.580 1193.860 2791.900 ;
        RECT 1411.580 2791.580 1411.900 2791.900 ;
        RECT 2236.820 2791.580 2237.140 2791.900 ;
        RECT 2392.300 2791.580 2392.620 2791.900 ;
        RECT 2404.260 2791.580 2404.580 2791.900 ;
        RECT 2442.900 2791.580 2443.220 2791.900 ;
        RECT 993.900 2790.900 994.220 2791.220 ;
        RECT 1417.100 2790.900 1417.420 2791.220 ;
        RECT 2242.340 2790.900 2242.660 2791.220 ;
        RECT 2420.820 2790.900 2421.140 2791.220 ;
        RECT 1191.700 2790.220 1192.020 2790.540 ;
        RECT 1613.980 2790.220 1614.300 2790.540 ;
        RECT 1620.420 2790.220 1620.740 2790.540 ;
        RECT 2428.180 2790.220 2428.500 2790.540 ;
        RECT 413.380 2789.540 413.700 2789.860 ;
        RECT 538.500 2789.540 538.820 2789.860 ;
        RECT 1648.940 2789.540 1649.260 2789.860 ;
        RECT 2417.140 2789.540 2417.460 2789.860 ;
        RECT 2434.620 2789.540 2434.940 2789.860 ;
        RECT 508.140 2788.860 508.460 2789.180 ;
        RECT 1581.780 2788.860 1582.100 2789.180 ;
        RECT 1661.820 2788.860 1662.140 2789.180 ;
        RECT 2249.700 2788.860 2250.020 2789.180 ;
        RECT 2418.060 2788.860 2418.380 2789.180 ;
        RECT 2439.220 2788.860 2439.540 2789.180 ;
        RECT 500.780 2788.180 501.100 2788.500 ;
        RECT 531.140 2788.180 531.460 2788.500 ;
        RECT 1007.700 2788.180 1008.020 2788.500 ;
        RECT 1035.300 2788.180 1035.620 2788.500 ;
        RECT 1051.860 2788.180 1052.180 2788.500 ;
        RECT 1086.820 2788.180 1087.140 2788.500 ;
        RECT 1626.860 2788.180 1627.180 2788.500 ;
        RECT 1724.380 2788.180 1724.700 2788.500 ;
        RECT 1765.780 2788.180 1766.100 2788.500 ;
        RECT 2303.980 2788.180 2304.300 2788.500 ;
        RECT 2445.660 2788.180 2445.980 2788.500 ;
        RECT 507.220 2787.500 507.540 2787.820 ;
        RECT 513.660 2787.500 513.980 2787.820 ;
        RECT 516.420 2787.500 516.740 2787.820 ;
        RECT 520.100 2787.500 520.420 2787.820 ;
        RECT 526.540 2787.500 526.860 2787.820 ;
        RECT 530.220 2787.500 530.540 2787.820 ;
        RECT 1034.380 2787.500 1034.700 2787.820 ;
        RECT 1039.900 2787.500 1040.220 2787.820 ;
        RECT 1046.340 2787.500 1046.660 2787.820 ;
        RECT 1061.980 2787.500 1062.300 2787.820 ;
        RECT 1067.500 2787.500 1067.820 2787.820 ;
        RECT 1073.940 2787.500 1074.260 2787.820 ;
        RECT 1081.300 2787.500 1081.620 2787.820 ;
        RECT 1089.580 2787.500 1089.900 2787.820 ;
        RECT 1096.020 2787.500 1096.340 2787.820 ;
        RECT 1103.380 2787.500 1103.700 2787.820 ;
        RECT 1109.820 2787.500 1110.140 2787.820 ;
        RECT 1116.260 2787.500 1116.580 2787.820 ;
        RECT 1121.780 2787.500 1122.100 2787.820 ;
        RECT 1754.740 2787.500 1755.060 2787.820 ;
        RECT 1772.220 2787.500 1772.540 2787.820 ;
        RECT 1778.660 2787.500 1778.980 2787.820 ;
        RECT 1783.260 2787.500 1783.580 2787.820 ;
        RECT 1789.700 2787.500 1790.020 2787.820 ;
        RECT 1761.180 2777.300 1761.500 2777.620 ;
        RECT 1796.140 2777.300 1796.460 2777.620 ;
        RECT 1841.220 2069.420 1841.540 2069.740 ;
        RECT 1844.900 2069.420 1845.220 2069.740 ;
        RECT 1851.340 2069.420 1851.660 2069.740 ;
        RECT 1859.620 2069.420 1859.940 2069.740 ;
        RECT 1865.140 2069.420 1865.460 2069.740 ;
        RECT 1901.020 2069.420 1901.340 2069.740 ;
        RECT 1923.100 2069.420 1923.420 2069.740 ;
        RECT 1941.500 2069.420 1941.820 2069.740 ;
        RECT 1953.460 2069.420 1953.780 2069.740 ;
        RECT 1964.500 2069.420 1964.820 2069.740 ;
        RECT 1947.020 2068.060 1947.340 2068.380 ;
        RECT 1960.820 2068.740 1961.140 2069.060 ;
        RECT 1989.340 2069.420 1989.660 2069.740 ;
        RECT 2015.100 2069.420 2015.420 2069.740 ;
        RECT 2039.020 2069.420 2039.340 2069.740 ;
        RECT 2052.820 2069.420 2053.140 2069.740 ;
        RECT 2354.580 2069.420 2354.900 2069.740 ;
        RECT 2373.900 2069.420 2374.220 2069.740 ;
        RECT 2391.380 2069.420 2391.700 2069.740 ;
        RECT 1980.140 2068.740 1980.460 2069.060 ;
        RECT 2381.260 2068.740 2381.580 2069.060 ;
        RECT 2387.700 2068.740 2388.020 2069.060 ;
        RECT 2528.460 2068.740 2528.780 2069.060 ;
        RECT 2396.900 2068.060 2397.220 2068.380 ;
        RECT 2534.900 2068.060 2535.220 2068.380 ;
        RECT 1932.300 2067.380 1932.620 2067.700 ;
        RECT 1946.100 2067.380 1946.420 2067.700 ;
        RECT 1907.460 2066.700 1907.780 2067.020 ;
        RECT 1912.060 2066.700 1912.380 2067.020 ;
        RECT 1871.580 2066.020 1871.900 2066.340 ;
        RECT 1877.100 2066.020 1877.420 2066.340 ;
        RECT 1879.860 2066.020 1880.180 2066.340 ;
        RECT 1889.060 2066.020 1889.380 2066.340 ;
        RECT 1894.580 2066.020 1894.900 2066.340 ;
        RECT 1935.980 2066.020 1936.300 2066.340 ;
        RECT 1973.700 2067.380 1974.020 2067.700 ;
        RECT 2007.740 2067.380 2008.060 2067.700 ;
        RECT 2021.540 2067.380 2021.860 2067.700 ;
        RECT 2403.340 2067.380 2403.660 2067.700 ;
        RECT 2429.100 2067.380 2429.420 2067.700 ;
        RECT 1987.500 2066.700 1987.820 2067.020 ;
        RECT 2011.420 2066.700 2011.740 2067.020 ;
        RECT 2409.780 2066.700 2410.100 2067.020 ;
        RECT 2417.140 2066.700 2417.460 2067.020 ;
        RECT 2023.380 2066.020 2023.700 2066.340 ;
        RECT 2422.660 2066.020 2422.980 2066.340 ;
        RECT 2442.900 2066.020 2443.220 2066.340 ;
        RECT 1847.660 2065.340 1847.980 2065.660 ;
        RECT 1854.100 2065.340 1854.420 2065.660 ;
        RECT 1882.620 2065.340 1882.940 2065.660 ;
        RECT 1911.140 2065.340 1911.460 2065.660 ;
        RECT 1913.900 2065.340 1914.220 2065.660 ;
        RECT 1925.860 2065.340 1926.180 2065.660 ;
        RECT 1958.980 2065.340 1959.300 2065.660 ;
        RECT 1990.260 2065.340 1990.580 2065.660 ;
        RECT 1999.460 2065.340 1999.780 2065.660 ;
        RECT 2436.460 2065.340 2436.780 2065.660 ;
        RECT 1948.860 2064.660 1949.180 2064.980 ;
        RECT 1955.300 2064.660 1955.620 2064.980 ;
        RECT 1967.260 2064.660 1967.580 2064.980 ;
        RECT 1981.980 2064.660 1982.300 2064.980 ;
        RECT 1993.020 2064.660 1993.340 2064.980 ;
        RECT 2450.260 2064.660 2450.580 2064.980 ;
        RECT 2456.700 2064.660 2457.020 2064.980 ;
        RECT 1869.740 2063.980 1870.060 2064.300 ;
        RECT 1886.300 2063.980 1886.620 2064.300 ;
        RECT 1890.900 2063.980 1891.220 2064.300 ;
        RECT 1898.260 2063.980 1898.580 2064.300 ;
        RECT 1976.460 2063.980 1976.780 2064.300 ;
        RECT 2002.220 2063.980 2002.540 2064.300 ;
        RECT 2016.940 2063.980 2017.260 2064.300 ;
        RECT 1838.460 2063.300 1838.780 2063.620 ;
        RECT 1856.860 2063.300 1857.180 2063.620 ;
        RECT 1863.300 2063.300 1863.620 2063.620 ;
        RECT 1873.420 2063.300 1873.740 2063.620 ;
        RECT 1904.700 2063.300 1905.020 2063.620 ;
        RECT 1917.580 2063.300 1917.900 2063.620 ;
        RECT 1920.340 2063.300 1920.660 2063.620 ;
        RECT 1929.540 2063.300 1929.860 2063.620 ;
        RECT 1940.580 2063.300 1940.900 2063.620 ;
        RECT 1970.940 2063.300 1971.260 2063.620 ;
        RECT 1995.780 2063.300 1996.100 2063.620 ;
        RECT 2005.900 2063.300 2006.220 2063.620 ;
        RECT 2340.780 2063.300 2341.100 2063.620 ;
        RECT 2347.220 2063.300 2347.540 2063.620 ;
        RECT 2360.100 2063.300 2360.420 2063.620 ;
        RECT 2459.460 2063.300 2459.780 2063.620 ;
        RECT 2465.900 2063.300 2466.220 2063.620 ;
        RECT 2472.340 2063.300 2472.660 2063.620 ;
        RECT 2478.780 2063.300 2479.100 2063.620 ;
        RECT 2484.300 2063.300 2484.620 2063.620 ;
        RECT 2491.660 2063.300 2491.980 2063.620 ;
        RECT 2498.100 2063.300 2498.420 2063.620 ;
        RECT 2505.460 2063.300 2505.780 2063.620 ;
        RECT 2513.740 2063.300 2514.060 2063.620 ;
        RECT 2518.340 2063.300 2518.660 2063.620 ;
        RECT 2522.020 2063.300 2522.340 2063.620 ;
        RECT 2590.100 2063.300 2590.420 2063.620 ;
        RECT 2028.800 2057.180 2029.120 2057.500 ;
        RECT 2367.230 2051.740 2367.550 2052.060 ;
        RECT 1417.100 1621.980 1417.420 1622.300 ;
        RECT 1411.580 1617.220 1411.900 1617.540 ;
        RECT 2103.420 1745.740 2103.740 1746.060 ;
        RECT 2099.740 1732.820 2100.060 1733.140 ;
        RECT 2103.420 1732.140 2103.740 1732.460 ;
        RECT 2114.460 1732.140 2114.780 1732.460 ;
        RECT 2139.300 1732.140 2139.620 1732.460 ;
        RECT 2234.060 1732.140 2234.380 1732.460 ;
        RECT 2238.660 1732.140 2238.980 1732.460 ;
        RECT 2189.900 1728.740 2190.220 1729.060 ;
        RECT 2235.900 1728.740 2236.220 1729.060 ;
        RECT 2188.980 1721.940 2189.300 1722.260 ;
        RECT 2103.420 1718.540 2103.740 1718.860 ;
        RECT 2188.060 1715.140 2188.380 1715.460 ;
        RECT 2240.500 1715.140 2240.820 1715.460 ;
        RECT 2247.860 1715.140 2248.180 1715.460 ;
        RECT 2253.380 1715.140 2253.700 1715.460 ;
        RECT 2102.500 1708.340 2102.820 1708.660 ;
        RECT 2139.300 1705.620 2139.620 1705.940 ;
        RECT 2197.260 1705.620 2197.580 1705.940 ;
        RECT 2102.500 1704.940 2102.820 1705.260 ;
        RECT 2222.100 1701.540 2222.420 1701.860 ;
        RECT 2227.620 1701.540 2227.940 1701.860 ;
        RECT 2637.940 1745.740 2638.260 1746.060 ;
        RECT 2639.780 1735.540 2640.100 1735.860 ;
        RECT 2637.940 1732.140 2638.260 1732.460 ;
        RECT 2637.940 1724.260 2638.260 1724.580 ;
        RECT 2639.780 1715.820 2640.100 1716.140 ;
        RECT 2637.940 1709.700 2638.260 1710.020 ;
        RECT 2637.940 1708.340 2638.260 1708.660 ;
      LAYER met4 ;
        RECT 1890.895 3264.175 1891.225 3264.505 ;
        RECT 1917.575 3264.175 1917.905 3264.505 ;
        RECT 2542.255 3264.175 2542.585 3264.505 ;
        RECT 2567.095 3264.175 2567.425 3264.505 ;
        RECT 1292.875 3258.055 1293.205 3258.385 ;
        RECT 1317.850 3258.055 1318.180 3258.385 ;
        RECT 394.025 3251.635 394.325 3256.235 ;
        RECT 400.265 3251.635 400.565 3256.235 ;
        RECT 406.505 3251.635 406.805 3256.235 ;
        RECT 412.745 3251.635 413.045 3256.235 ;
        RECT 418.985 3251.635 419.285 3256.235 ;
        RECT 425.225 3251.635 425.525 3256.235 ;
        RECT 431.465 3251.635 431.765 3256.235 ;
        RECT 437.705 3251.635 438.005 3256.235 ;
        RECT 443.945 3251.635 444.245 3256.235 ;
        RECT 450.185 3251.635 450.485 3256.235 ;
        RECT 456.425 3251.635 456.725 3256.235 ;
        RECT 462.665 3251.635 462.965 3256.235 ;
        RECT 468.905 3251.635 469.205 3256.235 ;
        RECT 475.145 3251.635 475.445 3256.235 ;
        RECT 481.385 3251.635 481.685 3256.235 ;
        RECT 487.625 3251.635 487.925 3256.235 ;
        RECT 493.865 3251.635 494.165 3256.235 ;
        RECT 500.105 3251.635 500.405 3256.235 ;
        RECT 506.345 3251.635 506.645 3256.235 ;
        RECT 512.585 3251.635 512.885 3256.235 ;
        RECT 518.825 3251.635 519.125 3256.235 ;
        RECT 525.065 3251.635 525.365 3256.235 ;
        RECT 531.305 3251.635 531.605 3256.235 ;
        RECT 537.545 3251.635 537.845 3256.235 ;
        RECT 543.785 3251.635 544.085 3256.235 ;
        RECT 550.025 3251.635 550.325 3256.235 ;
        RECT 556.265 3251.635 556.565 3256.235 ;
        RECT 562.505 3251.635 562.805 3256.235 ;
        RECT 568.745 3251.635 569.045 3256.235 ;
        RECT 574.985 3251.635 575.285 3256.235 ;
        RECT 581.225 3251.635 581.525 3256.235 ;
        RECT 587.465 3251.635 587.765 3256.235 ;
        RECT 642.890 3255.650 643.190 3256.235 ;
        RECT 646.135 3255.650 646.465 3255.665 ;
        RECT 642.890 3255.350 646.465 3255.650 ;
        RECT 642.890 3251.635 643.190 3255.350 ;
        RECT 646.135 3255.335 646.465 3255.350 ;
        RECT 667.865 3253.950 668.165 3256.235 ;
        RECT 669.135 3255.335 669.465 3255.665 ;
        RECT 669.150 3253.950 669.450 3255.335 ;
        RECT 667.865 3253.650 669.450 3253.950 ;
        RECT 667.865 3251.635 668.165 3253.650 ;
        RECT 1044.025 3251.635 1044.325 3256.235 ;
        RECT 1050.265 3251.635 1050.565 3256.235 ;
        RECT 1056.505 3251.635 1056.805 3256.235 ;
        RECT 1062.745 3251.635 1063.045 3256.235 ;
        RECT 1068.985 3251.635 1069.285 3256.235 ;
        RECT 1075.225 3251.635 1075.525 3256.235 ;
        RECT 1081.465 3251.635 1081.765 3256.235 ;
        RECT 1087.705 3251.635 1088.005 3256.235 ;
        RECT 1093.945 3251.635 1094.245 3256.235 ;
        RECT 1100.185 3251.635 1100.485 3256.235 ;
        RECT 1106.425 3251.635 1106.725 3256.235 ;
        RECT 1112.665 3251.635 1112.965 3256.235 ;
        RECT 1118.905 3251.635 1119.205 3256.235 ;
        RECT 1125.145 3251.635 1125.445 3256.235 ;
        RECT 1131.385 3251.635 1131.685 3256.235 ;
        RECT 1137.625 3251.635 1137.925 3256.235 ;
        RECT 1143.865 3251.635 1144.165 3256.235 ;
        RECT 1150.105 3251.635 1150.405 3256.235 ;
        RECT 1156.345 3251.635 1156.645 3256.235 ;
        RECT 1162.585 3251.635 1162.885 3256.235 ;
        RECT 1168.825 3251.635 1169.125 3256.235 ;
        RECT 1175.065 3251.635 1175.365 3256.235 ;
        RECT 1181.305 3251.635 1181.605 3256.235 ;
        RECT 1187.545 3251.635 1187.845 3256.235 ;
        RECT 1193.785 3251.635 1194.085 3256.235 ;
        RECT 1200.025 3251.635 1200.325 3256.235 ;
        RECT 1206.265 3251.635 1206.565 3256.235 ;
        RECT 1212.505 3251.635 1212.805 3256.235 ;
        RECT 1218.745 3251.635 1219.045 3256.235 ;
        RECT 1224.985 3251.635 1225.285 3256.235 ;
        RECT 1231.225 3251.635 1231.525 3256.235 ;
        RECT 1237.465 3251.635 1237.765 3256.235 ;
        RECT 1292.890 3251.635 1293.190 3258.055 ;
        RECT 1317.865 3251.635 1318.165 3258.055 ;
        RECT 1644.025 3251.635 1644.325 3256.235 ;
        RECT 1650.265 3251.635 1650.565 3256.235 ;
        RECT 1656.505 3251.635 1656.805 3256.235 ;
        RECT 1662.745 3251.635 1663.045 3256.235 ;
        RECT 1668.985 3251.635 1669.285 3256.235 ;
        RECT 1675.225 3251.635 1675.525 3256.235 ;
        RECT 1681.465 3251.635 1681.765 3256.235 ;
        RECT 1687.705 3251.635 1688.005 3256.235 ;
        RECT 1693.945 3251.635 1694.245 3256.235 ;
        RECT 1700.185 3251.635 1700.485 3256.235 ;
        RECT 1706.425 3251.635 1706.725 3256.235 ;
        RECT 1712.665 3251.635 1712.965 3256.235 ;
        RECT 1718.905 3251.635 1719.205 3256.235 ;
        RECT 1725.145 3251.635 1725.445 3256.235 ;
        RECT 1731.385 3251.635 1731.685 3256.235 ;
        RECT 1737.625 3251.635 1737.925 3256.235 ;
        RECT 1743.865 3251.635 1744.165 3256.235 ;
        RECT 1750.105 3251.635 1750.405 3256.235 ;
        RECT 1756.345 3251.635 1756.645 3256.235 ;
        RECT 1762.585 3251.635 1762.885 3256.235 ;
        RECT 1768.825 3251.635 1769.125 3256.235 ;
        RECT 1775.065 3251.635 1775.365 3256.235 ;
        RECT 1781.305 3251.635 1781.605 3256.235 ;
        RECT 1787.545 3251.635 1787.845 3256.235 ;
        RECT 1793.785 3251.635 1794.085 3256.235 ;
        RECT 1800.025 3251.635 1800.325 3256.235 ;
        RECT 1806.265 3251.635 1806.565 3256.235 ;
        RECT 1812.505 3251.635 1812.805 3256.235 ;
        RECT 1818.745 3251.635 1819.045 3256.235 ;
        RECT 1824.985 3251.635 1825.285 3256.235 ;
        RECT 1831.225 3251.635 1831.525 3256.235 ;
        RECT 1837.465 3251.635 1837.765 3256.235 ;
        RECT 1890.910 3255.650 1891.210 3264.175 ;
        RECT 1917.590 3256.235 1917.890 3264.175 ;
        RECT 1892.890 3255.650 1893.190 3256.235 ;
        RECT 1890.910 3255.350 1893.190 3255.650 ;
        RECT 1917.590 3255.350 1918.165 3256.235 ;
        RECT 1892.890 3251.635 1893.190 3255.350 ;
        RECT 1917.865 3251.635 1918.165 3255.350 ;
        RECT 2294.025 3251.635 2294.325 3256.235 ;
        RECT 2300.265 3251.635 2300.565 3256.235 ;
        RECT 2306.505 3251.635 2306.805 3256.235 ;
        RECT 2312.745 3251.635 2313.045 3256.235 ;
        RECT 2318.985 3251.635 2319.285 3256.235 ;
        RECT 2325.225 3251.635 2325.525 3256.235 ;
        RECT 2331.465 3251.635 2331.765 3256.235 ;
        RECT 2337.705 3251.635 2338.005 3256.235 ;
        RECT 2343.945 3251.635 2344.245 3256.235 ;
        RECT 2350.185 3251.635 2350.485 3256.235 ;
        RECT 2356.425 3251.635 2356.725 3256.235 ;
        RECT 2362.665 3251.635 2362.965 3256.235 ;
        RECT 2368.905 3251.635 2369.205 3256.235 ;
        RECT 2375.145 3251.635 2375.445 3256.235 ;
        RECT 2381.385 3251.635 2381.685 3256.235 ;
        RECT 2387.625 3251.635 2387.925 3256.235 ;
        RECT 2393.865 3251.635 2394.165 3256.235 ;
        RECT 2400.105 3251.635 2400.405 3256.235 ;
        RECT 2406.345 3251.635 2406.645 3256.235 ;
        RECT 2412.585 3251.635 2412.885 3256.235 ;
        RECT 2418.825 3251.635 2419.125 3256.235 ;
        RECT 2425.065 3251.635 2425.365 3256.235 ;
        RECT 2431.305 3251.635 2431.605 3256.235 ;
        RECT 2437.545 3251.635 2437.845 3256.235 ;
        RECT 2443.785 3251.635 2444.085 3256.235 ;
        RECT 2450.025 3251.635 2450.325 3256.235 ;
        RECT 2456.265 3251.635 2456.565 3256.235 ;
        RECT 2462.505 3251.635 2462.805 3256.235 ;
        RECT 2468.745 3251.635 2469.045 3256.235 ;
        RECT 2474.985 3251.635 2475.285 3256.235 ;
        RECT 2481.225 3251.635 2481.525 3256.235 ;
        RECT 2487.465 3251.635 2487.765 3256.235 ;
        RECT 2542.270 3255.650 2542.570 3264.175 ;
        RECT 2542.890 3255.650 2543.190 3256.235 ;
        RECT 2542.270 3255.350 2543.190 3255.650 ;
        RECT 2567.110 3255.650 2567.410 3264.175 ;
        RECT 2567.865 3255.650 2568.165 3256.235 ;
        RECT 2567.110 3255.350 2568.165 3255.650 ;
        RECT 2542.890 3251.635 2543.190 3255.350 ;
        RECT 2567.865 3251.635 2568.165 3255.350 ;
        RECT 302.550 2894.510 303.730 2895.690 ;
      LAYER met4 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met4 ;
        RECT 943.790 2894.510 944.970 2895.690 ;
      LAYER met4 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met4 ;
        RECT 1351.350 2935.310 1352.530 2936.490 ;
        RECT 1412.070 2894.510 1413.250 2895.690 ;
        RECT 1550.990 2894.510 1552.170 2895.690 ;
      LAYER met4 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met4 ;
        RECT 1937.390 2935.310 1938.570 2936.490 ;
        RECT 1946.095 2904.455 1946.425 2904.785 ;
        RECT 1946.110 2899.090 1946.410 2904.455 ;
        RECT 1945.670 2897.910 1946.850 2899.090 ;
        RECT 2186.710 2894.510 2187.890 2895.690 ;
      LAYER met4 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met4 ;
        RECT 2594.695 2904.455 2595.025 2904.785 ;
        RECT 2594.710 2899.090 2595.010 2904.455 ;
        RECT 2594.270 2897.910 2595.450 2899.090 ;
        RECT 334.010 2801.750 334.310 2804.600 ;
        RECT 339.850 2801.750 340.150 2804.600 ;
        RECT 345.690 2801.750 345.990 2804.600 ;
        RECT 351.530 2801.750 351.830 2804.600 ;
        RECT 334.010 2801.450 337.330 2801.750 ;
        RECT 334.010 2800.000 334.310 2801.450 ;
        RECT 337.030 2794.625 337.330 2801.450 ;
        RECT 339.850 2801.450 342.850 2801.750 ;
        RECT 339.850 2800.000 340.150 2801.450 ;
        RECT 342.550 2794.625 342.850 2801.450 ;
        RECT 345.690 2801.450 349.290 2801.750 ;
        RECT 345.690 2800.000 345.990 2801.450 ;
        RECT 337.015 2794.295 337.345 2794.625 ;
        RECT 342.535 2794.295 342.865 2794.625 ;
        RECT 348.990 2793.265 349.290 2801.450 ;
        RECT 350.830 2801.450 351.830 2801.750 ;
        RECT 350.830 2794.625 351.130 2801.450 ;
        RECT 351.530 2800.000 351.830 2801.450 ;
        RECT 357.370 2801.750 357.670 2804.600 ;
        RECT 363.210 2802.450 363.510 2804.600 ;
        RECT 361.870 2802.150 363.510 2802.450 ;
        RECT 357.370 2801.450 358.490 2801.750 ;
        RECT 357.370 2800.000 357.670 2801.450 ;
        RECT 358.190 2794.625 358.490 2801.450 ;
        RECT 361.870 2794.625 362.170 2802.150 ;
        RECT 363.210 2800.000 363.510 2802.150 ;
        RECT 363.830 2801.750 364.130 2804.600 ;
        RECT 369.050 2801.750 369.350 2804.600 ;
        RECT 363.830 2801.450 364.930 2801.750 ;
        RECT 363.830 2800.000 364.130 2801.450 ;
        RECT 364.630 2794.625 364.930 2801.450 ;
        RECT 368.310 2801.450 369.350 2801.750 ;
        RECT 368.310 2794.625 368.610 2801.450 ;
        RECT 369.050 2800.000 369.350 2801.450 ;
        RECT 369.670 2801.750 369.970 2804.600 ;
        RECT 374.890 2801.750 375.190 2804.600 ;
        RECT 369.670 2801.450 371.370 2801.750 ;
        RECT 369.670 2800.000 369.970 2801.450 ;
        RECT 371.070 2794.625 371.370 2801.450 ;
        RECT 374.750 2800.000 375.190 2801.750 ;
        RECT 375.510 2801.750 375.810 2804.600 ;
        RECT 380.730 2801.750 381.030 2804.600 ;
        RECT 375.510 2801.450 378.730 2801.750 ;
        RECT 375.510 2800.000 375.810 2801.450 ;
        RECT 374.750 2794.625 375.050 2800.000 ;
        RECT 378.430 2794.625 378.730 2801.450 ;
        RECT 379.350 2801.450 381.030 2801.750 ;
        RECT 350.815 2794.295 351.145 2794.625 ;
        RECT 358.175 2794.295 358.505 2794.625 ;
        RECT 361.855 2794.295 362.185 2794.625 ;
        RECT 364.615 2794.295 364.945 2794.625 ;
        RECT 368.295 2794.295 368.625 2794.625 ;
        RECT 371.055 2794.295 371.385 2794.625 ;
        RECT 374.735 2794.295 375.065 2794.625 ;
        RECT 378.415 2794.295 378.745 2794.625 ;
        RECT 379.350 2793.265 379.650 2801.450 ;
        RECT 380.730 2800.000 381.030 2801.450 ;
        RECT 381.350 2801.750 381.650 2804.600 ;
        RECT 381.350 2801.450 384.250 2801.750 ;
        RECT 381.350 2800.000 381.650 2801.450 ;
        RECT 383.950 2794.625 384.250 2801.450 ;
        RECT 386.570 2796.650 386.870 2804.600 ;
        RECT 387.190 2801.750 387.490 2804.600 ;
        RECT 392.410 2801.750 392.710 2804.600 ;
        RECT 387.190 2801.450 390.690 2801.750 ;
        RECT 387.190 2800.000 387.490 2801.450 ;
        RECT 386.570 2796.350 387.010 2796.650 ;
        RECT 386.710 2794.625 387.010 2796.350 ;
        RECT 390.390 2794.625 390.690 2801.450 ;
        RECT 392.230 2800.000 392.710 2801.750 ;
        RECT 393.030 2801.750 393.330 2804.600 ;
        RECT 398.250 2802.450 398.550 2804.600 ;
        RECT 396.830 2802.150 398.550 2802.450 ;
        RECT 393.030 2801.450 396.210 2801.750 ;
        RECT 393.030 2800.000 393.330 2801.450 ;
        RECT 383.935 2794.295 384.265 2794.625 ;
        RECT 386.695 2794.295 387.025 2794.625 ;
        RECT 390.375 2794.295 390.705 2794.625 ;
        RECT 392.230 2793.265 392.530 2800.000 ;
        RECT 395.910 2794.625 396.210 2801.450 ;
        RECT 395.895 2794.295 396.225 2794.625 ;
        RECT 396.830 2793.265 397.130 2802.150 ;
        RECT 398.250 2800.000 398.550 2802.150 ;
        RECT 398.870 2801.750 399.170 2804.600 ;
        RECT 404.090 2801.750 404.390 2804.600 ;
        RECT 398.870 2801.450 399.890 2801.750 ;
        RECT 398.870 2800.000 399.170 2801.450 ;
        RECT 399.590 2794.625 399.890 2801.450 ;
        RECT 403.270 2801.450 404.390 2801.750 ;
        RECT 403.270 2794.625 403.570 2801.450 ;
        RECT 404.090 2800.000 404.390 2801.450 ;
        RECT 404.710 2801.750 405.010 2804.600 ;
        RECT 409.930 2801.750 410.230 2804.600 ;
        RECT 404.710 2801.450 406.330 2801.750 ;
        RECT 404.710 2800.000 405.010 2801.450 ;
        RECT 406.030 2794.625 406.330 2801.450 ;
        RECT 409.710 2800.000 410.230 2801.750 ;
        RECT 410.550 2801.750 410.850 2804.600 ;
        RECT 415.770 2802.450 416.070 2804.600 ;
        RECT 414.310 2802.150 416.070 2802.450 ;
        RECT 410.550 2801.450 413.690 2801.750 ;
        RECT 410.550 2800.000 410.850 2801.450 ;
        RECT 409.710 2794.625 410.010 2800.000 ;
        RECT 399.575 2794.295 399.905 2794.625 ;
        RECT 403.255 2794.295 403.585 2794.625 ;
        RECT 406.015 2794.295 406.345 2794.625 ;
        RECT 409.695 2794.295 410.025 2794.625 ;
        RECT 348.975 2792.935 349.305 2793.265 ;
        RECT 379.335 2792.935 379.665 2793.265 ;
        RECT 392.215 2792.935 392.545 2793.265 ;
        RECT 396.815 2792.935 397.145 2793.265 ;
        RECT 413.390 2789.865 413.690 2801.450 ;
        RECT 414.310 2794.625 414.610 2802.150 ;
        RECT 415.770 2800.000 416.070 2802.150 ;
        RECT 416.390 2801.750 416.690 2804.600 ;
        RECT 421.610 2801.750 421.910 2804.600 ;
        RECT 416.390 2801.450 419.210 2801.750 ;
        RECT 416.390 2800.000 416.690 2801.450 ;
        RECT 418.910 2794.625 419.210 2801.450 ;
        RECT 420.750 2801.450 421.910 2801.750 ;
        RECT 420.750 2794.625 421.050 2801.450 ;
        RECT 421.610 2800.000 421.910 2801.450 ;
        RECT 422.230 2801.750 422.530 2804.600 ;
        RECT 427.450 2801.750 427.750 2804.600 ;
        RECT 422.230 2801.450 425.650 2801.750 ;
        RECT 422.230 2800.000 422.530 2801.450 ;
        RECT 425.350 2794.625 425.650 2801.450 ;
        RECT 427.190 2800.000 427.750 2801.750 ;
        RECT 428.070 2801.750 428.370 2804.600 ;
        RECT 433.290 2802.450 433.590 2804.600 ;
        RECT 431.790 2802.150 433.590 2802.450 ;
        RECT 428.070 2801.450 431.170 2801.750 ;
        RECT 428.070 2800.000 428.370 2801.450 ;
        RECT 414.295 2794.295 414.625 2794.625 ;
        RECT 418.895 2794.295 419.225 2794.625 ;
        RECT 420.735 2794.295 421.065 2794.625 ;
        RECT 425.335 2794.295 425.665 2794.625 ;
        RECT 427.190 2793.265 427.490 2800.000 ;
        RECT 430.870 2793.265 431.170 2801.450 ;
        RECT 431.790 2794.625 432.090 2802.150 ;
        RECT 433.290 2800.000 433.590 2802.150 ;
        RECT 433.910 2796.650 434.210 2804.600 ;
        RECT 439.130 2800.050 439.430 2804.600 ;
        RECT 439.750 2801.750 440.050 2804.600 ;
        RECT 444.970 2801.750 445.270 2804.600 ;
        RECT 439.750 2801.450 441.290 2801.750 ;
        RECT 439.130 2799.750 439.450 2800.050 ;
        RECT 439.750 2800.000 440.050 2801.450 ;
        RECT 433.630 2796.350 434.210 2796.650 ;
        RECT 433.630 2794.625 433.930 2796.350 ;
        RECT 439.150 2794.625 439.450 2799.750 ;
        RECT 440.990 2794.625 441.290 2801.450 ;
        RECT 444.670 2800.000 445.270 2801.750 ;
        RECT 444.670 2794.625 444.970 2800.000 ;
        RECT 445.590 2794.625 445.890 2804.600 ;
        RECT 450.810 2801.750 451.110 2804.600 ;
        RECT 449.270 2801.450 451.110 2801.750 ;
        RECT 449.270 2794.625 449.570 2801.450 ;
        RECT 450.810 2800.000 451.110 2801.450 ;
        RECT 451.430 2801.750 451.730 2804.600 ;
        RECT 456.650 2801.750 456.950 2804.600 ;
        RECT 451.430 2801.450 455.090 2801.750 ;
        RECT 451.430 2800.000 451.730 2801.450 ;
        RECT 454.790 2794.625 455.090 2801.450 ;
        RECT 455.710 2801.450 456.950 2801.750 ;
        RECT 431.775 2794.295 432.105 2794.625 ;
        RECT 433.615 2794.295 433.945 2794.625 ;
        RECT 439.135 2794.295 439.465 2794.625 ;
        RECT 440.975 2794.295 441.305 2794.625 ;
        RECT 444.655 2794.295 444.985 2794.625 ;
        RECT 445.575 2794.295 445.905 2794.625 ;
        RECT 449.255 2794.295 449.585 2794.625 ;
        RECT 454.775 2794.295 455.105 2794.625 ;
        RECT 455.710 2793.265 456.010 2801.450 ;
        RECT 456.650 2800.000 456.950 2801.450 ;
        RECT 457.270 2801.750 457.570 2804.600 ;
        RECT 457.270 2801.450 459.690 2801.750 ;
        RECT 457.270 2800.000 457.570 2801.450 ;
        RECT 459.390 2794.625 459.690 2801.450 ;
        RECT 462.490 2800.050 462.790 2804.600 ;
        RECT 462.150 2799.750 462.790 2800.050 ;
        RECT 463.110 2801.750 463.410 2804.600 ;
        RECT 468.330 2801.750 468.630 2804.600 ;
        RECT 463.110 2801.450 466.130 2801.750 ;
        RECT 463.110 2800.000 463.410 2801.450 ;
        RECT 462.150 2794.625 462.450 2799.750 ;
        RECT 459.375 2794.295 459.705 2794.625 ;
        RECT 462.135 2794.295 462.465 2794.625 ;
        RECT 465.830 2793.265 466.130 2801.450 ;
        RECT 466.750 2801.450 468.630 2801.750 ;
        RECT 466.750 2794.625 467.050 2801.450 ;
        RECT 468.330 2800.000 468.630 2801.450 ;
        RECT 468.950 2796.650 469.250 2804.600 ;
        RECT 474.170 2801.750 474.470 2804.600 ;
        RECT 468.590 2796.350 469.250 2796.650 ;
        RECT 474.110 2800.000 474.470 2801.750 ;
        RECT 474.790 2801.750 475.090 2804.600 ;
        RECT 480.010 2801.750 480.310 2804.600 ;
        RECT 474.790 2800.000 475.330 2801.750 ;
        RECT 468.590 2794.625 468.890 2796.350 ;
        RECT 466.735 2794.295 467.065 2794.625 ;
        RECT 468.575 2794.295 468.905 2794.625 ;
        RECT 474.110 2793.265 474.410 2800.000 ;
        RECT 475.030 2794.625 475.330 2800.000 ;
        RECT 478.710 2801.450 480.310 2801.750 ;
        RECT 478.710 2794.625 479.010 2801.450 ;
        RECT 480.010 2800.000 480.310 2801.450 ;
        RECT 480.630 2801.750 480.930 2804.600 ;
        RECT 485.850 2801.750 486.150 2804.600 ;
        RECT 480.630 2801.450 482.690 2801.750 ;
        RECT 480.630 2800.000 480.930 2801.450 ;
        RECT 482.390 2794.625 482.690 2801.450 ;
        RECT 485.150 2801.450 486.150 2801.750 ;
        RECT 485.150 2794.625 485.450 2801.450 ;
        RECT 485.850 2800.000 486.150 2801.450 ;
        RECT 486.470 2801.750 486.770 2804.600 ;
        RECT 491.690 2801.750 491.990 2804.600 ;
        RECT 486.470 2801.450 489.130 2801.750 ;
        RECT 486.470 2800.000 486.770 2801.450 ;
        RECT 488.830 2794.625 489.130 2801.450 ;
        RECT 491.590 2800.000 491.990 2801.750 ;
        RECT 492.310 2801.750 492.610 2804.600 ;
        RECT 492.310 2801.450 495.570 2801.750 ;
        RECT 492.310 2800.000 492.610 2801.450 ;
        RECT 491.590 2794.625 491.890 2800.000 ;
        RECT 495.270 2794.625 495.570 2801.450 ;
        RECT 497.530 2796.650 497.830 2804.600 ;
        RECT 498.150 2801.750 498.450 2804.600 ;
        RECT 503.370 2801.750 503.670 2804.600 ;
        RECT 498.150 2801.450 500.170 2801.750 ;
        RECT 498.150 2800.000 498.450 2801.450 ;
        RECT 497.530 2796.350 498.330 2796.650 ;
        RECT 475.015 2794.295 475.345 2794.625 ;
        RECT 478.695 2794.295 479.025 2794.625 ;
        RECT 482.375 2794.295 482.705 2794.625 ;
        RECT 485.135 2794.295 485.465 2794.625 ;
        RECT 488.815 2794.295 489.145 2794.625 ;
        RECT 491.575 2794.295 491.905 2794.625 ;
        RECT 495.255 2794.295 495.585 2794.625 ;
        RECT 427.175 2792.935 427.505 2793.265 ;
        RECT 430.855 2792.935 431.185 2793.265 ;
        RECT 455.695 2792.935 456.025 2793.265 ;
        RECT 465.815 2792.935 466.145 2793.265 ;
        RECT 474.095 2792.935 474.425 2793.265 ;
        RECT 498.030 2792.585 498.330 2796.350 ;
        RECT 499.870 2794.625 500.170 2801.450 ;
        RECT 500.790 2801.450 503.670 2801.750 ;
        RECT 499.855 2794.295 500.185 2794.625 ;
        RECT 498.015 2792.255 498.345 2792.585 ;
        RECT 413.375 2789.535 413.705 2789.865 ;
        RECT 500.790 2788.505 501.090 2801.450 ;
        RECT 503.370 2800.000 503.670 2801.450 ;
        RECT 503.990 2801.750 504.290 2804.600 ;
        RECT 509.210 2801.750 509.510 2804.600 ;
        RECT 503.990 2801.450 507.530 2801.750 ;
        RECT 503.990 2800.000 504.290 2801.450 ;
        RECT 500.775 2788.175 501.105 2788.505 ;
        RECT 507.230 2787.825 507.530 2801.450 ;
        RECT 508.150 2801.450 509.510 2801.750 ;
        RECT 508.150 2789.185 508.450 2801.450 ;
        RECT 509.210 2800.000 509.510 2801.450 ;
        RECT 509.830 2801.750 510.130 2804.600 ;
        RECT 515.050 2802.450 515.350 2804.600 ;
        RECT 513.670 2802.150 515.350 2802.450 ;
        RECT 509.830 2800.000 510.290 2801.750 ;
        RECT 509.990 2794.625 510.290 2800.000 ;
        RECT 509.975 2794.295 510.305 2794.625 ;
        RECT 508.135 2788.855 508.465 2789.185 ;
        RECT 513.670 2787.825 513.970 2802.150 ;
        RECT 515.050 2800.000 515.350 2802.150 ;
        RECT 515.670 2801.750 515.970 2804.600 ;
        RECT 520.890 2801.750 521.190 2804.600 ;
        RECT 515.670 2801.450 516.730 2801.750 ;
        RECT 515.670 2800.000 515.970 2801.450 ;
        RECT 516.430 2787.825 516.730 2801.450 ;
        RECT 520.110 2801.450 521.190 2801.750 ;
        RECT 520.110 2787.825 520.410 2801.450 ;
        RECT 520.890 2800.000 521.190 2801.450 ;
        RECT 521.510 2801.750 521.810 2804.600 ;
        RECT 526.730 2801.750 527.030 2804.600 ;
        RECT 521.510 2801.450 524.090 2801.750 ;
        RECT 521.510 2800.000 521.810 2801.450 ;
        RECT 523.790 2794.625 524.090 2801.450 ;
        RECT 526.550 2800.000 527.030 2801.750 ;
        RECT 527.350 2801.750 527.650 2804.600 ;
        RECT 532.570 2802.450 532.870 2804.600 ;
        RECT 531.150 2802.150 532.870 2802.450 ;
        RECT 527.350 2801.450 530.530 2801.750 ;
        RECT 527.350 2800.000 527.650 2801.450 ;
        RECT 523.775 2794.295 524.105 2794.625 ;
        RECT 526.550 2787.825 526.850 2800.000 ;
        RECT 530.230 2787.825 530.530 2801.450 ;
        RECT 531.150 2793.265 531.450 2802.150 ;
        RECT 532.570 2800.000 532.870 2802.150 ;
        RECT 533.190 2801.750 533.490 2804.600 ;
        RECT 533.190 2801.450 536.050 2801.750 ;
        RECT 533.190 2800.000 533.490 2801.450 ;
        RECT 535.750 2794.625 536.050 2801.450 ;
        RECT 538.410 2796.650 538.710 2804.600 ;
        RECT 539.030 2801.750 539.330 2804.600 ;
        RECT 544.250 2801.750 544.550 2804.600 ;
        RECT 539.030 2801.450 542.490 2801.750 ;
        RECT 539.030 2800.000 539.330 2801.450 ;
        RECT 538.410 2796.350 538.810 2796.650 ;
        RECT 535.735 2794.295 536.065 2794.625 ;
        RECT 531.135 2792.935 531.465 2793.265 ;
        RECT 531.150 2788.505 531.450 2792.935 ;
        RECT 538.510 2789.865 538.810 2796.350 ;
        RECT 542.190 2794.625 542.490 2801.450 ;
        RECT 543.110 2801.450 544.550 2801.750 ;
        RECT 542.175 2794.295 542.505 2794.625 ;
        RECT 543.110 2792.585 543.410 2801.450 ;
        RECT 544.250 2800.000 544.550 2801.450 ;
        RECT 544.870 2801.750 545.170 2804.600 ;
        RECT 984.010 2801.750 984.310 2804.600 ;
        RECT 989.850 2801.750 990.150 2804.600 ;
        RECT 995.690 2801.750 995.990 2804.600 ;
        RECT 1001.530 2801.750 1001.830 2804.600 ;
        RECT 544.870 2800.000 545.250 2801.750 ;
        RECT 544.950 2792.585 545.250 2800.000 ;
        RECT 981.030 2801.450 984.310 2801.750 ;
        RECT 981.030 2794.625 981.330 2801.450 ;
        RECT 984.010 2800.000 984.310 2801.450 ;
        RECT 986.550 2801.450 990.150 2801.750 ;
        RECT 981.015 2794.295 981.345 2794.625 ;
        RECT 543.095 2792.255 543.425 2792.585 ;
        RECT 544.935 2792.255 545.265 2792.585 ;
        RECT 986.550 2791.905 986.850 2801.450 ;
        RECT 989.850 2800.000 990.150 2801.450 ;
        RECT 993.910 2801.450 995.990 2801.750 ;
        RECT 986.535 2791.575 986.865 2791.905 ;
        RECT 993.910 2791.225 994.210 2801.450 ;
        RECT 995.690 2800.000 995.990 2801.450 ;
        RECT 1001.270 2800.000 1001.830 2801.750 ;
        RECT 1007.370 2800.050 1007.670 2804.600 ;
        RECT 1013.210 2801.750 1013.510 2804.600 ;
        RECT 1012.310 2801.450 1013.510 2801.750 ;
        RECT 1001.270 2794.625 1001.570 2800.000 ;
        RECT 1007.370 2799.750 1008.010 2800.050 ;
        RECT 1001.255 2794.295 1001.585 2794.625 ;
        RECT 993.895 2790.895 994.225 2791.225 ;
        RECT 538.495 2789.535 538.825 2789.865 ;
        RECT 1007.710 2788.505 1008.010 2799.750 ;
        RECT 1012.310 2793.265 1012.610 2801.450 ;
        RECT 1013.210 2800.000 1013.510 2801.450 ;
        RECT 1013.830 2796.650 1014.130 2804.600 ;
        RECT 1019.050 2801.750 1019.350 2804.600 ;
        RECT 1013.230 2796.350 1014.130 2796.650 ;
        RECT 1018.750 2800.000 1019.350 2801.750 ;
        RECT 1013.230 2794.625 1013.530 2796.350 ;
        RECT 1018.750 2794.625 1019.050 2800.000 ;
        RECT 1019.670 2794.625 1019.970 2804.600 ;
        RECT 1024.890 2801.750 1025.190 2804.600 ;
        RECT 1024.270 2801.450 1025.190 2801.750 ;
        RECT 1013.215 2794.295 1013.545 2794.625 ;
        RECT 1018.735 2794.295 1019.065 2794.625 ;
        RECT 1019.655 2794.295 1019.985 2794.625 ;
        RECT 1024.270 2793.265 1024.570 2801.450 ;
        RECT 1024.890 2800.000 1025.190 2801.450 ;
        RECT 1025.510 2801.750 1025.810 2804.600 ;
        RECT 1030.730 2801.750 1031.030 2804.600 ;
        RECT 1025.510 2801.450 1027.330 2801.750 ;
        RECT 1025.510 2800.000 1025.810 2801.450 ;
        RECT 1027.030 2794.625 1027.330 2801.450 ;
        RECT 1030.710 2800.000 1031.030 2801.750 ;
        RECT 1031.350 2801.750 1031.650 2804.600 ;
        RECT 1036.570 2802.450 1036.870 2804.600 ;
        RECT 1035.310 2802.150 1036.870 2802.450 ;
        RECT 1031.350 2801.450 1034.690 2801.750 ;
        RECT 1031.350 2800.000 1031.650 2801.450 ;
        RECT 1030.710 2794.625 1031.010 2800.000 ;
        RECT 1027.015 2794.295 1027.345 2794.625 ;
        RECT 1030.695 2794.295 1031.025 2794.625 ;
        RECT 1012.295 2792.935 1012.625 2793.265 ;
        RECT 1024.255 2792.935 1024.585 2793.265 ;
        RECT 531.135 2788.175 531.465 2788.505 ;
        RECT 1007.695 2788.175 1008.025 2788.505 ;
        RECT 1034.390 2787.825 1034.690 2801.450 ;
        RECT 1035.310 2788.505 1035.610 2802.150 ;
        RECT 1036.570 2800.000 1036.870 2802.150 ;
        RECT 1037.190 2801.750 1037.490 2804.600 ;
        RECT 1042.410 2801.750 1042.710 2804.600 ;
        RECT 1037.190 2801.450 1040.210 2801.750 ;
        RECT 1037.190 2800.000 1037.490 2801.450 ;
        RECT 1035.295 2788.175 1035.625 2788.505 ;
        RECT 1039.910 2787.825 1040.210 2801.450 ;
        RECT 1041.750 2801.450 1042.710 2801.750 ;
        RECT 1041.750 2794.625 1042.050 2801.450 ;
        RECT 1042.410 2800.000 1042.710 2801.450 ;
        RECT 1043.030 2801.750 1043.330 2804.600 ;
        RECT 1048.250 2801.750 1048.550 2804.600 ;
        RECT 1043.030 2801.450 1046.650 2801.750 ;
        RECT 1043.030 2800.000 1043.330 2801.450 ;
        RECT 1041.735 2794.295 1042.065 2794.625 ;
        RECT 1046.350 2787.825 1046.650 2801.450 ;
        RECT 1048.190 2800.000 1048.550 2801.750 ;
        RECT 1048.870 2801.750 1049.170 2804.600 ;
        RECT 1054.090 2801.750 1054.390 2804.600 ;
        RECT 1048.870 2801.450 1052.170 2801.750 ;
        RECT 1048.870 2800.000 1049.170 2801.450 ;
        RECT 1048.190 2793.265 1048.490 2800.000 ;
        RECT 1048.175 2792.935 1048.505 2793.265 ;
        RECT 1051.870 2788.505 1052.170 2801.450 ;
        RECT 1052.790 2801.450 1054.390 2801.750 ;
        RECT 1052.790 2794.625 1053.090 2801.450 ;
        RECT 1054.090 2800.000 1054.390 2801.450 ;
        RECT 1054.710 2800.050 1055.010 2804.600 ;
        RECT 1059.930 2801.750 1060.230 2804.600 ;
        RECT 1059.230 2801.450 1060.230 2801.750 ;
        RECT 1055.535 2800.050 1055.865 2800.065 ;
        RECT 1054.710 2799.750 1055.865 2800.050 ;
        RECT 1055.535 2799.735 1055.865 2799.750 ;
        RECT 1059.230 2794.625 1059.530 2801.450 ;
        RECT 1059.930 2800.000 1060.230 2801.450 ;
        RECT 1060.550 2801.750 1060.850 2804.600 ;
        RECT 1065.770 2801.750 1066.070 2804.600 ;
        RECT 1060.550 2801.450 1062.290 2801.750 ;
        RECT 1060.550 2800.000 1060.850 2801.450 ;
        RECT 1052.775 2794.295 1053.105 2794.625 ;
        RECT 1059.215 2794.295 1059.545 2794.625 ;
        RECT 1051.855 2788.175 1052.185 2788.505 ;
        RECT 1061.990 2787.825 1062.290 2801.450 ;
        RECT 1065.670 2800.000 1066.070 2801.750 ;
        RECT 1066.390 2801.750 1066.690 2804.600 ;
        RECT 1071.610 2802.450 1071.910 2804.600 ;
        RECT 1070.270 2802.150 1071.910 2802.450 ;
        RECT 1066.390 2801.450 1067.810 2801.750 ;
        RECT 1066.390 2800.000 1066.690 2801.450 ;
        RECT 1065.670 2794.625 1065.970 2800.000 ;
        RECT 1065.655 2794.295 1065.985 2794.625 ;
        RECT 1067.510 2787.825 1067.810 2801.450 ;
        RECT 1070.270 2794.625 1070.570 2802.150 ;
        RECT 1071.610 2800.000 1071.910 2802.150 ;
        RECT 1072.230 2801.750 1072.530 2804.600 ;
        RECT 1077.450 2801.750 1077.750 2804.600 ;
        RECT 1072.230 2801.450 1074.250 2801.750 ;
        RECT 1072.230 2800.000 1072.530 2801.450 ;
        RECT 1070.255 2794.295 1070.585 2794.625 ;
        RECT 1073.950 2787.825 1074.250 2801.450 ;
        RECT 1076.710 2801.450 1077.750 2801.750 ;
        RECT 1076.710 2794.625 1077.010 2801.450 ;
        RECT 1077.450 2800.000 1077.750 2801.450 ;
        RECT 1078.070 2801.750 1078.370 2804.600 ;
        RECT 1083.290 2801.750 1083.590 2804.600 ;
        RECT 1078.070 2801.450 1081.610 2801.750 ;
        RECT 1078.070 2800.000 1078.370 2801.450 ;
        RECT 1076.695 2794.295 1077.025 2794.625 ;
        RECT 1081.310 2787.825 1081.610 2801.450 ;
        RECT 1083.150 2800.000 1083.590 2801.750 ;
        RECT 1083.910 2801.750 1084.210 2804.600 ;
        RECT 1089.130 2802.450 1089.430 2804.600 ;
        RECT 1087.750 2802.150 1089.430 2802.450 ;
        RECT 1083.910 2801.450 1087.130 2801.750 ;
        RECT 1083.910 2800.000 1084.210 2801.450 ;
        RECT 1083.150 2794.625 1083.450 2800.000 ;
        RECT 1083.135 2794.295 1083.465 2794.625 ;
        RECT 1086.830 2788.505 1087.130 2801.450 ;
        RECT 1087.750 2793.945 1088.050 2802.150 ;
        RECT 1089.130 2800.000 1089.430 2802.150 ;
        RECT 1089.750 2796.650 1090.050 2804.600 ;
        RECT 1094.970 2801.750 1095.270 2804.600 ;
        RECT 1089.590 2796.350 1090.050 2796.650 ;
        RECT 1094.190 2801.450 1095.270 2801.750 ;
        RECT 1087.735 2793.615 1088.065 2793.945 ;
        RECT 1086.815 2788.175 1087.145 2788.505 ;
        RECT 1089.590 2787.825 1089.890 2796.350 ;
        RECT 1094.190 2794.625 1094.490 2801.450 ;
        RECT 1094.970 2800.000 1095.270 2801.450 ;
        RECT 1095.590 2800.050 1095.890 2804.600 ;
        RECT 1100.810 2801.750 1101.110 2804.600 ;
        RECT 1095.590 2799.750 1096.330 2800.050 ;
        RECT 1094.175 2794.295 1094.505 2794.625 ;
        RECT 1096.030 2787.825 1096.330 2799.750 ;
        RECT 1100.630 2800.000 1101.110 2801.750 ;
        RECT 1101.430 2801.750 1101.730 2804.600 ;
        RECT 1106.650 2802.450 1106.950 2804.600 ;
        RECT 1105.230 2802.150 1106.950 2802.450 ;
        RECT 1101.430 2801.450 1103.690 2801.750 ;
        RECT 1101.430 2800.000 1101.730 2801.450 ;
        RECT 1100.630 2794.625 1100.930 2800.000 ;
        RECT 1100.615 2794.295 1100.945 2794.625 ;
        RECT 1103.390 2787.825 1103.690 2801.450 ;
        RECT 1105.230 2794.625 1105.530 2802.150 ;
        RECT 1106.650 2800.000 1106.950 2802.150 ;
        RECT 1107.270 2801.750 1107.570 2804.600 ;
        RECT 1112.490 2801.750 1112.790 2804.600 ;
        RECT 1107.270 2801.450 1110.130 2801.750 ;
        RECT 1107.270 2800.000 1107.570 2801.450 ;
        RECT 1105.215 2794.295 1105.545 2794.625 ;
        RECT 1109.830 2787.825 1110.130 2801.450 ;
        RECT 1111.670 2801.450 1112.790 2801.750 ;
        RECT 1111.670 2794.625 1111.970 2801.450 ;
        RECT 1112.490 2800.000 1112.790 2801.450 ;
        RECT 1113.110 2801.750 1113.410 2804.600 ;
        RECT 1118.330 2801.750 1118.630 2804.600 ;
        RECT 1113.110 2801.450 1116.570 2801.750 ;
        RECT 1113.110 2800.000 1113.410 2801.450 ;
        RECT 1111.655 2794.295 1111.985 2794.625 ;
        RECT 1116.270 2787.825 1116.570 2801.450 ;
        RECT 1118.110 2800.000 1118.630 2801.750 ;
        RECT 1118.950 2801.750 1119.250 2804.600 ;
        RECT 1124.170 2801.750 1124.470 2804.600 ;
        RECT 1118.950 2801.450 1122.090 2801.750 ;
        RECT 1118.950 2800.000 1119.250 2801.450 ;
        RECT 1118.110 2793.945 1118.410 2800.000 ;
        RECT 1118.095 2793.615 1118.425 2793.945 ;
        RECT 1121.790 2787.825 1122.090 2801.450 ;
        RECT 1122.710 2801.450 1124.470 2801.750 ;
        RECT 1122.710 2794.625 1123.010 2801.450 ;
        RECT 1124.170 2800.000 1124.470 2801.450 ;
        RECT 1124.790 2801.750 1125.090 2804.600 ;
        RECT 1130.010 2801.750 1130.310 2804.600 ;
        RECT 1124.790 2801.450 1128.530 2801.750 ;
        RECT 1124.790 2800.000 1125.090 2801.450 ;
        RECT 1122.695 2794.295 1123.025 2794.625 ;
        RECT 1128.230 2793.945 1128.530 2801.450 ;
        RECT 1129.150 2801.450 1130.310 2801.750 ;
        RECT 1129.150 2794.625 1129.450 2801.450 ;
        RECT 1130.010 2800.000 1130.310 2801.450 ;
        RECT 1130.630 2800.050 1130.930 2804.600 ;
        RECT 1135.850 2801.750 1136.150 2804.600 ;
        RECT 1130.630 2799.750 1131.290 2800.050 ;
        RECT 1130.990 2794.625 1131.290 2799.750 ;
        RECT 1135.590 2800.000 1136.150 2801.750 ;
        RECT 1136.470 2801.750 1136.770 2804.600 ;
        RECT 1141.690 2802.450 1141.990 2804.600 ;
        RECT 1140.190 2802.150 1141.990 2802.450 ;
        RECT 1136.470 2801.450 1137.730 2801.750 ;
        RECT 1136.470 2800.000 1136.770 2801.450 ;
        RECT 1135.590 2794.625 1135.890 2800.000 ;
        RECT 1137.430 2794.625 1137.730 2801.450 ;
        RECT 1140.190 2794.625 1140.490 2802.150 ;
        RECT 1141.690 2800.000 1141.990 2802.150 ;
        RECT 1142.310 2801.750 1142.610 2804.600 ;
        RECT 1142.310 2801.450 1144.170 2801.750 ;
        RECT 1142.310 2800.000 1142.610 2801.450 ;
        RECT 1143.870 2794.625 1144.170 2801.450 ;
        RECT 1147.530 2800.050 1147.830 2804.600 ;
        RECT 1148.150 2801.750 1148.450 2804.600 ;
        RECT 1153.370 2801.750 1153.670 2804.600 ;
        RECT 1148.150 2801.450 1151.530 2801.750 ;
        RECT 1147.530 2799.750 1147.850 2800.050 ;
        RECT 1148.150 2800.000 1148.450 2801.450 ;
        RECT 1147.550 2794.625 1147.850 2799.750 ;
        RECT 1151.230 2794.625 1151.530 2801.450 ;
        RECT 1153.070 2800.000 1153.670 2801.750 ;
        RECT 1129.135 2794.295 1129.465 2794.625 ;
        RECT 1130.975 2794.295 1131.305 2794.625 ;
        RECT 1135.575 2794.295 1135.905 2794.625 ;
        RECT 1137.415 2794.295 1137.745 2794.625 ;
        RECT 1140.175 2794.295 1140.505 2794.625 ;
        RECT 1143.855 2794.295 1144.185 2794.625 ;
        RECT 1147.535 2794.295 1147.865 2794.625 ;
        RECT 1151.215 2794.295 1151.545 2794.625 ;
        RECT 1128.215 2793.615 1128.545 2793.945 ;
        RECT 1153.070 2791.905 1153.370 2800.000 ;
        RECT 1153.990 2794.625 1154.290 2804.600 ;
        RECT 1159.210 2796.650 1159.510 2804.600 ;
        RECT 1159.830 2801.750 1160.130 2804.600 ;
        RECT 1165.050 2801.750 1165.350 2804.600 ;
        RECT 1159.830 2801.450 1163.490 2801.750 ;
        RECT 1159.830 2800.000 1160.130 2801.450 ;
        RECT 1159.210 2796.350 1159.810 2796.650 ;
        RECT 1153.975 2794.295 1154.305 2794.625 ;
        RECT 1159.510 2793.945 1159.810 2796.350 ;
        RECT 1163.190 2793.945 1163.490 2801.450 ;
        RECT 1164.110 2801.450 1165.350 2801.750 ;
        RECT 1159.495 2793.615 1159.825 2793.945 ;
        RECT 1163.175 2793.615 1163.505 2793.945 ;
        RECT 1164.110 2792.585 1164.410 2801.450 ;
        RECT 1165.050 2800.000 1165.350 2801.450 ;
        RECT 1165.670 2796.650 1165.970 2804.600 ;
        RECT 1170.890 2801.750 1171.190 2804.600 ;
        RECT 1165.030 2796.350 1165.970 2796.650 ;
        RECT 1167.790 2801.450 1171.190 2801.750 ;
        RECT 1165.030 2794.625 1165.330 2796.350 ;
        RECT 1167.790 2794.625 1168.090 2801.450 ;
        RECT 1170.890 2800.000 1171.190 2801.450 ;
        RECT 1171.510 2801.750 1171.810 2804.600 ;
        RECT 1176.730 2801.750 1177.030 2804.600 ;
        RECT 1171.510 2801.450 1172.690 2801.750 ;
        RECT 1171.510 2800.000 1171.810 2801.450 ;
        RECT 1172.390 2794.625 1172.690 2801.450 ;
        RECT 1173.310 2801.450 1177.030 2801.750 ;
        RECT 1165.015 2794.295 1165.345 2794.625 ;
        RECT 1167.775 2794.295 1168.105 2794.625 ;
        RECT 1172.375 2794.295 1172.705 2794.625 ;
        RECT 1173.310 2793.945 1173.610 2801.450 ;
        RECT 1176.730 2800.000 1177.030 2801.450 ;
        RECT 1177.350 2801.750 1177.650 2804.600 ;
        RECT 1182.570 2801.750 1182.870 2804.600 ;
        RECT 1177.350 2801.450 1179.130 2801.750 ;
        RECT 1177.350 2800.000 1177.650 2801.450 ;
        RECT 1178.830 2794.625 1179.130 2801.450 ;
        RECT 1180.670 2801.450 1182.870 2801.750 ;
        RECT 1178.815 2794.295 1179.145 2794.625 ;
        RECT 1180.670 2793.945 1180.970 2801.450 ;
        RECT 1182.570 2800.000 1182.870 2801.450 ;
        RECT 1183.190 2801.750 1183.490 2804.600 ;
        RECT 1188.410 2801.750 1188.710 2804.600 ;
        RECT 1183.190 2801.450 1186.490 2801.750 ;
        RECT 1183.190 2800.000 1183.490 2801.450 ;
        RECT 1186.190 2794.625 1186.490 2801.450 ;
        RECT 1187.110 2801.450 1188.710 2801.750 ;
        RECT 1186.175 2794.295 1186.505 2794.625 ;
        RECT 1187.110 2793.945 1187.410 2801.450 ;
        RECT 1188.410 2800.000 1188.710 2801.450 ;
        RECT 1189.030 2801.750 1189.330 2804.600 ;
        RECT 1194.250 2801.750 1194.550 2804.600 ;
        RECT 1189.030 2801.450 1192.010 2801.750 ;
        RECT 1189.030 2800.000 1189.330 2801.450 ;
        RECT 1173.295 2793.615 1173.625 2793.945 ;
        RECT 1180.655 2793.615 1180.985 2793.945 ;
        RECT 1187.095 2793.615 1187.425 2793.945 ;
        RECT 1164.095 2792.255 1164.425 2792.585 ;
        RECT 1153.055 2791.575 1153.385 2791.905 ;
        RECT 1191.710 2790.545 1192.010 2801.450 ;
        RECT 1193.550 2801.450 1194.550 2801.750 ;
        RECT 1193.550 2791.905 1193.850 2801.450 ;
        RECT 1194.250 2800.000 1194.550 2801.450 ;
        RECT 1194.870 2801.750 1195.170 2804.600 ;
        RECT 1584.010 2801.750 1584.310 2804.600 ;
        RECT 1589.850 2801.750 1590.150 2804.600 ;
        RECT 1595.690 2801.750 1595.990 2804.600 ;
        RECT 1194.870 2801.450 1198.450 2801.750 ;
        RECT 1194.870 2800.000 1195.170 2801.450 ;
        RECT 1198.150 2794.625 1198.450 2801.450 ;
        RECT 1581.790 2801.450 1584.310 2801.750 ;
        RECT 1198.135 2794.295 1198.465 2794.625 ;
        RECT 1193.535 2791.575 1193.865 2791.905 ;
        RECT 1411.575 2791.575 1411.905 2791.905 ;
        RECT 1191.695 2790.215 1192.025 2790.545 ;
        RECT 507.215 2787.495 507.545 2787.825 ;
        RECT 513.655 2787.495 513.985 2787.825 ;
        RECT 516.415 2787.495 516.745 2787.825 ;
        RECT 520.095 2787.495 520.425 2787.825 ;
        RECT 526.535 2787.495 526.865 2787.825 ;
        RECT 530.215 2787.495 530.545 2787.825 ;
        RECT 1034.375 2787.495 1034.705 2787.825 ;
        RECT 1039.895 2787.495 1040.225 2787.825 ;
        RECT 1046.335 2787.495 1046.665 2787.825 ;
        RECT 1061.975 2787.495 1062.305 2787.825 ;
        RECT 1067.495 2787.495 1067.825 2787.825 ;
        RECT 1073.935 2787.495 1074.265 2787.825 ;
        RECT 1081.295 2787.495 1081.625 2787.825 ;
        RECT 1089.575 2787.495 1089.905 2787.825 ;
        RECT 1096.015 2787.495 1096.345 2787.825 ;
        RECT 1103.375 2787.495 1103.705 2787.825 ;
        RECT 1109.815 2787.495 1110.145 2787.825 ;
        RECT 1116.255 2787.495 1116.585 2787.825 ;
        RECT 1121.775 2787.495 1122.105 2787.825 ;
        RECT 292.020 2715.000 295.020 2785.000 ;
        RECT 310.020 2715.000 313.020 2785.000 ;
        RECT 328.020 2715.000 331.020 2785.000 ;
        RECT 364.020 2715.000 367.020 2785.000 ;
        RECT 454.020 2715.000 457.020 2785.000 ;
        RECT 472.020 2715.000 475.020 2785.000 ;
        RECT 490.020 2715.000 493.020 2785.000 ;
        RECT 508.020 2715.000 511.020 2785.000 ;
        RECT 544.020 2715.000 547.020 2785.000 ;
        RECT 634.020 2715.000 637.020 2785.000 ;
        RECT 652.020 2715.000 655.020 2785.000 ;
        RECT 670.020 2715.000 673.020 2785.000 ;
        RECT 688.020 2715.000 691.020 2785.000 ;
        RECT 994.020 2715.000 997.020 2785.000 ;
        RECT 1012.020 2715.000 1015.020 2785.000 ;
        RECT 1030.020 2715.000 1033.020 2785.000 ;
        RECT 1048.020 2715.000 1051.020 2785.000 ;
        RECT 1084.020 2715.000 1087.020 2785.000 ;
        RECT 1174.020 2715.000 1177.020 2785.000 ;
        RECT 1192.020 2715.000 1195.020 2785.000 ;
        RECT 1210.020 2715.000 1213.020 2785.000 ;
        RECT 1228.020 2715.000 1231.020 2785.000 ;
        RECT 1264.020 2715.000 1267.020 2785.000 ;
      LAYER met4 ;
        RECT 323.295 2688.640 1389.905 2697.345 ;
        RECT 323.295 1610.240 397.440 2688.640 ;
        RECT 399.840 1610.240 1389.905 2688.640 ;
      LAYER met4 ;
        RECT 1411.590 1617.545 1411.890 2791.575 ;
        RECT 1417.095 2790.895 1417.425 2791.225 ;
        RECT 1417.110 1622.305 1417.410 2790.895 ;
        RECT 1581.790 2789.185 1582.090 2801.450 ;
        RECT 1584.010 2800.000 1584.310 2801.450 ;
        RECT 1587.310 2801.450 1590.150 2801.750 ;
        RECT 1587.310 2794.625 1587.610 2801.450 ;
        RECT 1589.850 2800.000 1590.150 2801.450 ;
        RECT 1594.670 2801.450 1595.990 2801.750 ;
        RECT 1594.670 2794.625 1594.970 2801.450 ;
        RECT 1595.690 2800.000 1595.990 2801.450 ;
        RECT 1601.530 2800.050 1601.830 2804.600 ;
        RECT 1607.370 2801.750 1607.670 2804.600 ;
        RECT 1613.210 2801.750 1613.510 2804.600 ;
        RECT 1601.110 2799.750 1601.830 2800.050 ;
        RECT 1604.790 2801.450 1607.670 2801.750 ;
        RECT 1601.110 2794.625 1601.410 2799.750 ;
        RECT 1587.295 2794.295 1587.625 2794.625 ;
        RECT 1594.655 2794.295 1594.985 2794.625 ;
        RECT 1601.095 2794.295 1601.425 2794.625 ;
        RECT 1604.790 2793.945 1605.090 2801.450 ;
        RECT 1607.370 2800.000 1607.670 2801.450 ;
        RECT 1613.070 2800.000 1613.510 2801.750 ;
        RECT 1613.830 2801.750 1614.130 2804.600 ;
        RECT 1619.050 2802.450 1619.350 2804.600 ;
        RECT 1617.670 2802.150 1619.350 2802.450 ;
        RECT 1613.830 2800.000 1614.290 2801.750 ;
        RECT 1613.070 2793.945 1613.370 2800.000 ;
        RECT 1604.775 2793.615 1605.105 2793.945 ;
        RECT 1613.055 2793.615 1613.385 2793.945 ;
        RECT 1613.990 2790.545 1614.290 2800.000 ;
        RECT 1617.670 2793.265 1617.970 2802.150 ;
        RECT 1619.050 2800.000 1619.350 2802.150 ;
        RECT 1619.670 2801.750 1619.970 2804.600 ;
        RECT 1624.890 2801.750 1625.190 2804.600 ;
        RECT 1619.670 2801.450 1620.730 2801.750 ;
        RECT 1619.670 2800.000 1619.970 2801.450 ;
        RECT 1617.655 2792.935 1617.985 2793.265 ;
        RECT 1620.430 2790.545 1620.730 2801.450 ;
        RECT 1624.110 2801.450 1625.190 2801.750 ;
        RECT 1624.110 2793.265 1624.410 2801.450 ;
        RECT 1624.890 2800.000 1625.190 2801.450 ;
        RECT 1625.510 2802.450 1625.810 2804.600 ;
        RECT 1625.510 2802.150 1627.170 2802.450 ;
        RECT 1625.510 2800.000 1625.810 2802.150 ;
        RECT 1624.095 2792.935 1624.425 2793.265 ;
        RECT 1613.975 2790.215 1614.305 2790.545 ;
        RECT 1620.415 2790.215 1620.745 2790.545 ;
        RECT 1581.775 2788.855 1582.105 2789.185 ;
        RECT 1626.870 2788.505 1627.170 2802.150 ;
        RECT 1630.730 2801.750 1631.030 2804.600 ;
        RECT 1630.550 2800.000 1631.030 2801.750 ;
        RECT 1631.350 2801.750 1631.650 2804.600 ;
        RECT 1636.570 2802.450 1636.870 2804.600 ;
        RECT 1635.150 2802.150 1636.870 2802.450 ;
        RECT 1631.350 2800.000 1631.770 2801.750 ;
        RECT 1630.550 2793.945 1630.850 2800.000 ;
        RECT 1631.470 2794.625 1631.770 2800.000 ;
        RECT 1631.455 2794.295 1631.785 2794.625 ;
        RECT 1630.535 2793.615 1630.865 2793.945 ;
        RECT 1635.150 2793.265 1635.450 2802.150 ;
        RECT 1636.570 2800.000 1636.870 2802.150 ;
        RECT 1637.190 2801.750 1637.490 2804.600 ;
        RECT 1637.190 2801.450 1638.210 2801.750 ;
        RECT 1637.190 2800.000 1637.490 2801.450 ;
        RECT 1637.910 2794.625 1638.210 2801.450 ;
        RECT 1642.410 2796.650 1642.710 2804.600 ;
        RECT 1643.030 2802.450 1643.330 2804.600 ;
        RECT 1643.030 2802.150 1644.650 2802.450 ;
        RECT 1643.030 2800.000 1643.330 2802.150 ;
        RECT 1642.410 2796.350 1642.810 2796.650 ;
        RECT 1637.895 2794.295 1638.225 2794.625 ;
        RECT 1642.510 2793.265 1642.810 2796.350 ;
        RECT 1644.350 2793.945 1644.650 2802.150 ;
        RECT 1648.250 2801.750 1648.550 2804.600 ;
        RECT 1648.030 2800.000 1648.550 2801.750 ;
        RECT 1648.870 2801.750 1649.170 2804.600 ;
        RECT 1654.090 2802.450 1654.390 2804.600 ;
        RECT 1652.630 2802.150 1654.390 2802.450 ;
        RECT 1648.870 2800.000 1649.250 2801.750 ;
        RECT 1648.030 2794.625 1648.330 2800.000 ;
        RECT 1648.015 2794.295 1648.345 2794.625 ;
        RECT 1644.335 2793.615 1644.665 2793.945 ;
        RECT 1635.135 2792.935 1635.465 2793.265 ;
        RECT 1642.495 2792.935 1642.825 2793.265 ;
        RECT 1648.950 2789.865 1649.250 2800.000 ;
        RECT 1652.630 2793.945 1652.930 2802.150 ;
        RECT 1654.090 2800.000 1654.390 2802.150 ;
        RECT 1654.710 2801.750 1655.010 2804.600 ;
        RECT 1659.930 2801.750 1660.230 2804.600 ;
        RECT 1654.710 2801.450 1655.690 2801.750 ;
        RECT 1654.710 2800.000 1655.010 2801.450 ;
        RECT 1655.390 2794.625 1655.690 2801.450 ;
        RECT 1659.070 2801.450 1660.230 2801.750 ;
        RECT 1659.070 2794.625 1659.370 2801.450 ;
        RECT 1659.930 2800.000 1660.230 2801.450 ;
        RECT 1660.550 2802.450 1660.850 2804.600 ;
        RECT 1660.550 2802.150 1662.130 2802.450 ;
        RECT 1660.550 2800.000 1660.850 2802.150 ;
        RECT 1655.375 2794.295 1655.705 2794.625 ;
        RECT 1659.055 2794.295 1659.385 2794.625 ;
        RECT 1652.615 2793.615 1652.945 2793.945 ;
        RECT 1648.935 2789.535 1649.265 2789.865 ;
        RECT 1661.830 2789.185 1662.130 2802.150 ;
        RECT 1665.770 2801.750 1666.070 2804.600 ;
        RECT 1665.510 2800.000 1666.070 2801.750 ;
        RECT 1666.390 2801.750 1666.690 2804.600 ;
        RECT 1671.610 2802.450 1671.910 2804.600 ;
        RECT 1670.110 2802.150 1671.910 2802.450 ;
        RECT 1666.390 2800.000 1666.730 2801.750 ;
        RECT 1665.510 2793.945 1665.810 2800.000 ;
        RECT 1666.430 2794.625 1666.730 2800.000 ;
        RECT 1666.415 2794.295 1666.745 2794.625 ;
        RECT 1670.110 2793.945 1670.410 2802.150 ;
        RECT 1671.610 2800.000 1671.910 2802.150 ;
        RECT 1672.230 2801.750 1672.530 2804.600 ;
        RECT 1672.230 2801.450 1673.170 2801.750 ;
        RECT 1672.230 2800.000 1672.530 2801.450 ;
        RECT 1672.870 2794.625 1673.170 2801.450 ;
        RECT 1677.450 2800.050 1677.750 2804.600 ;
        RECT 1678.070 2802.450 1678.370 2804.600 ;
        RECT 1678.070 2802.150 1679.610 2802.450 ;
        RECT 1677.450 2799.750 1677.770 2800.050 ;
        RECT 1678.070 2800.000 1678.370 2802.150 ;
        RECT 1672.855 2794.295 1673.185 2794.625 ;
        RECT 1677.470 2793.945 1677.770 2799.750 ;
        RECT 1679.310 2794.625 1679.610 2802.150 ;
        RECT 1683.290 2801.750 1683.590 2804.600 ;
        RECT 1682.990 2800.000 1683.590 2801.750 ;
        RECT 1679.295 2794.295 1679.625 2794.625 ;
        RECT 1682.990 2793.945 1683.290 2800.000 ;
        RECT 1683.910 2794.625 1684.210 2804.600 ;
        RECT 1689.130 2801.750 1689.430 2804.600 ;
        RECT 1688.510 2801.450 1689.430 2801.750 ;
        RECT 1688.510 2794.625 1688.810 2801.450 ;
        RECT 1689.130 2800.000 1689.430 2801.450 ;
        RECT 1689.750 2796.650 1690.050 2804.600 ;
        RECT 1694.970 2801.750 1695.270 2804.600 ;
        RECT 1689.430 2796.350 1690.050 2796.650 ;
        RECT 1694.950 2800.000 1695.270 2801.750 ;
        RECT 1695.590 2801.750 1695.890 2804.600 ;
        RECT 1700.810 2802.450 1701.110 2804.600 ;
        RECT 1699.550 2802.150 1701.110 2802.450 ;
        RECT 1695.590 2800.000 1696.170 2801.750 ;
        RECT 1683.895 2794.295 1684.225 2794.625 ;
        RECT 1688.495 2794.295 1688.825 2794.625 ;
        RECT 1689.430 2793.945 1689.730 2796.350 ;
        RECT 1694.950 2793.945 1695.250 2800.000 ;
        RECT 1695.870 2794.625 1696.170 2800.000 ;
        RECT 1695.855 2794.295 1696.185 2794.625 ;
        RECT 1699.550 2793.945 1699.850 2802.150 ;
        RECT 1700.810 2800.000 1701.110 2802.150 ;
        RECT 1701.430 2801.750 1701.730 2804.600 ;
        RECT 1706.650 2801.750 1706.950 2804.600 ;
        RECT 1701.430 2801.450 1702.610 2801.750 ;
        RECT 1701.430 2800.000 1701.730 2801.450 ;
        RECT 1702.310 2794.625 1702.610 2801.450 ;
        RECT 1705.990 2801.450 1706.950 2801.750 ;
        RECT 1702.295 2794.295 1702.625 2794.625 ;
        RECT 1705.990 2793.945 1706.290 2801.450 ;
        RECT 1706.650 2800.000 1706.950 2801.450 ;
        RECT 1707.270 2802.450 1707.570 2804.600 ;
        RECT 1707.270 2802.150 1709.050 2802.450 ;
        RECT 1707.270 2800.000 1707.570 2802.150 ;
        RECT 1708.750 2794.625 1709.050 2802.150 ;
        RECT 1712.490 2801.750 1712.790 2804.600 ;
        RECT 1712.430 2800.000 1712.790 2801.750 ;
        RECT 1713.110 2801.750 1713.410 2804.600 ;
        RECT 1713.110 2800.000 1713.650 2801.750 ;
        RECT 1718.330 2800.050 1718.630 2804.600 ;
        RECT 1708.735 2794.295 1709.065 2794.625 ;
        RECT 1712.430 2793.945 1712.730 2800.000 ;
        RECT 1713.350 2794.625 1713.650 2800.000 ;
        RECT 1717.950 2799.750 1718.630 2800.050 ;
        RECT 1718.950 2801.750 1719.250 2804.600 ;
        RECT 1724.170 2801.750 1724.470 2804.600 ;
        RECT 1718.950 2801.450 1720.090 2801.750 ;
        RECT 1718.950 2800.000 1719.250 2801.450 ;
        RECT 1713.335 2794.295 1713.665 2794.625 ;
        RECT 1717.950 2793.945 1718.250 2799.750 ;
        RECT 1719.790 2794.625 1720.090 2801.450 ;
        RECT 1721.630 2801.450 1724.470 2801.750 ;
        RECT 1721.630 2794.625 1721.930 2801.450 ;
        RECT 1724.170 2800.000 1724.470 2801.450 ;
        RECT 1724.790 2796.650 1725.090 2804.600 ;
        RECT 1730.010 2801.750 1730.310 2804.600 ;
        RECT 1724.390 2796.350 1725.090 2796.650 ;
        RECT 1729.910 2800.000 1730.310 2801.750 ;
        RECT 1730.630 2801.750 1730.930 2804.600 ;
        RECT 1735.850 2801.750 1736.150 2804.600 ;
        RECT 1730.630 2800.000 1731.130 2801.750 ;
        RECT 1719.775 2794.295 1720.105 2794.625 ;
        RECT 1721.615 2794.295 1721.945 2794.625 ;
        RECT 1665.495 2793.615 1665.825 2793.945 ;
        RECT 1670.095 2793.615 1670.425 2793.945 ;
        RECT 1677.455 2793.615 1677.785 2793.945 ;
        RECT 1682.975 2793.615 1683.305 2793.945 ;
        RECT 1689.415 2793.615 1689.745 2793.945 ;
        RECT 1694.935 2793.615 1695.265 2793.945 ;
        RECT 1699.535 2793.615 1699.865 2793.945 ;
        RECT 1705.975 2793.615 1706.305 2793.945 ;
        RECT 1712.415 2793.615 1712.745 2793.945 ;
        RECT 1717.935 2793.615 1718.265 2793.945 ;
        RECT 1661.815 2788.855 1662.145 2789.185 ;
        RECT 1724.390 2788.505 1724.690 2796.350 ;
        RECT 1729.910 2793.945 1730.210 2800.000 ;
        RECT 1730.830 2794.625 1731.130 2800.000 ;
        RECT 1734.510 2801.450 1736.150 2801.750 ;
        RECT 1730.815 2794.295 1731.145 2794.625 ;
        RECT 1734.510 2793.945 1734.810 2801.450 ;
        RECT 1735.850 2800.000 1736.150 2801.450 ;
        RECT 1736.470 2801.750 1736.770 2804.600 ;
        RECT 1741.690 2801.750 1741.990 2804.600 ;
        RECT 1736.470 2801.450 1737.570 2801.750 ;
        RECT 1736.470 2800.000 1736.770 2801.450 ;
        RECT 1737.270 2794.625 1737.570 2801.450 ;
        RECT 1740.950 2801.450 1741.990 2801.750 ;
        RECT 1737.255 2794.295 1737.585 2794.625 ;
        RECT 1740.950 2793.945 1741.250 2801.450 ;
        RECT 1741.690 2800.000 1741.990 2801.450 ;
        RECT 1742.310 2802.450 1742.610 2804.600 ;
        RECT 1742.310 2802.150 1744.010 2802.450 ;
        RECT 1742.310 2800.000 1742.610 2802.150 ;
        RECT 1743.710 2794.625 1744.010 2802.150 ;
        RECT 1747.530 2801.750 1747.830 2804.600 ;
        RECT 1747.390 2800.000 1747.830 2801.750 ;
        RECT 1748.150 2801.750 1748.450 2804.600 ;
        RECT 1748.150 2800.000 1748.610 2801.750 ;
        RECT 1753.370 2800.050 1753.670 2804.600 ;
        RECT 1743.695 2794.295 1744.025 2794.625 ;
        RECT 1747.390 2793.945 1747.690 2800.000 ;
        RECT 1748.310 2794.625 1748.610 2800.000 ;
        RECT 1752.910 2799.750 1753.670 2800.050 ;
        RECT 1753.990 2801.750 1754.290 2804.600 ;
        RECT 1753.990 2801.450 1755.050 2801.750 ;
        RECT 1753.990 2800.000 1754.290 2801.450 ;
        RECT 1748.295 2794.295 1748.625 2794.625 ;
        RECT 1729.895 2793.615 1730.225 2793.945 ;
        RECT 1734.495 2793.615 1734.825 2793.945 ;
        RECT 1740.935 2793.615 1741.265 2793.945 ;
        RECT 1747.375 2793.615 1747.705 2793.945 ;
        RECT 1752.910 2792.585 1753.210 2799.750 ;
        RECT 1752.895 2792.255 1753.225 2792.585 ;
        RECT 1626.855 2788.175 1627.185 2788.505 ;
        RECT 1724.375 2788.175 1724.705 2788.505 ;
        RECT 1754.750 2787.825 1755.050 2801.450 ;
        RECT 1759.210 2796.665 1759.510 2804.600 ;
        RECT 1759.830 2802.450 1760.130 2804.600 ;
        RECT 1759.830 2802.150 1761.490 2802.450 ;
        RECT 1759.830 2800.000 1760.130 2802.150 ;
        RECT 1759.210 2796.350 1759.665 2796.665 ;
        RECT 1759.335 2796.335 1759.665 2796.350 ;
        RECT 1754.735 2787.495 1755.065 2787.825 ;
        RECT 1761.190 2777.625 1761.490 2802.150 ;
        RECT 1765.050 2801.750 1765.350 2804.600 ;
        RECT 1762.110 2801.450 1765.350 2801.750 ;
        RECT 1762.110 2794.625 1762.410 2801.450 ;
        RECT 1765.050 2800.000 1765.350 2801.450 ;
        RECT 1765.670 2801.750 1765.970 2804.600 ;
        RECT 1770.890 2801.750 1771.190 2804.600 ;
        RECT 1765.670 2800.000 1766.090 2801.750 ;
        RECT 1762.095 2794.295 1762.425 2794.625 ;
        RECT 1765.790 2788.505 1766.090 2800.000 ;
        RECT 1767.630 2801.450 1771.190 2801.750 ;
        RECT 1767.630 2793.945 1767.930 2801.450 ;
        RECT 1770.890 2800.000 1771.190 2801.450 ;
        RECT 1771.510 2801.750 1771.810 2804.600 ;
        RECT 1776.730 2801.750 1777.030 2804.600 ;
        RECT 1771.510 2801.450 1772.530 2801.750 ;
        RECT 1771.510 2800.000 1771.810 2801.450 ;
        RECT 1767.615 2793.615 1767.945 2793.945 ;
        RECT 1765.775 2788.175 1766.105 2788.505 ;
        RECT 1772.230 2787.825 1772.530 2801.450 ;
        RECT 1774.070 2801.450 1777.030 2801.750 ;
        RECT 1774.070 2793.945 1774.370 2801.450 ;
        RECT 1776.730 2800.000 1777.030 2801.450 ;
        RECT 1777.350 2802.450 1777.650 2804.600 ;
        RECT 1777.350 2802.150 1778.970 2802.450 ;
        RECT 1777.350 2800.000 1777.650 2802.150 ;
        RECT 1774.055 2793.615 1774.385 2793.945 ;
        RECT 1778.670 2787.825 1778.970 2802.150 ;
        RECT 1782.570 2801.750 1782.870 2804.600 ;
        RECT 1780.510 2801.450 1782.870 2801.750 ;
        RECT 1780.510 2794.625 1780.810 2801.450 ;
        RECT 1782.570 2800.000 1782.870 2801.450 ;
        RECT 1783.190 2801.750 1783.490 2804.600 ;
        RECT 1783.190 2800.000 1783.570 2801.750 ;
        RECT 1788.410 2800.050 1788.710 2804.600 ;
        RECT 1780.495 2794.295 1780.825 2794.625 ;
        RECT 1783.270 2787.825 1783.570 2800.000 ;
        RECT 1787.870 2799.750 1788.710 2800.050 ;
        RECT 1789.030 2801.750 1789.330 2804.600 ;
        RECT 1789.030 2801.450 1790.010 2801.750 ;
        RECT 1789.030 2800.000 1789.330 2801.450 ;
        RECT 1787.870 2792.585 1788.170 2799.750 ;
        RECT 1787.855 2792.255 1788.185 2792.585 ;
        RECT 1789.710 2787.825 1790.010 2801.450 ;
        RECT 1794.250 2796.665 1794.550 2804.600 ;
        RECT 1794.870 2802.450 1795.170 2804.600 ;
        RECT 1794.870 2802.150 1796.450 2802.450 ;
        RECT 1794.870 2800.000 1795.170 2802.150 ;
        RECT 1794.250 2796.350 1794.625 2796.665 ;
        RECT 1794.295 2796.335 1794.625 2796.350 ;
        RECT 1772.215 2787.495 1772.545 2787.825 ;
        RECT 1778.655 2787.495 1778.985 2787.825 ;
        RECT 1783.255 2787.495 1783.585 2787.825 ;
        RECT 1789.695 2787.495 1790.025 2787.825 ;
        RECT 1796.150 2777.625 1796.450 2802.150 ;
        RECT 2234.010 2801.750 2234.310 2804.600 ;
        RECT 2239.850 2801.750 2240.150 2804.600 ;
        RECT 2245.690 2801.750 2245.990 2804.600 ;
        RECT 2251.530 2801.750 2251.830 2804.600 ;
        RECT 2257.370 2801.750 2257.670 2804.600 ;
        RECT 2231.310 2801.450 2234.310 2801.750 ;
        RECT 2231.310 2794.625 2231.610 2801.450 ;
        RECT 2234.010 2800.000 2234.310 2801.450 ;
        RECT 2236.830 2801.450 2240.150 2801.750 ;
        RECT 2231.295 2794.295 2231.625 2794.625 ;
        RECT 2236.830 2791.905 2237.130 2801.450 ;
        RECT 2239.850 2800.000 2240.150 2801.450 ;
        RECT 2242.350 2801.450 2245.990 2801.750 ;
        RECT 2236.815 2791.575 2237.145 2791.905 ;
        RECT 2242.350 2791.225 2242.650 2801.450 ;
        RECT 2245.690 2800.000 2245.990 2801.450 ;
        RECT 2249.710 2801.450 2251.830 2801.750 ;
        RECT 2242.335 2790.895 2242.665 2791.225 ;
        RECT 2249.710 2789.185 2250.010 2801.450 ;
        RECT 2251.530 2800.000 2251.830 2801.450 ;
        RECT 2257.070 2800.000 2257.670 2801.750 ;
        RECT 2257.070 2794.625 2257.370 2800.000 ;
        RECT 2263.210 2796.650 2263.510 2804.600 ;
        RECT 2263.830 2801.750 2264.130 2804.600 ;
        RECT 2269.050 2801.750 2269.350 2804.600 ;
        RECT 2263.830 2801.450 2264.730 2801.750 ;
        RECT 2263.830 2800.000 2264.130 2801.450 ;
        RECT 2263.210 2796.350 2263.810 2796.650 ;
        RECT 2257.055 2794.295 2257.385 2794.625 ;
        RECT 2263.510 2793.265 2263.810 2796.350 ;
        RECT 2264.430 2794.625 2264.730 2801.450 ;
        RECT 2268.110 2801.450 2269.350 2801.750 ;
        RECT 2268.110 2794.625 2268.410 2801.450 ;
        RECT 2269.050 2800.000 2269.350 2801.450 ;
        RECT 2269.670 2796.650 2269.970 2804.600 ;
        RECT 2274.890 2802.450 2275.190 2804.600 ;
        RECT 2269.030 2796.350 2269.970 2796.650 ;
        RECT 2273.630 2802.150 2275.190 2802.450 ;
        RECT 2264.415 2794.295 2264.745 2794.625 ;
        RECT 2268.095 2794.295 2268.425 2794.625 ;
        RECT 2269.030 2793.945 2269.330 2796.350 ;
        RECT 2273.630 2793.945 2273.930 2802.150 ;
        RECT 2274.890 2800.000 2275.190 2802.150 ;
        RECT 2275.510 2801.750 2275.810 2804.600 ;
        RECT 2280.730 2801.750 2281.030 2804.600 ;
        RECT 2275.510 2801.450 2276.690 2801.750 ;
        RECT 2275.510 2800.000 2275.810 2801.450 ;
        RECT 2276.390 2794.625 2276.690 2801.450 ;
        RECT 2280.070 2801.450 2281.030 2801.750 ;
        RECT 2276.375 2794.295 2276.705 2794.625 ;
        RECT 2280.070 2793.945 2280.370 2801.450 ;
        RECT 2280.730 2800.000 2281.030 2801.450 ;
        RECT 2281.350 2802.450 2281.650 2804.600 ;
        RECT 2281.350 2802.150 2283.130 2802.450 ;
        RECT 2281.350 2800.000 2281.650 2802.150 ;
        RECT 2282.830 2794.625 2283.130 2802.150 ;
        RECT 2286.570 2801.750 2286.870 2804.600 ;
        RECT 2286.510 2800.000 2286.870 2801.750 ;
        RECT 2287.190 2801.750 2287.490 2804.600 ;
        RECT 2287.190 2800.000 2287.730 2801.750 ;
        RECT 2292.410 2800.050 2292.710 2804.600 ;
        RECT 2282.815 2794.295 2283.145 2794.625 ;
        RECT 2286.510 2793.945 2286.810 2800.000 ;
        RECT 2287.430 2794.625 2287.730 2800.000 ;
        RECT 2292.030 2799.750 2292.710 2800.050 ;
        RECT 2293.030 2801.750 2293.330 2804.600 ;
        RECT 2298.250 2801.750 2298.550 2804.600 ;
        RECT 2293.030 2801.450 2294.170 2801.750 ;
        RECT 2293.030 2800.000 2293.330 2801.450 ;
        RECT 2287.415 2794.295 2287.745 2794.625 ;
        RECT 2292.030 2793.945 2292.330 2799.750 ;
        RECT 2293.870 2794.625 2294.170 2801.450 ;
        RECT 2297.550 2801.450 2298.550 2801.750 ;
        RECT 2293.855 2794.295 2294.185 2794.625 ;
        RECT 2269.015 2793.615 2269.345 2793.945 ;
        RECT 2273.615 2793.615 2273.945 2793.945 ;
        RECT 2280.055 2793.615 2280.385 2793.945 ;
        RECT 2286.495 2793.615 2286.825 2793.945 ;
        RECT 2292.015 2793.615 2292.345 2793.945 ;
        RECT 2297.550 2793.265 2297.850 2801.450 ;
        RECT 2298.250 2800.000 2298.550 2801.450 ;
        RECT 2298.870 2802.450 2299.170 2804.600 ;
        RECT 2298.870 2802.150 2300.610 2802.450 ;
        RECT 2298.870 2800.000 2299.170 2802.150 ;
        RECT 2300.310 2794.625 2300.610 2802.150 ;
        RECT 2304.090 2801.750 2304.390 2804.600 ;
        RECT 2303.990 2800.000 2304.390 2801.750 ;
        RECT 2304.710 2801.750 2305.010 2804.600 ;
        RECT 2309.930 2801.750 2310.230 2804.600 ;
        RECT 2304.710 2800.000 2305.210 2801.750 ;
        RECT 2300.295 2794.295 2300.625 2794.625 ;
        RECT 2263.495 2792.935 2263.825 2793.265 ;
        RECT 2297.535 2792.935 2297.865 2793.265 ;
        RECT 2249.695 2788.855 2250.025 2789.185 ;
        RECT 2303.990 2788.505 2304.290 2800.000 ;
        RECT 2304.910 2794.625 2305.210 2800.000 ;
        RECT 2308.590 2801.450 2310.230 2801.750 ;
        RECT 2308.590 2794.625 2308.890 2801.450 ;
        RECT 2309.930 2800.000 2310.230 2801.450 ;
        RECT 2310.550 2796.650 2310.850 2804.600 ;
        RECT 2315.770 2801.750 2316.070 2804.600 ;
        RECT 2310.430 2796.350 2310.850 2796.650 ;
        RECT 2315.030 2801.450 2316.070 2801.750 ;
        RECT 2304.895 2794.295 2305.225 2794.625 ;
        RECT 2308.575 2794.295 2308.905 2794.625 ;
        RECT 2310.430 2793.945 2310.730 2796.350 ;
        RECT 2315.030 2793.945 2315.330 2801.450 ;
        RECT 2315.770 2800.000 2316.070 2801.450 ;
        RECT 2316.390 2800.050 2316.690 2804.600 ;
        RECT 2321.610 2801.750 2321.910 2804.600 ;
        RECT 2316.390 2799.750 2317.170 2800.050 ;
        RECT 2316.870 2794.625 2317.170 2799.750 ;
        RECT 2321.470 2800.000 2321.910 2801.750 ;
        RECT 2322.230 2801.750 2322.530 2804.600 ;
        RECT 2327.450 2801.750 2327.750 2804.600 ;
        RECT 2322.230 2800.000 2322.690 2801.750 ;
        RECT 2316.855 2794.295 2317.185 2794.625 ;
        RECT 2321.470 2793.945 2321.770 2800.000 ;
        RECT 2322.390 2794.625 2322.690 2800.000 ;
        RECT 2326.070 2801.450 2327.750 2801.750 ;
        RECT 2322.375 2794.295 2322.705 2794.625 ;
        RECT 2326.070 2793.945 2326.370 2801.450 ;
        RECT 2327.450 2800.000 2327.750 2801.450 ;
        RECT 2328.070 2801.750 2328.370 2804.600 ;
        RECT 2333.290 2801.750 2333.590 2804.600 ;
        RECT 2328.070 2801.450 2329.130 2801.750 ;
        RECT 2328.070 2800.000 2328.370 2801.450 ;
        RECT 2328.830 2794.625 2329.130 2801.450 ;
        RECT 2332.510 2801.450 2333.590 2801.750 ;
        RECT 2328.815 2794.295 2329.145 2794.625 ;
        RECT 2332.510 2793.945 2332.810 2801.450 ;
        RECT 2333.290 2800.000 2333.590 2801.450 ;
        RECT 2333.910 2800.050 2334.210 2804.600 ;
        RECT 2339.130 2801.750 2339.430 2804.600 ;
        RECT 2333.910 2799.750 2334.650 2800.050 ;
        RECT 2334.350 2794.625 2334.650 2799.750 ;
        RECT 2338.950 2800.000 2339.430 2801.750 ;
        RECT 2339.750 2801.750 2340.050 2804.600 ;
        RECT 2344.970 2802.450 2345.270 2804.600 ;
        RECT 2343.550 2802.150 2345.270 2802.450 ;
        RECT 2339.750 2800.000 2340.170 2801.750 ;
        RECT 2334.335 2794.295 2334.665 2794.625 ;
        RECT 2310.415 2793.615 2310.745 2793.945 ;
        RECT 2315.015 2793.615 2315.345 2793.945 ;
        RECT 2321.455 2793.615 2321.785 2793.945 ;
        RECT 2326.055 2793.615 2326.385 2793.945 ;
        RECT 2332.495 2793.615 2332.825 2793.945 ;
        RECT 2338.950 2793.265 2339.250 2800.000 ;
        RECT 2339.870 2794.625 2340.170 2800.000 ;
        RECT 2343.550 2794.625 2343.850 2802.150 ;
        RECT 2344.970 2800.000 2345.270 2802.150 ;
        RECT 2345.590 2796.650 2345.890 2804.600 ;
        RECT 2350.810 2801.750 2351.110 2804.600 ;
        RECT 2345.390 2796.350 2345.890 2796.650 ;
        RECT 2349.990 2801.450 2351.110 2801.750 ;
        RECT 2339.855 2794.295 2340.185 2794.625 ;
        RECT 2343.535 2794.295 2343.865 2794.625 ;
        RECT 2345.390 2793.945 2345.690 2796.350 ;
        RECT 2345.375 2793.615 2345.705 2793.945 ;
        RECT 2349.990 2793.265 2350.290 2801.450 ;
        RECT 2350.810 2800.000 2351.110 2801.450 ;
        RECT 2351.430 2800.050 2351.730 2804.600 ;
        RECT 2356.650 2801.750 2356.950 2804.600 ;
        RECT 2351.430 2799.750 2352.130 2800.050 ;
        RECT 2351.830 2794.625 2352.130 2799.750 ;
        RECT 2356.430 2800.000 2356.950 2801.750 ;
        RECT 2357.270 2801.750 2357.570 2804.600 ;
        RECT 2362.490 2802.450 2362.790 2804.600 ;
        RECT 2361.030 2802.150 2362.790 2802.450 ;
        RECT 2357.270 2800.000 2357.650 2801.750 ;
        RECT 2351.815 2794.295 2352.145 2794.625 ;
        RECT 2356.430 2793.945 2356.730 2800.000 ;
        RECT 2357.350 2794.625 2357.650 2800.000 ;
        RECT 2357.335 2794.295 2357.665 2794.625 ;
        RECT 2361.030 2793.945 2361.330 2802.150 ;
        RECT 2362.490 2800.000 2362.790 2802.150 ;
        RECT 2363.110 2801.750 2363.410 2804.600 ;
        RECT 2368.330 2801.750 2368.630 2804.600 ;
        RECT 2363.110 2801.450 2364.090 2801.750 ;
        RECT 2363.110 2800.000 2363.410 2801.450 ;
        RECT 2363.790 2794.625 2364.090 2801.450 ;
        RECT 2367.470 2801.450 2368.630 2801.750 ;
        RECT 2363.775 2794.295 2364.105 2794.625 ;
        RECT 2367.470 2793.945 2367.770 2801.450 ;
        RECT 2368.330 2800.000 2368.630 2801.450 ;
        RECT 2368.950 2802.450 2369.250 2804.600 ;
        RECT 2368.950 2802.150 2370.530 2802.450 ;
        RECT 2368.950 2800.000 2369.250 2802.150 ;
        RECT 2370.230 2794.625 2370.530 2802.150 ;
        RECT 2374.170 2801.750 2374.470 2804.600 ;
        RECT 2373.910 2800.000 2374.470 2801.750 ;
        RECT 2374.790 2801.750 2375.090 2804.600 ;
        RECT 2380.010 2801.750 2380.310 2804.600 ;
        RECT 2374.790 2800.000 2375.130 2801.750 ;
        RECT 2370.215 2794.295 2370.545 2794.625 ;
        RECT 2373.910 2793.945 2374.210 2800.000 ;
        RECT 2374.830 2794.625 2375.130 2800.000 ;
        RECT 2377.590 2801.450 2380.310 2801.750 ;
        RECT 2377.590 2794.625 2377.890 2801.450 ;
        RECT 2380.010 2800.000 2380.310 2801.450 ;
        RECT 2380.630 2801.750 2380.930 2804.600 ;
        RECT 2385.850 2801.750 2386.150 2804.600 ;
        RECT 2380.630 2801.450 2381.570 2801.750 ;
        RECT 2380.630 2800.000 2380.930 2801.450 ;
        RECT 2381.270 2794.625 2381.570 2801.450 ;
        RECT 2383.110 2801.450 2386.150 2801.750 ;
        RECT 2383.110 2794.625 2383.410 2801.450 ;
        RECT 2385.850 2800.000 2386.150 2801.450 ;
        RECT 2386.470 2800.050 2386.770 2804.600 ;
        RECT 2391.690 2801.750 2391.990 2804.600 ;
        RECT 2389.550 2801.450 2391.990 2801.750 ;
        RECT 2386.470 2799.750 2387.090 2800.050 ;
        RECT 2374.815 2794.295 2375.145 2794.625 ;
        RECT 2377.575 2794.295 2377.905 2794.625 ;
        RECT 2381.255 2794.295 2381.585 2794.625 ;
        RECT 2383.095 2794.295 2383.425 2794.625 ;
        RECT 2356.415 2793.615 2356.745 2793.945 ;
        RECT 2361.015 2793.615 2361.345 2793.945 ;
        RECT 2367.455 2793.615 2367.785 2793.945 ;
        RECT 2373.895 2793.615 2374.225 2793.945 ;
        RECT 2386.790 2793.265 2387.090 2799.750 ;
        RECT 2389.550 2794.625 2389.850 2801.450 ;
        RECT 2391.690 2800.000 2391.990 2801.450 ;
        RECT 2389.535 2794.295 2389.865 2794.625 ;
        RECT 2338.935 2792.935 2339.265 2793.265 ;
        RECT 2349.975 2792.935 2350.305 2793.265 ;
        RECT 2386.775 2792.935 2387.105 2793.265 ;
        RECT 2392.310 2791.905 2392.610 2804.600 ;
        RECT 2397.530 2801.750 2397.830 2804.600 ;
        RECT 2395.070 2801.450 2397.830 2801.750 ;
        RECT 2395.070 2794.625 2395.370 2801.450 ;
        RECT 2397.530 2800.000 2397.830 2801.450 ;
        RECT 2398.150 2801.750 2398.450 2804.600 ;
        RECT 2403.370 2801.750 2403.670 2804.600 ;
        RECT 2398.150 2801.450 2399.050 2801.750 ;
        RECT 2398.150 2800.000 2398.450 2801.450 ;
        RECT 2395.055 2794.295 2395.385 2794.625 ;
        RECT 2398.750 2792.585 2399.050 2801.450 ;
        RECT 2402.430 2801.450 2403.670 2801.750 ;
        RECT 2402.430 2794.625 2402.730 2801.450 ;
        RECT 2403.370 2800.000 2403.670 2801.450 ;
        RECT 2403.990 2801.750 2404.290 2804.600 ;
        RECT 2409.210 2802.450 2409.510 2804.600 ;
        RECT 2407.950 2802.150 2409.510 2802.450 ;
        RECT 2403.990 2800.000 2404.570 2801.750 ;
        RECT 2402.415 2794.295 2402.745 2794.625 ;
        RECT 2398.735 2792.255 2399.065 2792.585 ;
        RECT 2404.270 2791.905 2404.570 2800.000 ;
        RECT 2407.950 2793.265 2408.250 2802.150 ;
        RECT 2409.210 2800.000 2409.510 2802.150 ;
        RECT 2409.830 2801.750 2410.130 2804.600 ;
        RECT 2409.830 2801.450 2411.010 2801.750 ;
        RECT 2409.830 2800.000 2410.130 2801.450 ;
        RECT 2407.935 2792.935 2408.265 2793.265 ;
        RECT 2410.710 2792.585 2411.010 2801.450 ;
        RECT 2415.050 2796.650 2415.350 2804.600 ;
        RECT 2415.670 2802.450 2415.970 2804.600 ;
        RECT 2415.670 2802.150 2417.450 2802.450 ;
        RECT 2415.670 2800.000 2415.970 2802.150 ;
        RECT 2415.050 2796.350 2415.610 2796.650 ;
        RECT 2415.310 2792.585 2415.610 2796.350 ;
        RECT 2410.695 2792.255 2411.025 2792.585 ;
        RECT 2415.295 2792.255 2415.625 2792.585 ;
        RECT 2392.295 2791.575 2392.625 2791.905 ;
        RECT 2404.255 2791.575 2404.585 2791.905 ;
        RECT 2417.150 2789.865 2417.450 2802.150 ;
        RECT 2420.890 2801.750 2421.190 2804.600 ;
        RECT 2418.070 2801.450 2421.190 2801.750 ;
        RECT 2417.135 2789.535 2417.465 2789.865 ;
        RECT 2418.070 2789.185 2418.370 2801.450 ;
        RECT 2420.890 2800.000 2421.190 2801.450 ;
        RECT 2421.510 2796.650 2421.810 2804.600 ;
        RECT 2426.730 2801.750 2427.030 2804.600 ;
        RECT 2420.830 2796.350 2421.810 2796.650 ;
        RECT 2423.590 2801.450 2427.030 2801.750 ;
        RECT 2420.830 2791.225 2421.130 2796.350 ;
        RECT 2423.590 2793.945 2423.890 2801.450 ;
        RECT 2426.730 2800.000 2427.030 2801.450 ;
        RECT 2427.350 2801.750 2427.650 2804.600 ;
        RECT 2432.570 2801.750 2432.870 2804.600 ;
        RECT 2427.350 2801.450 2428.490 2801.750 ;
        RECT 2427.350 2800.000 2427.650 2801.450 ;
        RECT 2423.575 2793.615 2423.905 2793.945 ;
        RECT 2420.815 2790.895 2421.145 2791.225 ;
        RECT 2428.190 2790.545 2428.490 2801.450 ;
        RECT 2430.030 2801.450 2432.870 2801.750 ;
        RECT 2430.030 2792.585 2430.330 2801.450 ;
        RECT 2432.570 2800.000 2432.870 2801.450 ;
        RECT 2433.190 2802.450 2433.490 2804.600 ;
        RECT 2433.190 2802.150 2434.930 2802.450 ;
        RECT 2433.190 2800.000 2433.490 2802.150 ;
        RECT 2430.015 2792.255 2430.345 2792.585 ;
        RECT 2428.175 2790.215 2428.505 2790.545 ;
        RECT 2434.630 2789.865 2434.930 2802.150 ;
        RECT 2438.410 2801.750 2438.710 2804.600 ;
        RECT 2436.470 2801.450 2438.710 2801.750 ;
        RECT 2436.470 2792.585 2436.770 2801.450 ;
        RECT 2438.410 2800.000 2438.710 2801.450 ;
        RECT 2439.030 2801.750 2439.330 2804.600 ;
        RECT 2444.250 2801.750 2444.550 2804.600 ;
        RECT 2439.030 2800.000 2439.530 2801.750 ;
        RECT 2436.455 2792.255 2436.785 2792.585 ;
        RECT 2434.615 2789.535 2434.945 2789.865 ;
        RECT 2439.230 2789.185 2439.530 2800.000 ;
        RECT 2442.910 2801.450 2444.550 2801.750 ;
        RECT 2442.910 2791.905 2443.210 2801.450 ;
        RECT 2444.250 2800.000 2444.550 2801.450 ;
        RECT 2444.870 2801.750 2445.170 2804.600 ;
        RECT 2444.870 2801.450 2445.970 2801.750 ;
        RECT 2444.870 2800.000 2445.170 2801.450 ;
        RECT 2442.895 2791.575 2443.225 2791.905 ;
        RECT 2418.055 2788.855 2418.385 2789.185 ;
        RECT 2439.215 2788.855 2439.545 2789.185 ;
        RECT 2445.670 2788.505 2445.970 2801.450 ;
        RECT 2303.975 2788.175 2304.305 2788.505 ;
        RECT 2445.655 2788.175 2445.985 2788.505 ;
        RECT 1761.175 2777.295 1761.505 2777.625 ;
        RECT 1796.135 2777.295 1796.465 2777.625 ;
        RECT 1841.215 2069.415 1841.545 2069.745 ;
        RECT 1844.895 2069.415 1845.225 2069.745 ;
        RECT 1851.335 2069.415 1851.665 2069.745 ;
        RECT 1859.615 2069.415 1859.945 2069.745 ;
        RECT 1865.135 2069.415 1865.465 2069.745 ;
        RECT 1901.015 2069.415 1901.345 2069.745 ;
        RECT 1923.095 2069.415 1923.425 2069.745 ;
        RECT 1941.495 2069.415 1941.825 2069.745 ;
        RECT 1953.455 2069.415 1953.785 2069.745 ;
        RECT 1964.495 2069.415 1964.825 2069.745 ;
        RECT 1989.335 2069.415 1989.665 2069.745 ;
        RECT 2015.095 2069.415 2015.425 2069.745 ;
        RECT 2039.015 2069.415 2039.345 2069.745 ;
        RECT 2052.815 2069.415 2053.145 2069.745 ;
        RECT 2354.575 2069.415 2354.905 2069.745 ;
        RECT 2373.895 2069.415 2374.225 2069.745 ;
        RECT 2391.375 2069.415 2391.705 2069.745 ;
        RECT 1838.455 2063.295 1838.785 2063.625 ;
        RECT 1838.470 2055.450 1838.770 2063.295 ;
        RECT 1841.230 2058.850 1841.530 2069.415 ;
        RECT 1841.230 2058.550 1842.230 2058.850 ;
        RECT 1841.310 2055.450 1841.610 2056.235 ;
        RECT 1838.470 2055.150 1841.610 2055.450 ;
        RECT 1841.310 2051.635 1841.610 2055.150 ;
        RECT 1841.930 2051.635 1842.230 2058.550 ;
        RECT 1844.910 2055.450 1845.210 2069.415 ;
        RECT 1847.655 2065.335 1847.985 2065.665 ;
        RECT 1847.670 2058.850 1847.970 2065.335 ;
        RECT 1847.670 2058.550 1848.070 2058.850 ;
        RECT 1847.150 2055.450 1847.450 2056.235 ;
        RECT 1844.910 2055.150 1847.450 2055.450 ;
        RECT 1847.150 2051.635 1847.450 2055.150 ;
        RECT 1847.770 2051.635 1848.070 2058.550 ;
        RECT 1851.350 2055.450 1851.650 2069.415 ;
        RECT 1854.095 2065.335 1854.425 2065.665 ;
        RECT 1854.110 2058.850 1854.410 2065.335 ;
        RECT 1856.855 2063.295 1857.185 2063.625 ;
        RECT 1853.610 2058.550 1854.410 2058.850 ;
        RECT 1852.990 2055.450 1853.290 2056.235 ;
        RECT 1851.350 2055.150 1853.290 2055.450 ;
        RECT 1852.990 2051.635 1853.290 2055.150 ;
        RECT 1853.610 2051.635 1853.910 2058.550 ;
        RECT 1856.870 2055.450 1857.170 2063.295 ;
        RECT 1859.630 2056.235 1859.930 2069.415 ;
        RECT 1863.295 2063.295 1863.625 2063.625 ;
        RECT 1858.830 2055.450 1859.130 2056.235 ;
        RECT 1856.870 2055.150 1859.130 2055.450 ;
        RECT 1858.830 2051.635 1859.130 2055.150 ;
        RECT 1859.450 2055.150 1859.930 2056.235 ;
        RECT 1859.450 2051.635 1859.750 2055.150 ;
        RECT 1863.310 2053.750 1863.610 2063.295 ;
        RECT 1865.150 2058.850 1865.450 2069.415 ;
        RECT 1871.575 2066.015 1871.905 2066.345 ;
        RECT 1877.095 2066.015 1877.425 2066.345 ;
        RECT 1879.855 2066.015 1880.185 2066.345 ;
        RECT 1889.055 2066.015 1889.385 2066.345 ;
        RECT 1894.575 2066.015 1894.905 2066.345 ;
        RECT 1869.735 2063.975 1870.065 2064.305 ;
        RECT 1865.150 2058.550 1865.590 2058.850 ;
        RECT 1864.670 2053.750 1864.970 2056.235 ;
        RECT 1863.310 2053.450 1864.970 2053.750 ;
        RECT 1864.670 2051.635 1864.970 2053.450 ;
        RECT 1865.290 2051.635 1865.590 2058.550 ;
        RECT 1869.750 2055.450 1870.050 2063.975 ;
        RECT 1871.590 2058.850 1871.890 2066.015 ;
        RECT 1873.415 2063.295 1873.745 2063.625 ;
        RECT 1871.130 2058.550 1871.890 2058.850 ;
        RECT 1870.510 2055.450 1870.810 2056.235 ;
        RECT 1869.750 2055.150 1870.810 2055.450 ;
        RECT 1870.510 2051.635 1870.810 2055.150 ;
        RECT 1871.130 2051.635 1871.430 2058.550 ;
        RECT 1873.430 2055.450 1873.730 2063.295 ;
        RECT 1877.110 2056.235 1877.410 2066.015 ;
        RECT 1876.350 2055.450 1876.650 2056.235 ;
        RECT 1873.430 2055.150 1876.650 2055.450 ;
        RECT 1876.350 2051.635 1876.650 2055.150 ;
        RECT 1876.970 2055.150 1877.410 2056.235 ;
        RECT 1879.870 2055.450 1880.170 2066.015 ;
        RECT 1882.615 2065.335 1882.945 2065.665 ;
        RECT 1882.630 2058.850 1882.930 2065.335 ;
        RECT 1886.295 2063.975 1886.625 2064.305 ;
        RECT 1882.630 2058.550 1883.110 2058.850 ;
        RECT 1882.190 2055.450 1882.490 2056.235 ;
        RECT 1879.870 2055.150 1882.490 2055.450 ;
        RECT 1876.970 2051.635 1877.270 2055.150 ;
        RECT 1882.190 2051.635 1882.490 2055.150 ;
        RECT 1882.810 2051.635 1883.110 2058.550 ;
        RECT 1886.310 2055.450 1886.610 2063.975 ;
        RECT 1889.070 2058.850 1889.370 2066.015 ;
        RECT 1890.895 2063.975 1891.225 2064.305 ;
        RECT 1888.650 2058.550 1889.370 2058.850 ;
        RECT 1888.030 2055.450 1888.330 2056.235 ;
        RECT 1886.310 2055.150 1888.330 2055.450 ;
        RECT 1888.030 2051.635 1888.330 2055.150 ;
        RECT 1888.650 2051.635 1888.950 2058.550 ;
        RECT 1890.910 2055.450 1891.210 2063.975 ;
        RECT 1894.590 2056.235 1894.890 2066.015 ;
        RECT 1898.255 2063.975 1898.585 2064.305 ;
        RECT 1893.870 2055.450 1894.170 2056.235 ;
        RECT 1890.910 2055.150 1894.170 2055.450 ;
        RECT 1893.870 2051.635 1894.170 2055.150 ;
        RECT 1894.490 2055.150 1894.890 2056.235 ;
        RECT 1894.490 2051.635 1894.790 2055.150 ;
        RECT 1898.270 2053.750 1898.570 2063.975 ;
        RECT 1899.710 2053.750 1900.010 2056.235 ;
        RECT 1898.270 2053.450 1900.010 2053.750 ;
        RECT 1899.710 2051.635 1900.010 2053.450 ;
        RECT 1900.330 2055.450 1900.630 2056.235 ;
        RECT 1901.030 2055.450 1901.330 2069.415 ;
        RECT 1907.455 2066.695 1907.785 2067.025 ;
        RECT 1912.055 2066.695 1912.385 2067.025 ;
        RECT 1904.695 2063.295 1905.025 2063.625 ;
        RECT 1900.330 2055.150 1901.330 2055.450 ;
        RECT 1904.710 2055.450 1905.010 2063.295 ;
        RECT 1905.550 2055.450 1905.850 2056.235 ;
        RECT 1904.710 2055.150 1905.850 2055.450 ;
        RECT 1900.330 2051.635 1900.630 2055.150 ;
        RECT 1905.550 2051.635 1905.850 2055.150 ;
        RECT 1906.170 2053.750 1906.470 2056.235 ;
        RECT 1907.470 2053.750 1907.770 2066.695 ;
        RECT 1911.135 2065.335 1911.465 2065.665 ;
        RECT 1911.150 2056.235 1911.450 2065.335 ;
        RECT 1912.070 2056.235 1912.370 2066.695 ;
        RECT 1913.895 2065.335 1914.225 2065.665 ;
        RECT 1911.150 2055.150 1911.690 2056.235 ;
        RECT 1906.170 2053.450 1907.770 2053.750 ;
        RECT 1906.170 2051.635 1906.470 2053.450 ;
        RECT 1911.390 2051.635 1911.690 2055.150 ;
        RECT 1912.010 2055.150 1912.370 2056.235 ;
        RECT 1913.910 2055.450 1914.210 2065.335 ;
        RECT 1917.575 2063.295 1917.905 2063.625 ;
        RECT 1920.335 2063.295 1920.665 2063.625 ;
        RECT 1917.590 2058.850 1917.890 2063.295 ;
        RECT 1917.590 2058.550 1918.150 2058.850 ;
        RECT 1917.230 2055.450 1917.530 2056.235 ;
        RECT 1913.910 2055.150 1917.530 2055.450 ;
        RECT 1912.010 2051.635 1912.310 2055.150 ;
        RECT 1917.230 2051.635 1917.530 2055.150 ;
        RECT 1917.850 2051.635 1918.150 2058.550 ;
        RECT 1920.350 2055.450 1920.650 2063.295 ;
        RECT 1923.110 2058.850 1923.410 2069.415 ;
        RECT 1932.295 2067.375 1932.625 2067.705 ;
        RECT 1925.855 2065.335 1926.185 2065.665 ;
        RECT 1923.110 2058.550 1923.990 2058.850 ;
        RECT 1923.070 2055.450 1923.370 2056.235 ;
        RECT 1920.350 2055.150 1923.370 2055.450 ;
        RECT 1923.070 2051.635 1923.370 2055.150 ;
        RECT 1923.690 2051.635 1923.990 2058.550 ;
        RECT 1925.870 2055.450 1926.170 2065.335 ;
        RECT 1929.535 2063.295 1929.865 2063.625 ;
        RECT 1929.550 2056.235 1929.850 2063.295 ;
        RECT 1928.910 2055.450 1929.210 2056.235 ;
        RECT 1925.870 2055.150 1929.210 2055.450 ;
        RECT 1928.910 2051.635 1929.210 2055.150 ;
        RECT 1929.530 2055.150 1929.850 2056.235 ;
        RECT 1932.310 2055.450 1932.610 2067.375 ;
        RECT 1935.975 2066.015 1936.305 2066.345 ;
        RECT 1934.750 2055.450 1935.050 2056.235 ;
        RECT 1932.310 2055.150 1935.050 2055.450 ;
        RECT 1929.530 2051.635 1929.830 2055.150 ;
        RECT 1934.750 2051.635 1935.050 2055.150 ;
        RECT 1935.370 2055.450 1935.670 2056.235 ;
        RECT 1935.990 2055.450 1936.290 2066.015 ;
        RECT 1940.575 2063.295 1940.905 2063.625 ;
        RECT 1935.370 2055.150 1936.290 2055.450 ;
        RECT 1935.370 2051.635 1935.670 2055.150 ;
        RECT 1940.590 2051.635 1940.890 2063.295 ;
        RECT 1941.510 2056.235 1941.810 2069.415 ;
        RECT 1947.015 2068.055 1947.345 2068.385 ;
        RECT 1946.095 2067.375 1946.425 2067.705 ;
        RECT 1946.110 2058.850 1946.410 2067.375 ;
        RECT 1947.030 2058.850 1947.330 2068.055 ;
        RECT 1948.855 2064.655 1949.185 2064.985 ;
        RECT 1946.110 2058.550 1946.730 2058.850 ;
        RECT 1947.030 2058.550 1947.350 2058.850 ;
        RECT 1941.210 2055.150 1941.810 2056.235 ;
        RECT 1941.210 2051.635 1941.510 2055.150 ;
        RECT 1946.430 2051.635 1946.730 2058.550 ;
        RECT 1947.050 2051.635 1947.350 2058.550 ;
        RECT 1948.870 2055.450 1949.170 2064.655 ;
        RECT 1953.470 2058.850 1953.770 2069.415 ;
        RECT 1960.815 2068.735 1961.145 2069.065 ;
        RECT 1958.975 2065.335 1959.305 2065.665 ;
        RECT 1955.295 2064.655 1955.625 2064.985 ;
        RECT 1952.890 2058.550 1953.770 2058.850 ;
        RECT 1952.270 2055.450 1952.570 2056.235 ;
        RECT 1948.870 2055.150 1952.570 2055.450 ;
        RECT 1952.270 2051.635 1952.570 2055.150 ;
        RECT 1952.890 2051.635 1953.190 2058.550 ;
        RECT 1955.310 2055.450 1955.610 2064.655 ;
        RECT 1958.990 2056.235 1959.290 2065.335 ;
        RECT 1958.110 2055.450 1958.410 2056.235 ;
        RECT 1955.310 2055.150 1958.410 2055.450 ;
        RECT 1958.110 2051.635 1958.410 2055.150 ;
        RECT 1958.730 2055.150 1959.290 2056.235 ;
        RECT 1960.830 2055.450 1961.130 2068.735 ;
        RECT 1964.510 2058.850 1964.810 2069.415 ;
        RECT 1980.135 2068.735 1980.465 2069.065 ;
        RECT 1973.695 2067.375 1974.025 2067.705 ;
        RECT 1967.255 2064.655 1967.585 2064.985 ;
        RECT 1964.510 2058.550 1964.870 2058.850 ;
        RECT 1963.950 2055.450 1964.250 2056.235 ;
        RECT 1960.830 2055.150 1964.250 2055.450 ;
        RECT 1958.730 2051.635 1959.030 2055.150 ;
        RECT 1963.950 2051.635 1964.250 2055.150 ;
        RECT 1964.570 2051.635 1964.870 2058.550 ;
        RECT 1967.270 2055.450 1967.570 2064.655 ;
        RECT 1970.935 2063.295 1971.265 2063.625 ;
        RECT 1970.950 2058.850 1971.250 2063.295 ;
        RECT 1970.410 2058.550 1971.250 2058.850 ;
        RECT 1969.790 2055.450 1970.090 2056.235 ;
        RECT 1967.270 2055.150 1970.090 2055.450 ;
        RECT 1969.790 2051.635 1970.090 2055.150 ;
        RECT 1970.410 2051.635 1970.710 2058.550 ;
        RECT 1973.710 2055.450 1974.010 2067.375 ;
        RECT 1976.455 2063.975 1976.785 2064.305 ;
        RECT 1976.470 2056.235 1976.770 2063.975 ;
        RECT 1975.630 2055.450 1975.930 2056.235 ;
        RECT 1973.710 2055.150 1975.930 2055.450 ;
        RECT 1975.630 2051.635 1975.930 2055.150 ;
        RECT 1976.250 2055.150 1976.770 2056.235 ;
        RECT 1976.250 2051.635 1976.550 2055.150 ;
        RECT 1980.150 2053.750 1980.450 2068.735 ;
        RECT 1987.495 2066.695 1987.825 2067.025 ;
        RECT 1981.975 2064.655 1982.305 2064.985 ;
        RECT 1981.990 2058.850 1982.290 2064.655 ;
        RECT 1987.510 2058.850 1987.810 2066.695 ;
        RECT 1981.990 2058.550 1982.390 2058.850 ;
        RECT 1981.470 2053.750 1981.770 2056.235 ;
        RECT 1980.150 2053.450 1981.770 2053.750 ;
        RECT 1981.470 2051.635 1981.770 2053.450 ;
        RECT 1982.090 2051.635 1982.390 2058.550 ;
        RECT 1987.310 2058.550 1987.810 2058.850 ;
        RECT 1987.310 2051.635 1987.610 2058.550 ;
        RECT 1987.930 2053.750 1988.230 2056.235 ;
        RECT 1989.350 2053.750 1989.650 2069.415 ;
        RECT 2007.735 2067.375 2008.065 2067.705 ;
        RECT 1990.255 2065.335 1990.585 2065.665 ;
        RECT 1999.455 2065.335 1999.785 2065.665 ;
        RECT 1990.270 2055.450 1990.570 2065.335 ;
        RECT 1993.015 2064.655 1993.345 2064.985 ;
        RECT 1993.030 2058.850 1993.330 2064.655 ;
        RECT 1995.775 2063.295 1996.105 2063.625 ;
        RECT 1993.030 2058.550 1994.070 2058.850 ;
        RECT 1993.150 2055.450 1993.450 2056.235 ;
        RECT 1990.270 2055.150 1993.450 2055.450 ;
        RECT 1987.930 2053.450 1989.650 2053.750 ;
        RECT 1987.930 2051.635 1988.230 2053.450 ;
        RECT 1993.150 2051.635 1993.450 2055.150 ;
        RECT 1993.770 2051.635 1994.070 2058.550 ;
        RECT 1995.790 2055.450 1996.090 2063.295 ;
        RECT 1999.470 2058.850 1999.770 2065.335 ;
        RECT 2002.215 2063.975 2002.545 2064.305 ;
        RECT 1999.470 2058.550 1999.910 2058.850 ;
        RECT 1998.990 2055.450 1999.290 2056.235 ;
        RECT 1995.790 2055.150 1999.290 2055.450 ;
        RECT 1998.990 2051.635 1999.290 2055.150 ;
        RECT 1999.610 2051.635 1999.910 2058.550 ;
        RECT 2002.230 2055.450 2002.530 2063.975 ;
        RECT 2005.895 2063.295 2006.225 2063.625 ;
        RECT 2005.910 2058.850 2006.210 2063.295 ;
        RECT 2005.450 2058.550 2006.210 2058.850 ;
        RECT 2004.830 2055.450 2005.130 2056.235 ;
        RECT 2002.230 2055.150 2005.130 2055.450 ;
        RECT 2004.830 2051.635 2005.130 2055.150 ;
        RECT 2005.450 2051.635 2005.750 2058.550 ;
        RECT 2007.750 2055.450 2008.050 2067.375 ;
        RECT 2011.415 2066.695 2011.745 2067.025 ;
        RECT 2011.430 2056.235 2011.730 2066.695 ;
        RECT 2010.670 2055.450 2010.970 2056.235 ;
        RECT 2007.750 2055.150 2010.970 2055.450 ;
        RECT 2010.670 2051.635 2010.970 2055.150 ;
        RECT 2011.290 2055.150 2011.730 2056.235 ;
        RECT 2015.110 2055.450 2015.410 2069.415 ;
        RECT 2021.535 2067.375 2021.865 2067.705 ;
        RECT 2016.935 2063.975 2017.265 2064.305 ;
        RECT 2016.950 2058.850 2017.250 2063.975 ;
        RECT 2016.950 2058.550 2017.430 2058.850 ;
        RECT 2016.510 2055.450 2016.810 2056.235 ;
        RECT 2015.110 2055.150 2016.810 2055.450 ;
        RECT 2011.290 2051.635 2011.590 2055.150 ;
        RECT 2016.510 2051.635 2016.810 2055.150 ;
        RECT 2017.130 2051.635 2017.430 2058.550 ;
        RECT 2021.550 2055.450 2021.850 2067.375 ;
        RECT 2023.375 2066.015 2023.705 2066.345 ;
        RECT 2023.390 2058.850 2023.690 2066.015 ;
        RECT 2022.970 2058.550 2023.690 2058.850 ;
        RECT 2022.350 2055.450 2022.650 2056.235 ;
        RECT 2021.550 2055.150 2022.650 2055.450 ;
        RECT 2022.350 2051.635 2022.650 2055.150 ;
        RECT 2022.970 2051.635 2023.270 2058.550 ;
        RECT 2028.795 2057.175 2029.125 2057.505 ;
        RECT 2028.810 2055.450 2029.110 2057.175 ;
        RECT 2034.650 2055.450 2034.950 2056.235 ;
        RECT 2039.030 2055.450 2039.330 2069.415 ;
        RECT 2040.490 2055.450 2040.790 2056.235 ;
        RECT 2046.330 2055.450 2046.630 2056.235 ;
        RECT 2028.810 2055.150 2046.630 2055.450 ;
        RECT 2028.810 2051.635 2029.110 2055.150 ;
        RECT 2034.650 2051.635 2034.950 2055.150 ;
        RECT 2040.490 2051.635 2040.790 2055.150 ;
        RECT 2046.330 2051.635 2046.630 2055.150 ;
        RECT 2052.170 2055.450 2052.470 2056.235 ;
        RECT 2052.830 2055.450 2053.130 2069.415 ;
        RECT 2340.775 2063.295 2341.105 2063.625 ;
        RECT 2347.215 2063.295 2347.545 2063.625 ;
        RECT 2052.170 2055.150 2053.130 2055.450 ;
        RECT 2340.790 2055.450 2341.090 2063.295 ;
        RECT 2344.025 2055.450 2344.325 2056.235 ;
        RECT 2340.790 2055.150 2344.325 2055.450 ;
        RECT 2347.230 2055.450 2347.530 2063.295 ;
        RECT 2350.265 2055.450 2350.565 2056.235 ;
        RECT 2347.230 2055.150 2350.565 2055.450 ;
        RECT 2354.590 2055.450 2354.890 2069.415 ;
        RECT 2360.095 2063.295 2360.425 2063.625 ;
        RECT 2356.505 2055.450 2356.805 2056.235 ;
        RECT 2354.590 2055.150 2356.805 2055.450 ;
        RECT 2360.110 2055.450 2360.410 2063.295 ;
        RECT 2362.745 2055.450 2363.045 2056.235 ;
        RECT 2360.110 2055.150 2363.045 2055.450 ;
        RECT 2052.170 2051.635 2052.470 2055.150 ;
        RECT 2344.025 2051.635 2344.325 2055.150 ;
        RECT 2350.265 2051.635 2350.565 2055.150 ;
        RECT 2356.505 2051.635 2356.805 2055.150 ;
        RECT 2362.745 2051.635 2363.045 2055.150 ;
        RECT 2367.225 2052.050 2367.555 2052.065 ;
        RECT 2368.985 2052.050 2369.285 2056.235 ;
        RECT 2373.910 2053.750 2374.210 2069.415 ;
        RECT 2381.255 2068.735 2381.585 2069.065 ;
        RECT 2387.695 2068.735 2388.025 2069.065 ;
        RECT 2381.270 2056.235 2381.570 2068.735 ;
        RECT 2387.710 2056.235 2388.010 2068.735 ;
        RECT 2375.225 2053.750 2375.525 2056.235 ;
        RECT 2381.270 2055.150 2381.765 2056.235 ;
        RECT 2373.910 2053.450 2375.525 2053.750 ;
        RECT 2367.225 2051.750 2369.285 2052.050 ;
        RECT 2367.225 2051.735 2367.555 2051.750 ;
        RECT 2368.985 2051.635 2369.285 2051.750 ;
        RECT 2375.225 2051.635 2375.525 2053.450 ;
        RECT 2381.465 2051.635 2381.765 2055.150 ;
        RECT 2387.705 2055.150 2388.010 2056.235 ;
        RECT 2391.390 2055.450 2391.690 2069.415 ;
        RECT 2528.455 2068.735 2528.785 2069.065 ;
        RECT 2396.895 2068.055 2397.225 2068.385 ;
        RECT 2393.945 2055.450 2394.245 2056.235 ;
        RECT 2391.390 2055.150 2394.245 2055.450 ;
        RECT 2396.910 2055.450 2397.210 2068.055 ;
        RECT 2403.335 2067.375 2403.665 2067.705 ;
        RECT 2429.095 2067.375 2429.425 2067.705 ;
        RECT 2400.185 2055.450 2400.485 2056.235 ;
        RECT 2396.910 2055.150 2400.485 2055.450 ;
        RECT 2403.350 2055.450 2403.650 2067.375 ;
        RECT 2409.775 2066.695 2410.105 2067.025 ;
        RECT 2417.135 2066.695 2417.465 2067.025 ;
        RECT 2406.425 2055.450 2406.725 2056.235 ;
        RECT 2403.350 2055.150 2406.725 2055.450 ;
        RECT 2409.790 2055.450 2410.090 2066.695 ;
        RECT 2412.665 2055.450 2412.965 2056.235 ;
        RECT 2409.790 2055.150 2412.965 2055.450 ;
        RECT 2417.150 2055.450 2417.450 2066.695 ;
        RECT 2422.655 2066.015 2422.985 2066.345 ;
        RECT 2418.905 2055.450 2419.205 2056.235 ;
        RECT 2417.150 2055.150 2419.205 2055.450 ;
        RECT 2422.670 2055.450 2422.970 2066.015 ;
        RECT 2425.145 2055.450 2425.445 2056.235 ;
        RECT 2422.670 2055.150 2425.445 2055.450 ;
        RECT 2429.110 2055.450 2429.410 2067.375 ;
        RECT 2442.895 2066.015 2443.225 2066.345 ;
        RECT 2436.455 2065.335 2436.785 2065.665 ;
        RECT 2431.385 2055.450 2431.685 2056.235 ;
        RECT 2429.110 2055.150 2431.685 2055.450 ;
        RECT 2436.470 2055.450 2436.770 2065.335 ;
        RECT 2437.625 2055.450 2437.925 2056.235 ;
        RECT 2436.470 2055.150 2437.925 2055.450 ;
        RECT 2442.910 2055.450 2443.210 2066.015 ;
        RECT 2450.255 2064.655 2450.585 2064.985 ;
        RECT 2456.695 2064.655 2457.025 2064.985 ;
        RECT 2450.270 2056.235 2450.570 2064.655 ;
        RECT 2456.710 2058.850 2457.010 2064.655 ;
        RECT 2459.455 2063.295 2459.785 2063.625 ;
        RECT 2465.895 2063.295 2466.225 2063.625 ;
        RECT 2472.335 2063.295 2472.665 2063.625 ;
        RECT 2478.775 2063.295 2479.105 2063.625 ;
        RECT 2484.295 2063.295 2484.625 2063.625 ;
        RECT 2491.655 2063.295 2491.985 2063.625 ;
        RECT 2498.095 2063.295 2498.425 2063.625 ;
        RECT 2505.455 2063.295 2505.785 2063.625 ;
        RECT 2513.735 2063.295 2514.065 2063.625 ;
        RECT 2518.335 2063.295 2518.665 2063.625 ;
        RECT 2522.015 2063.295 2522.345 2063.625 ;
        RECT 2443.865 2055.450 2444.165 2056.235 ;
        RECT 2442.910 2055.150 2444.165 2055.450 ;
        RECT 2387.705 2051.635 2388.005 2055.150 ;
        RECT 2393.945 2051.635 2394.245 2055.150 ;
        RECT 2400.185 2051.635 2400.485 2055.150 ;
        RECT 2406.425 2051.635 2406.725 2055.150 ;
        RECT 2412.665 2051.635 2412.965 2055.150 ;
        RECT 2418.905 2051.635 2419.205 2055.150 ;
        RECT 2425.145 2051.635 2425.445 2055.150 ;
        RECT 2431.385 2051.635 2431.685 2055.150 ;
        RECT 2437.625 2051.635 2437.925 2055.150 ;
        RECT 2443.865 2051.635 2444.165 2055.150 ;
        RECT 2450.105 2055.150 2450.570 2056.235 ;
        RECT 2456.345 2058.550 2457.010 2058.850 ;
        RECT 2450.105 2051.635 2450.405 2055.150 ;
        RECT 2456.345 2051.635 2456.645 2058.550 ;
        RECT 2459.470 2055.450 2459.770 2063.295 ;
        RECT 2462.585 2055.450 2462.885 2056.235 ;
        RECT 2459.470 2055.150 2462.885 2055.450 ;
        RECT 2465.910 2055.450 2466.210 2063.295 ;
        RECT 2468.825 2055.450 2469.125 2056.235 ;
        RECT 2465.910 2055.150 2469.125 2055.450 ;
        RECT 2472.350 2055.450 2472.650 2063.295 ;
        RECT 2475.065 2055.450 2475.365 2056.235 ;
        RECT 2472.350 2055.150 2475.365 2055.450 ;
        RECT 2478.790 2055.450 2479.090 2063.295 ;
        RECT 2481.305 2055.450 2481.605 2056.235 ;
        RECT 2478.790 2055.150 2481.605 2055.450 ;
        RECT 2484.310 2055.450 2484.610 2063.295 ;
        RECT 2487.545 2055.450 2487.845 2056.235 ;
        RECT 2484.310 2055.150 2487.845 2055.450 ;
        RECT 2491.670 2055.450 2491.970 2063.295 ;
        RECT 2493.785 2055.450 2494.085 2056.235 ;
        RECT 2491.670 2055.150 2494.085 2055.450 ;
        RECT 2498.110 2055.450 2498.410 2063.295 ;
        RECT 2500.025 2055.450 2500.325 2056.235 ;
        RECT 2498.110 2055.150 2500.325 2055.450 ;
        RECT 2505.470 2055.450 2505.770 2063.295 ;
        RECT 2506.265 2055.450 2506.565 2056.235 ;
        RECT 2505.470 2055.150 2506.565 2055.450 ;
        RECT 2462.585 2051.635 2462.885 2055.150 ;
        RECT 2468.825 2051.635 2469.125 2055.150 ;
        RECT 2475.065 2051.635 2475.365 2055.150 ;
        RECT 2481.305 2051.635 2481.605 2055.150 ;
        RECT 2487.545 2051.635 2487.845 2055.150 ;
        RECT 2493.785 2051.635 2494.085 2055.150 ;
        RECT 2500.025 2051.635 2500.325 2055.150 ;
        RECT 2506.265 2051.635 2506.565 2055.150 ;
        RECT 2512.505 2053.750 2512.805 2056.235 ;
        RECT 2513.750 2053.750 2514.050 2063.295 ;
        RECT 2518.350 2058.850 2518.650 2063.295 ;
        RECT 2518.350 2058.550 2519.045 2058.850 ;
        RECT 2512.505 2053.450 2514.050 2053.750 ;
        RECT 2512.505 2051.635 2512.805 2053.450 ;
        RECT 2518.745 2051.635 2519.045 2058.550 ;
        RECT 2522.030 2055.450 2522.330 2063.295 ;
        RECT 2524.985 2055.450 2525.285 2056.235 ;
        RECT 2522.030 2055.150 2525.285 2055.450 ;
        RECT 2528.470 2055.450 2528.770 2068.735 ;
        RECT 2534.895 2068.055 2535.225 2068.385 ;
        RECT 2531.225 2055.450 2531.525 2056.235 ;
        RECT 2528.470 2055.150 2531.525 2055.450 ;
        RECT 2534.910 2055.450 2535.210 2068.055 ;
        RECT 2590.095 2063.295 2590.425 2063.625 ;
        RECT 2537.465 2055.450 2537.765 2056.235 ;
        RECT 2534.910 2055.150 2537.765 2055.450 ;
        RECT 2590.110 2055.450 2590.410 2063.295 ;
        RECT 2592.890 2055.450 2593.190 2056.235 ;
        RECT 2590.110 2055.150 2593.190 2055.450 ;
        RECT 2524.985 2051.635 2525.285 2055.150 ;
        RECT 2531.225 2051.635 2531.525 2055.150 ;
        RECT 2537.465 2051.635 2537.765 2055.150 ;
        RECT 2592.890 2051.635 2593.190 2055.150 ;
        RECT 1417.095 1621.975 1417.425 1622.305 ;
        RECT 1411.575 1617.215 1411.905 1617.545 ;
      LAYER met4 ;
        RECT 323.295 1606.975 1389.905 1610.240 ;
        RECT 1705.000 1605.000 2081.480 2051.235 ;
      LAYER met4 ;
        RECT 2102.990 1745.310 2104.170 1746.490 ;
        RECT 2099.735 1732.890 2100.065 1733.145 ;
        RECT 2099.310 1731.710 2100.490 1732.890 ;
        RECT 2102.990 1731.710 2104.170 1732.890 ;
        RECT 2114.030 1731.710 2115.210 1732.890 ;
        RECT 2138.870 1731.710 2140.050 1732.890 ;
        RECT 2233.630 1731.710 2234.810 1732.890 ;
        RECT 2238.230 1731.710 2239.410 1732.890 ;
        RECT 2189.470 1728.310 2190.650 1729.490 ;
        RECT 2235.470 1728.310 2236.650 1729.490 ;
        RECT 2188.550 1724.910 2189.730 1726.090 ;
        RECT 2188.990 1722.265 2189.290 1724.910 ;
        RECT 2188.975 1721.935 2189.305 1722.265 ;
        RECT 2103.415 1718.535 2103.745 1718.865 ;
        RECT 2103.430 1715.890 2103.730 1718.535 ;
        RECT 2102.990 1714.710 2104.170 1715.890 ;
        RECT 2187.630 1714.710 2188.810 1715.890 ;
        RECT 2240.070 1714.710 2241.250 1715.890 ;
        RECT 2247.430 1714.710 2248.610 1715.890 ;
        RECT 2253.375 1715.135 2253.705 1715.465 ;
        RECT 2227.190 1711.310 2228.370 1712.490 ;
        RECT 2102.070 1707.910 2103.250 1709.090 ;
        RECT 2221.670 1708.650 2222.850 1709.090 ;
        RECT 2225.350 1708.650 2226.530 1709.090 ;
        RECT 2221.670 1708.350 2226.530 1708.650 ;
        RECT 2221.670 1707.910 2222.850 1708.350 ;
        RECT 2225.350 1707.910 2226.530 1708.350 ;
        RECT 2139.295 1705.690 2139.625 1705.945 ;
        RECT 2102.070 1704.510 2103.250 1705.690 ;
        RECT 2138.870 1704.510 2140.050 1705.690 ;
        RECT 2197.255 1705.615 2197.585 1705.945 ;
        RECT 2197.270 1698.890 2197.570 1705.615 ;
        RECT 2221.670 1701.110 2222.850 1702.290 ;
        RECT 2227.630 1701.865 2227.930 1711.310 ;
        RECT 2227.615 1701.535 2227.945 1701.865 ;
        RECT 2196.830 1697.710 2198.010 1698.890 ;
        RECT 2253.390 1692.090 2253.690 1715.135 ;
        RECT 2252.950 1690.910 2254.130 1692.090 ;
      LAYER met4 ;
        RECT 2255.000 1605.000 2631.480 2051.235 ;
      LAYER met4 ;
        RECT 2637.510 1745.310 2638.690 1746.490 ;
        RECT 2639.775 1735.535 2640.105 1735.865 ;
        RECT 2639.790 1732.890 2640.090 1735.535 ;
        RECT 2637.935 1732.135 2638.265 1732.465 ;
        RECT 2637.950 1729.490 2638.250 1732.135 ;
        RECT 2639.350 1731.710 2640.530 1732.890 ;
        RECT 2637.510 1728.310 2638.690 1729.490 ;
        RECT 2637.510 1724.910 2638.690 1726.090 ;
        RECT 2637.950 1724.585 2638.250 1724.910 ;
        RECT 2637.935 1724.255 2638.265 1724.585 ;
        RECT 2637.510 1714.710 2638.690 1715.890 ;
        RECT 2639.775 1715.815 2640.105 1716.145 ;
        RECT 2637.950 1710.025 2638.250 1714.710 ;
        RECT 2637.935 1709.695 2638.265 1710.025 ;
        RECT 2637.510 1707.910 2638.690 1709.090 ;
        RECT 2639.790 1702.290 2640.090 1715.815 ;
        RECT 2639.350 1701.110 2640.530 1702.290 ;
        RECT 1743.290 1600.000 1743.590 1604.600 ;
        RECT 1798.715 1600.000 1799.015 1604.600 ;
        RECT 1804.955 1600.000 1805.255 1604.600 ;
        RECT 1811.195 1600.000 1811.495 1604.600 ;
        RECT 1817.435 1600.000 1817.735 1604.600 ;
        RECT 1823.675 1600.000 1823.975 1604.600 ;
        RECT 1829.915 1600.000 1830.215 1604.600 ;
        RECT 1836.155 1600.000 1836.455 1604.600 ;
        RECT 1842.395 1600.000 1842.695 1604.600 ;
        RECT 1848.635 1600.000 1848.935 1604.600 ;
        RECT 1854.875 1600.000 1855.175 1604.600 ;
        RECT 1861.115 1600.000 1861.415 1604.600 ;
        RECT 1867.355 1600.000 1867.655 1604.600 ;
        RECT 1873.595 1600.000 1873.895 1604.600 ;
        RECT 1879.835 1600.000 1880.135 1604.600 ;
        RECT 1886.075 1600.000 1886.375 1604.600 ;
        RECT 1892.315 1600.000 1892.615 1604.600 ;
        RECT 1898.555 1600.000 1898.855 1604.600 ;
        RECT 1904.795 1600.000 1905.095 1604.600 ;
        RECT 1911.035 1600.000 1911.335 1604.600 ;
        RECT 1917.275 1600.000 1917.575 1604.600 ;
        RECT 1923.515 1600.000 1923.815 1604.600 ;
        RECT 1929.755 1600.000 1930.055 1604.600 ;
        RECT 1935.995 1600.000 1936.295 1604.600 ;
        RECT 1942.235 1600.000 1942.535 1604.600 ;
        RECT 1948.475 1600.000 1948.775 1604.600 ;
        RECT 1954.715 1600.000 1955.015 1604.600 ;
        RECT 1960.955 1600.000 1961.255 1604.600 ;
        RECT 1967.195 1600.000 1967.495 1604.600 ;
        RECT 1973.435 1600.000 1973.735 1604.600 ;
        RECT 1979.675 1600.000 1979.975 1604.600 ;
        RECT 1985.915 1600.000 1986.215 1604.600 ;
        RECT 1992.155 1600.000 1992.455 1604.600 ;
        RECT 2284.010 1600.000 2284.310 1604.600 ;
        RECT 2289.850 1600.000 2290.150 1604.600 ;
        RECT 2295.690 1600.000 2295.990 1604.600 ;
        RECT 2301.530 1600.000 2301.830 1604.600 ;
        RECT 2307.370 1600.000 2307.670 1604.600 ;
        RECT 2313.210 1600.000 2313.510 1604.600 ;
        RECT 2313.830 1600.000 2314.130 1604.600 ;
        RECT 2319.050 1600.000 2319.350 1604.600 ;
        RECT 2319.670 1600.000 2319.970 1604.600 ;
        RECT 2324.890 1600.000 2325.190 1604.600 ;
        RECT 2325.510 1600.000 2325.810 1604.600 ;
        RECT 2330.730 1600.000 2331.030 1604.600 ;
        RECT 2331.350 1600.000 2331.650 1604.600 ;
        RECT 2336.570 1600.000 2336.870 1604.600 ;
        RECT 2337.190 1600.000 2337.490 1604.600 ;
        RECT 2342.410 1600.000 2342.710 1604.600 ;
        RECT 2343.030 1600.000 2343.330 1604.600 ;
        RECT 2348.250 1600.000 2348.550 1604.600 ;
        RECT 2348.870 1600.000 2349.170 1604.600 ;
        RECT 2354.090 1600.000 2354.390 1604.600 ;
        RECT 2354.710 1600.000 2355.010 1604.600 ;
        RECT 2359.930 1600.000 2360.230 1604.600 ;
        RECT 2360.550 1600.000 2360.850 1604.600 ;
        RECT 2365.770 1600.000 2366.070 1604.600 ;
        RECT 2366.390 1600.000 2366.690 1604.600 ;
        RECT 2371.610 1600.000 2371.910 1604.600 ;
        RECT 2372.230 1600.000 2372.530 1604.600 ;
        RECT 2377.450 1600.000 2377.750 1604.600 ;
        RECT 2378.070 1600.000 2378.370 1604.600 ;
        RECT 2383.290 1600.000 2383.590 1604.600 ;
        RECT 2383.910 1600.000 2384.210 1604.600 ;
        RECT 2389.130 1600.000 2389.430 1604.600 ;
        RECT 2389.750 1600.000 2390.050 1604.600 ;
        RECT 2394.970 1600.000 2395.270 1604.600 ;
        RECT 2395.590 1600.000 2395.890 1604.600 ;
        RECT 2400.810 1600.000 2401.110 1604.600 ;
        RECT 2401.430 1600.000 2401.730 1604.600 ;
        RECT 2406.650 1600.000 2406.950 1604.600 ;
        RECT 2407.270 1600.000 2407.570 1604.600 ;
        RECT 2412.490 1600.000 2412.790 1604.600 ;
        RECT 2413.110 1600.000 2413.410 1604.600 ;
        RECT 2418.330 1600.000 2418.630 1604.600 ;
        RECT 2418.950 1600.000 2419.250 1604.600 ;
        RECT 2424.170 1600.000 2424.470 1604.600 ;
        RECT 2424.790 1600.000 2425.090 1604.600 ;
        RECT 2430.010 1600.000 2430.310 1604.600 ;
        RECT 2430.630 1600.000 2430.930 1604.600 ;
        RECT 2435.850 1600.000 2436.150 1604.600 ;
        RECT 2436.470 1600.000 2436.770 1604.600 ;
        RECT 2441.690 1600.000 2441.990 1604.600 ;
        RECT 2442.310 1600.000 2442.610 1604.600 ;
        RECT 2447.530 1600.000 2447.830 1604.600 ;
        RECT 2448.150 1600.000 2448.450 1604.600 ;
        RECT 2453.370 1600.000 2453.670 1604.600 ;
        RECT 2453.990 1600.000 2454.290 1604.600 ;
        RECT 2459.210 1600.000 2459.510 1604.600 ;
        RECT 2459.830 1600.000 2460.130 1604.600 ;
        RECT 2465.050 1600.000 2465.350 1604.600 ;
        RECT 2465.670 1600.000 2465.970 1604.600 ;
        RECT 2470.890 1600.000 2471.190 1604.600 ;
        RECT 2471.510 1600.000 2471.810 1604.600 ;
        RECT 2476.730 1600.000 2477.030 1604.600 ;
        RECT 2477.350 1600.000 2477.650 1604.600 ;
        RECT 2482.570 1600.000 2482.870 1604.600 ;
        RECT 2483.190 1600.000 2483.490 1604.600 ;
        RECT 2488.410 1600.000 2488.710 1604.600 ;
        RECT 2489.030 1600.000 2489.330 1604.600 ;
        RECT 2494.250 1600.000 2494.550 1604.600 ;
        RECT 2494.870 1600.000 2495.170 1604.600 ;
        RECT 1768.020 1515.000 1771.020 1585.000 ;
        RECT 1804.020 1515.000 1807.020 1585.000 ;
        RECT 1822.020 1515.000 1825.020 1585.000 ;
        RECT 1840.020 1515.000 1843.020 1585.000 ;
        RECT 1858.020 1515.000 1861.020 1585.000 ;
        RECT 1948.020 1515.000 1951.020 1585.000 ;
        RECT 1984.020 1515.000 1987.020 1585.000 ;
        RECT 2002.020 1515.000 2005.020 1585.000 ;
        RECT 2020.020 1515.000 2023.020 1585.000 ;
        RECT 2038.020 1515.000 2041.020 1585.000 ;
        RECT 2308.020 1515.000 2311.020 1585.000 ;
        RECT 2344.020 1515.000 2347.020 1585.000 ;
        RECT 2362.020 1515.000 2365.020 1585.000 ;
        RECT 2380.020 1515.000 2383.020 1585.000 ;
        RECT 2398.020 1515.000 2401.020 1585.000 ;
        RECT 2488.020 1515.000 2491.020 1585.000 ;
        RECT 2524.020 1515.000 2527.020 1585.000 ;
        RECT 2542.020 1515.000 2545.020 1585.000 ;
        RECT 2560.020 1515.000 2563.020 1585.000 ;
        RECT 2578.020 1515.000 2581.020 1585.000 ;
      LAYER met4 ;
        RECT 1573.295 1488.640 2639.905 1497.345 ;
        RECT 1573.295 410.240 1647.440 1488.640 ;
        RECT 1649.840 410.240 2639.905 1488.640 ;
        RECT 1573.295 406.975 2639.905 410.240 ;
      LAYER met5 ;
        RECT 1351.140 2935.100 1938.780 2936.700 ;
        RECT 1945.460 2897.700 2595.660 2899.300 ;
        RECT 302.340 2894.300 2188.100 2895.900 ;
        RECT 2102.780 1745.100 2638.900 1746.700 ;
        RECT 2099.100 1729.700 2100.700 1733.100 ;
        RECT 2102.780 1731.500 2115.420 1733.100 ;
        RECT 2138.660 1731.500 2235.020 1733.100 ;
        RECT 2238.020 1731.500 2640.740 1733.100 ;
        RECT 2099.100 1728.100 2190.860 1729.700 ;
        RECT 2235.260 1728.100 2638.900 1729.700 ;
        RECT 2188.340 1724.700 2638.900 1726.300 ;
        RECT 2102.780 1714.500 2189.020 1716.100 ;
        RECT 2239.860 1714.500 2248.820 1716.100 ;
        RECT 2267.460 1714.500 2349.100 1716.100 ;
        RECT 2267.460 1712.700 2269.060 1714.500 ;
        RECT 2226.980 1711.100 2269.060 1712.700 ;
        RECT 2347.500 1712.700 2349.100 1714.500 ;
        RECT 2394.420 1714.500 2430.060 1716.100 ;
        RECT 2394.420 1712.700 2396.020 1714.500 ;
        RECT 2347.500 1711.100 2356.460 1712.700 ;
        RECT 2354.860 1709.300 2356.460 1711.100 ;
        RECT 2359.460 1711.100 2396.020 1712.700 ;
        RECT 2428.460 1712.700 2430.060 1714.500 ;
        RECT 2443.180 1714.500 2512.860 1716.100 ;
        RECT 2443.180 1712.700 2444.780 1714.500 ;
        RECT 2511.260 1712.700 2512.860 1714.500 ;
        RECT 2606.940 1714.500 2638.900 1716.100 ;
        RECT 2428.460 1711.100 2444.780 1712.700 ;
        RECT 2475.380 1711.100 2490.780 1712.700 ;
        RECT 2511.260 1711.100 2577.260 1712.700 ;
        RECT 2359.460 1709.300 2361.060 1711.100 ;
        RECT 2101.860 1707.700 2223.060 1709.300 ;
        RECT 2225.140 1707.700 2250.660 1709.300 ;
        RECT 2249.060 1705.900 2250.660 1707.700 ;
        RECT 2301.500 1707.700 2352.780 1709.300 ;
        RECT 2354.860 1707.700 2361.060 1709.300 ;
        RECT 2363.140 1707.700 2388.660 1709.300 ;
        RECT 2301.500 1705.900 2303.100 1707.700 ;
        RECT 2101.860 1704.300 2140.260 1705.900 ;
        RECT 2220.540 1700.900 2223.060 1705.900 ;
        RECT 2249.060 1704.300 2297.580 1705.900 ;
        RECT 2295.980 1702.500 2297.580 1704.300 ;
        RECT 2300.580 1704.300 2303.100 1705.900 ;
        RECT 2351.180 1705.900 2352.780 1707.700 ;
        RECT 2363.140 1705.900 2364.740 1707.700 ;
        RECT 2351.180 1704.300 2364.740 1705.900 ;
        RECT 2300.580 1702.500 2302.180 1704.300 ;
        RECT 2387.060 1702.500 2388.660 1707.700 ;
        RECT 2475.380 1705.900 2476.980 1711.100 ;
        RECT 2489.180 1709.300 2490.780 1711.100 ;
        RECT 2575.660 1709.300 2577.260 1711.100 ;
        RECT 2606.940 1709.300 2608.540 1714.500 ;
        RECT 2489.180 1707.700 2540.460 1709.300 ;
        RECT 2575.660 1707.700 2608.540 1709.300 ;
        RECT 2610.620 1707.700 2638.900 1709.300 ;
        RECT 2431.220 1704.300 2476.980 1705.900 ;
        RECT 2431.220 1702.500 2432.820 1704.300 ;
        RECT 2295.980 1700.900 2302.180 1702.500 ;
        RECT 2339.220 1700.900 2349.100 1702.500 ;
        RECT 2387.060 1700.900 2432.820 1702.500 ;
        RECT 2538.860 1702.500 2540.460 1707.700 ;
        RECT 2610.620 1705.900 2612.220 1707.700 ;
        RECT 2609.700 1704.300 2612.220 1705.900 ;
        RECT 2538.860 1700.900 2574.500 1702.500 ;
        RECT 2220.540 1699.100 2222.140 1700.900 ;
        RECT 2196.620 1697.500 2222.140 1699.100 ;
        RECT 2295.980 1694.100 2298.500 1700.900 ;
        RECT 2339.220 1699.100 2340.820 1700.900 ;
        RECT 2320.820 1697.500 2340.820 1699.100 ;
        RECT 2320.820 1692.300 2322.420 1697.500 ;
        RECT 2347.500 1695.700 2349.100 1700.900 ;
        RECT 2572.900 1699.100 2574.500 1700.900 ;
        RECT 2609.700 1699.100 2611.300 1704.300 ;
        RECT 2434.900 1697.500 2487.100 1699.100 ;
        RECT 2434.900 1695.700 2436.500 1697.500 ;
        RECT 2347.500 1694.100 2350.020 1695.700 ;
        RECT 2252.740 1690.700 2322.420 1692.300 ;
        RECT 2348.420 1692.300 2350.020 1694.100 ;
        RECT 2390.740 1694.100 2436.500 1695.700 ;
        RECT 2390.740 1692.300 2392.340 1694.100 ;
        RECT 2348.420 1690.700 2392.340 1692.300 ;
        RECT 2485.500 1692.300 2487.100 1697.500 ;
        RECT 2489.180 1697.500 2534.940 1699.100 ;
        RECT 2572.900 1697.500 2611.300 1699.100 ;
        RECT 2614.300 1700.900 2640.740 1702.500 ;
        RECT 2489.180 1692.300 2490.780 1697.500 ;
        RECT 2533.340 1695.700 2534.940 1697.500 ;
        RECT 2533.340 1694.100 2537.700 1695.700 ;
        RECT 2485.500 1690.700 2490.780 1692.300 ;
        RECT 2536.100 1692.300 2537.700 1694.100 ;
        RECT 2539.780 1694.100 2549.660 1695.700 ;
        RECT 2539.780 1692.300 2541.380 1694.100 ;
        RECT 2536.100 1690.700 2541.380 1692.300 ;
        RECT 2548.060 1692.300 2549.660 1694.100 ;
        RECT 2614.300 1692.300 2615.900 1700.900 ;
        RECT 2548.060 1690.700 2615.900 1692.300 ;
  END
END user_project_wrapper
END LIBRARY

