magic
tech sky130A
magscale 1 2
timestamp 1608587418
<< obsli1 >>
rect 1104 2159 218868 237745
<< obsm1 >>
rect 1026 892 218946 237856
<< metal2 >>
rect 1030 239200 1086 240000
rect 3054 239200 3110 240000
rect 5170 239200 5226 240000
rect 7194 239200 7250 240000
rect 9310 239200 9366 240000
rect 11334 239200 11390 240000
rect 13450 239200 13506 240000
rect 15474 239200 15530 240000
rect 17590 239200 17646 240000
rect 19706 239200 19762 240000
rect 21730 239200 21786 240000
rect 23846 239200 23902 240000
rect 25870 239200 25926 240000
rect 27986 239200 28042 240000
rect 30010 239200 30066 240000
rect 32126 239200 32182 240000
rect 34150 239200 34206 240000
rect 36266 239200 36322 240000
rect 38382 239200 38438 240000
rect 40406 239200 40462 240000
rect 42522 239200 42578 240000
rect 44546 239200 44602 240000
rect 46662 239200 46718 240000
rect 48686 239200 48742 240000
rect 50802 239200 50858 240000
rect 52826 239200 52882 240000
rect 54942 239200 54998 240000
rect 57058 239200 57114 240000
rect 59082 239200 59138 240000
rect 61198 239200 61254 240000
rect 63222 239200 63278 240000
rect 65338 239200 65394 240000
rect 67362 239200 67418 240000
rect 69478 239200 69534 240000
rect 71502 239200 71558 240000
rect 73618 239200 73674 240000
rect 75734 239200 75790 240000
rect 77758 239200 77814 240000
rect 79874 239200 79930 240000
rect 81898 239200 81954 240000
rect 84014 239200 84070 240000
rect 86038 239200 86094 240000
rect 88154 239200 88210 240000
rect 90178 239200 90234 240000
rect 92294 239200 92350 240000
rect 94410 239200 94466 240000
rect 96434 239200 96490 240000
rect 98550 239200 98606 240000
rect 100574 239200 100630 240000
rect 102690 239200 102746 240000
rect 104714 239200 104770 240000
rect 106830 239200 106886 240000
rect 108854 239200 108910 240000
rect 110970 239200 111026 240000
rect 113086 239200 113142 240000
rect 115110 239200 115166 240000
rect 117226 239200 117282 240000
rect 119250 239200 119306 240000
rect 121366 239200 121422 240000
rect 123390 239200 123446 240000
rect 125506 239200 125562 240000
rect 127530 239200 127586 240000
rect 129646 239200 129702 240000
rect 131762 239200 131818 240000
rect 133786 239200 133842 240000
rect 135902 239200 135958 240000
rect 137926 239200 137982 240000
rect 140042 239200 140098 240000
rect 142066 239200 142122 240000
rect 144182 239200 144238 240000
rect 146206 239200 146262 240000
rect 148322 239200 148378 240000
rect 150438 239200 150494 240000
rect 152462 239200 152518 240000
rect 154578 239200 154634 240000
rect 156602 239200 156658 240000
rect 158718 239200 158774 240000
rect 160742 239200 160798 240000
rect 162858 239200 162914 240000
rect 164882 239200 164938 240000
rect 166998 239200 167054 240000
rect 169114 239200 169170 240000
rect 171138 239200 171194 240000
rect 173254 239200 173310 240000
rect 175278 239200 175334 240000
rect 177394 239200 177450 240000
rect 179418 239200 179474 240000
rect 181534 239200 181590 240000
rect 183558 239200 183614 240000
rect 185674 239200 185730 240000
rect 187790 239200 187846 240000
rect 189814 239200 189870 240000
rect 191930 239200 191986 240000
rect 193954 239200 194010 240000
rect 196070 239200 196126 240000
rect 198094 239200 198150 240000
rect 200210 239200 200266 240000
rect 202234 239200 202290 240000
rect 204350 239200 204406 240000
rect 206466 239200 206522 240000
rect 208490 239200 208546 240000
rect 210606 239200 210662 240000
rect 212630 239200 212686 240000
rect 214746 239200 214802 240000
rect 216770 239200 216826 240000
rect 218886 239200 218942 240000
rect 938 0 994 800
rect 2870 0 2926 800
rect 4802 0 4858 800
rect 6734 0 6790 800
rect 8666 0 8722 800
rect 10598 0 10654 800
rect 12530 0 12586 800
rect 14554 0 14610 800
rect 16486 0 16542 800
rect 18418 0 18474 800
rect 20350 0 20406 800
rect 22282 0 22338 800
rect 24214 0 24270 800
rect 26238 0 26294 800
rect 28170 0 28226 800
rect 30102 0 30158 800
rect 32034 0 32090 800
rect 33966 0 34022 800
rect 35898 0 35954 800
rect 37922 0 37978 800
rect 39854 0 39910 800
rect 41786 0 41842 800
rect 43718 0 43774 800
rect 45650 0 45706 800
rect 47582 0 47638 800
rect 49514 0 49570 800
rect 51538 0 51594 800
rect 53470 0 53526 800
rect 55402 0 55458 800
rect 57334 0 57390 800
rect 59266 0 59322 800
rect 61198 0 61254 800
rect 63222 0 63278 800
rect 65154 0 65210 800
rect 67086 0 67142 800
rect 69018 0 69074 800
rect 70950 0 71006 800
rect 72882 0 72938 800
rect 74906 0 74962 800
rect 76838 0 76894 800
rect 78770 0 78826 800
rect 80702 0 80758 800
rect 82634 0 82690 800
rect 84566 0 84622 800
rect 86590 0 86646 800
rect 88522 0 88578 800
rect 90454 0 90510 800
rect 92386 0 92442 800
rect 94318 0 94374 800
rect 96250 0 96306 800
rect 98182 0 98238 800
rect 100206 0 100262 800
rect 102138 0 102194 800
rect 104070 0 104126 800
rect 106002 0 106058 800
rect 107934 0 107990 800
rect 109866 0 109922 800
rect 111890 0 111946 800
rect 113822 0 113878 800
rect 115754 0 115810 800
rect 117686 0 117742 800
rect 119618 0 119674 800
rect 121550 0 121606 800
rect 123574 0 123630 800
rect 125506 0 125562 800
rect 127438 0 127494 800
rect 129370 0 129426 800
rect 131302 0 131358 800
rect 133234 0 133290 800
rect 135166 0 135222 800
rect 137190 0 137246 800
rect 139122 0 139178 800
rect 141054 0 141110 800
rect 142986 0 143042 800
rect 144918 0 144974 800
rect 146850 0 146906 800
rect 148874 0 148930 800
rect 150806 0 150862 800
rect 152738 0 152794 800
rect 154670 0 154726 800
rect 156602 0 156658 800
rect 158534 0 158590 800
rect 160558 0 160614 800
rect 162490 0 162546 800
rect 164422 0 164478 800
rect 166354 0 166410 800
rect 168286 0 168342 800
rect 170218 0 170274 800
rect 172242 0 172298 800
rect 174174 0 174230 800
rect 176106 0 176162 800
rect 178038 0 178094 800
rect 179970 0 180026 800
rect 181902 0 181958 800
rect 183834 0 183890 800
rect 185858 0 185914 800
rect 187790 0 187846 800
rect 189722 0 189778 800
rect 191654 0 191710 800
rect 193586 0 193642 800
rect 195518 0 195574 800
rect 197542 0 197598 800
rect 199474 0 199530 800
rect 201406 0 201462 800
rect 203338 0 203394 800
rect 205270 0 205326 800
rect 207202 0 207258 800
rect 209226 0 209282 800
rect 211158 0 211214 800
rect 213090 0 213146 800
rect 215022 0 215078 800
rect 216954 0 217010 800
rect 218886 0 218942 800
<< obsm2 >>
rect 952 239144 974 239200
rect 1142 239144 2998 239200
rect 3166 239144 5114 239200
rect 5282 239144 7138 239200
rect 7306 239144 9254 239200
rect 9422 239144 11278 239200
rect 11446 239144 13394 239200
rect 13562 239144 15418 239200
rect 15586 239144 17534 239200
rect 17702 239144 19650 239200
rect 19818 239144 21674 239200
rect 21842 239144 23790 239200
rect 23958 239144 25814 239200
rect 25982 239144 27930 239200
rect 28098 239144 29954 239200
rect 30122 239144 32070 239200
rect 32238 239144 34094 239200
rect 34262 239144 36210 239200
rect 36378 239144 38326 239200
rect 38494 239144 40350 239200
rect 40518 239144 42466 239200
rect 42634 239144 44490 239200
rect 44658 239144 46606 239200
rect 46774 239144 48630 239200
rect 48798 239144 50746 239200
rect 50914 239144 52770 239200
rect 52938 239144 54886 239200
rect 55054 239144 57002 239200
rect 57170 239144 59026 239200
rect 59194 239144 61142 239200
rect 61310 239144 63166 239200
rect 63334 239144 65282 239200
rect 65450 239144 67306 239200
rect 67474 239144 69422 239200
rect 69590 239144 71446 239200
rect 71614 239144 73562 239200
rect 73730 239144 75678 239200
rect 75846 239144 77702 239200
rect 77870 239144 79818 239200
rect 79986 239144 81842 239200
rect 82010 239144 83958 239200
rect 84126 239144 85982 239200
rect 86150 239144 88098 239200
rect 88266 239144 90122 239200
rect 90290 239144 92238 239200
rect 92406 239144 94354 239200
rect 94522 239144 96378 239200
rect 96546 239144 98494 239200
rect 98662 239144 100518 239200
rect 100686 239144 102634 239200
rect 102802 239144 104658 239200
rect 104826 239144 106774 239200
rect 106942 239144 108798 239200
rect 108966 239144 110914 239200
rect 111082 239144 113030 239200
rect 113198 239144 115054 239200
rect 115222 239144 117170 239200
rect 117338 239144 119194 239200
rect 119362 239144 121310 239200
rect 121478 239144 123334 239200
rect 123502 239144 125450 239200
rect 125618 239144 127474 239200
rect 127642 239144 129590 239200
rect 129758 239144 131706 239200
rect 131874 239144 133730 239200
rect 133898 239144 135846 239200
rect 136014 239144 137870 239200
rect 138038 239144 139986 239200
rect 140154 239144 142010 239200
rect 142178 239144 144126 239200
rect 144294 239144 146150 239200
rect 146318 239144 148266 239200
rect 148434 239144 150382 239200
rect 150550 239144 152406 239200
rect 152574 239144 154522 239200
rect 154690 239144 156546 239200
rect 156714 239144 158662 239200
rect 158830 239144 160686 239200
rect 160854 239144 162802 239200
rect 162970 239144 164826 239200
rect 164994 239144 166942 239200
rect 167110 239144 169058 239200
rect 169226 239144 171082 239200
rect 171250 239144 173198 239200
rect 173366 239144 175222 239200
rect 175390 239144 177338 239200
rect 177506 239144 179362 239200
rect 179530 239144 181478 239200
rect 181646 239144 183502 239200
rect 183670 239144 185618 239200
rect 185786 239144 187734 239200
rect 187902 239144 189758 239200
rect 189926 239144 191874 239200
rect 192042 239144 193898 239200
rect 194066 239144 196014 239200
rect 196182 239144 198038 239200
rect 198206 239144 200154 239200
rect 200322 239144 202178 239200
rect 202346 239144 204294 239200
rect 204462 239144 206410 239200
rect 206578 239144 208434 239200
rect 208602 239144 210550 239200
rect 210718 239144 212574 239200
rect 212742 239144 214690 239200
rect 214858 239144 216714 239200
rect 216882 239144 218830 239200
rect 218998 239144 219126 239200
rect 952 856 219126 239144
rect 1050 800 2814 856
rect 2982 800 4746 856
rect 4914 800 6678 856
rect 6846 800 8610 856
rect 8778 800 10542 856
rect 10710 800 12474 856
rect 12642 800 14498 856
rect 14666 800 16430 856
rect 16598 800 18362 856
rect 18530 800 20294 856
rect 20462 800 22226 856
rect 22394 800 24158 856
rect 24326 800 26182 856
rect 26350 800 28114 856
rect 28282 800 30046 856
rect 30214 800 31978 856
rect 32146 800 33910 856
rect 34078 800 35842 856
rect 36010 800 37866 856
rect 38034 800 39798 856
rect 39966 800 41730 856
rect 41898 800 43662 856
rect 43830 800 45594 856
rect 45762 800 47526 856
rect 47694 800 49458 856
rect 49626 800 51482 856
rect 51650 800 53414 856
rect 53582 800 55346 856
rect 55514 800 57278 856
rect 57446 800 59210 856
rect 59378 800 61142 856
rect 61310 800 63166 856
rect 63334 800 65098 856
rect 65266 800 67030 856
rect 67198 800 68962 856
rect 69130 800 70894 856
rect 71062 800 72826 856
rect 72994 800 74850 856
rect 75018 800 76782 856
rect 76950 800 78714 856
rect 78882 800 80646 856
rect 80814 800 82578 856
rect 82746 800 84510 856
rect 84678 800 86534 856
rect 86702 800 88466 856
rect 88634 800 90398 856
rect 90566 800 92330 856
rect 92498 800 94262 856
rect 94430 800 96194 856
rect 96362 800 98126 856
rect 98294 800 100150 856
rect 100318 800 102082 856
rect 102250 800 104014 856
rect 104182 800 105946 856
rect 106114 800 107878 856
rect 108046 800 109810 856
rect 109978 800 111834 856
rect 112002 800 113766 856
rect 113934 800 115698 856
rect 115866 800 117630 856
rect 117798 800 119562 856
rect 119730 800 121494 856
rect 121662 800 123518 856
rect 123686 800 125450 856
rect 125618 800 127382 856
rect 127550 800 129314 856
rect 129482 800 131246 856
rect 131414 800 133178 856
rect 133346 800 135110 856
rect 135278 800 137134 856
rect 137302 800 139066 856
rect 139234 800 140998 856
rect 141166 800 142930 856
rect 143098 800 144862 856
rect 145030 800 146794 856
rect 146962 800 148818 856
rect 148986 800 150750 856
rect 150918 800 152682 856
rect 152850 800 154614 856
rect 154782 800 156546 856
rect 156714 800 158478 856
rect 158646 800 160502 856
rect 160670 800 162434 856
rect 162602 800 164366 856
rect 164534 800 166298 856
rect 166466 800 168230 856
rect 168398 800 170162 856
rect 170330 800 172186 856
rect 172354 800 174118 856
rect 174286 800 176050 856
rect 176218 800 177982 856
rect 178150 800 179914 856
rect 180082 800 181846 856
rect 182014 800 183778 856
rect 183946 800 185802 856
rect 185970 800 187734 856
rect 187902 800 189666 856
rect 189834 800 191598 856
rect 191766 800 193530 856
rect 193698 800 195462 856
rect 195630 800 197486 856
rect 197654 800 199418 856
rect 199586 800 201350 856
rect 201518 800 203282 856
rect 203450 800 205214 856
rect 205382 800 207146 856
rect 207314 800 209170 856
rect 209338 800 211102 856
rect 211270 800 213034 856
rect 213202 800 214966 856
rect 215134 800 216898 856
rect 217066 800 218830 856
rect 218998 800 219126 856
<< metal3 >>
rect 0 238824 800 238944
rect 219200 238824 220000 238944
rect 0 236784 800 236904
rect 219200 236648 220000 236768
rect 0 234608 800 234728
rect 219200 234472 220000 234592
rect 0 232568 800 232688
rect 219200 232296 220000 232416
rect 0 230392 800 230512
rect 219200 230120 220000 230240
rect 0 228352 800 228472
rect 219200 227808 220000 227928
rect 0 226176 800 226296
rect 219200 225632 220000 225752
rect 0 224136 800 224256
rect 219200 223456 220000 223576
rect 0 221960 800 222080
rect 219200 221280 220000 221400
rect 0 219920 800 220040
rect 219200 219104 220000 219224
rect 0 217744 800 217864
rect 219200 216792 220000 216912
rect 0 215704 800 215824
rect 219200 214616 220000 214736
rect 0 213528 800 213648
rect 219200 212440 220000 212560
rect 0 211488 800 211608
rect 219200 210264 220000 210384
rect 0 209312 800 209432
rect 219200 208088 220000 208208
rect 0 207272 800 207392
rect 219200 205776 220000 205896
rect 0 205096 800 205216
rect 219200 203600 220000 203720
rect 0 203056 800 203176
rect 219200 201424 220000 201544
rect 0 200880 800 201000
rect 219200 199248 220000 199368
rect 0 198840 800 198960
rect 219200 197072 220000 197192
rect 0 196664 800 196784
rect 0 194624 800 194744
rect 219200 194760 220000 194880
rect 0 192448 800 192568
rect 219200 192584 220000 192704
rect 0 190408 800 190528
rect 219200 190408 220000 190528
rect 0 188232 800 188352
rect 219200 188232 220000 188352
rect 0 186192 800 186312
rect 219200 186056 220000 186176
rect 0 184016 800 184136
rect 219200 183744 220000 183864
rect 0 181976 800 182096
rect 219200 181568 220000 181688
rect 0 179936 800 180056
rect 219200 179392 220000 179512
rect 0 177760 800 177880
rect 219200 177216 220000 177336
rect 0 175720 800 175840
rect 219200 175040 220000 175160
rect 0 173544 800 173664
rect 219200 172864 220000 172984
rect 0 171504 800 171624
rect 219200 170552 220000 170672
rect 0 169328 800 169448
rect 219200 168376 220000 168496
rect 0 167288 800 167408
rect 219200 166200 220000 166320
rect 0 165112 800 165232
rect 219200 164024 220000 164144
rect 0 163072 800 163192
rect 219200 161848 220000 161968
rect 0 160896 800 161016
rect 219200 159536 220000 159656
rect 0 158856 800 158976
rect 219200 157360 220000 157480
rect 0 156680 800 156800
rect 219200 155184 220000 155304
rect 0 154640 800 154760
rect 219200 153008 220000 153128
rect 0 152464 800 152584
rect 219200 150832 220000 150952
rect 0 150424 800 150544
rect 219200 148520 220000 148640
rect 0 148248 800 148368
rect 0 146208 800 146328
rect 219200 146344 220000 146464
rect 0 144032 800 144152
rect 219200 144168 220000 144288
rect 0 141992 800 142112
rect 219200 141992 220000 142112
rect 0 139816 800 139936
rect 219200 139816 220000 139936
rect 0 137776 800 137896
rect 219200 137504 220000 137624
rect 0 135600 800 135720
rect 219200 135328 220000 135448
rect 0 133560 800 133680
rect 219200 133152 220000 133272
rect 0 131384 800 131504
rect 219200 130976 220000 131096
rect 0 129344 800 129464
rect 219200 128800 220000 128920
rect 0 127168 800 127288
rect 219200 126488 220000 126608
rect 0 125128 800 125248
rect 219200 124312 220000 124432
rect 0 122952 800 123072
rect 219200 122136 220000 122256
rect 0 120912 800 121032
rect 219200 119960 220000 120080
rect 0 118872 800 118992
rect 219200 117784 220000 117904
rect 0 116696 800 116816
rect 219200 115608 220000 115728
rect 0 114656 800 114776
rect 219200 113296 220000 113416
rect 0 112480 800 112600
rect 219200 111120 220000 111240
rect 0 110440 800 110560
rect 219200 108944 220000 109064
rect 0 108264 800 108384
rect 219200 106768 220000 106888
rect 0 106224 800 106344
rect 219200 104592 220000 104712
rect 0 104048 800 104168
rect 219200 102280 220000 102400
rect 0 102008 800 102128
rect 219200 100104 220000 100224
rect 0 99832 800 99952
rect 0 97792 800 97912
rect 219200 97928 220000 98048
rect 0 95616 800 95736
rect 219200 95752 220000 95872
rect 0 93576 800 93696
rect 219200 93576 220000 93696
rect 0 91400 800 91520
rect 219200 91264 220000 91384
rect 0 89360 800 89480
rect 219200 89088 220000 89208
rect 0 87184 800 87304
rect 219200 86912 220000 87032
rect 0 85144 800 85264
rect 219200 84736 220000 84856
rect 0 82968 800 83088
rect 219200 82560 220000 82680
rect 0 80928 800 81048
rect 219200 80248 220000 80368
rect 0 78752 800 78872
rect 219200 78072 220000 78192
rect 0 76712 800 76832
rect 219200 75896 220000 76016
rect 0 74536 800 74656
rect 219200 73720 220000 73840
rect 0 72496 800 72616
rect 219200 71544 220000 71664
rect 0 70320 800 70440
rect 219200 69232 220000 69352
rect 0 68280 800 68400
rect 219200 67056 220000 67176
rect 0 66104 800 66224
rect 219200 64880 220000 65000
rect 0 64064 800 64184
rect 219200 62704 220000 62824
rect 0 61888 800 62008
rect 219200 60528 220000 60648
rect 0 59848 800 59968
rect 219200 58352 220000 58472
rect 0 57808 800 57928
rect 219200 56040 220000 56160
rect 0 55632 800 55752
rect 219200 53864 220000 53984
rect 0 53592 800 53712
rect 219200 51688 220000 51808
rect 0 51416 800 51536
rect 0 49376 800 49496
rect 219200 49512 220000 49632
rect 0 47200 800 47320
rect 219200 47336 220000 47456
rect 0 45160 800 45280
rect 219200 45024 220000 45144
rect 0 42984 800 43104
rect 219200 42848 220000 42968
rect 0 40944 800 41064
rect 219200 40672 220000 40792
rect 0 38768 800 38888
rect 219200 38496 220000 38616
rect 0 36728 800 36848
rect 219200 36320 220000 36440
rect 0 34552 800 34672
rect 219200 34008 220000 34128
rect 0 32512 800 32632
rect 219200 31832 220000 31952
rect 0 30336 800 30456
rect 219200 29656 220000 29776
rect 0 28296 800 28416
rect 219200 27480 220000 27600
rect 0 26120 800 26240
rect 219200 25304 220000 25424
rect 0 24080 800 24200
rect 219200 22992 220000 23112
rect 0 21904 800 22024
rect 219200 20816 220000 20936
rect 0 19864 800 19984
rect 219200 18640 220000 18760
rect 0 17688 800 17808
rect 219200 16464 220000 16584
rect 0 15648 800 15768
rect 219200 14288 220000 14408
rect 0 13472 800 13592
rect 219200 11976 220000 12096
rect 0 11432 800 11552
rect 219200 9800 220000 9920
rect 0 9256 800 9376
rect 219200 7624 220000 7744
rect 0 7216 800 7336
rect 219200 5448 220000 5568
rect 0 5040 800 5160
rect 219200 3272 220000 3392
rect 0 3000 800 3120
rect 0 960 800 1080
rect 219200 1096 220000 1216
<< obsm3 >>
rect 880 238744 219120 238917
rect 798 236984 219200 238744
rect 880 236848 219200 236984
rect 880 236704 219120 236848
rect 798 236568 219120 236704
rect 798 234808 219200 236568
rect 880 234672 219200 234808
rect 880 234528 219120 234672
rect 798 234392 219120 234528
rect 798 232768 219200 234392
rect 880 232496 219200 232768
rect 880 232488 219120 232496
rect 798 232216 219120 232488
rect 798 230592 219200 232216
rect 880 230320 219200 230592
rect 880 230312 219120 230320
rect 798 230040 219120 230312
rect 798 228552 219200 230040
rect 880 228272 219200 228552
rect 798 228008 219200 228272
rect 798 227728 219120 228008
rect 798 226376 219200 227728
rect 880 226096 219200 226376
rect 798 225832 219200 226096
rect 798 225552 219120 225832
rect 798 224336 219200 225552
rect 880 224056 219200 224336
rect 798 223656 219200 224056
rect 798 223376 219120 223656
rect 798 222160 219200 223376
rect 880 221880 219200 222160
rect 798 221480 219200 221880
rect 798 221200 219120 221480
rect 798 220120 219200 221200
rect 880 219840 219200 220120
rect 798 219304 219200 219840
rect 798 219024 219120 219304
rect 798 217944 219200 219024
rect 880 217664 219200 217944
rect 798 216992 219200 217664
rect 798 216712 219120 216992
rect 798 215904 219200 216712
rect 880 215624 219200 215904
rect 798 214816 219200 215624
rect 798 214536 219120 214816
rect 798 213728 219200 214536
rect 880 213448 219200 213728
rect 798 212640 219200 213448
rect 798 212360 219120 212640
rect 798 211688 219200 212360
rect 880 211408 219200 211688
rect 798 210464 219200 211408
rect 798 210184 219120 210464
rect 798 209512 219200 210184
rect 880 209232 219200 209512
rect 798 208288 219200 209232
rect 798 208008 219120 208288
rect 798 207472 219200 208008
rect 880 207192 219200 207472
rect 798 205976 219200 207192
rect 798 205696 219120 205976
rect 798 205296 219200 205696
rect 880 205016 219200 205296
rect 798 203800 219200 205016
rect 798 203520 219120 203800
rect 798 203256 219200 203520
rect 880 202976 219200 203256
rect 798 201624 219200 202976
rect 798 201344 219120 201624
rect 798 201080 219200 201344
rect 880 200800 219200 201080
rect 798 199448 219200 200800
rect 798 199168 219120 199448
rect 798 199040 219200 199168
rect 880 198760 219200 199040
rect 798 197272 219200 198760
rect 798 196992 219120 197272
rect 798 196864 219200 196992
rect 880 196584 219200 196864
rect 798 194960 219200 196584
rect 798 194824 219120 194960
rect 880 194680 219120 194824
rect 880 194544 219200 194680
rect 798 192784 219200 194544
rect 798 192648 219120 192784
rect 880 192504 219120 192648
rect 880 192368 219200 192504
rect 798 190608 219200 192368
rect 880 190328 219120 190608
rect 798 188432 219200 190328
rect 880 188152 219120 188432
rect 798 186392 219200 188152
rect 880 186256 219200 186392
rect 880 186112 219120 186256
rect 798 185976 219120 186112
rect 798 184216 219200 185976
rect 880 183944 219200 184216
rect 880 183936 219120 183944
rect 798 183664 219120 183936
rect 798 182176 219200 183664
rect 880 181896 219200 182176
rect 798 181768 219200 181896
rect 798 181488 219120 181768
rect 798 180136 219200 181488
rect 880 179856 219200 180136
rect 798 179592 219200 179856
rect 798 179312 219120 179592
rect 798 177960 219200 179312
rect 880 177680 219200 177960
rect 798 177416 219200 177680
rect 798 177136 219120 177416
rect 798 175920 219200 177136
rect 880 175640 219200 175920
rect 798 175240 219200 175640
rect 798 174960 219120 175240
rect 798 173744 219200 174960
rect 880 173464 219200 173744
rect 798 173064 219200 173464
rect 798 172784 219120 173064
rect 798 171704 219200 172784
rect 880 171424 219200 171704
rect 798 170752 219200 171424
rect 798 170472 219120 170752
rect 798 169528 219200 170472
rect 880 169248 219200 169528
rect 798 168576 219200 169248
rect 798 168296 219120 168576
rect 798 167488 219200 168296
rect 880 167208 219200 167488
rect 798 166400 219200 167208
rect 798 166120 219120 166400
rect 798 165312 219200 166120
rect 880 165032 219200 165312
rect 798 164224 219200 165032
rect 798 163944 219120 164224
rect 798 163272 219200 163944
rect 880 162992 219200 163272
rect 798 162048 219200 162992
rect 798 161768 219120 162048
rect 798 161096 219200 161768
rect 880 160816 219200 161096
rect 798 159736 219200 160816
rect 798 159456 219120 159736
rect 798 159056 219200 159456
rect 880 158776 219200 159056
rect 798 157560 219200 158776
rect 798 157280 219120 157560
rect 798 156880 219200 157280
rect 880 156600 219200 156880
rect 798 155384 219200 156600
rect 798 155104 219120 155384
rect 798 154840 219200 155104
rect 880 154560 219200 154840
rect 798 153208 219200 154560
rect 798 152928 219120 153208
rect 798 152664 219200 152928
rect 880 152384 219200 152664
rect 798 151032 219200 152384
rect 798 150752 219120 151032
rect 798 150624 219200 150752
rect 880 150344 219200 150624
rect 798 148720 219200 150344
rect 798 148448 219120 148720
rect 880 148440 219120 148448
rect 880 148168 219200 148440
rect 798 146544 219200 148168
rect 798 146408 219120 146544
rect 880 146264 219120 146408
rect 880 146128 219200 146264
rect 798 144368 219200 146128
rect 798 144232 219120 144368
rect 880 144088 219120 144232
rect 880 143952 219200 144088
rect 798 142192 219200 143952
rect 880 141912 219120 142192
rect 798 140016 219200 141912
rect 880 139736 219120 140016
rect 798 137976 219200 139736
rect 880 137704 219200 137976
rect 880 137696 219120 137704
rect 798 137424 219120 137696
rect 798 135800 219200 137424
rect 880 135528 219200 135800
rect 880 135520 219120 135528
rect 798 135248 219120 135520
rect 798 133760 219200 135248
rect 880 133480 219200 133760
rect 798 133352 219200 133480
rect 798 133072 219120 133352
rect 798 131584 219200 133072
rect 880 131304 219200 131584
rect 798 131176 219200 131304
rect 798 130896 219120 131176
rect 798 129544 219200 130896
rect 880 129264 219200 129544
rect 798 129000 219200 129264
rect 798 128720 219120 129000
rect 798 127368 219200 128720
rect 880 127088 219200 127368
rect 798 126688 219200 127088
rect 798 126408 219120 126688
rect 798 125328 219200 126408
rect 880 125048 219200 125328
rect 798 124512 219200 125048
rect 798 124232 219120 124512
rect 798 123152 219200 124232
rect 880 122872 219200 123152
rect 798 122336 219200 122872
rect 798 122056 219120 122336
rect 798 121112 219200 122056
rect 880 120832 219200 121112
rect 798 120160 219200 120832
rect 798 119880 219120 120160
rect 798 119072 219200 119880
rect 880 118792 219200 119072
rect 798 117984 219200 118792
rect 798 117704 219120 117984
rect 798 116896 219200 117704
rect 880 116616 219200 116896
rect 798 115808 219200 116616
rect 798 115528 219120 115808
rect 798 114856 219200 115528
rect 880 114576 219200 114856
rect 798 113496 219200 114576
rect 798 113216 219120 113496
rect 798 112680 219200 113216
rect 880 112400 219200 112680
rect 798 111320 219200 112400
rect 798 111040 219120 111320
rect 798 110640 219200 111040
rect 880 110360 219200 110640
rect 798 109144 219200 110360
rect 798 108864 219120 109144
rect 798 108464 219200 108864
rect 880 108184 219200 108464
rect 798 106968 219200 108184
rect 798 106688 219120 106968
rect 798 106424 219200 106688
rect 880 106144 219200 106424
rect 798 104792 219200 106144
rect 798 104512 219120 104792
rect 798 104248 219200 104512
rect 880 103968 219200 104248
rect 798 102480 219200 103968
rect 798 102208 219120 102480
rect 880 102200 219120 102208
rect 880 101928 219200 102200
rect 798 100304 219200 101928
rect 798 100032 219120 100304
rect 880 100024 219120 100032
rect 880 99752 219200 100024
rect 798 98128 219200 99752
rect 798 97992 219120 98128
rect 880 97848 219120 97992
rect 880 97712 219200 97848
rect 798 95952 219200 97712
rect 798 95816 219120 95952
rect 880 95672 219120 95816
rect 880 95536 219200 95672
rect 798 93776 219200 95536
rect 880 93496 219120 93776
rect 798 91600 219200 93496
rect 880 91464 219200 91600
rect 880 91320 219120 91464
rect 798 91184 219120 91320
rect 798 89560 219200 91184
rect 880 89288 219200 89560
rect 880 89280 219120 89288
rect 798 89008 219120 89280
rect 798 87384 219200 89008
rect 880 87112 219200 87384
rect 880 87104 219120 87112
rect 798 86832 219120 87104
rect 798 85344 219200 86832
rect 880 85064 219200 85344
rect 798 84936 219200 85064
rect 798 84656 219120 84936
rect 798 83168 219200 84656
rect 880 82888 219200 83168
rect 798 82760 219200 82888
rect 798 82480 219120 82760
rect 798 81128 219200 82480
rect 880 80848 219200 81128
rect 798 80448 219200 80848
rect 798 80168 219120 80448
rect 798 78952 219200 80168
rect 880 78672 219200 78952
rect 798 78272 219200 78672
rect 798 77992 219120 78272
rect 798 76912 219200 77992
rect 880 76632 219200 76912
rect 798 76096 219200 76632
rect 798 75816 219120 76096
rect 798 74736 219200 75816
rect 880 74456 219200 74736
rect 798 73920 219200 74456
rect 798 73640 219120 73920
rect 798 72696 219200 73640
rect 880 72416 219200 72696
rect 798 71744 219200 72416
rect 798 71464 219120 71744
rect 798 70520 219200 71464
rect 880 70240 219200 70520
rect 798 69432 219200 70240
rect 798 69152 219120 69432
rect 798 68480 219200 69152
rect 880 68200 219200 68480
rect 798 67256 219200 68200
rect 798 66976 219120 67256
rect 798 66304 219200 66976
rect 880 66024 219200 66304
rect 798 65080 219200 66024
rect 798 64800 219120 65080
rect 798 64264 219200 64800
rect 880 63984 219200 64264
rect 798 62904 219200 63984
rect 798 62624 219120 62904
rect 798 62088 219200 62624
rect 880 61808 219200 62088
rect 798 60728 219200 61808
rect 798 60448 219120 60728
rect 798 60048 219200 60448
rect 880 59768 219200 60048
rect 798 58552 219200 59768
rect 798 58272 219120 58552
rect 798 58008 219200 58272
rect 880 57728 219200 58008
rect 798 56240 219200 57728
rect 798 55960 219120 56240
rect 798 55832 219200 55960
rect 880 55552 219200 55832
rect 798 54064 219200 55552
rect 798 53792 219120 54064
rect 880 53784 219120 53792
rect 880 53512 219200 53784
rect 798 51888 219200 53512
rect 798 51616 219120 51888
rect 880 51608 219120 51616
rect 880 51336 219200 51608
rect 798 49712 219200 51336
rect 798 49576 219120 49712
rect 880 49432 219120 49576
rect 880 49296 219200 49432
rect 798 47536 219200 49296
rect 798 47400 219120 47536
rect 880 47256 219120 47400
rect 880 47120 219200 47256
rect 798 45360 219200 47120
rect 880 45224 219200 45360
rect 880 45080 219120 45224
rect 798 44944 219120 45080
rect 798 43184 219200 44944
rect 880 43048 219200 43184
rect 880 42904 219120 43048
rect 798 42768 219120 42904
rect 798 41144 219200 42768
rect 880 40872 219200 41144
rect 880 40864 219120 40872
rect 798 40592 219120 40864
rect 798 38968 219200 40592
rect 880 38696 219200 38968
rect 880 38688 219120 38696
rect 798 38416 219120 38688
rect 798 36928 219200 38416
rect 880 36648 219200 36928
rect 798 36520 219200 36648
rect 798 36240 219120 36520
rect 798 34752 219200 36240
rect 880 34472 219200 34752
rect 798 34208 219200 34472
rect 798 33928 219120 34208
rect 798 32712 219200 33928
rect 880 32432 219200 32712
rect 798 32032 219200 32432
rect 798 31752 219120 32032
rect 798 30536 219200 31752
rect 880 30256 219200 30536
rect 798 29856 219200 30256
rect 798 29576 219120 29856
rect 798 28496 219200 29576
rect 880 28216 219200 28496
rect 798 27680 219200 28216
rect 798 27400 219120 27680
rect 798 26320 219200 27400
rect 880 26040 219200 26320
rect 798 25504 219200 26040
rect 798 25224 219120 25504
rect 798 24280 219200 25224
rect 880 24000 219200 24280
rect 798 23192 219200 24000
rect 798 22912 219120 23192
rect 798 22104 219200 22912
rect 880 21824 219200 22104
rect 798 21016 219200 21824
rect 798 20736 219120 21016
rect 798 20064 219200 20736
rect 880 19784 219200 20064
rect 798 18840 219200 19784
rect 798 18560 219120 18840
rect 798 17888 219200 18560
rect 880 17608 219200 17888
rect 798 16664 219200 17608
rect 798 16384 219120 16664
rect 798 15848 219200 16384
rect 880 15568 219200 15848
rect 798 14488 219200 15568
rect 798 14208 219120 14488
rect 798 13672 219200 14208
rect 880 13392 219200 13672
rect 798 12176 219200 13392
rect 798 11896 219120 12176
rect 798 11632 219200 11896
rect 880 11352 219200 11632
rect 798 10000 219200 11352
rect 798 9720 219120 10000
rect 798 9456 219200 9720
rect 880 9176 219200 9456
rect 798 7824 219200 9176
rect 798 7544 219120 7824
rect 798 7416 219200 7544
rect 880 7136 219200 7416
rect 798 5648 219200 7136
rect 798 5368 219120 5648
rect 798 5240 219200 5368
rect 880 4960 219200 5240
rect 798 3472 219200 4960
rect 798 3200 219120 3472
rect 880 3192 219120 3200
rect 880 2920 219200 3192
rect 798 1296 219200 2920
rect 798 1160 219120 1296
rect 880 1016 219120 1160
rect 880 880 219200 1016
rect 798 851 219200 880
<< metal4 >>
rect 4208 2128 4528 237776
rect 19568 2128 19888 237776
<< obsm4 >>
rect 2819 2128 4128 237776
rect 4608 2128 19488 237776
rect 19968 2128 217613 237776
<< labels >>
rlabel metal3 s 219200 97928 220000 98048 6 cpu_addr_e[0]
port 1 nsew default output
rlabel metal3 s 219200 119960 220000 120080 6 cpu_addr_e[10]
port 2 nsew default output
rlabel metal3 s 219200 122136 220000 122256 6 cpu_addr_e[11]
port 3 nsew default output
rlabel metal3 s 219200 124312 220000 124432 6 cpu_addr_e[12]
port 4 nsew default output
rlabel metal3 s 219200 126488 220000 126608 6 cpu_addr_e[13]
port 5 nsew default output
rlabel metal3 s 219200 128800 220000 128920 6 cpu_addr_e[14]
port 6 nsew default output
rlabel metal3 s 219200 130976 220000 131096 6 cpu_addr_e[15]
port 7 nsew default output
rlabel metal3 s 219200 100104 220000 100224 6 cpu_addr_e[1]
port 8 nsew default output
rlabel metal3 s 219200 102280 220000 102400 6 cpu_addr_e[2]
port 9 nsew default output
rlabel metal3 s 219200 104592 220000 104712 6 cpu_addr_e[3]
port 10 nsew default output
rlabel metal3 s 219200 106768 220000 106888 6 cpu_addr_e[4]
port 11 nsew default output
rlabel metal3 s 219200 108944 220000 109064 6 cpu_addr_e[5]
port 12 nsew default output
rlabel metal3 s 219200 111120 220000 111240 6 cpu_addr_e[6]
port 13 nsew default output
rlabel metal3 s 219200 113296 220000 113416 6 cpu_addr_e[7]
port 14 nsew default output
rlabel metal3 s 219200 115608 220000 115728 6 cpu_addr_e[8]
port 15 nsew default output
rlabel metal3 s 219200 117784 220000 117904 6 cpu_addr_e[9]
port 16 nsew default output
rlabel metal2 s 67362 239200 67418 240000 6 cpu_addr_n[0]
port 17 nsew default output
rlabel metal2 s 88154 239200 88210 240000 6 cpu_addr_n[10]
port 18 nsew default output
rlabel metal2 s 90178 239200 90234 240000 6 cpu_addr_n[11]
port 19 nsew default output
rlabel metal2 s 92294 239200 92350 240000 6 cpu_addr_n[12]
port 20 nsew default output
rlabel metal2 s 94410 239200 94466 240000 6 cpu_addr_n[13]
port 21 nsew default output
rlabel metal2 s 96434 239200 96490 240000 6 cpu_addr_n[14]
port 22 nsew default output
rlabel metal2 s 98550 239200 98606 240000 6 cpu_addr_n[15]
port 23 nsew default output
rlabel metal2 s 69478 239200 69534 240000 6 cpu_addr_n[1]
port 24 nsew default output
rlabel metal2 s 71502 239200 71558 240000 6 cpu_addr_n[2]
port 25 nsew default output
rlabel metal2 s 73618 239200 73674 240000 6 cpu_addr_n[3]
port 26 nsew default output
rlabel metal2 s 75734 239200 75790 240000 6 cpu_addr_n[4]
port 27 nsew default output
rlabel metal2 s 77758 239200 77814 240000 6 cpu_addr_n[5]
port 28 nsew default output
rlabel metal2 s 79874 239200 79930 240000 6 cpu_addr_n[6]
port 29 nsew default output
rlabel metal2 s 81898 239200 81954 240000 6 cpu_addr_n[7]
port 30 nsew default output
rlabel metal2 s 84014 239200 84070 240000 6 cpu_addr_n[8]
port 31 nsew default output
rlabel metal2 s 86038 239200 86094 240000 6 cpu_addr_n[9]
port 32 nsew default output
rlabel metal3 s 219200 5448 220000 5568 6 cpu_dtr_e0[0]
port 33 nsew default input
rlabel metal3 s 219200 27480 220000 27600 6 cpu_dtr_e0[10]
port 34 nsew default input
rlabel metal3 s 219200 29656 220000 29776 6 cpu_dtr_e0[11]
port 35 nsew default input
rlabel metal3 s 219200 31832 220000 31952 6 cpu_dtr_e0[12]
port 36 nsew default input
rlabel metal3 s 219200 34008 220000 34128 6 cpu_dtr_e0[13]
port 37 nsew default input
rlabel metal3 s 219200 36320 220000 36440 6 cpu_dtr_e0[14]
port 38 nsew default input
rlabel metal3 s 219200 38496 220000 38616 6 cpu_dtr_e0[15]
port 39 nsew default input
rlabel metal3 s 219200 40672 220000 40792 6 cpu_dtr_e0[16]
port 40 nsew default input
rlabel metal3 s 219200 42848 220000 42968 6 cpu_dtr_e0[17]
port 41 nsew default input
rlabel metal3 s 219200 45024 220000 45144 6 cpu_dtr_e0[18]
port 42 nsew default input
rlabel metal3 s 219200 47336 220000 47456 6 cpu_dtr_e0[19]
port 43 nsew default input
rlabel metal3 s 219200 7624 220000 7744 6 cpu_dtr_e0[1]
port 44 nsew default input
rlabel metal3 s 219200 49512 220000 49632 6 cpu_dtr_e0[20]
port 45 nsew default input
rlabel metal3 s 219200 51688 220000 51808 6 cpu_dtr_e0[21]
port 46 nsew default input
rlabel metal3 s 219200 53864 220000 53984 6 cpu_dtr_e0[22]
port 47 nsew default input
rlabel metal3 s 219200 56040 220000 56160 6 cpu_dtr_e0[23]
port 48 nsew default input
rlabel metal3 s 219200 58352 220000 58472 6 cpu_dtr_e0[24]
port 49 nsew default input
rlabel metal3 s 219200 60528 220000 60648 6 cpu_dtr_e0[25]
port 50 nsew default input
rlabel metal3 s 219200 62704 220000 62824 6 cpu_dtr_e0[26]
port 51 nsew default input
rlabel metal3 s 219200 64880 220000 65000 6 cpu_dtr_e0[27]
port 52 nsew default input
rlabel metal3 s 219200 67056 220000 67176 6 cpu_dtr_e0[28]
port 53 nsew default input
rlabel metal3 s 219200 69232 220000 69352 6 cpu_dtr_e0[29]
port 54 nsew default input
rlabel metal3 s 219200 9800 220000 9920 6 cpu_dtr_e0[2]
port 55 nsew default input
rlabel metal3 s 219200 71544 220000 71664 6 cpu_dtr_e0[30]
port 56 nsew default input
rlabel metal3 s 219200 73720 220000 73840 6 cpu_dtr_e0[31]
port 57 nsew default input
rlabel metal3 s 219200 11976 220000 12096 6 cpu_dtr_e0[3]
port 58 nsew default input
rlabel metal3 s 219200 14288 220000 14408 6 cpu_dtr_e0[4]
port 59 nsew default input
rlabel metal3 s 219200 16464 220000 16584 6 cpu_dtr_e0[5]
port 60 nsew default input
rlabel metal3 s 219200 18640 220000 18760 6 cpu_dtr_e0[6]
port 61 nsew default input
rlabel metal3 s 219200 20816 220000 20936 6 cpu_dtr_e0[7]
port 62 nsew default input
rlabel metal3 s 219200 22992 220000 23112 6 cpu_dtr_e0[8]
port 63 nsew default input
rlabel metal3 s 219200 25304 220000 25424 6 cpu_dtr_e0[9]
port 64 nsew default input
rlabel metal3 s 219200 168376 220000 168496 6 cpu_dtr_e1[0]
port 65 nsew default input
rlabel metal3 s 219200 190408 220000 190528 6 cpu_dtr_e1[10]
port 66 nsew default input
rlabel metal3 s 219200 192584 220000 192704 6 cpu_dtr_e1[11]
port 67 nsew default input
rlabel metal3 s 219200 194760 220000 194880 6 cpu_dtr_e1[12]
port 68 nsew default input
rlabel metal3 s 219200 197072 220000 197192 6 cpu_dtr_e1[13]
port 69 nsew default input
rlabel metal3 s 219200 199248 220000 199368 6 cpu_dtr_e1[14]
port 70 nsew default input
rlabel metal3 s 219200 201424 220000 201544 6 cpu_dtr_e1[15]
port 71 nsew default input
rlabel metal3 s 219200 203600 220000 203720 6 cpu_dtr_e1[16]
port 72 nsew default input
rlabel metal3 s 219200 205776 220000 205896 6 cpu_dtr_e1[17]
port 73 nsew default input
rlabel metal3 s 219200 208088 220000 208208 6 cpu_dtr_e1[18]
port 74 nsew default input
rlabel metal3 s 219200 210264 220000 210384 6 cpu_dtr_e1[19]
port 75 nsew default input
rlabel metal3 s 219200 170552 220000 170672 6 cpu_dtr_e1[1]
port 76 nsew default input
rlabel metal3 s 219200 212440 220000 212560 6 cpu_dtr_e1[20]
port 77 nsew default input
rlabel metal3 s 219200 214616 220000 214736 6 cpu_dtr_e1[21]
port 78 nsew default input
rlabel metal3 s 219200 216792 220000 216912 6 cpu_dtr_e1[22]
port 79 nsew default input
rlabel metal3 s 219200 219104 220000 219224 6 cpu_dtr_e1[23]
port 80 nsew default input
rlabel metal3 s 219200 221280 220000 221400 6 cpu_dtr_e1[24]
port 81 nsew default input
rlabel metal3 s 219200 223456 220000 223576 6 cpu_dtr_e1[25]
port 82 nsew default input
rlabel metal3 s 219200 225632 220000 225752 6 cpu_dtr_e1[26]
port 83 nsew default input
rlabel metal3 s 219200 227808 220000 227928 6 cpu_dtr_e1[27]
port 84 nsew default input
rlabel metal3 s 219200 230120 220000 230240 6 cpu_dtr_e1[28]
port 85 nsew default input
rlabel metal3 s 219200 232296 220000 232416 6 cpu_dtr_e1[29]
port 86 nsew default input
rlabel metal3 s 219200 172864 220000 172984 6 cpu_dtr_e1[2]
port 87 nsew default input
rlabel metal3 s 219200 234472 220000 234592 6 cpu_dtr_e1[30]
port 88 nsew default input
rlabel metal3 s 219200 236648 220000 236768 6 cpu_dtr_e1[31]
port 89 nsew default input
rlabel metal3 s 219200 175040 220000 175160 6 cpu_dtr_e1[3]
port 90 nsew default input
rlabel metal3 s 219200 177216 220000 177336 6 cpu_dtr_e1[4]
port 91 nsew default input
rlabel metal3 s 219200 179392 220000 179512 6 cpu_dtr_e1[5]
port 92 nsew default input
rlabel metal3 s 219200 181568 220000 181688 6 cpu_dtr_e1[6]
port 93 nsew default input
rlabel metal3 s 219200 183744 220000 183864 6 cpu_dtr_e1[7]
port 94 nsew default input
rlabel metal3 s 219200 186056 220000 186176 6 cpu_dtr_e1[8]
port 95 nsew default input
rlabel metal3 s 219200 188232 220000 188352 6 cpu_dtr_e1[9]
port 96 nsew default input
rlabel metal2 s 1030 239200 1086 240000 6 cpu_dtr_n0[0]
port 97 nsew default input
rlabel metal2 s 21730 239200 21786 240000 6 cpu_dtr_n0[10]
port 98 nsew default input
rlabel metal2 s 23846 239200 23902 240000 6 cpu_dtr_n0[11]
port 99 nsew default input
rlabel metal2 s 25870 239200 25926 240000 6 cpu_dtr_n0[12]
port 100 nsew default input
rlabel metal2 s 27986 239200 28042 240000 6 cpu_dtr_n0[13]
port 101 nsew default input
rlabel metal2 s 30010 239200 30066 240000 6 cpu_dtr_n0[14]
port 102 nsew default input
rlabel metal2 s 32126 239200 32182 240000 6 cpu_dtr_n0[15]
port 103 nsew default input
rlabel metal2 s 34150 239200 34206 240000 6 cpu_dtr_n0[16]
port 104 nsew default input
rlabel metal2 s 36266 239200 36322 240000 6 cpu_dtr_n0[17]
port 105 nsew default input
rlabel metal2 s 38382 239200 38438 240000 6 cpu_dtr_n0[18]
port 106 nsew default input
rlabel metal2 s 40406 239200 40462 240000 6 cpu_dtr_n0[19]
port 107 nsew default input
rlabel metal2 s 3054 239200 3110 240000 6 cpu_dtr_n0[1]
port 108 nsew default input
rlabel metal2 s 42522 239200 42578 240000 6 cpu_dtr_n0[20]
port 109 nsew default input
rlabel metal2 s 44546 239200 44602 240000 6 cpu_dtr_n0[21]
port 110 nsew default input
rlabel metal2 s 46662 239200 46718 240000 6 cpu_dtr_n0[22]
port 111 nsew default input
rlabel metal2 s 48686 239200 48742 240000 6 cpu_dtr_n0[23]
port 112 nsew default input
rlabel metal2 s 50802 239200 50858 240000 6 cpu_dtr_n0[24]
port 113 nsew default input
rlabel metal2 s 52826 239200 52882 240000 6 cpu_dtr_n0[25]
port 114 nsew default input
rlabel metal2 s 54942 239200 54998 240000 6 cpu_dtr_n0[26]
port 115 nsew default input
rlabel metal2 s 57058 239200 57114 240000 6 cpu_dtr_n0[27]
port 116 nsew default input
rlabel metal2 s 59082 239200 59138 240000 6 cpu_dtr_n0[28]
port 117 nsew default input
rlabel metal2 s 61198 239200 61254 240000 6 cpu_dtr_n0[29]
port 118 nsew default input
rlabel metal2 s 5170 239200 5226 240000 6 cpu_dtr_n0[2]
port 119 nsew default input
rlabel metal2 s 63222 239200 63278 240000 6 cpu_dtr_n0[30]
port 120 nsew default input
rlabel metal2 s 65338 239200 65394 240000 6 cpu_dtr_n0[31]
port 121 nsew default input
rlabel metal2 s 7194 239200 7250 240000 6 cpu_dtr_n0[3]
port 122 nsew default input
rlabel metal2 s 9310 239200 9366 240000 6 cpu_dtr_n0[4]
port 123 nsew default input
rlabel metal2 s 11334 239200 11390 240000 6 cpu_dtr_n0[5]
port 124 nsew default input
rlabel metal2 s 13450 239200 13506 240000 6 cpu_dtr_n0[6]
port 125 nsew default input
rlabel metal2 s 15474 239200 15530 240000 6 cpu_dtr_n0[7]
port 126 nsew default input
rlabel metal2 s 17590 239200 17646 240000 6 cpu_dtr_n0[8]
port 127 nsew default input
rlabel metal2 s 19706 239200 19762 240000 6 cpu_dtr_n0[9]
port 128 nsew default input
rlabel metal2 s 154578 239200 154634 240000 6 cpu_dtr_n1[0]
port 129 nsew default input
rlabel metal2 s 175278 239200 175334 240000 6 cpu_dtr_n1[10]
port 130 nsew default input
rlabel metal2 s 177394 239200 177450 240000 6 cpu_dtr_n1[11]
port 131 nsew default input
rlabel metal2 s 179418 239200 179474 240000 6 cpu_dtr_n1[12]
port 132 nsew default input
rlabel metal2 s 181534 239200 181590 240000 6 cpu_dtr_n1[13]
port 133 nsew default input
rlabel metal2 s 183558 239200 183614 240000 6 cpu_dtr_n1[14]
port 134 nsew default input
rlabel metal2 s 185674 239200 185730 240000 6 cpu_dtr_n1[15]
port 135 nsew default input
rlabel metal2 s 187790 239200 187846 240000 6 cpu_dtr_n1[16]
port 136 nsew default input
rlabel metal2 s 189814 239200 189870 240000 6 cpu_dtr_n1[17]
port 137 nsew default input
rlabel metal2 s 191930 239200 191986 240000 6 cpu_dtr_n1[18]
port 138 nsew default input
rlabel metal2 s 193954 239200 194010 240000 6 cpu_dtr_n1[19]
port 139 nsew default input
rlabel metal2 s 156602 239200 156658 240000 6 cpu_dtr_n1[1]
port 140 nsew default input
rlabel metal2 s 196070 239200 196126 240000 6 cpu_dtr_n1[20]
port 141 nsew default input
rlabel metal2 s 198094 239200 198150 240000 6 cpu_dtr_n1[21]
port 142 nsew default input
rlabel metal2 s 200210 239200 200266 240000 6 cpu_dtr_n1[22]
port 143 nsew default input
rlabel metal2 s 202234 239200 202290 240000 6 cpu_dtr_n1[23]
port 144 nsew default input
rlabel metal2 s 204350 239200 204406 240000 6 cpu_dtr_n1[24]
port 145 nsew default input
rlabel metal2 s 206466 239200 206522 240000 6 cpu_dtr_n1[25]
port 146 nsew default input
rlabel metal2 s 208490 239200 208546 240000 6 cpu_dtr_n1[26]
port 147 nsew default input
rlabel metal2 s 210606 239200 210662 240000 6 cpu_dtr_n1[27]
port 148 nsew default input
rlabel metal2 s 212630 239200 212686 240000 6 cpu_dtr_n1[28]
port 149 nsew default input
rlabel metal2 s 214746 239200 214802 240000 6 cpu_dtr_n1[29]
port 150 nsew default input
rlabel metal2 s 158718 239200 158774 240000 6 cpu_dtr_n1[2]
port 151 nsew default input
rlabel metal2 s 216770 239200 216826 240000 6 cpu_dtr_n1[30]
port 152 nsew default input
rlabel metal2 s 218886 239200 218942 240000 6 cpu_dtr_n1[31]
port 153 nsew default input
rlabel metal2 s 160742 239200 160798 240000 6 cpu_dtr_n1[3]
port 154 nsew default input
rlabel metal2 s 162858 239200 162914 240000 6 cpu_dtr_n1[4]
port 155 nsew default input
rlabel metal2 s 164882 239200 164938 240000 6 cpu_dtr_n1[5]
port 156 nsew default input
rlabel metal2 s 166998 239200 167054 240000 6 cpu_dtr_n1[6]
port 157 nsew default input
rlabel metal2 s 169114 239200 169170 240000 6 cpu_dtr_n1[7]
port 158 nsew default input
rlabel metal2 s 171138 239200 171194 240000 6 cpu_dtr_n1[8]
port 159 nsew default input
rlabel metal2 s 173254 239200 173310 240000 6 cpu_dtr_n1[9]
port 160 nsew default input
rlabel metal3 s 219200 133152 220000 133272 6 cpu_dtw_e[0]
port 161 nsew default output
rlabel metal3 s 219200 155184 220000 155304 6 cpu_dtw_e[10]
port 162 nsew default output
rlabel metal3 s 219200 157360 220000 157480 6 cpu_dtw_e[11]
port 163 nsew default output
rlabel metal3 s 219200 159536 220000 159656 6 cpu_dtw_e[12]
port 164 nsew default output
rlabel metal3 s 219200 161848 220000 161968 6 cpu_dtw_e[13]
port 165 nsew default output
rlabel metal3 s 219200 164024 220000 164144 6 cpu_dtw_e[14]
port 166 nsew default output
rlabel metal3 s 219200 166200 220000 166320 6 cpu_dtw_e[15]
port 167 nsew default output
rlabel metal3 s 219200 135328 220000 135448 6 cpu_dtw_e[1]
port 168 nsew default output
rlabel metal3 s 219200 137504 220000 137624 6 cpu_dtw_e[2]
port 169 nsew default output
rlabel metal3 s 219200 139816 220000 139936 6 cpu_dtw_e[3]
port 170 nsew default output
rlabel metal3 s 219200 141992 220000 142112 6 cpu_dtw_e[4]
port 171 nsew default output
rlabel metal3 s 219200 144168 220000 144288 6 cpu_dtw_e[5]
port 172 nsew default output
rlabel metal3 s 219200 146344 220000 146464 6 cpu_dtw_e[6]
port 173 nsew default output
rlabel metal3 s 219200 148520 220000 148640 6 cpu_dtw_e[7]
port 174 nsew default output
rlabel metal3 s 219200 150832 220000 150952 6 cpu_dtw_e[8]
port 175 nsew default output
rlabel metal3 s 219200 153008 220000 153128 6 cpu_dtw_e[9]
port 176 nsew default output
rlabel metal2 s 121366 239200 121422 240000 6 cpu_dtw_n[0]
port 177 nsew default output
rlabel metal2 s 142066 239200 142122 240000 6 cpu_dtw_n[10]
port 178 nsew default output
rlabel metal2 s 144182 239200 144238 240000 6 cpu_dtw_n[11]
port 179 nsew default output
rlabel metal2 s 146206 239200 146262 240000 6 cpu_dtw_n[12]
port 180 nsew default output
rlabel metal2 s 148322 239200 148378 240000 6 cpu_dtw_n[13]
port 181 nsew default output
rlabel metal2 s 150438 239200 150494 240000 6 cpu_dtw_n[14]
port 182 nsew default output
rlabel metal2 s 152462 239200 152518 240000 6 cpu_dtw_n[15]
port 183 nsew default output
rlabel metal2 s 123390 239200 123446 240000 6 cpu_dtw_n[1]
port 184 nsew default output
rlabel metal2 s 125506 239200 125562 240000 6 cpu_dtw_n[2]
port 185 nsew default output
rlabel metal2 s 127530 239200 127586 240000 6 cpu_dtw_n[3]
port 186 nsew default output
rlabel metal2 s 129646 239200 129702 240000 6 cpu_dtw_n[4]
port 187 nsew default output
rlabel metal2 s 131762 239200 131818 240000 6 cpu_dtw_n[5]
port 188 nsew default output
rlabel metal2 s 133786 239200 133842 240000 6 cpu_dtw_n[6]
port 189 nsew default output
rlabel metal2 s 135902 239200 135958 240000 6 cpu_dtw_n[7]
port 190 nsew default output
rlabel metal2 s 137926 239200 137982 240000 6 cpu_dtw_n[8]
port 191 nsew default output
rlabel metal2 s 140042 239200 140098 240000 6 cpu_dtw_n[9]
port 192 nsew default output
rlabel metal3 s 219200 75896 220000 76016 6 cpu_mask_e[0]
port 193 nsew default output
rlabel metal3 s 219200 78072 220000 78192 6 cpu_mask_e[1]
port 194 nsew default output
rlabel metal3 s 219200 80248 220000 80368 6 cpu_mask_e[2]
port 195 nsew default output
rlabel metal3 s 219200 82560 220000 82680 6 cpu_mask_e[3]
port 196 nsew default output
rlabel metal3 s 219200 84736 220000 84856 6 cpu_mask_e[4]
port 197 nsew default output
rlabel metal3 s 219200 86912 220000 87032 6 cpu_mask_e[5]
port 198 nsew default output
rlabel metal3 s 219200 89088 220000 89208 6 cpu_mask_e[6]
port 199 nsew default output
rlabel metal3 s 219200 91264 220000 91384 6 cpu_mask_e[7]
port 200 nsew default output
rlabel metal2 s 100574 239200 100630 240000 6 cpu_mask_n[0]
port 201 nsew default output
rlabel metal2 s 102690 239200 102746 240000 6 cpu_mask_n[1]
port 202 nsew default output
rlabel metal2 s 104714 239200 104770 240000 6 cpu_mask_n[2]
port 203 nsew default output
rlabel metal2 s 106830 239200 106886 240000 6 cpu_mask_n[3]
port 204 nsew default output
rlabel metal2 s 108854 239200 108910 240000 6 cpu_mask_n[4]
port 205 nsew default output
rlabel metal2 s 110970 239200 111026 240000 6 cpu_mask_n[5]
port 206 nsew default output
rlabel metal2 s 113086 239200 113142 240000 6 cpu_mask_n[6]
port 207 nsew default output
rlabel metal2 s 115110 239200 115166 240000 6 cpu_mask_n[7]
port 208 nsew default output
rlabel metal3 s 219200 93576 220000 93696 6 cpu_wen_e[0]
port 209 nsew default output
rlabel metal3 s 219200 95752 220000 95872 6 cpu_wen_e[1]
port 210 nsew default output
rlabel metal2 s 117226 239200 117282 240000 6 cpu_wen_n[0]
port 211 nsew default output
rlabel metal2 s 119250 239200 119306 240000 6 cpu_wen_n[1]
port 212 nsew default output
rlabel metal3 s 0 960 800 1080 6 io_in[0]
port 213 nsew default input
rlabel metal3 s 0 64064 800 64184 6 io_in[10]
port 214 nsew default input
rlabel metal3 s 0 70320 800 70440 6 io_in[11]
port 215 nsew default input
rlabel metal3 s 0 76712 800 76832 6 io_in[12]
port 216 nsew default input
rlabel metal3 s 0 82968 800 83088 6 io_in[13]
port 217 nsew default input
rlabel metal3 s 0 89360 800 89480 6 io_in[14]
port 218 nsew default input
rlabel metal3 s 0 95616 800 95736 6 io_in[15]
port 219 nsew default input
rlabel metal3 s 0 102008 800 102128 6 io_in[16]
port 220 nsew default input
rlabel metal3 s 0 108264 800 108384 6 io_in[17]
port 221 nsew default input
rlabel metal3 s 0 114656 800 114776 6 io_in[18]
port 222 nsew default input
rlabel metal3 s 0 120912 800 121032 6 io_in[19]
port 223 nsew default input
rlabel metal3 s 0 7216 800 7336 6 io_in[1]
port 224 nsew default input
rlabel metal3 s 0 127168 800 127288 6 io_in[20]
port 225 nsew default input
rlabel metal3 s 0 133560 800 133680 6 io_in[21]
port 226 nsew default input
rlabel metal3 s 0 139816 800 139936 6 io_in[22]
port 227 nsew default input
rlabel metal3 s 0 146208 800 146328 6 io_in[23]
port 228 nsew default input
rlabel metal3 s 0 152464 800 152584 6 io_in[24]
port 229 nsew default input
rlabel metal3 s 0 158856 800 158976 6 io_in[25]
port 230 nsew default input
rlabel metal3 s 0 165112 800 165232 6 io_in[26]
port 231 nsew default input
rlabel metal3 s 0 171504 800 171624 6 io_in[27]
port 232 nsew default input
rlabel metal3 s 0 177760 800 177880 6 io_in[28]
port 233 nsew default input
rlabel metal3 s 0 184016 800 184136 6 io_in[29]
port 234 nsew default input
rlabel metal3 s 0 13472 800 13592 6 io_in[2]
port 235 nsew default input
rlabel metal3 s 0 190408 800 190528 6 io_in[30]
port 236 nsew default input
rlabel metal3 s 0 196664 800 196784 6 io_in[31]
port 237 nsew default input
rlabel metal3 s 0 203056 800 203176 6 io_in[32]
port 238 nsew default input
rlabel metal3 s 0 209312 800 209432 6 io_in[33]
port 239 nsew default input
rlabel metal3 s 0 215704 800 215824 6 io_in[34]
port 240 nsew default input
rlabel metal3 s 0 221960 800 222080 6 io_in[35]
port 241 nsew default input
rlabel metal3 s 0 228352 800 228472 6 io_in[36]
port 242 nsew default input
rlabel metal3 s 0 234608 800 234728 6 io_in[37]
port 243 nsew default input
rlabel metal3 s 0 19864 800 19984 6 io_in[3]
port 244 nsew default input
rlabel metal3 s 0 26120 800 26240 6 io_in[4]
port 245 nsew default input
rlabel metal3 s 0 32512 800 32632 6 io_in[5]
port 246 nsew default input
rlabel metal3 s 0 38768 800 38888 6 io_in[6]
port 247 nsew default input
rlabel metal3 s 0 45160 800 45280 6 io_in[7]
port 248 nsew default input
rlabel metal3 s 0 51416 800 51536 6 io_in[8]
port 249 nsew default input
rlabel metal3 s 0 57808 800 57928 6 io_in[9]
port 250 nsew default input
rlabel metal3 s 0 3000 800 3120 6 io_oeb[0]
port 251 nsew default output
rlabel metal3 s 0 66104 800 66224 6 io_oeb[10]
port 252 nsew default output
rlabel metal3 s 0 72496 800 72616 6 io_oeb[11]
port 253 nsew default output
rlabel metal3 s 0 78752 800 78872 6 io_oeb[12]
port 254 nsew default output
rlabel metal3 s 0 85144 800 85264 6 io_oeb[13]
port 255 nsew default output
rlabel metal3 s 0 91400 800 91520 6 io_oeb[14]
port 256 nsew default output
rlabel metal3 s 0 97792 800 97912 6 io_oeb[15]
port 257 nsew default output
rlabel metal3 s 0 104048 800 104168 6 io_oeb[16]
port 258 nsew default output
rlabel metal3 s 0 110440 800 110560 6 io_oeb[17]
port 259 nsew default output
rlabel metal3 s 0 116696 800 116816 6 io_oeb[18]
port 260 nsew default output
rlabel metal3 s 0 122952 800 123072 6 io_oeb[19]
port 261 nsew default output
rlabel metal3 s 0 9256 800 9376 6 io_oeb[1]
port 262 nsew default output
rlabel metal3 s 0 129344 800 129464 6 io_oeb[20]
port 263 nsew default output
rlabel metal3 s 0 135600 800 135720 6 io_oeb[21]
port 264 nsew default output
rlabel metal3 s 0 141992 800 142112 6 io_oeb[22]
port 265 nsew default output
rlabel metal3 s 0 148248 800 148368 6 io_oeb[23]
port 266 nsew default output
rlabel metal3 s 0 154640 800 154760 6 io_oeb[24]
port 267 nsew default output
rlabel metal3 s 0 160896 800 161016 6 io_oeb[25]
port 268 nsew default output
rlabel metal3 s 0 167288 800 167408 6 io_oeb[26]
port 269 nsew default output
rlabel metal3 s 0 173544 800 173664 6 io_oeb[27]
port 270 nsew default output
rlabel metal3 s 0 179936 800 180056 6 io_oeb[28]
port 271 nsew default output
rlabel metal3 s 0 186192 800 186312 6 io_oeb[29]
port 272 nsew default output
rlabel metal3 s 0 15648 800 15768 6 io_oeb[2]
port 273 nsew default output
rlabel metal3 s 0 192448 800 192568 6 io_oeb[30]
port 274 nsew default output
rlabel metal3 s 0 198840 800 198960 6 io_oeb[31]
port 275 nsew default output
rlabel metal3 s 0 205096 800 205216 6 io_oeb[32]
port 276 nsew default output
rlabel metal3 s 0 211488 800 211608 6 io_oeb[33]
port 277 nsew default output
rlabel metal3 s 0 217744 800 217864 6 io_oeb[34]
port 278 nsew default output
rlabel metal3 s 0 224136 800 224256 6 io_oeb[35]
port 279 nsew default output
rlabel metal3 s 0 230392 800 230512 6 io_oeb[36]
port 280 nsew default output
rlabel metal3 s 0 236784 800 236904 6 io_oeb[37]
port 281 nsew default output
rlabel metal3 s 0 21904 800 22024 6 io_oeb[3]
port 282 nsew default output
rlabel metal3 s 0 28296 800 28416 6 io_oeb[4]
port 283 nsew default output
rlabel metal3 s 0 34552 800 34672 6 io_oeb[5]
port 284 nsew default output
rlabel metal3 s 0 40944 800 41064 6 io_oeb[6]
port 285 nsew default output
rlabel metal3 s 0 47200 800 47320 6 io_oeb[7]
port 286 nsew default output
rlabel metal3 s 0 53592 800 53712 6 io_oeb[8]
port 287 nsew default output
rlabel metal3 s 0 59848 800 59968 6 io_oeb[9]
port 288 nsew default output
rlabel metal3 s 0 5040 800 5160 6 io_out[0]
port 289 nsew default output
rlabel metal3 s 0 68280 800 68400 6 io_out[10]
port 290 nsew default output
rlabel metal3 s 0 74536 800 74656 6 io_out[11]
port 291 nsew default output
rlabel metal3 s 0 80928 800 81048 6 io_out[12]
port 292 nsew default output
rlabel metal3 s 0 87184 800 87304 6 io_out[13]
port 293 nsew default output
rlabel metal3 s 0 93576 800 93696 6 io_out[14]
port 294 nsew default output
rlabel metal3 s 0 99832 800 99952 6 io_out[15]
port 295 nsew default output
rlabel metal3 s 0 106224 800 106344 6 io_out[16]
port 296 nsew default output
rlabel metal3 s 0 112480 800 112600 6 io_out[17]
port 297 nsew default output
rlabel metal3 s 0 118872 800 118992 6 io_out[18]
port 298 nsew default output
rlabel metal3 s 0 125128 800 125248 6 io_out[19]
port 299 nsew default output
rlabel metal3 s 0 11432 800 11552 6 io_out[1]
port 300 nsew default output
rlabel metal3 s 0 131384 800 131504 6 io_out[20]
port 301 nsew default output
rlabel metal3 s 0 137776 800 137896 6 io_out[21]
port 302 nsew default output
rlabel metal3 s 0 144032 800 144152 6 io_out[22]
port 303 nsew default output
rlabel metal3 s 0 150424 800 150544 6 io_out[23]
port 304 nsew default output
rlabel metal3 s 0 156680 800 156800 6 io_out[24]
port 305 nsew default output
rlabel metal3 s 0 163072 800 163192 6 io_out[25]
port 306 nsew default output
rlabel metal3 s 0 169328 800 169448 6 io_out[26]
port 307 nsew default output
rlabel metal3 s 0 175720 800 175840 6 io_out[27]
port 308 nsew default output
rlabel metal3 s 0 181976 800 182096 6 io_out[28]
port 309 nsew default output
rlabel metal3 s 0 188232 800 188352 6 io_out[29]
port 310 nsew default output
rlabel metal3 s 0 17688 800 17808 6 io_out[2]
port 311 nsew default output
rlabel metal3 s 0 194624 800 194744 6 io_out[30]
port 312 nsew default output
rlabel metal3 s 0 200880 800 201000 6 io_out[31]
port 313 nsew default output
rlabel metal3 s 0 207272 800 207392 6 io_out[32]
port 314 nsew default output
rlabel metal3 s 0 213528 800 213648 6 io_out[33]
port 315 nsew default output
rlabel metal3 s 0 219920 800 220040 6 io_out[34]
port 316 nsew default output
rlabel metal3 s 0 226176 800 226296 6 io_out[35]
port 317 nsew default output
rlabel metal3 s 0 232568 800 232688 6 io_out[36]
port 318 nsew default output
rlabel metal3 s 0 238824 800 238944 6 io_out[37]
port 319 nsew default output
rlabel metal3 s 0 24080 800 24200 6 io_out[3]
port 320 nsew default output
rlabel metal3 s 0 30336 800 30456 6 io_out[4]
port 321 nsew default output
rlabel metal3 s 0 36728 800 36848 6 io_out[5]
port 322 nsew default output
rlabel metal3 s 0 42984 800 43104 6 io_out[6]
port 323 nsew default output
rlabel metal3 s 0 49376 800 49496 6 io_out[7]
port 324 nsew default output
rlabel metal3 s 0 55632 800 55752 6 io_out[8]
port 325 nsew default output
rlabel metal3 s 0 61888 800 62008 6 io_out[9]
port 326 nsew default output
rlabel metal2 s 207202 0 207258 800 6 la_data_in[0]
port 327 nsew default input
rlabel metal2 s 213090 0 213146 800 6 la_data_in[1]
port 328 nsew default input
rlabel metal2 s 209226 0 209282 800 6 la_data_out[0]
port 329 nsew default output
rlabel metal2 s 215022 0 215078 800 6 la_data_out[1]
port 330 nsew default output
rlabel metal2 s 218886 0 218942 800 6 la_data_out[2]
port 331 nsew default output
rlabel metal2 s 211158 0 211214 800 6 la_oen[0]
port 332 nsew default input
rlabel metal2 s 216954 0 217010 800 6 la_oen[1]
port 333 nsew default input
rlabel metal3 s 219200 3272 220000 3392 6 one
port 334 nsew default output
rlabel metal3 s 219200 238824 220000 238944 6 ram_ce
port 335 nsew default output
rlabel metal2 s 938 0 994 800 6 wb_clk_i
port 336 nsew default input
rlabel metal2 s 2870 0 2926 800 6 wb_rst_i
port 337 nsew default input
rlabel metal2 s 4802 0 4858 800 6 wbs_ack_o
port 338 nsew default output
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[0]
port 339 nsew default input
rlabel metal2 s 78770 0 78826 800 6 wbs_adr_i[10]
port 340 nsew default input
rlabel metal2 s 84566 0 84622 800 6 wbs_adr_i[11]
port 341 nsew default input
rlabel metal2 s 90454 0 90510 800 6 wbs_adr_i[12]
port 342 nsew default input
rlabel metal2 s 96250 0 96306 800 6 wbs_adr_i[13]
port 343 nsew default input
rlabel metal2 s 102138 0 102194 800 6 wbs_adr_i[14]
port 344 nsew default input
rlabel metal2 s 107934 0 107990 800 6 wbs_adr_i[15]
port 345 nsew default input
rlabel metal2 s 113822 0 113878 800 6 wbs_adr_i[16]
port 346 nsew default input
rlabel metal2 s 119618 0 119674 800 6 wbs_adr_i[17]
port 347 nsew default input
rlabel metal2 s 125506 0 125562 800 6 wbs_adr_i[18]
port 348 nsew default input
rlabel metal2 s 131302 0 131358 800 6 wbs_adr_i[19]
port 349 nsew default input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[1]
port 350 nsew default input
rlabel metal2 s 137190 0 137246 800 6 wbs_adr_i[20]
port 351 nsew default input
rlabel metal2 s 142986 0 143042 800 6 wbs_adr_i[21]
port 352 nsew default input
rlabel metal2 s 148874 0 148930 800 6 wbs_adr_i[22]
port 353 nsew default input
rlabel metal2 s 154670 0 154726 800 6 wbs_adr_i[23]
port 354 nsew default input
rlabel metal2 s 160558 0 160614 800 6 wbs_adr_i[24]
port 355 nsew default input
rlabel metal2 s 166354 0 166410 800 6 wbs_adr_i[25]
port 356 nsew default input
rlabel metal2 s 172242 0 172298 800 6 wbs_adr_i[26]
port 357 nsew default input
rlabel metal2 s 178038 0 178094 800 6 wbs_adr_i[27]
port 358 nsew default input
rlabel metal2 s 183834 0 183890 800 6 wbs_adr_i[28]
port 359 nsew default input
rlabel metal2 s 189722 0 189778 800 6 wbs_adr_i[29]
port 360 nsew default input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[2]
port 361 nsew default input
rlabel metal2 s 195518 0 195574 800 6 wbs_adr_i[30]
port 362 nsew default input
rlabel metal2 s 201406 0 201462 800 6 wbs_adr_i[31]
port 363 nsew default input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[3]
port 364 nsew default input
rlabel metal2 s 43718 0 43774 800 6 wbs_adr_i[4]
port 365 nsew default input
rlabel metal2 s 49514 0 49570 800 6 wbs_adr_i[5]
port 366 nsew default input
rlabel metal2 s 55402 0 55458 800 6 wbs_adr_i[6]
port 367 nsew default input
rlabel metal2 s 61198 0 61254 800 6 wbs_adr_i[7]
port 368 nsew default input
rlabel metal2 s 67086 0 67142 800 6 wbs_adr_i[8]
port 369 nsew default input
rlabel metal2 s 72882 0 72938 800 6 wbs_adr_i[9]
port 370 nsew default input
rlabel metal2 s 6734 0 6790 800 6 wbs_cyc_i
port 371 nsew default input
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_i[0]
port 372 nsew default input
rlabel metal2 s 80702 0 80758 800 6 wbs_dat_i[10]
port 373 nsew default input
rlabel metal2 s 86590 0 86646 800 6 wbs_dat_i[11]
port 374 nsew default input
rlabel metal2 s 92386 0 92442 800 6 wbs_dat_i[12]
port 375 nsew default input
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_i[13]
port 376 nsew default input
rlabel metal2 s 104070 0 104126 800 6 wbs_dat_i[14]
port 377 nsew default input
rlabel metal2 s 109866 0 109922 800 6 wbs_dat_i[15]
port 378 nsew default input
rlabel metal2 s 115754 0 115810 800 6 wbs_dat_i[16]
port 379 nsew default input
rlabel metal2 s 121550 0 121606 800 6 wbs_dat_i[17]
port 380 nsew default input
rlabel metal2 s 127438 0 127494 800 6 wbs_dat_i[18]
port 381 nsew default input
rlabel metal2 s 133234 0 133290 800 6 wbs_dat_i[19]
port 382 nsew default input
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_i[1]
port 383 nsew default input
rlabel metal2 s 139122 0 139178 800 6 wbs_dat_i[20]
port 384 nsew default input
rlabel metal2 s 144918 0 144974 800 6 wbs_dat_i[21]
port 385 nsew default input
rlabel metal2 s 150806 0 150862 800 6 wbs_dat_i[22]
port 386 nsew default input
rlabel metal2 s 156602 0 156658 800 6 wbs_dat_i[23]
port 387 nsew default input
rlabel metal2 s 162490 0 162546 800 6 wbs_dat_i[24]
port 388 nsew default input
rlabel metal2 s 168286 0 168342 800 6 wbs_dat_i[25]
port 389 nsew default input
rlabel metal2 s 174174 0 174230 800 6 wbs_dat_i[26]
port 390 nsew default input
rlabel metal2 s 179970 0 180026 800 6 wbs_dat_i[27]
port 391 nsew default input
rlabel metal2 s 185858 0 185914 800 6 wbs_dat_i[28]
port 392 nsew default input
rlabel metal2 s 191654 0 191710 800 6 wbs_dat_i[29]
port 393 nsew default input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[2]
port 394 nsew default input
rlabel metal2 s 197542 0 197598 800 6 wbs_dat_i[30]
port 395 nsew default input
rlabel metal2 s 203338 0 203394 800 6 wbs_dat_i[31]
port 396 nsew default input
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_i[3]
port 397 nsew default input
rlabel metal2 s 45650 0 45706 800 6 wbs_dat_i[4]
port 398 nsew default input
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_i[5]
port 399 nsew default input
rlabel metal2 s 57334 0 57390 800 6 wbs_dat_i[6]
port 400 nsew default input
rlabel metal2 s 63222 0 63278 800 6 wbs_dat_i[7]
port 401 nsew default input
rlabel metal2 s 69018 0 69074 800 6 wbs_dat_i[8]
port 402 nsew default input
rlabel metal2 s 74906 0 74962 800 6 wbs_dat_i[9]
port 403 nsew default input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[0]
port 404 nsew default output
rlabel metal2 s 82634 0 82690 800 6 wbs_dat_o[10]
port 405 nsew default output
rlabel metal2 s 88522 0 88578 800 6 wbs_dat_o[11]
port 406 nsew default output
rlabel metal2 s 94318 0 94374 800 6 wbs_dat_o[12]
port 407 nsew default output
rlabel metal2 s 100206 0 100262 800 6 wbs_dat_o[13]
port 408 nsew default output
rlabel metal2 s 106002 0 106058 800 6 wbs_dat_o[14]
port 409 nsew default output
rlabel metal2 s 111890 0 111946 800 6 wbs_dat_o[15]
port 410 nsew default output
rlabel metal2 s 117686 0 117742 800 6 wbs_dat_o[16]
port 411 nsew default output
rlabel metal2 s 123574 0 123630 800 6 wbs_dat_o[17]
port 412 nsew default output
rlabel metal2 s 129370 0 129426 800 6 wbs_dat_o[18]
port 413 nsew default output
rlabel metal2 s 135166 0 135222 800 6 wbs_dat_o[19]
port 414 nsew default output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[1]
port 415 nsew default output
rlabel metal2 s 141054 0 141110 800 6 wbs_dat_o[20]
port 416 nsew default output
rlabel metal2 s 146850 0 146906 800 6 wbs_dat_o[21]
port 417 nsew default output
rlabel metal2 s 152738 0 152794 800 6 wbs_dat_o[22]
port 418 nsew default output
rlabel metal2 s 158534 0 158590 800 6 wbs_dat_o[23]
port 419 nsew default output
rlabel metal2 s 164422 0 164478 800 6 wbs_dat_o[24]
port 420 nsew default output
rlabel metal2 s 170218 0 170274 800 6 wbs_dat_o[25]
port 421 nsew default output
rlabel metal2 s 176106 0 176162 800 6 wbs_dat_o[26]
port 422 nsew default output
rlabel metal2 s 181902 0 181958 800 6 wbs_dat_o[27]
port 423 nsew default output
rlabel metal2 s 187790 0 187846 800 6 wbs_dat_o[28]
port 424 nsew default output
rlabel metal2 s 193586 0 193642 800 6 wbs_dat_o[29]
port 425 nsew default output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[2]
port 426 nsew default output
rlabel metal2 s 199474 0 199530 800 6 wbs_dat_o[30]
port 427 nsew default output
rlabel metal2 s 205270 0 205326 800 6 wbs_dat_o[31]
port 428 nsew default output
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_o[3]
port 429 nsew default output
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_o[4]
port 430 nsew default output
rlabel metal2 s 53470 0 53526 800 6 wbs_dat_o[5]
port 431 nsew default output
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_o[6]
port 432 nsew default output
rlabel metal2 s 65154 0 65210 800 6 wbs_dat_o[7]
port 433 nsew default output
rlabel metal2 s 70950 0 71006 800 6 wbs_dat_o[8]
port 434 nsew default output
rlabel metal2 s 76838 0 76894 800 6 wbs_dat_o[9]
port 435 nsew default output
rlabel metal2 s 18418 0 18474 800 6 wbs_sel_i[0]
port 436 nsew default input
rlabel metal2 s 26238 0 26294 800 6 wbs_sel_i[1]
port 437 nsew default input
rlabel metal2 s 33966 0 34022 800 6 wbs_sel_i[2]
port 438 nsew default input
rlabel metal2 s 41786 0 41842 800 6 wbs_sel_i[3]
port 439 nsew default input
rlabel metal2 s 8666 0 8722 800 6 wbs_stb_i
port 440 nsew default input
rlabel metal2 s 10598 0 10654 800 6 wbs_we_i
port 441 nsew default input
rlabel metal3 s 219200 1096 220000 1216 6 zero
port 442 nsew default output
rlabel metal4 s 4208 2128 4528 237776 6 VPWR
port 443 nsew power input
rlabel metal4 s 19568 2128 19888 237776 6 VGND
port 444 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 220000 240000
string LEFview TRUE
<< end >>
