VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hs32_core1
  CLASS BLOCK ;
  FOREIGN hs32_core1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1400.000 BY 1200.000 ;
  PIN cpu_addr_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END cpu_addr_e[0]
  PIN cpu_addr_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 673.530 0.000 673.810 4.000 ;
    END
  END cpu_addr_e[10]
  PIN cpu_addr_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 686.410 0.000 686.690 4.000 ;
    END
  END cpu_addr_e[11]
  PIN cpu_addr_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END cpu_addr_e[12]
  PIN cpu_addr_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END cpu_addr_e[13]
  PIN cpu_addr_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END cpu_addr_e[14]
  PIN cpu_addr_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 737.930 0.000 738.210 4.000 ;
    END
  END cpu_addr_e[15]
  PIN cpu_addr_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.070 0.000 558.350 4.000 ;
    END
  END cpu_addr_e[1]
  PIN cpu_addr_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END cpu_addr_e[2]
  PIN cpu_addr_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END cpu_addr_e[3]
  PIN cpu_addr_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END cpu_addr_e[4]
  PIN cpu_addr_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END cpu_addr_e[5]
  PIN cpu_addr_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END cpu_addr_e[6]
  PIN cpu_addr_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 4.000 ;
    END
  END cpu_addr_e[7]
  PIN cpu_addr_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 647.770 0.000 648.050 4.000 ;
    END
  END cpu_addr_e[8]
  PIN cpu_addr_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END cpu_addr_e[9]
  PIN cpu_addr_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 545.190 1196.000 545.470 1200.000 ;
    END
  END cpu_addr_n[0]
  PIN cpu_addr_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 673.530 1196.000 673.810 1200.000 ;
    END
  END cpu_addr_n[10]
  PIN cpu_addr_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 686.410 1196.000 686.690 1200.000 ;
    END
  END cpu_addr_n[11]
  PIN cpu_addr_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 699.290 1196.000 699.570 1200.000 ;
    END
  END cpu_addr_n[12]
  PIN cpu_addr_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 712.170 1196.000 712.450 1200.000 ;
    END
  END cpu_addr_n[13]
  PIN cpu_addr_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 725.050 1196.000 725.330 1200.000 ;
    END
  END cpu_addr_n[14]
  PIN cpu_addr_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 737.930 1196.000 738.210 1200.000 ;
    END
  END cpu_addr_n[15]
  PIN cpu_addr_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.070 1196.000 558.350 1200.000 ;
    END
  END cpu_addr_n[1]
  PIN cpu_addr_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.950 1196.000 571.230 1200.000 ;
    END
  END cpu_addr_n[2]
  PIN cpu_addr_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 583.830 1196.000 584.110 1200.000 ;
    END
  END cpu_addr_n[3]
  PIN cpu_addr_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 596.710 1196.000 596.990 1200.000 ;
    END
  END cpu_addr_n[4]
  PIN cpu_addr_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 609.590 1196.000 609.870 1200.000 ;
    END
  END cpu_addr_n[5]
  PIN cpu_addr_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 622.470 1196.000 622.750 1200.000 ;
    END
  END cpu_addr_n[6]
  PIN cpu_addr_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 634.890 1196.000 635.170 1200.000 ;
    END
  END cpu_addr_n[7]
  PIN cpu_addr_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 647.770 1196.000 648.050 1200.000 ;
    END
  END cpu_addr_n[8]
  PIN cpu_addr_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 660.650 1196.000 660.930 1200.000 ;
    END
  END cpu_addr_n[9]
  PIN cpu_dtr_e0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END cpu_dtr_e0[0]
  PIN cpu_dtr_e0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END cpu_dtr_e0[10]
  PIN cpu_dtr_e0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END cpu_dtr_e0[11]
  PIN cpu_dtr_e0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END cpu_dtr_e0[12]
  PIN cpu_dtr_e0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END cpu_dtr_e0[13]
  PIN cpu_dtr_e0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END cpu_dtr_e0[14]
  PIN cpu_dtr_e0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END cpu_dtr_e0[15]
  PIN cpu_dtr_e0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END cpu_dtr_e0[16]
  PIN cpu_dtr_e0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END cpu_dtr_e0[17]
  PIN cpu_dtr_e0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END cpu_dtr_e0[18]
  PIN cpu_dtr_e0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END cpu_dtr_e0[19]
  PIN cpu_dtr_e0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END cpu_dtr_e0[1]
  PIN cpu_dtr_e0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END cpu_dtr_e0[20]
  PIN cpu_dtr_e0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END cpu_dtr_e0[21]
  PIN cpu_dtr_e0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END cpu_dtr_e0[22]
  PIN cpu_dtr_e0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END cpu_dtr_e0[23]
  PIN cpu_dtr_e0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END cpu_dtr_e0[24]
  PIN cpu_dtr_e0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END cpu_dtr_e0[25]
  PIN cpu_dtr_e0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END cpu_dtr_e0[26]
  PIN cpu_dtr_e0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END cpu_dtr_e0[27]
  PIN cpu_dtr_e0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END cpu_dtr_e0[28]
  PIN cpu_dtr_e0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END cpu_dtr_e0[29]
  PIN cpu_dtr_e0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END cpu_dtr_e0[2]
  PIN cpu_dtr_e0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END cpu_dtr_e0[30]
  PIN cpu_dtr_e0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END cpu_dtr_e0[31]
  PIN cpu_dtr_e0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END cpu_dtr_e0[3]
  PIN cpu_dtr_e0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END cpu_dtr_e0[4]
  PIN cpu_dtr_e0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END cpu_dtr_e0[5]
  PIN cpu_dtr_e0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END cpu_dtr_e0[6]
  PIN cpu_dtr_e0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END cpu_dtr_e0[7]
  PIN cpu_dtr_e0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END cpu_dtr_e0[8]
  PIN cpu_dtr_e0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END cpu_dtr_e0[9]
  PIN cpu_dtr_e1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 994.610 0.000 994.890 4.000 ;
    END
  END cpu_dtr_e1[0]
  PIN cpu_dtr_e1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1122.950 0.000 1123.230 4.000 ;
    END
  END cpu_dtr_e1[10]
  PIN cpu_dtr_e1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1135.830 0.000 1136.110 4.000 ;
    END
  END cpu_dtr_e1[11]
  PIN cpu_dtr_e1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1148.710 0.000 1148.990 4.000 ;
    END
  END cpu_dtr_e1[12]
  PIN cpu_dtr_e1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1161.590 0.000 1161.870 4.000 ;
    END
  END cpu_dtr_e1[13]
  PIN cpu_dtr_e1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1174.470 0.000 1174.750 4.000 ;
    END
  END cpu_dtr_e1[14]
  PIN cpu_dtr_e1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1187.350 0.000 1187.630 4.000 ;
    END
  END cpu_dtr_e1[15]
  PIN cpu_dtr_e1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1200.230 0.000 1200.510 4.000 ;
    END
  END cpu_dtr_e1[16]
  PIN cpu_dtr_e1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1213.110 0.000 1213.390 4.000 ;
    END
  END cpu_dtr_e1[17]
  PIN cpu_dtr_e1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1225.990 0.000 1226.270 4.000 ;
    END
  END cpu_dtr_e1[18]
  PIN cpu_dtr_e1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1238.870 0.000 1239.150 4.000 ;
    END
  END cpu_dtr_e1[19]
  PIN cpu_dtr_e1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.490 0.000 1007.770 4.000 ;
    END
  END cpu_dtr_e1[1]
  PIN cpu_dtr_e1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.290 0.000 1251.570 4.000 ;
    END
  END cpu_dtr_e1[20]
  PIN cpu_dtr_e1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1264.170 0.000 1264.450 4.000 ;
    END
  END cpu_dtr_e1[21]
  PIN cpu_dtr_e1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.050 0.000 1277.330 4.000 ;
    END
  END cpu_dtr_e1[22]
  PIN cpu_dtr_e1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1289.930 0.000 1290.210 4.000 ;
    END
  END cpu_dtr_e1[23]
  PIN cpu_dtr_e1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1302.810 0.000 1303.090 4.000 ;
    END
  END cpu_dtr_e1[24]
  PIN cpu_dtr_e1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1315.690 0.000 1315.970 4.000 ;
    END
  END cpu_dtr_e1[25]
  PIN cpu_dtr_e1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.570 0.000 1328.850 4.000 ;
    END
  END cpu_dtr_e1[26]
  PIN cpu_dtr_e1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1341.450 0.000 1341.730 4.000 ;
    END
  END cpu_dtr_e1[27]
  PIN cpu_dtr_e1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1354.330 0.000 1354.610 4.000 ;
    END
  END cpu_dtr_e1[28]
  PIN cpu_dtr_e1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1367.210 0.000 1367.490 4.000 ;
    END
  END cpu_dtr_e1[29]
  PIN cpu_dtr_e1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.370 0.000 1020.650 4.000 ;
    END
  END cpu_dtr_e1[2]
  PIN cpu_dtr_e1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1380.090 0.000 1380.370 4.000 ;
    END
  END cpu_dtr_e1[30]
  PIN cpu_dtr_e1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1392.970 0.000 1393.250 4.000 ;
    END
  END cpu_dtr_e1[31]
  PIN cpu_dtr_e1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1033.250 0.000 1033.530 4.000 ;
    END
  END cpu_dtr_e1[3]
  PIN cpu_dtr_e1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END cpu_dtr_e1[4]
  PIN cpu_dtr_e1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1059.010 0.000 1059.290 4.000 ;
    END
  END cpu_dtr_e1[5]
  PIN cpu_dtr_e1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1071.890 0.000 1072.170 4.000 ;
    END
  END cpu_dtr_e1[6]
  PIN cpu_dtr_e1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1084.770 0.000 1085.050 4.000 ;
    END
  END cpu_dtr_e1[7]
  PIN cpu_dtr_e1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.190 0.000 1097.470 4.000 ;
    END
  END cpu_dtr_e1[8]
  PIN cpu_dtr_e1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.070 0.000 1110.350 4.000 ;
    END
  END cpu_dtr_e1[9]
  PIN cpu_dtr_n0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 1196.000 31.650 1200.000 ;
    END
  END cpu_dtr_n0[0]
  PIN cpu_dtr_n0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.170 1196.000 160.450 1200.000 ;
    END
  END cpu_dtr_n0[10]
  PIN cpu_dtr_n0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.590 1196.000 172.870 1200.000 ;
    END
  END cpu_dtr_n0[11]
  PIN cpu_dtr_n0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.470 1196.000 185.750 1200.000 ;
    END
  END cpu_dtr_n0[12]
  PIN cpu_dtr_n0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 198.350 1196.000 198.630 1200.000 ;
    END
  END cpu_dtr_n0[13]
  PIN cpu_dtr_n0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.230 1196.000 211.510 1200.000 ;
    END
  END cpu_dtr_n0[14]
  PIN cpu_dtr_n0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.110 1196.000 224.390 1200.000 ;
    END
  END cpu_dtr_n0[15]
  PIN cpu_dtr_n0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.990 1196.000 237.270 1200.000 ;
    END
  END cpu_dtr_n0[16]
  PIN cpu_dtr_n0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 249.870 1196.000 250.150 1200.000 ;
    END
  END cpu_dtr_n0[17]
  PIN cpu_dtr_n0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 262.750 1196.000 263.030 1200.000 ;
    END
  END cpu_dtr_n0[18]
  PIN cpu_dtr_n0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.630 1196.000 275.910 1200.000 ;
    END
  END cpu_dtr_n0[19]
  PIN cpu_dtr_n0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 1196.000 44.530 1200.000 ;
    END
  END cpu_dtr_n0[1]
  PIN cpu_dtr_n0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.510 1196.000 288.790 1200.000 ;
    END
  END cpu_dtr_n0[20]
  PIN cpu_dtr_n0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.390 1196.000 301.670 1200.000 ;
    END
  END cpu_dtr_n0[21]
  PIN cpu_dtr_n0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 314.270 1196.000 314.550 1200.000 ;
    END
  END cpu_dtr_n0[22]
  PIN cpu_dtr_n0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 326.690 1196.000 326.970 1200.000 ;
    END
  END cpu_dtr_n0[23]
  PIN cpu_dtr_n0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 339.570 1196.000 339.850 1200.000 ;
    END
  END cpu_dtr_n0[24]
  PIN cpu_dtr_n0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 352.450 1196.000 352.730 1200.000 ;
    END
  END cpu_dtr_n0[25]
  PIN cpu_dtr_n0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.330 1196.000 365.610 1200.000 ;
    END
  END cpu_dtr_n0[26]
  PIN cpu_dtr_n0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 378.210 1196.000 378.490 1200.000 ;
    END
  END cpu_dtr_n0[27]
  PIN cpu_dtr_n0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 391.090 1196.000 391.370 1200.000 ;
    END
  END cpu_dtr_n0[28]
  PIN cpu_dtr_n0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.970 1196.000 404.250 1200.000 ;
    END
  END cpu_dtr_n0[29]
  PIN cpu_dtr_n0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 1196.000 57.410 1200.000 ;
    END
  END cpu_dtr_n0[2]
  PIN cpu_dtr_n0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 416.850 1196.000 417.130 1200.000 ;
    END
  END cpu_dtr_n0[30]
  PIN cpu_dtr_n0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 429.730 1196.000 430.010 1200.000 ;
    END
  END cpu_dtr_n0[31]
  PIN cpu_dtr_n0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.010 1196.000 70.290 1200.000 ;
    END
  END cpu_dtr_n0[3]
  PIN cpu_dtr_n0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.890 1196.000 83.170 1200.000 ;
    END
  END cpu_dtr_n0[4]
  PIN cpu_dtr_n0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.770 1196.000 96.050 1200.000 ;
    END
  END cpu_dtr_n0[5]
  PIN cpu_dtr_n0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.650 1196.000 108.930 1200.000 ;
    END
  END cpu_dtr_n0[6]
  PIN cpu_dtr_n0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.530 1196.000 121.810 1200.000 ;
    END
  END cpu_dtr_n0[7]
  PIN cpu_dtr_n0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.410 1196.000 134.690 1200.000 ;
    END
  END cpu_dtr_n0[8]
  PIN cpu_dtr_n0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 147.290 1196.000 147.570 1200.000 ;
    END
  END cpu_dtr_n0[9]
  PIN cpu_dtr_n1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 994.610 1196.000 994.890 1200.000 ;
    END
  END cpu_dtr_n1[0]
  PIN cpu_dtr_n1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1122.950 1196.000 1123.230 1200.000 ;
    END
  END cpu_dtr_n1[10]
  PIN cpu_dtr_n1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1135.830 1196.000 1136.110 1200.000 ;
    END
  END cpu_dtr_n1[11]
  PIN cpu_dtr_n1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1148.710 1196.000 1148.990 1200.000 ;
    END
  END cpu_dtr_n1[12]
  PIN cpu_dtr_n1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1161.590 1196.000 1161.870 1200.000 ;
    END
  END cpu_dtr_n1[13]
  PIN cpu_dtr_n1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1174.470 1196.000 1174.750 1200.000 ;
    END
  END cpu_dtr_n1[14]
  PIN cpu_dtr_n1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1187.350 1196.000 1187.630 1200.000 ;
    END
  END cpu_dtr_n1[15]
  PIN cpu_dtr_n1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1200.230 1196.000 1200.510 1200.000 ;
    END
  END cpu_dtr_n1[16]
  PIN cpu_dtr_n1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1213.110 1196.000 1213.390 1200.000 ;
    END
  END cpu_dtr_n1[17]
  PIN cpu_dtr_n1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1225.990 1196.000 1226.270 1200.000 ;
    END
  END cpu_dtr_n1[18]
  PIN cpu_dtr_n1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1238.870 1196.000 1239.150 1200.000 ;
    END
  END cpu_dtr_n1[19]
  PIN cpu_dtr_n1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.490 1196.000 1007.770 1200.000 ;
    END
  END cpu_dtr_n1[1]
  PIN cpu_dtr_n1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.290 1196.000 1251.570 1200.000 ;
    END
  END cpu_dtr_n1[20]
  PIN cpu_dtr_n1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1264.170 1196.000 1264.450 1200.000 ;
    END
  END cpu_dtr_n1[21]
  PIN cpu_dtr_n1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.050 1196.000 1277.330 1200.000 ;
    END
  END cpu_dtr_n1[22]
  PIN cpu_dtr_n1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1289.930 1196.000 1290.210 1200.000 ;
    END
  END cpu_dtr_n1[23]
  PIN cpu_dtr_n1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1302.810 1196.000 1303.090 1200.000 ;
    END
  END cpu_dtr_n1[24]
  PIN cpu_dtr_n1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1315.690 1196.000 1315.970 1200.000 ;
    END
  END cpu_dtr_n1[25]
  PIN cpu_dtr_n1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.570 1196.000 1328.850 1200.000 ;
    END
  END cpu_dtr_n1[26]
  PIN cpu_dtr_n1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1341.450 1196.000 1341.730 1200.000 ;
    END
  END cpu_dtr_n1[27]
  PIN cpu_dtr_n1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1354.330 1196.000 1354.610 1200.000 ;
    END
  END cpu_dtr_n1[28]
  PIN cpu_dtr_n1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1367.210 1196.000 1367.490 1200.000 ;
    END
  END cpu_dtr_n1[29]
  PIN cpu_dtr_n1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.370 1196.000 1020.650 1200.000 ;
    END
  END cpu_dtr_n1[2]
  PIN cpu_dtr_n1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1380.090 1196.000 1380.370 1200.000 ;
    END
  END cpu_dtr_n1[30]
  PIN cpu_dtr_n1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1392.970 1196.000 1393.250 1200.000 ;
    END
  END cpu_dtr_n1[31]
  PIN cpu_dtr_n1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1033.250 1196.000 1033.530 1200.000 ;
    END
  END cpu_dtr_n1[3]
  PIN cpu_dtr_n1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1046.130 1196.000 1046.410 1200.000 ;
    END
  END cpu_dtr_n1[4]
  PIN cpu_dtr_n1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1059.010 1196.000 1059.290 1200.000 ;
    END
  END cpu_dtr_n1[5]
  PIN cpu_dtr_n1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1071.890 1196.000 1072.170 1200.000 ;
    END
  END cpu_dtr_n1[6]
  PIN cpu_dtr_n1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1084.770 1196.000 1085.050 1200.000 ;
    END
  END cpu_dtr_n1[7]
  PIN cpu_dtr_n1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.190 1196.000 1097.470 1200.000 ;
    END
  END cpu_dtr_n1[8]
  PIN cpu_dtr_n1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.070 1196.000 1110.350 1200.000 ;
    END
  END cpu_dtr_n1[9]
  PIN cpu_dtw_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END cpu_dtw_e[0]
  PIN cpu_dtw_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END cpu_dtw_e[10]
  PIN cpu_dtw_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 930.670 0.000 930.950 4.000 ;
    END
  END cpu_dtw_e[11]
  PIN cpu_dtw_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 943.090 0.000 943.370 4.000 ;
    END
  END cpu_dtw_e[12]
  PIN cpu_dtw_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 955.970 0.000 956.250 4.000 ;
    END
  END cpu_dtw_e[13]
  PIN cpu_dtw_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 968.850 0.000 969.130 4.000 ;
    END
  END cpu_dtw_e[14]
  PIN cpu_dtw_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 981.730 0.000 982.010 4.000 ;
    END
  END cpu_dtw_e[15]
  PIN cpu_dtw_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END cpu_dtw_e[1]
  PIN cpu_dtw_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END cpu_dtw_e[2]
  PIN cpu_dtw_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END cpu_dtw_e[3]
  PIN cpu_dtw_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END cpu_dtw_e[4]
  PIN cpu_dtw_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END cpu_dtw_e[5]
  PIN cpu_dtw_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END cpu_dtw_e[6]
  PIN cpu_dtw_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END cpu_dtw_e[7]
  PIN cpu_dtw_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END cpu_dtw_e[8]
  PIN cpu_dtw_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END cpu_dtw_e[9]
  PIN cpu_dtw_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 788.990 1196.000 789.270 1200.000 ;
    END
  END cpu_dtw_n[0]
  PIN cpu_dtw_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 917.790 1196.000 918.070 1200.000 ;
    END
  END cpu_dtw_n[10]
  PIN cpu_dtw_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 930.670 1196.000 930.950 1200.000 ;
    END
  END cpu_dtw_n[11]
  PIN cpu_dtw_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 943.090 1196.000 943.370 1200.000 ;
    END
  END cpu_dtw_n[12]
  PIN cpu_dtw_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 955.970 1196.000 956.250 1200.000 ;
    END
  END cpu_dtw_n[13]
  PIN cpu_dtw_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 968.850 1196.000 969.130 1200.000 ;
    END
  END cpu_dtw_n[14]
  PIN cpu_dtw_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 981.730 1196.000 982.010 1200.000 ;
    END
  END cpu_dtw_n[15]
  PIN cpu_dtw_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 801.870 1196.000 802.150 1200.000 ;
    END
  END cpu_dtw_n[1]
  PIN cpu_dtw_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 814.750 1196.000 815.030 1200.000 ;
    END
  END cpu_dtw_n[2]
  PIN cpu_dtw_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 827.630 1196.000 827.910 1200.000 ;
    END
  END cpu_dtw_n[3]
  PIN cpu_dtw_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 840.510 1196.000 840.790 1200.000 ;
    END
  END cpu_dtw_n[4]
  PIN cpu_dtw_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 853.390 1196.000 853.670 1200.000 ;
    END
  END cpu_dtw_n[5]
  PIN cpu_dtw_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 866.270 1196.000 866.550 1200.000 ;
    END
  END cpu_dtw_n[6]
  PIN cpu_dtw_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 879.150 1196.000 879.430 1200.000 ;
    END
  END cpu_dtw_n[7]
  PIN cpu_dtw_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 892.030 1196.000 892.310 1200.000 ;
    END
  END cpu_dtw_n[8]
  PIN cpu_dtw_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 904.910 1196.000 905.190 1200.000 ;
    END
  END cpu_dtw_n[9]
  PIN cpu_mask_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END cpu_mask_e[0]
  PIN cpu_mask_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END cpu_mask_e[1]
  PIN cpu_mask_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END cpu_mask_e[2]
  PIN cpu_mask_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END cpu_mask_e[3]
  PIN cpu_mask_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 493.670 0.000 493.950 4.000 ;
    END
  END cpu_mask_e[4]
  PIN cpu_mask_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 4.000 ;
    END
  END cpu_mask_e[5]
  PIN cpu_mask_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END cpu_mask_e[6]
  PIN cpu_mask_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END cpu_mask_e[7]
  PIN cpu_mask_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 442.610 1196.000 442.890 1200.000 ;
    END
  END cpu_mask_n[0]
  PIN cpu_mask_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.490 1196.000 455.770 1200.000 ;
    END
  END cpu_mask_n[1]
  PIN cpu_mask_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 468.370 1196.000 468.650 1200.000 ;
    END
  END cpu_mask_n[2]
  PIN cpu_mask_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 480.790 1196.000 481.070 1200.000 ;
    END
  END cpu_mask_n[3]
  PIN cpu_mask_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 493.670 1196.000 493.950 1200.000 ;
    END
  END cpu_mask_n[4]
  PIN cpu_mask_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 506.550 1196.000 506.830 1200.000 ;
    END
  END cpu_mask_n[5]
  PIN cpu_mask_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.430 1196.000 519.710 1200.000 ;
    END
  END cpu_mask_n[6]
  PIN cpu_mask_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 532.310 1196.000 532.590 1200.000 ;
    END
  END cpu_mask_n[7]
  PIN cpu_wen_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END cpu_wen_e[0]
  PIN cpu_wen_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END cpu_wen_e[1]
  PIN cpu_wen_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.690 1196.000 763.970 1200.000 ;
    END
  END cpu_wen_n[0]
  PIN cpu_wen_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 776.570 1196.000 776.850 1200.000 ;
    END
  END cpu_wen_n[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 4.800 1400.000 5.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 320.320 1400.000 320.920 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 351.600 1400.000 352.200 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 383.560 1400.000 384.160 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 414.840 1400.000 415.440 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 446.800 1400.000 447.400 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 478.080 1400.000 478.680 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 510.040 1400.000 510.640 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 541.320 1400.000 541.920 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 573.280 1400.000 573.880 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 604.560 1400.000 605.160 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 36.080 1400.000 36.680 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 635.840 1400.000 636.440 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 667.800 1400.000 668.400 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 699.080 1400.000 699.680 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 731.040 1400.000 731.640 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 762.320 1400.000 762.920 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 794.280 1400.000 794.880 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 825.560 1400.000 826.160 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 857.520 1400.000 858.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 888.800 1400.000 889.400 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 920.080 1400.000 920.680 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 67.360 1400.000 67.960 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 952.040 1400.000 952.640 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 983.320 1400.000 983.920 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1015.280 1400.000 1015.880 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1046.560 1400.000 1047.160 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1078.520 1400.000 1079.120 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1109.800 1400.000 1110.400 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1141.760 1400.000 1142.360 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1173.040 1400.000 1173.640 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 99.320 1400.000 99.920 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 130.600 1400.000 131.200 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 162.560 1400.000 163.160 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 193.840 1400.000 194.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 225.800 1400.000 226.400 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 257.080 1400.000 257.680 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1396.000 289.040 1400.000 289.640 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 15.000 1400.000 15.600 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 330.520 1400.000 331.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 362.480 1400.000 363.080 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 393.760 1400.000 394.360 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 425.720 1400.000 426.320 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 457.000 1400.000 457.600 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 488.960 1400.000 489.560 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 520.240 1400.000 520.840 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 552.200 1400.000 552.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 583.480 1400.000 584.080 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 614.760 1400.000 615.360 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 46.280 1400.000 46.880 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 646.720 1400.000 647.320 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 678.000 1400.000 678.600 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 709.960 1400.000 710.560 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 741.240 1400.000 741.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 773.200 1400.000 773.800 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 804.480 1400.000 805.080 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 836.440 1400.000 837.040 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 867.720 1400.000 868.320 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 899.680 1400.000 900.280 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 930.960 1400.000 931.560 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 78.240 1400.000 78.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 962.240 1400.000 962.840 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 994.200 1400.000 994.800 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1025.480 1400.000 1026.080 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1057.440 1400.000 1058.040 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1088.720 1400.000 1089.320 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1120.680 1400.000 1121.280 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1151.960 1400.000 1152.560 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1183.920 1400.000 1184.520 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 109.520 1400.000 110.120 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 141.480 1400.000 142.080 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 172.760 1400.000 173.360 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 204.720 1400.000 205.320 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 236.000 1400.000 236.600 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 267.960 1400.000 268.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 299.240 1400.000 299.840 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 25.200 1400.000 25.800 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 341.400 1400.000 342.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 372.680 1400.000 373.280 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 404.640 1400.000 405.240 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 435.920 1400.000 436.520 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 467.880 1400.000 468.480 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 499.160 1400.000 499.760 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 531.120 1400.000 531.720 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 562.400 1400.000 563.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 594.360 1400.000 594.960 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 625.640 1400.000 626.240 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 57.160 1400.000 57.760 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 656.920 1400.000 657.520 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 688.880 1400.000 689.480 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 720.160 1400.000 720.760 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 752.120 1400.000 752.720 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 783.400 1400.000 784.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 815.360 1400.000 815.960 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 846.640 1400.000 847.240 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 878.600 1400.000 879.200 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 909.880 1400.000 910.480 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 941.160 1400.000 941.760 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 88.440 1400.000 89.040 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 973.120 1400.000 973.720 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1004.400 1400.000 1005.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1036.360 1400.000 1036.960 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1067.640 1400.000 1068.240 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1099.600 1400.000 1100.200 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1130.880 1400.000 1131.480 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1162.840 1400.000 1163.440 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 1194.120 1400.000 1194.720 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 120.400 1400.000 121.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 151.680 1400.000 152.280 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 183.640 1400.000 184.240 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 214.920 1400.000 215.520 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 246.880 1400.000 247.480 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 278.160 1400.000 278.760 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1396.000 309.440 1400.000 310.040 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1130.200 4.000 1130.800 ;
    END
  END la_data_in[0]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.160 4.000 1162.760 ;
    END
  END la_data_in[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.080 4.000 1141.680 ;
    END
  END la_data_out[0]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END la_data_out[1]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.120 4.000 1194.720 ;
    END
  END la_data_out[2]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1151.280 4.000 1151.880 ;
    END
  END la_oen[0]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.240 4.000 1183.840 ;
    END
  END la_oen[1]
  PIN one_e
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END one_e
  PIN one_n
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 1196.000 18.770 1200.000 ;
    END
  END one_n
  PIN ram_ce_e
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 750.810 0.000 751.090 4.000 ;
    END
  END ram_ce_e
  PIN ram_ce_n
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 750.810 1196.000 751.090 1200.000 ;
    END
  END ram_ce_n
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.000 4.000 780.600 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.960 4.000 812.560 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.200 4.000 875.800 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.160 4.000 907.760 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.120 4.000 939.720 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.080 4.000 971.680 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1035.000 4.000 1035.600 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.280 4.000 1066.880 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.920 4.000 504.520 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.960 4.000 727.560 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.200 4.000 790.800 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.160 4.000 822.760 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.120 4.000 854.720 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.080 4.000 886.680 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.000 4.000 950.600 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 981.280 4.000 981.880 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.200 4.000 1045.800 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.160 4.000 1077.760 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.120 4.000 1109.720 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.080 4.000 376.680 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.880 4.000 451.480 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.160 4.000 482.760 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.080 4.000 546.680 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.000 4.000 610.600 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.920 4.000 674.520 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.200 4.000 705.800 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 4.000 737.760 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.120 4.000 769.720 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.080 4.000 801.680 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.960 4.000 897.560 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.200 4.000 960.800 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.160 4.000 992.760 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.120 4.000 1024.720 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.080 4.000 1056.680 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.000 4.000 1120.600 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wbs_we_i
  PIN zero_e
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END zero_e
  PIN zero_n
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 1196.000 6.350 1200.000 ;
    END
  END zero_n
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1188.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 5.865 1394.260 1188.725 ;
      LAYER met1 ;
        RECT 5.520 5.820 1394.260 1189.620 ;
      LAYER met2 ;
        RECT 6.630 1195.720 18.210 1196.000 ;
        RECT 19.050 1195.720 31.090 1196.000 ;
        RECT 31.930 1195.720 43.970 1196.000 ;
        RECT 44.810 1195.720 56.850 1196.000 ;
        RECT 57.690 1195.720 69.730 1196.000 ;
        RECT 70.570 1195.720 82.610 1196.000 ;
        RECT 83.450 1195.720 95.490 1196.000 ;
        RECT 96.330 1195.720 108.370 1196.000 ;
        RECT 109.210 1195.720 121.250 1196.000 ;
        RECT 122.090 1195.720 134.130 1196.000 ;
        RECT 134.970 1195.720 147.010 1196.000 ;
        RECT 147.850 1195.720 159.890 1196.000 ;
        RECT 160.730 1195.720 172.310 1196.000 ;
        RECT 173.150 1195.720 185.190 1196.000 ;
        RECT 186.030 1195.720 198.070 1196.000 ;
        RECT 198.910 1195.720 210.950 1196.000 ;
        RECT 211.790 1195.720 223.830 1196.000 ;
        RECT 224.670 1195.720 236.710 1196.000 ;
        RECT 237.550 1195.720 249.590 1196.000 ;
        RECT 250.430 1195.720 262.470 1196.000 ;
        RECT 263.310 1195.720 275.350 1196.000 ;
        RECT 276.190 1195.720 288.230 1196.000 ;
        RECT 289.070 1195.720 301.110 1196.000 ;
        RECT 301.950 1195.720 313.990 1196.000 ;
        RECT 314.830 1195.720 326.410 1196.000 ;
        RECT 327.250 1195.720 339.290 1196.000 ;
        RECT 340.130 1195.720 352.170 1196.000 ;
        RECT 353.010 1195.720 365.050 1196.000 ;
        RECT 365.890 1195.720 377.930 1196.000 ;
        RECT 378.770 1195.720 390.810 1196.000 ;
        RECT 391.650 1195.720 403.690 1196.000 ;
        RECT 404.530 1195.720 416.570 1196.000 ;
        RECT 417.410 1195.720 429.450 1196.000 ;
        RECT 430.290 1195.720 442.330 1196.000 ;
        RECT 443.170 1195.720 455.210 1196.000 ;
        RECT 456.050 1195.720 468.090 1196.000 ;
        RECT 468.930 1195.720 480.510 1196.000 ;
        RECT 481.350 1195.720 493.390 1196.000 ;
        RECT 494.230 1195.720 506.270 1196.000 ;
        RECT 507.110 1195.720 519.150 1196.000 ;
        RECT 519.990 1195.720 532.030 1196.000 ;
        RECT 532.870 1195.720 544.910 1196.000 ;
        RECT 545.750 1195.720 557.790 1196.000 ;
        RECT 558.630 1195.720 570.670 1196.000 ;
        RECT 571.510 1195.720 583.550 1196.000 ;
        RECT 584.390 1195.720 596.430 1196.000 ;
        RECT 597.270 1195.720 609.310 1196.000 ;
        RECT 610.150 1195.720 622.190 1196.000 ;
        RECT 623.030 1195.720 634.610 1196.000 ;
        RECT 635.450 1195.720 647.490 1196.000 ;
        RECT 648.330 1195.720 660.370 1196.000 ;
        RECT 661.210 1195.720 673.250 1196.000 ;
        RECT 674.090 1195.720 686.130 1196.000 ;
        RECT 686.970 1195.720 699.010 1196.000 ;
        RECT 699.850 1195.720 711.890 1196.000 ;
        RECT 712.730 1195.720 724.770 1196.000 ;
        RECT 725.610 1195.720 737.650 1196.000 ;
        RECT 738.490 1195.720 750.530 1196.000 ;
        RECT 751.370 1195.720 763.410 1196.000 ;
        RECT 764.250 1195.720 776.290 1196.000 ;
        RECT 777.130 1195.720 788.710 1196.000 ;
        RECT 789.550 1195.720 801.590 1196.000 ;
        RECT 802.430 1195.720 814.470 1196.000 ;
        RECT 815.310 1195.720 827.350 1196.000 ;
        RECT 828.190 1195.720 840.230 1196.000 ;
        RECT 841.070 1195.720 853.110 1196.000 ;
        RECT 853.950 1195.720 865.990 1196.000 ;
        RECT 866.830 1195.720 878.870 1196.000 ;
        RECT 879.710 1195.720 891.750 1196.000 ;
        RECT 892.590 1195.720 904.630 1196.000 ;
        RECT 905.470 1195.720 917.510 1196.000 ;
        RECT 918.350 1195.720 930.390 1196.000 ;
        RECT 931.230 1195.720 942.810 1196.000 ;
        RECT 943.650 1195.720 955.690 1196.000 ;
        RECT 956.530 1195.720 968.570 1196.000 ;
        RECT 969.410 1195.720 981.450 1196.000 ;
        RECT 982.290 1195.720 994.330 1196.000 ;
        RECT 995.170 1195.720 1007.210 1196.000 ;
        RECT 1008.050 1195.720 1020.090 1196.000 ;
        RECT 1020.930 1195.720 1032.970 1196.000 ;
        RECT 1033.810 1195.720 1045.850 1196.000 ;
        RECT 1046.690 1195.720 1058.730 1196.000 ;
        RECT 1059.570 1195.720 1071.610 1196.000 ;
        RECT 1072.450 1195.720 1084.490 1196.000 ;
        RECT 1085.330 1195.720 1096.910 1196.000 ;
        RECT 1097.750 1195.720 1109.790 1196.000 ;
        RECT 1110.630 1195.720 1122.670 1196.000 ;
        RECT 1123.510 1195.720 1135.550 1196.000 ;
        RECT 1136.390 1195.720 1148.430 1196.000 ;
        RECT 1149.270 1195.720 1161.310 1196.000 ;
        RECT 1162.150 1195.720 1174.190 1196.000 ;
        RECT 1175.030 1195.720 1187.070 1196.000 ;
        RECT 1187.910 1195.720 1199.950 1196.000 ;
        RECT 1200.790 1195.720 1212.830 1196.000 ;
        RECT 1213.670 1195.720 1225.710 1196.000 ;
        RECT 1226.550 1195.720 1238.590 1196.000 ;
        RECT 1239.430 1195.720 1251.010 1196.000 ;
        RECT 1251.850 1195.720 1263.890 1196.000 ;
        RECT 1264.730 1195.720 1276.770 1196.000 ;
        RECT 1277.610 1195.720 1289.650 1196.000 ;
        RECT 1290.490 1195.720 1302.530 1196.000 ;
        RECT 1303.370 1195.720 1315.410 1196.000 ;
        RECT 1316.250 1195.720 1328.290 1196.000 ;
        RECT 1329.130 1195.720 1341.170 1196.000 ;
        RECT 1342.010 1195.720 1354.050 1196.000 ;
        RECT 1354.890 1195.720 1366.930 1196.000 ;
        RECT 1367.770 1195.720 1379.810 1196.000 ;
        RECT 1380.650 1195.720 1392.690 1196.000 ;
        RECT 1393.530 1195.720 1395.550 1196.000 ;
        RECT 6.080 4.280 1395.550 1195.720 ;
        RECT 6.630 4.000 18.210 4.280 ;
        RECT 19.050 4.000 31.090 4.280 ;
        RECT 31.930 4.000 43.970 4.280 ;
        RECT 44.810 4.000 56.850 4.280 ;
        RECT 57.690 4.000 69.730 4.280 ;
        RECT 70.570 4.000 82.610 4.280 ;
        RECT 83.450 4.000 95.490 4.280 ;
        RECT 96.330 4.000 108.370 4.280 ;
        RECT 109.210 4.000 121.250 4.280 ;
        RECT 122.090 4.000 134.130 4.280 ;
        RECT 134.970 4.000 147.010 4.280 ;
        RECT 147.850 4.000 159.890 4.280 ;
        RECT 160.730 4.000 172.310 4.280 ;
        RECT 173.150 4.000 185.190 4.280 ;
        RECT 186.030 4.000 198.070 4.280 ;
        RECT 198.910 4.000 210.950 4.280 ;
        RECT 211.790 4.000 223.830 4.280 ;
        RECT 224.670 4.000 236.710 4.280 ;
        RECT 237.550 4.000 249.590 4.280 ;
        RECT 250.430 4.000 262.470 4.280 ;
        RECT 263.310 4.000 275.350 4.280 ;
        RECT 276.190 4.000 288.230 4.280 ;
        RECT 289.070 4.000 301.110 4.280 ;
        RECT 301.950 4.000 313.990 4.280 ;
        RECT 314.830 4.000 326.410 4.280 ;
        RECT 327.250 4.000 339.290 4.280 ;
        RECT 340.130 4.000 352.170 4.280 ;
        RECT 353.010 4.000 365.050 4.280 ;
        RECT 365.890 4.000 377.930 4.280 ;
        RECT 378.770 4.000 390.810 4.280 ;
        RECT 391.650 4.000 403.690 4.280 ;
        RECT 404.530 4.000 416.570 4.280 ;
        RECT 417.410 4.000 429.450 4.280 ;
        RECT 430.290 4.000 442.330 4.280 ;
        RECT 443.170 4.000 455.210 4.280 ;
        RECT 456.050 4.000 468.090 4.280 ;
        RECT 468.930 4.000 480.510 4.280 ;
        RECT 481.350 4.000 493.390 4.280 ;
        RECT 494.230 4.000 506.270 4.280 ;
        RECT 507.110 4.000 519.150 4.280 ;
        RECT 519.990 4.000 532.030 4.280 ;
        RECT 532.870 4.000 544.910 4.280 ;
        RECT 545.750 4.000 557.790 4.280 ;
        RECT 558.630 4.000 570.670 4.280 ;
        RECT 571.510 4.000 583.550 4.280 ;
        RECT 584.390 4.000 596.430 4.280 ;
        RECT 597.270 4.000 609.310 4.280 ;
        RECT 610.150 4.000 622.190 4.280 ;
        RECT 623.030 4.000 634.610 4.280 ;
        RECT 635.450 4.000 647.490 4.280 ;
        RECT 648.330 4.000 660.370 4.280 ;
        RECT 661.210 4.000 673.250 4.280 ;
        RECT 674.090 4.000 686.130 4.280 ;
        RECT 686.970 4.000 699.010 4.280 ;
        RECT 699.850 4.000 711.890 4.280 ;
        RECT 712.730 4.000 724.770 4.280 ;
        RECT 725.610 4.000 737.650 4.280 ;
        RECT 738.490 4.000 750.530 4.280 ;
        RECT 751.370 4.000 763.410 4.280 ;
        RECT 764.250 4.000 776.290 4.280 ;
        RECT 777.130 4.000 788.710 4.280 ;
        RECT 789.550 4.000 801.590 4.280 ;
        RECT 802.430 4.000 814.470 4.280 ;
        RECT 815.310 4.000 827.350 4.280 ;
        RECT 828.190 4.000 840.230 4.280 ;
        RECT 841.070 4.000 853.110 4.280 ;
        RECT 853.950 4.000 865.990 4.280 ;
        RECT 866.830 4.000 878.870 4.280 ;
        RECT 879.710 4.000 891.750 4.280 ;
        RECT 892.590 4.000 904.630 4.280 ;
        RECT 905.470 4.000 917.510 4.280 ;
        RECT 918.350 4.000 930.390 4.280 ;
        RECT 931.230 4.000 942.810 4.280 ;
        RECT 943.650 4.000 955.690 4.280 ;
        RECT 956.530 4.000 968.570 4.280 ;
        RECT 969.410 4.000 981.450 4.280 ;
        RECT 982.290 4.000 994.330 4.280 ;
        RECT 995.170 4.000 1007.210 4.280 ;
        RECT 1008.050 4.000 1020.090 4.280 ;
        RECT 1020.930 4.000 1032.970 4.280 ;
        RECT 1033.810 4.000 1045.850 4.280 ;
        RECT 1046.690 4.000 1058.730 4.280 ;
        RECT 1059.570 4.000 1071.610 4.280 ;
        RECT 1072.450 4.000 1084.490 4.280 ;
        RECT 1085.330 4.000 1096.910 4.280 ;
        RECT 1097.750 4.000 1109.790 4.280 ;
        RECT 1110.630 4.000 1122.670 4.280 ;
        RECT 1123.510 4.000 1135.550 4.280 ;
        RECT 1136.390 4.000 1148.430 4.280 ;
        RECT 1149.270 4.000 1161.310 4.280 ;
        RECT 1162.150 4.000 1174.190 4.280 ;
        RECT 1175.030 4.000 1187.070 4.280 ;
        RECT 1187.910 4.000 1199.950 4.280 ;
        RECT 1200.790 4.000 1212.830 4.280 ;
        RECT 1213.670 4.000 1225.710 4.280 ;
        RECT 1226.550 4.000 1238.590 4.280 ;
        RECT 1239.430 4.000 1251.010 4.280 ;
        RECT 1251.850 4.000 1263.890 4.280 ;
        RECT 1264.730 4.000 1276.770 4.280 ;
        RECT 1277.610 4.000 1289.650 4.280 ;
        RECT 1290.490 4.000 1302.530 4.280 ;
        RECT 1303.370 4.000 1315.410 4.280 ;
        RECT 1316.250 4.000 1328.290 4.280 ;
        RECT 1329.130 4.000 1341.170 4.280 ;
        RECT 1342.010 4.000 1354.050 4.280 ;
        RECT 1354.890 4.000 1366.930 4.280 ;
        RECT 1367.770 4.000 1379.810 4.280 ;
        RECT 1380.650 4.000 1392.690 4.280 ;
        RECT 1393.530 4.000 1395.550 4.280 ;
      LAYER met3 ;
        RECT 4.400 1193.720 1395.600 1194.585 ;
        RECT 3.990 1184.920 1396.000 1193.720 ;
        RECT 3.990 1184.240 1395.600 1184.920 ;
        RECT 4.400 1183.520 1395.600 1184.240 ;
        RECT 4.400 1182.840 1396.000 1183.520 ;
        RECT 3.990 1174.040 1396.000 1182.840 ;
        RECT 4.400 1172.640 1395.600 1174.040 ;
        RECT 3.990 1163.840 1396.000 1172.640 ;
        RECT 3.990 1163.160 1395.600 1163.840 ;
        RECT 4.400 1162.440 1395.600 1163.160 ;
        RECT 4.400 1161.760 1396.000 1162.440 ;
        RECT 3.990 1152.960 1396.000 1161.760 ;
        RECT 3.990 1152.280 1395.600 1152.960 ;
        RECT 4.400 1151.560 1395.600 1152.280 ;
        RECT 4.400 1150.880 1396.000 1151.560 ;
        RECT 3.990 1142.760 1396.000 1150.880 ;
        RECT 3.990 1142.080 1395.600 1142.760 ;
        RECT 4.400 1141.360 1395.600 1142.080 ;
        RECT 4.400 1140.680 1396.000 1141.360 ;
        RECT 3.990 1131.880 1396.000 1140.680 ;
        RECT 3.990 1131.200 1395.600 1131.880 ;
        RECT 4.400 1130.480 1395.600 1131.200 ;
        RECT 4.400 1129.800 1396.000 1130.480 ;
        RECT 3.990 1121.680 1396.000 1129.800 ;
        RECT 3.990 1121.000 1395.600 1121.680 ;
        RECT 4.400 1120.280 1395.600 1121.000 ;
        RECT 4.400 1119.600 1396.000 1120.280 ;
        RECT 3.990 1110.800 1396.000 1119.600 ;
        RECT 3.990 1110.120 1395.600 1110.800 ;
        RECT 4.400 1109.400 1395.600 1110.120 ;
        RECT 4.400 1108.720 1396.000 1109.400 ;
        RECT 3.990 1100.600 1396.000 1108.720 ;
        RECT 3.990 1099.240 1395.600 1100.600 ;
        RECT 4.400 1099.200 1395.600 1099.240 ;
        RECT 4.400 1097.840 1396.000 1099.200 ;
        RECT 3.990 1089.720 1396.000 1097.840 ;
        RECT 3.990 1089.040 1395.600 1089.720 ;
        RECT 4.400 1088.320 1395.600 1089.040 ;
        RECT 4.400 1087.640 1396.000 1088.320 ;
        RECT 3.990 1079.520 1396.000 1087.640 ;
        RECT 3.990 1078.160 1395.600 1079.520 ;
        RECT 4.400 1078.120 1395.600 1078.160 ;
        RECT 4.400 1076.760 1396.000 1078.120 ;
        RECT 3.990 1068.640 1396.000 1076.760 ;
        RECT 3.990 1067.280 1395.600 1068.640 ;
        RECT 4.400 1067.240 1395.600 1067.280 ;
        RECT 4.400 1065.880 1396.000 1067.240 ;
        RECT 3.990 1058.440 1396.000 1065.880 ;
        RECT 3.990 1057.080 1395.600 1058.440 ;
        RECT 4.400 1057.040 1395.600 1057.080 ;
        RECT 4.400 1055.680 1396.000 1057.040 ;
        RECT 3.990 1047.560 1396.000 1055.680 ;
        RECT 3.990 1046.200 1395.600 1047.560 ;
        RECT 4.400 1046.160 1395.600 1046.200 ;
        RECT 4.400 1044.800 1396.000 1046.160 ;
        RECT 3.990 1037.360 1396.000 1044.800 ;
        RECT 3.990 1036.000 1395.600 1037.360 ;
        RECT 4.400 1035.960 1395.600 1036.000 ;
        RECT 4.400 1034.600 1396.000 1035.960 ;
        RECT 3.990 1026.480 1396.000 1034.600 ;
        RECT 3.990 1025.120 1395.600 1026.480 ;
        RECT 4.400 1025.080 1395.600 1025.120 ;
        RECT 4.400 1023.720 1396.000 1025.080 ;
        RECT 3.990 1016.280 1396.000 1023.720 ;
        RECT 3.990 1014.880 1395.600 1016.280 ;
        RECT 3.990 1014.240 1396.000 1014.880 ;
        RECT 4.400 1012.840 1396.000 1014.240 ;
        RECT 3.990 1005.400 1396.000 1012.840 ;
        RECT 3.990 1004.040 1395.600 1005.400 ;
        RECT 4.400 1004.000 1395.600 1004.040 ;
        RECT 4.400 1002.640 1396.000 1004.000 ;
        RECT 3.990 995.200 1396.000 1002.640 ;
        RECT 3.990 993.800 1395.600 995.200 ;
        RECT 3.990 993.160 1396.000 993.800 ;
        RECT 4.400 991.760 1396.000 993.160 ;
        RECT 3.990 984.320 1396.000 991.760 ;
        RECT 3.990 982.920 1395.600 984.320 ;
        RECT 3.990 982.280 1396.000 982.920 ;
        RECT 4.400 980.880 1396.000 982.280 ;
        RECT 3.990 974.120 1396.000 980.880 ;
        RECT 3.990 972.720 1395.600 974.120 ;
        RECT 3.990 972.080 1396.000 972.720 ;
        RECT 4.400 970.680 1396.000 972.080 ;
        RECT 3.990 963.240 1396.000 970.680 ;
        RECT 3.990 961.840 1395.600 963.240 ;
        RECT 3.990 961.200 1396.000 961.840 ;
        RECT 4.400 959.800 1396.000 961.200 ;
        RECT 3.990 953.040 1396.000 959.800 ;
        RECT 3.990 951.640 1395.600 953.040 ;
        RECT 3.990 951.000 1396.000 951.640 ;
        RECT 4.400 949.600 1396.000 951.000 ;
        RECT 3.990 942.160 1396.000 949.600 ;
        RECT 3.990 940.760 1395.600 942.160 ;
        RECT 3.990 940.120 1396.000 940.760 ;
        RECT 4.400 938.720 1396.000 940.120 ;
        RECT 3.990 931.960 1396.000 938.720 ;
        RECT 3.990 930.560 1395.600 931.960 ;
        RECT 3.990 929.240 1396.000 930.560 ;
        RECT 4.400 927.840 1396.000 929.240 ;
        RECT 3.990 921.080 1396.000 927.840 ;
        RECT 3.990 919.680 1395.600 921.080 ;
        RECT 3.990 919.040 1396.000 919.680 ;
        RECT 4.400 917.640 1396.000 919.040 ;
        RECT 3.990 910.880 1396.000 917.640 ;
        RECT 3.990 909.480 1395.600 910.880 ;
        RECT 3.990 908.160 1396.000 909.480 ;
        RECT 4.400 906.760 1396.000 908.160 ;
        RECT 3.990 900.680 1396.000 906.760 ;
        RECT 3.990 899.280 1395.600 900.680 ;
        RECT 3.990 897.960 1396.000 899.280 ;
        RECT 4.400 896.560 1396.000 897.960 ;
        RECT 3.990 889.800 1396.000 896.560 ;
        RECT 3.990 888.400 1395.600 889.800 ;
        RECT 3.990 887.080 1396.000 888.400 ;
        RECT 4.400 885.680 1396.000 887.080 ;
        RECT 3.990 879.600 1396.000 885.680 ;
        RECT 3.990 878.200 1395.600 879.600 ;
        RECT 3.990 876.200 1396.000 878.200 ;
        RECT 4.400 874.800 1396.000 876.200 ;
        RECT 3.990 868.720 1396.000 874.800 ;
        RECT 3.990 867.320 1395.600 868.720 ;
        RECT 3.990 866.000 1396.000 867.320 ;
        RECT 4.400 864.600 1396.000 866.000 ;
        RECT 3.990 858.520 1396.000 864.600 ;
        RECT 3.990 857.120 1395.600 858.520 ;
        RECT 3.990 855.120 1396.000 857.120 ;
        RECT 4.400 853.720 1396.000 855.120 ;
        RECT 3.990 847.640 1396.000 853.720 ;
        RECT 3.990 846.240 1395.600 847.640 ;
        RECT 3.990 844.240 1396.000 846.240 ;
        RECT 4.400 842.840 1396.000 844.240 ;
        RECT 3.990 837.440 1396.000 842.840 ;
        RECT 3.990 836.040 1395.600 837.440 ;
        RECT 3.990 834.040 1396.000 836.040 ;
        RECT 4.400 832.640 1396.000 834.040 ;
        RECT 3.990 826.560 1396.000 832.640 ;
        RECT 3.990 825.160 1395.600 826.560 ;
        RECT 3.990 823.160 1396.000 825.160 ;
        RECT 4.400 821.760 1396.000 823.160 ;
        RECT 3.990 816.360 1396.000 821.760 ;
        RECT 3.990 814.960 1395.600 816.360 ;
        RECT 3.990 812.960 1396.000 814.960 ;
        RECT 4.400 811.560 1396.000 812.960 ;
        RECT 3.990 805.480 1396.000 811.560 ;
        RECT 3.990 804.080 1395.600 805.480 ;
        RECT 3.990 802.080 1396.000 804.080 ;
        RECT 4.400 800.680 1396.000 802.080 ;
        RECT 3.990 795.280 1396.000 800.680 ;
        RECT 3.990 793.880 1395.600 795.280 ;
        RECT 3.990 791.200 1396.000 793.880 ;
        RECT 4.400 789.800 1396.000 791.200 ;
        RECT 3.990 784.400 1396.000 789.800 ;
        RECT 3.990 783.000 1395.600 784.400 ;
        RECT 3.990 781.000 1396.000 783.000 ;
        RECT 4.400 779.600 1396.000 781.000 ;
        RECT 3.990 774.200 1396.000 779.600 ;
        RECT 3.990 772.800 1395.600 774.200 ;
        RECT 3.990 770.120 1396.000 772.800 ;
        RECT 4.400 768.720 1396.000 770.120 ;
        RECT 3.990 763.320 1396.000 768.720 ;
        RECT 3.990 761.920 1395.600 763.320 ;
        RECT 3.990 759.240 1396.000 761.920 ;
        RECT 4.400 757.840 1396.000 759.240 ;
        RECT 3.990 753.120 1396.000 757.840 ;
        RECT 3.990 751.720 1395.600 753.120 ;
        RECT 3.990 749.040 1396.000 751.720 ;
        RECT 4.400 747.640 1396.000 749.040 ;
        RECT 3.990 742.240 1396.000 747.640 ;
        RECT 3.990 740.840 1395.600 742.240 ;
        RECT 3.990 738.160 1396.000 740.840 ;
        RECT 4.400 736.760 1396.000 738.160 ;
        RECT 3.990 732.040 1396.000 736.760 ;
        RECT 3.990 730.640 1395.600 732.040 ;
        RECT 3.990 727.960 1396.000 730.640 ;
        RECT 4.400 726.560 1396.000 727.960 ;
        RECT 3.990 721.160 1396.000 726.560 ;
        RECT 3.990 719.760 1395.600 721.160 ;
        RECT 3.990 717.080 1396.000 719.760 ;
        RECT 4.400 715.680 1396.000 717.080 ;
        RECT 3.990 710.960 1396.000 715.680 ;
        RECT 3.990 709.560 1395.600 710.960 ;
        RECT 3.990 706.200 1396.000 709.560 ;
        RECT 4.400 704.800 1396.000 706.200 ;
        RECT 3.990 700.080 1396.000 704.800 ;
        RECT 3.990 698.680 1395.600 700.080 ;
        RECT 3.990 696.000 1396.000 698.680 ;
        RECT 4.400 694.600 1396.000 696.000 ;
        RECT 3.990 689.880 1396.000 694.600 ;
        RECT 3.990 688.480 1395.600 689.880 ;
        RECT 3.990 685.120 1396.000 688.480 ;
        RECT 4.400 683.720 1396.000 685.120 ;
        RECT 3.990 679.000 1396.000 683.720 ;
        RECT 3.990 677.600 1395.600 679.000 ;
        RECT 3.990 674.920 1396.000 677.600 ;
        RECT 4.400 673.520 1396.000 674.920 ;
        RECT 3.990 668.800 1396.000 673.520 ;
        RECT 3.990 667.400 1395.600 668.800 ;
        RECT 3.990 664.040 1396.000 667.400 ;
        RECT 4.400 662.640 1396.000 664.040 ;
        RECT 3.990 657.920 1396.000 662.640 ;
        RECT 3.990 656.520 1395.600 657.920 ;
        RECT 3.990 653.160 1396.000 656.520 ;
        RECT 4.400 651.760 1396.000 653.160 ;
        RECT 3.990 647.720 1396.000 651.760 ;
        RECT 3.990 646.320 1395.600 647.720 ;
        RECT 3.990 642.960 1396.000 646.320 ;
        RECT 4.400 641.560 1396.000 642.960 ;
        RECT 3.990 636.840 1396.000 641.560 ;
        RECT 3.990 635.440 1395.600 636.840 ;
        RECT 3.990 632.080 1396.000 635.440 ;
        RECT 4.400 630.680 1396.000 632.080 ;
        RECT 3.990 626.640 1396.000 630.680 ;
        RECT 3.990 625.240 1395.600 626.640 ;
        RECT 3.990 621.200 1396.000 625.240 ;
        RECT 4.400 619.800 1396.000 621.200 ;
        RECT 3.990 615.760 1396.000 619.800 ;
        RECT 3.990 614.360 1395.600 615.760 ;
        RECT 3.990 611.000 1396.000 614.360 ;
        RECT 4.400 609.600 1396.000 611.000 ;
        RECT 3.990 605.560 1396.000 609.600 ;
        RECT 3.990 604.160 1395.600 605.560 ;
        RECT 3.990 600.120 1396.000 604.160 ;
        RECT 4.400 598.720 1396.000 600.120 ;
        RECT 3.990 595.360 1396.000 598.720 ;
        RECT 3.990 593.960 1395.600 595.360 ;
        RECT 3.990 589.920 1396.000 593.960 ;
        RECT 4.400 588.520 1396.000 589.920 ;
        RECT 3.990 584.480 1396.000 588.520 ;
        RECT 3.990 583.080 1395.600 584.480 ;
        RECT 3.990 579.040 1396.000 583.080 ;
        RECT 4.400 577.640 1396.000 579.040 ;
        RECT 3.990 574.280 1396.000 577.640 ;
        RECT 3.990 572.880 1395.600 574.280 ;
        RECT 3.990 568.160 1396.000 572.880 ;
        RECT 4.400 566.760 1396.000 568.160 ;
        RECT 3.990 563.400 1396.000 566.760 ;
        RECT 3.990 562.000 1395.600 563.400 ;
        RECT 3.990 557.960 1396.000 562.000 ;
        RECT 4.400 556.560 1396.000 557.960 ;
        RECT 3.990 553.200 1396.000 556.560 ;
        RECT 3.990 551.800 1395.600 553.200 ;
        RECT 3.990 547.080 1396.000 551.800 ;
        RECT 4.400 545.680 1396.000 547.080 ;
        RECT 3.990 542.320 1396.000 545.680 ;
        RECT 3.990 540.920 1395.600 542.320 ;
        RECT 3.990 536.200 1396.000 540.920 ;
        RECT 4.400 534.800 1396.000 536.200 ;
        RECT 3.990 532.120 1396.000 534.800 ;
        RECT 3.990 530.720 1395.600 532.120 ;
        RECT 3.990 526.000 1396.000 530.720 ;
        RECT 4.400 524.600 1396.000 526.000 ;
        RECT 3.990 521.240 1396.000 524.600 ;
        RECT 3.990 519.840 1395.600 521.240 ;
        RECT 3.990 515.120 1396.000 519.840 ;
        RECT 4.400 513.720 1396.000 515.120 ;
        RECT 3.990 511.040 1396.000 513.720 ;
        RECT 3.990 509.640 1395.600 511.040 ;
        RECT 3.990 504.920 1396.000 509.640 ;
        RECT 4.400 503.520 1396.000 504.920 ;
        RECT 3.990 500.160 1396.000 503.520 ;
        RECT 3.990 498.760 1395.600 500.160 ;
        RECT 3.990 494.040 1396.000 498.760 ;
        RECT 4.400 492.640 1396.000 494.040 ;
        RECT 3.990 489.960 1396.000 492.640 ;
        RECT 3.990 488.560 1395.600 489.960 ;
        RECT 3.990 483.160 1396.000 488.560 ;
        RECT 4.400 481.760 1396.000 483.160 ;
        RECT 3.990 479.080 1396.000 481.760 ;
        RECT 3.990 477.680 1395.600 479.080 ;
        RECT 3.990 472.960 1396.000 477.680 ;
        RECT 4.400 471.560 1396.000 472.960 ;
        RECT 3.990 468.880 1396.000 471.560 ;
        RECT 3.990 467.480 1395.600 468.880 ;
        RECT 3.990 462.080 1396.000 467.480 ;
        RECT 4.400 460.680 1396.000 462.080 ;
        RECT 3.990 458.000 1396.000 460.680 ;
        RECT 3.990 456.600 1395.600 458.000 ;
        RECT 3.990 451.880 1396.000 456.600 ;
        RECT 4.400 450.480 1396.000 451.880 ;
        RECT 3.990 447.800 1396.000 450.480 ;
        RECT 3.990 446.400 1395.600 447.800 ;
        RECT 3.990 441.000 1396.000 446.400 ;
        RECT 4.400 439.600 1396.000 441.000 ;
        RECT 3.990 436.920 1396.000 439.600 ;
        RECT 3.990 435.520 1395.600 436.920 ;
        RECT 3.990 430.120 1396.000 435.520 ;
        RECT 4.400 428.720 1396.000 430.120 ;
        RECT 3.990 426.720 1396.000 428.720 ;
        RECT 3.990 425.320 1395.600 426.720 ;
        RECT 3.990 419.920 1396.000 425.320 ;
        RECT 4.400 418.520 1396.000 419.920 ;
        RECT 3.990 415.840 1396.000 418.520 ;
        RECT 3.990 414.440 1395.600 415.840 ;
        RECT 3.990 409.040 1396.000 414.440 ;
        RECT 4.400 407.640 1396.000 409.040 ;
        RECT 3.990 405.640 1396.000 407.640 ;
        RECT 3.990 404.240 1395.600 405.640 ;
        RECT 3.990 398.160 1396.000 404.240 ;
        RECT 4.400 396.760 1396.000 398.160 ;
        RECT 3.990 394.760 1396.000 396.760 ;
        RECT 3.990 393.360 1395.600 394.760 ;
        RECT 3.990 387.960 1396.000 393.360 ;
        RECT 4.400 386.560 1396.000 387.960 ;
        RECT 3.990 384.560 1396.000 386.560 ;
        RECT 3.990 383.160 1395.600 384.560 ;
        RECT 3.990 377.080 1396.000 383.160 ;
        RECT 4.400 375.680 1396.000 377.080 ;
        RECT 3.990 373.680 1396.000 375.680 ;
        RECT 3.990 372.280 1395.600 373.680 ;
        RECT 3.990 366.880 1396.000 372.280 ;
        RECT 4.400 365.480 1396.000 366.880 ;
        RECT 3.990 363.480 1396.000 365.480 ;
        RECT 3.990 362.080 1395.600 363.480 ;
        RECT 3.990 356.000 1396.000 362.080 ;
        RECT 4.400 354.600 1396.000 356.000 ;
        RECT 3.990 352.600 1396.000 354.600 ;
        RECT 3.990 351.200 1395.600 352.600 ;
        RECT 3.990 345.120 1396.000 351.200 ;
        RECT 4.400 343.720 1396.000 345.120 ;
        RECT 3.990 342.400 1396.000 343.720 ;
        RECT 3.990 341.000 1395.600 342.400 ;
        RECT 3.990 334.920 1396.000 341.000 ;
        RECT 4.400 333.520 1396.000 334.920 ;
        RECT 3.990 331.520 1396.000 333.520 ;
        RECT 3.990 330.120 1395.600 331.520 ;
        RECT 3.990 324.040 1396.000 330.120 ;
        RECT 4.400 322.640 1396.000 324.040 ;
        RECT 3.990 321.320 1396.000 322.640 ;
        RECT 3.990 319.920 1395.600 321.320 ;
        RECT 3.990 313.160 1396.000 319.920 ;
        RECT 4.400 311.760 1396.000 313.160 ;
        RECT 3.990 310.440 1396.000 311.760 ;
        RECT 3.990 309.040 1395.600 310.440 ;
        RECT 3.990 302.960 1396.000 309.040 ;
        RECT 4.400 301.560 1396.000 302.960 ;
        RECT 3.990 300.240 1396.000 301.560 ;
        RECT 3.990 298.840 1395.600 300.240 ;
        RECT 3.990 292.080 1396.000 298.840 ;
        RECT 4.400 290.680 1396.000 292.080 ;
        RECT 3.990 290.040 1396.000 290.680 ;
        RECT 3.990 288.640 1395.600 290.040 ;
        RECT 3.990 281.880 1396.000 288.640 ;
        RECT 4.400 280.480 1396.000 281.880 ;
        RECT 3.990 279.160 1396.000 280.480 ;
        RECT 3.990 277.760 1395.600 279.160 ;
        RECT 3.990 271.000 1396.000 277.760 ;
        RECT 4.400 269.600 1396.000 271.000 ;
        RECT 3.990 268.960 1396.000 269.600 ;
        RECT 3.990 267.560 1395.600 268.960 ;
        RECT 3.990 260.120 1396.000 267.560 ;
        RECT 4.400 258.720 1396.000 260.120 ;
        RECT 3.990 258.080 1396.000 258.720 ;
        RECT 3.990 256.680 1395.600 258.080 ;
        RECT 3.990 249.920 1396.000 256.680 ;
        RECT 4.400 248.520 1396.000 249.920 ;
        RECT 3.990 247.880 1396.000 248.520 ;
        RECT 3.990 246.480 1395.600 247.880 ;
        RECT 3.990 239.040 1396.000 246.480 ;
        RECT 4.400 237.640 1396.000 239.040 ;
        RECT 3.990 237.000 1396.000 237.640 ;
        RECT 3.990 235.600 1395.600 237.000 ;
        RECT 3.990 228.840 1396.000 235.600 ;
        RECT 4.400 227.440 1396.000 228.840 ;
        RECT 3.990 226.800 1396.000 227.440 ;
        RECT 3.990 225.400 1395.600 226.800 ;
        RECT 3.990 217.960 1396.000 225.400 ;
        RECT 4.400 216.560 1396.000 217.960 ;
        RECT 3.990 215.920 1396.000 216.560 ;
        RECT 3.990 214.520 1395.600 215.920 ;
        RECT 3.990 207.080 1396.000 214.520 ;
        RECT 4.400 205.720 1396.000 207.080 ;
        RECT 4.400 205.680 1395.600 205.720 ;
        RECT 3.990 204.320 1395.600 205.680 ;
        RECT 3.990 196.880 1396.000 204.320 ;
        RECT 4.400 195.480 1396.000 196.880 ;
        RECT 3.990 194.840 1396.000 195.480 ;
        RECT 3.990 193.440 1395.600 194.840 ;
        RECT 3.990 186.000 1396.000 193.440 ;
        RECT 4.400 184.640 1396.000 186.000 ;
        RECT 4.400 184.600 1395.600 184.640 ;
        RECT 3.990 183.240 1395.600 184.600 ;
        RECT 3.990 175.120 1396.000 183.240 ;
        RECT 4.400 173.760 1396.000 175.120 ;
        RECT 4.400 173.720 1395.600 173.760 ;
        RECT 3.990 172.360 1395.600 173.720 ;
        RECT 3.990 164.920 1396.000 172.360 ;
        RECT 4.400 163.560 1396.000 164.920 ;
        RECT 4.400 163.520 1395.600 163.560 ;
        RECT 3.990 162.160 1395.600 163.520 ;
        RECT 3.990 154.040 1396.000 162.160 ;
        RECT 4.400 152.680 1396.000 154.040 ;
        RECT 4.400 152.640 1395.600 152.680 ;
        RECT 3.990 151.280 1395.600 152.640 ;
        RECT 3.990 143.840 1396.000 151.280 ;
        RECT 4.400 142.480 1396.000 143.840 ;
        RECT 4.400 142.440 1395.600 142.480 ;
        RECT 3.990 141.080 1395.600 142.440 ;
        RECT 3.990 132.960 1396.000 141.080 ;
        RECT 4.400 131.600 1396.000 132.960 ;
        RECT 4.400 131.560 1395.600 131.600 ;
        RECT 3.990 130.200 1395.600 131.560 ;
        RECT 3.990 122.080 1396.000 130.200 ;
        RECT 4.400 121.400 1396.000 122.080 ;
        RECT 4.400 120.680 1395.600 121.400 ;
        RECT 3.990 120.000 1395.600 120.680 ;
        RECT 3.990 111.880 1396.000 120.000 ;
        RECT 4.400 110.520 1396.000 111.880 ;
        RECT 4.400 110.480 1395.600 110.520 ;
        RECT 3.990 109.120 1395.600 110.480 ;
        RECT 3.990 101.000 1396.000 109.120 ;
        RECT 4.400 100.320 1396.000 101.000 ;
        RECT 4.400 99.600 1395.600 100.320 ;
        RECT 3.990 98.920 1395.600 99.600 ;
        RECT 3.990 90.120 1396.000 98.920 ;
        RECT 4.400 89.440 1396.000 90.120 ;
        RECT 4.400 88.720 1395.600 89.440 ;
        RECT 3.990 88.040 1395.600 88.720 ;
        RECT 3.990 79.920 1396.000 88.040 ;
        RECT 4.400 79.240 1396.000 79.920 ;
        RECT 4.400 78.520 1395.600 79.240 ;
        RECT 3.990 77.840 1395.600 78.520 ;
        RECT 3.990 69.040 1396.000 77.840 ;
        RECT 4.400 68.360 1396.000 69.040 ;
        RECT 4.400 67.640 1395.600 68.360 ;
        RECT 3.990 66.960 1395.600 67.640 ;
        RECT 3.990 58.840 1396.000 66.960 ;
        RECT 4.400 58.160 1396.000 58.840 ;
        RECT 4.400 57.440 1395.600 58.160 ;
        RECT 3.990 56.760 1395.600 57.440 ;
        RECT 3.990 47.960 1396.000 56.760 ;
        RECT 4.400 47.280 1396.000 47.960 ;
        RECT 4.400 46.560 1395.600 47.280 ;
        RECT 3.990 45.880 1395.600 46.560 ;
        RECT 3.990 37.080 1396.000 45.880 ;
        RECT 4.400 35.680 1395.600 37.080 ;
        RECT 3.990 26.880 1396.000 35.680 ;
        RECT 4.400 26.200 1396.000 26.880 ;
        RECT 4.400 25.480 1395.600 26.200 ;
        RECT 3.990 24.800 1395.600 25.480 ;
        RECT 3.990 16.000 1396.000 24.800 ;
        RECT 4.400 14.600 1395.600 16.000 ;
        RECT 3.990 5.800 1396.000 14.600 ;
        RECT 4.400 4.950 1395.600 5.800 ;
      LAYER met4 ;
        RECT 16.855 10.240 20.640 1188.880 ;
        RECT 23.040 10.240 97.440 1188.880 ;
        RECT 99.840 10.240 1378.785 1188.880 ;
        RECT 16.855 6.295 1378.785 10.240 ;
  END
END hs32_core1
END LIBRARY

