VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hs32_core1
  CLASS BLOCK ;
  FOREIGN hs32_core1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1200.000 ;
  PIN cpu_addr_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END cpu_addr_e[0]
  PIN cpu_addr_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END cpu_addr_e[10]
  PIN cpu_addr_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END cpu_addr_e[11]
  PIN cpu_addr_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END cpu_addr_e[12]
  PIN cpu_addr_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 632.590 0.000 632.870 4.000 ;
    END
  END cpu_addr_e[13]
  PIN cpu_addr_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END cpu_addr_e[14]
  PIN cpu_addr_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 654.670 0.000 654.950 4.000 ;
    END
  END cpu_addr_e[15]
  PIN cpu_addr_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END cpu_addr_e[1]
  PIN cpu_addr_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END cpu_addr_e[2]
  PIN cpu_addr_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END cpu_addr_e[3]
  PIN cpu_addr_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END cpu_addr_e[4]
  PIN cpu_addr_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END cpu_addr_e[5]
  PIN cpu_addr_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END cpu_addr_e[6]
  PIN cpu_addr_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END cpu_addr_e[7]
  PIN cpu_addr_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END cpu_addr_e[8]
  PIN cpu_addr_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END cpu_addr_e[9]
  PIN cpu_addr_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.130 1196.000 379.410 1200.000 ;
    END
  END cpu_addr_n[0]
  PIN cpu_addr_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.530 1196.000 489.810 1200.000 ;
    END
  END cpu_addr_n[10]
  PIN cpu_addr_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 500.570 1196.000 500.850 1200.000 ;
    END
  END cpu_addr_n[11]
  PIN cpu_addr_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 511.610 1196.000 511.890 1200.000 ;
    END
  END cpu_addr_n[12]
  PIN cpu_addr_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 522.190 1196.000 522.470 1200.000 ;
    END
  END cpu_addr_n[13]
  PIN cpu_addr_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 533.230 1196.000 533.510 1200.000 ;
    END
  END cpu_addr_n[14]
  PIN cpu_addr_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 544.270 1196.000 544.550 1200.000 ;
    END
  END cpu_addr_n[15]
  PIN cpu_addr_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 390.170 1196.000 390.450 1200.000 ;
    END
  END cpu_addr_n[1]
  PIN cpu_addr_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.210 1196.000 401.490 1200.000 ;
    END
  END cpu_addr_n[2]
  PIN cpu_addr_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 412.250 1196.000 412.530 1200.000 ;
    END
  END cpu_addr_n[3]
  PIN cpu_addr_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.290 1196.000 423.570 1200.000 ;
    END
  END cpu_addr_n[4]
  PIN cpu_addr_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 434.330 1196.000 434.610 1200.000 ;
    END
  END cpu_addr_n[5]
  PIN cpu_addr_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.370 1196.000 445.650 1200.000 ;
    END
  END cpu_addr_n[6]
  PIN cpu_addr_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.410 1196.000 456.690 1200.000 ;
    END
  END cpu_addr_n[7]
  PIN cpu_addr_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 467.450 1196.000 467.730 1200.000 ;
    END
  END cpu_addr_n[8]
  PIN cpu_addr_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 478.490 1196.000 478.770 1200.000 ;
    END
  END cpu_addr_n[9]
  PIN cpu_dtr_e0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END cpu_dtr_e0[0]
  PIN cpu_dtr_e0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END cpu_dtr_e0[10]
  PIN cpu_dtr_e0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END cpu_dtr_e0[11]
  PIN cpu_dtr_e0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END cpu_dtr_e0[12]
  PIN cpu_dtr_e0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END cpu_dtr_e0[13]
  PIN cpu_dtr_e0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END cpu_dtr_e0[14]
  PIN cpu_dtr_e0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END cpu_dtr_e0[15]
  PIN cpu_dtr_e0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END cpu_dtr_e0[16]
  PIN cpu_dtr_e0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END cpu_dtr_e0[17]
  PIN cpu_dtr_e0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END cpu_dtr_e0[18]
  PIN cpu_dtr_e0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END cpu_dtr_e0[19]
  PIN cpu_dtr_e0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END cpu_dtr_e0[1]
  PIN cpu_dtr_e0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END cpu_dtr_e0[20]
  PIN cpu_dtr_e0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END cpu_dtr_e0[21]
  PIN cpu_dtr_e0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END cpu_dtr_e0[22]
  PIN cpu_dtr_e0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END cpu_dtr_e0[23]
  PIN cpu_dtr_e0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END cpu_dtr_e0[24]
  PIN cpu_dtr_e0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END cpu_dtr_e0[25]
  PIN cpu_dtr_e0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END cpu_dtr_e0[26]
  PIN cpu_dtr_e0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END cpu_dtr_e0[27]
  PIN cpu_dtr_e0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END cpu_dtr_e0[28]
  PIN cpu_dtr_e0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END cpu_dtr_e0[29]
  PIN cpu_dtr_e0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END cpu_dtr_e0[2]
  PIN cpu_dtr_e0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END cpu_dtr_e0[30]
  PIN cpu_dtr_e0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END cpu_dtr_e0[31]
  PIN cpu_dtr_e0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END cpu_dtr_e0[3]
  PIN cpu_dtr_e0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END cpu_dtr_e0[4]
  PIN cpu_dtr_e0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END cpu_dtr_e0[5]
  PIN cpu_dtr_e0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END cpu_dtr_e0[6]
  PIN cpu_dtr_e0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END cpu_dtr_e0[7]
  PIN cpu_dtr_e0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END cpu_dtr_e0[8]
  PIN cpu_dtr_e0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END cpu_dtr_e0[9]
  PIN cpu_dtr_e1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END cpu_dtr_e1[0]
  PIN cpu_dtr_e1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 951.830 0.000 952.110 4.000 ;
    END
  END cpu_dtr_e1[10]
  PIN cpu_dtr_e1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END cpu_dtr_e1[11]
  PIN cpu_dtr_e1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 973.910 0.000 974.190 4.000 ;
    END
  END cpu_dtr_e1[12]
  PIN cpu_dtr_e1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.950 0.000 985.230 4.000 ;
    END
  END cpu_dtr_e1[13]
  PIN cpu_dtr_e1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 995.990 0.000 996.270 4.000 ;
    END
  END cpu_dtr_e1[14]
  PIN cpu_dtr_e1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.030 0.000 1007.310 4.000 ;
    END
  END cpu_dtr_e1[15]
  PIN cpu_dtr_e1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1018.070 0.000 1018.350 4.000 ;
    END
  END cpu_dtr_e1[16]
  PIN cpu_dtr_e1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1029.110 0.000 1029.390 4.000 ;
    END
  END cpu_dtr_e1[17]
  PIN cpu_dtr_e1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1039.690 0.000 1039.970 4.000 ;
    END
  END cpu_dtr_e1[18]
  PIN cpu_dtr_e1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1050.730 0.000 1051.010 4.000 ;
    END
  END cpu_dtr_e1[19]
  PIN cpu_dtr_e1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 852.930 0.000 853.210 4.000 ;
    END
  END cpu_dtr_e1[1]
  PIN cpu_dtr_e1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.770 0.000 1062.050 4.000 ;
    END
  END cpu_dtr_e1[20]
  PIN cpu_dtr_e1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1072.810 0.000 1073.090 4.000 ;
    END
  END cpu_dtr_e1[21]
  PIN cpu_dtr_e1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.850 0.000 1084.130 4.000 ;
    END
  END cpu_dtr_e1[22]
  PIN cpu_dtr_e1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.890 0.000 1095.170 4.000 ;
    END
  END cpu_dtr_e1[23]
  PIN cpu_dtr_e1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1105.930 0.000 1106.210 4.000 ;
    END
  END cpu_dtr_e1[24]
  PIN cpu_dtr_e1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1116.970 0.000 1117.250 4.000 ;
    END
  END cpu_dtr_e1[25]
  PIN cpu_dtr_e1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1128.010 0.000 1128.290 4.000 ;
    END
  END cpu_dtr_e1[26]
  PIN cpu_dtr_e1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1139.050 0.000 1139.330 4.000 ;
    END
  END cpu_dtr_e1[27]
  PIN cpu_dtr_e1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.090 0.000 1150.370 4.000 ;
    END
  END cpu_dtr_e1[28]
  PIN cpu_dtr_e1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1161.130 0.000 1161.410 4.000 ;
    END
  END cpu_dtr_e1[29]
  PIN cpu_dtr_e1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 863.510 0.000 863.790 4.000 ;
    END
  END cpu_dtr_e1[2]
  PIN cpu_dtr_e1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1172.170 0.000 1172.450 4.000 ;
    END
  END cpu_dtr_e1[30]
  PIN cpu_dtr_e1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1183.210 0.000 1183.490 4.000 ;
    END
  END cpu_dtr_e1[31]
  PIN cpu_dtr_e1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 874.550 0.000 874.830 4.000 ;
    END
  END cpu_dtr_e1[3]
  PIN cpu_dtr_e1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END cpu_dtr_e1[4]
  PIN cpu_dtr_e1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.630 0.000 896.910 4.000 ;
    END
  END cpu_dtr_e1[5]
  PIN cpu_dtr_e1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 907.670 0.000 907.950 4.000 ;
    END
  END cpu_dtr_e1[6]
  PIN cpu_dtr_e1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.710 0.000 918.990 4.000 ;
    END
  END cpu_dtr_e1[7]
  PIN cpu_dtr_e1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.750 0.000 930.030 4.000 ;
    END
  END cpu_dtr_e1[8]
  PIN cpu_dtr_e1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 940.790 0.000 941.070 4.000 ;
    END
  END cpu_dtr_e1[9]
  PIN cpu_dtr_n0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 1196.000 27.050 1200.000 ;
    END
  END cpu_dtr_n0[0]
  PIN cpu_dtr_n0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.170 1196.000 137.450 1200.000 ;
    END
  END cpu_dtr_n0[10]
  PIN cpu_dtr_n0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.210 1196.000 148.490 1200.000 ;
    END
  END cpu_dtr_n0[11]
  PIN cpu_dtr_n0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 1196.000 159.530 1200.000 ;
    END
  END cpu_dtr_n0[12]
  PIN cpu_dtr_n0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 1196.000 170.570 1200.000 ;
    END
  END cpu_dtr_n0[13]
  PIN cpu_dtr_n0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.870 1196.000 181.150 1200.000 ;
    END
  END cpu_dtr_n0[14]
  PIN cpu_dtr_n0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.910 1196.000 192.190 1200.000 ;
    END
  END cpu_dtr_n0[15]
  PIN cpu_dtr_n0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.950 1196.000 203.230 1200.000 ;
    END
  END cpu_dtr_n0[16]
  PIN cpu_dtr_n0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.990 1196.000 214.270 1200.000 ;
    END
  END cpu_dtr_n0[17]
  PIN cpu_dtr_n0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 225.030 1196.000 225.310 1200.000 ;
    END
  END cpu_dtr_n0[18]
  PIN cpu_dtr_n0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.070 1196.000 236.350 1200.000 ;
    END
  END cpu_dtr_n0[19]
  PIN cpu_dtr_n0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 1196.000 38.090 1200.000 ;
    END
  END cpu_dtr_n0[1]
  PIN cpu_dtr_n0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.110 1196.000 247.390 1200.000 ;
    END
  END cpu_dtr_n0[20]
  PIN cpu_dtr_n0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.150 1196.000 258.430 1200.000 ;
    END
  END cpu_dtr_n0[21]
  PIN cpu_dtr_n0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.190 1196.000 269.470 1200.000 ;
    END
  END cpu_dtr_n0[22]
  PIN cpu_dtr_n0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 280.230 1196.000 280.510 1200.000 ;
    END
  END cpu_dtr_n0[23]
  PIN cpu_dtr_n0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.270 1196.000 291.550 1200.000 ;
    END
  END cpu_dtr_n0[24]
  PIN cpu_dtr_n0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.310 1196.000 302.590 1200.000 ;
    END
  END cpu_dtr_n0[25]
  PIN cpu_dtr_n0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 313.350 1196.000 313.630 1200.000 ;
    END
  END cpu_dtr_n0[26]
  PIN cpu_dtr_n0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 324.390 1196.000 324.670 1200.000 ;
    END
  END cpu_dtr_n0[27]
  PIN cpu_dtr_n0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.430 1196.000 335.710 1200.000 ;
    END
  END cpu_dtr_n0[28]
  PIN cpu_dtr_n0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 346.470 1196.000 346.750 1200.000 ;
    END
  END cpu_dtr_n0[29]
  PIN cpu_dtr_n0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 1196.000 49.130 1200.000 ;
    END
  END cpu_dtr_n0[2]
  PIN cpu_dtr_n0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.050 1196.000 357.330 1200.000 ;
    END
  END cpu_dtr_n0[30]
  PIN cpu_dtr_n0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 368.090 1196.000 368.370 1200.000 ;
    END
  END cpu_dtr_n0[31]
  PIN cpu_dtr_n0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 1196.000 60.170 1200.000 ;
    END
  END cpu_dtr_n0[3]
  PIN cpu_dtr_n0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 1196.000 71.210 1200.000 ;
    END
  END cpu_dtr_n0[4]
  PIN cpu_dtr_n0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.970 1196.000 82.250 1200.000 ;
    END
  END cpu_dtr_n0[5]
  PIN cpu_dtr_n0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.010 1196.000 93.290 1200.000 ;
    END
  END cpu_dtr_n0[6]
  PIN cpu_dtr_n0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.050 1196.000 104.330 1200.000 ;
    END
  END cpu_dtr_n0[7]
  PIN cpu_dtr_n0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 1196.000 115.370 1200.000 ;
    END
  END cpu_dtr_n0[8]
  PIN cpu_dtr_n0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.130 1196.000 126.410 1200.000 ;
    END
  END cpu_dtr_n0[9]
  PIN cpu_dtr_n1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 841.890 1196.000 842.170 1200.000 ;
    END
  END cpu_dtr_n1[0]
  PIN cpu_dtr_n1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 951.830 1196.000 952.110 1200.000 ;
    END
  END cpu_dtr_n1[10]
  PIN cpu_dtr_n1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 962.870 1196.000 963.150 1200.000 ;
    END
  END cpu_dtr_n1[11]
  PIN cpu_dtr_n1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 973.910 1196.000 974.190 1200.000 ;
    END
  END cpu_dtr_n1[12]
  PIN cpu_dtr_n1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.950 1196.000 985.230 1200.000 ;
    END
  END cpu_dtr_n1[13]
  PIN cpu_dtr_n1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 995.990 1196.000 996.270 1200.000 ;
    END
  END cpu_dtr_n1[14]
  PIN cpu_dtr_n1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.030 1196.000 1007.310 1200.000 ;
    END
  END cpu_dtr_n1[15]
  PIN cpu_dtr_n1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1018.070 1196.000 1018.350 1200.000 ;
    END
  END cpu_dtr_n1[16]
  PIN cpu_dtr_n1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1029.110 1196.000 1029.390 1200.000 ;
    END
  END cpu_dtr_n1[17]
  PIN cpu_dtr_n1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1039.690 1196.000 1039.970 1200.000 ;
    END
  END cpu_dtr_n1[18]
  PIN cpu_dtr_n1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1050.730 1196.000 1051.010 1200.000 ;
    END
  END cpu_dtr_n1[19]
  PIN cpu_dtr_n1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 852.930 1196.000 853.210 1200.000 ;
    END
  END cpu_dtr_n1[1]
  PIN cpu_dtr_n1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.770 1196.000 1062.050 1200.000 ;
    END
  END cpu_dtr_n1[20]
  PIN cpu_dtr_n1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1072.810 1196.000 1073.090 1200.000 ;
    END
  END cpu_dtr_n1[21]
  PIN cpu_dtr_n1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.850 1196.000 1084.130 1200.000 ;
    END
  END cpu_dtr_n1[22]
  PIN cpu_dtr_n1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.890 1196.000 1095.170 1200.000 ;
    END
  END cpu_dtr_n1[23]
  PIN cpu_dtr_n1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1105.930 1196.000 1106.210 1200.000 ;
    END
  END cpu_dtr_n1[24]
  PIN cpu_dtr_n1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1116.970 1196.000 1117.250 1200.000 ;
    END
  END cpu_dtr_n1[25]
  PIN cpu_dtr_n1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1128.010 1196.000 1128.290 1200.000 ;
    END
  END cpu_dtr_n1[26]
  PIN cpu_dtr_n1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1139.050 1196.000 1139.330 1200.000 ;
    END
  END cpu_dtr_n1[27]
  PIN cpu_dtr_n1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.090 1196.000 1150.370 1200.000 ;
    END
  END cpu_dtr_n1[28]
  PIN cpu_dtr_n1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1161.130 1196.000 1161.410 1200.000 ;
    END
  END cpu_dtr_n1[29]
  PIN cpu_dtr_n1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 863.510 1196.000 863.790 1200.000 ;
    END
  END cpu_dtr_n1[2]
  PIN cpu_dtr_n1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1172.170 1196.000 1172.450 1200.000 ;
    END
  END cpu_dtr_n1[30]
  PIN cpu_dtr_n1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1183.210 1196.000 1183.490 1200.000 ;
    END
  END cpu_dtr_n1[31]
  PIN cpu_dtr_n1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 874.550 1196.000 874.830 1200.000 ;
    END
  END cpu_dtr_n1[3]
  PIN cpu_dtr_n1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 885.590 1196.000 885.870 1200.000 ;
    END
  END cpu_dtr_n1[4]
  PIN cpu_dtr_n1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.630 1196.000 896.910 1200.000 ;
    END
  END cpu_dtr_n1[5]
  PIN cpu_dtr_n1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 907.670 1196.000 907.950 1200.000 ;
    END
  END cpu_dtr_n1[6]
  PIN cpu_dtr_n1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.710 1196.000 918.990 1200.000 ;
    END
  END cpu_dtr_n1[7]
  PIN cpu_dtr_n1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.750 1196.000 930.030 1200.000 ;
    END
  END cpu_dtr_n1[8]
  PIN cpu_dtr_n1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 940.790 1196.000 941.070 1200.000 ;
    END
  END cpu_dtr_n1[9]
  PIN cpu_dtw_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END cpu_dtw_e[0]
  PIN cpu_dtw_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END cpu_dtw_e[10]
  PIN cpu_dtw_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END cpu_dtw_e[11]
  PIN cpu_dtw_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END cpu_dtw_e[12]
  PIN cpu_dtw_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 808.770 0.000 809.050 4.000 ;
    END
  END cpu_dtw_e[13]
  PIN cpu_dtw_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END cpu_dtw_e[14]
  PIN cpu_dtw_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END cpu_dtw_e[15]
  PIN cpu_dtw_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END cpu_dtw_e[1]
  PIN cpu_dtw_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 687.790 0.000 688.070 4.000 ;
    END
  END cpu_dtw_e[2]
  PIN cpu_dtw_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END cpu_dtw_e[3]
  PIN cpu_dtw_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END cpu_dtw_e[4]
  PIN cpu_dtw_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END cpu_dtw_e[5]
  PIN cpu_dtw_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END cpu_dtw_e[6]
  PIN cpu_dtw_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 742.530 0.000 742.810 4.000 ;
    END
  END cpu_dtw_e[7]
  PIN cpu_dtw_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END cpu_dtw_e[8]
  PIN cpu_dtw_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END cpu_dtw_e[9]
  PIN cpu_dtw_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 665.710 1196.000 665.990 1200.000 ;
    END
  END cpu_dtw_n[0]
  PIN cpu_dtw_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 775.650 1196.000 775.930 1200.000 ;
    END
  END cpu_dtw_n[10]
  PIN cpu_dtw_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.690 1196.000 786.970 1200.000 ;
    END
  END cpu_dtw_n[11]
  PIN cpu_dtw_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 797.730 1196.000 798.010 1200.000 ;
    END
  END cpu_dtw_n[12]
  PIN cpu_dtw_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 808.770 1196.000 809.050 1200.000 ;
    END
  END cpu_dtw_n[13]
  PIN cpu_dtw_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 819.810 1196.000 820.090 1200.000 ;
    END
  END cpu_dtw_n[14]
  PIN cpu_dtw_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 830.850 1196.000 831.130 1200.000 ;
    END
  END cpu_dtw_n[15]
  PIN cpu_dtw_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 676.750 1196.000 677.030 1200.000 ;
    END
  END cpu_dtw_n[1]
  PIN cpu_dtw_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 687.790 1196.000 688.070 1200.000 ;
    END
  END cpu_dtw_n[2]
  PIN cpu_dtw_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 698.370 1196.000 698.650 1200.000 ;
    END
  END cpu_dtw_n[3]
  PIN cpu_dtw_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 709.410 1196.000 709.690 1200.000 ;
    END
  END cpu_dtw_n[4]
  PIN cpu_dtw_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 720.450 1196.000 720.730 1200.000 ;
    END
  END cpu_dtw_n[5]
  PIN cpu_dtw_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.490 1196.000 731.770 1200.000 ;
    END
  END cpu_dtw_n[6]
  PIN cpu_dtw_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 742.530 1196.000 742.810 1200.000 ;
    END
  END cpu_dtw_n[7]
  PIN cpu_dtw_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 753.570 1196.000 753.850 1200.000 ;
    END
  END cpu_dtw_n[8]
  PIN cpu_dtw_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 764.610 1196.000 764.890 1200.000 ;
    END
  END cpu_dtw_n[9]
  PIN cpu_mask_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END cpu_mask_e[0]
  PIN cpu_mask_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END cpu_mask_e[1]
  PIN cpu_mask_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END cpu_mask_e[2]
  PIN cpu_mask_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END cpu_mask_e[3]
  PIN cpu_mask_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END cpu_mask_e[4]
  PIN cpu_mask_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END cpu_mask_e[5]
  PIN cpu_mask_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END cpu_mask_e[6]
  PIN cpu_mask_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END cpu_mask_e[7]
  PIN cpu_mask_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.310 1196.000 555.590 1200.000 ;
    END
  END cpu_mask_n[0]
  PIN cpu_mask_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 566.350 1196.000 566.630 1200.000 ;
    END
  END cpu_mask_n[1]
  PIN cpu_mask_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 577.390 1196.000 577.670 1200.000 ;
    END
  END cpu_mask_n[2]
  PIN cpu_mask_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 588.430 1196.000 588.710 1200.000 ;
    END
  END cpu_mask_n[3]
  PIN cpu_mask_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 599.470 1196.000 599.750 1200.000 ;
    END
  END cpu_mask_n[4]
  PIN cpu_mask_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 610.510 1196.000 610.790 1200.000 ;
    END
  END cpu_mask_n[5]
  PIN cpu_mask_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 621.550 1196.000 621.830 1200.000 ;
    END
  END cpu_mask_n[6]
  PIN cpu_mask_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 632.590 1196.000 632.870 1200.000 ;
    END
  END cpu_mask_n[7]
  PIN cpu_wen_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END cpu_wen_e[0]
  PIN cpu_wen_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END cpu_wen_e[1]
  PIN cpu_wen_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 643.630 1196.000 643.910 1200.000 ;
    END
  END cpu_wen_n[0]
  PIN cpu_wen_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 654.670 1196.000 654.950 1200.000 ;
    END
  END cpu_wen_n[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 4.800 1200.000 5.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 320.320 1200.000 320.920 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 351.600 1200.000 352.200 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 383.560 1200.000 384.160 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 414.840 1200.000 415.440 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 446.800 1200.000 447.400 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 478.080 1200.000 478.680 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 510.040 1200.000 510.640 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 541.320 1200.000 541.920 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 573.280 1200.000 573.880 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 604.560 1200.000 605.160 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 36.080 1200.000 36.680 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 635.840 1200.000 636.440 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 667.800 1200.000 668.400 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 699.080 1200.000 699.680 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 731.040 1200.000 731.640 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 762.320 1200.000 762.920 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 794.280 1200.000 794.880 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 825.560 1200.000 826.160 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 857.520 1200.000 858.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 888.800 1200.000 889.400 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 920.080 1200.000 920.680 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 67.360 1200.000 67.960 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 952.040 1200.000 952.640 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 983.320 1200.000 983.920 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1015.280 1200.000 1015.880 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1046.560 1200.000 1047.160 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1078.520 1200.000 1079.120 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1109.800 1200.000 1110.400 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1141.760 1200.000 1142.360 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1173.040 1200.000 1173.640 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 99.320 1200.000 99.920 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 130.600 1200.000 131.200 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 162.560 1200.000 163.160 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 193.840 1200.000 194.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 225.800 1200.000 226.400 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 257.080 1200.000 257.680 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 289.040 1200.000 289.640 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 15.000 1200.000 15.600 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 330.520 1200.000 331.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 362.480 1200.000 363.080 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 393.760 1200.000 394.360 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 425.720 1200.000 426.320 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 457.000 1200.000 457.600 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 488.960 1200.000 489.560 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 520.240 1200.000 520.840 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 552.200 1200.000 552.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 583.480 1200.000 584.080 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 614.760 1200.000 615.360 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 46.280 1200.000 46.880 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 646.720 1200.000 647.320 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 678.000 1200.000 678.600 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 709.960 1200.000 710.560 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 741.240 1200.000 741.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 773.200 1200.000 773.800 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 804.480 1200.000 805.080 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 836.440 1200.000 837.040 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 867.720 1200.000 868.320 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 899.680 1200.000 900.280 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 930.960 1200.000 931.560 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 78.240 1200.000 78.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 962.240 1200.000 962.840 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 994.200 1200.000 994.800 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1025.480 1200.000 1026.080 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1057.440 1200.000 1058.040 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1088.720 1200.000 1089.320 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1120.680 1200.000 1121.280 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1151.960 1200.000 1152.560 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1183.920 1200.000 1184.520 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 109.520 1200.000 110.120 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 141.480 1200.000 142.080 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 172.760 1200.000 173.360 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 204.720 1200.000 205.320 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 236.000 1200.000 236.600 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 267.960 1200.000 268.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 299.240 1200.000 299.840 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 25.200 1200.000 25.800 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 341.400 1200.000 342.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 372.680 1200.000 373.280 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 404.640 1200.000 405.240 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 435.920 1200.000 436.520 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 467.880 1200.000 468.480 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 499.160 1200.000 499.760 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 531.120 1200.000 531.720 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 562.400 1200.000 563.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 594.360 1200.000 594.960 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 625.640 1200.000 626.240 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 57.160 1200.000 57.760 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 656.920 1200.000 657.520 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 688.880 1200.000 689.480 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 720.160 1200.000 720.760 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 752.120 1200.000 752.720 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 783.400 1200.000 784.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 815.360 1200.000 815.960 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 846.640 1200.000 847.240 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 878.600 1200.000 879.200 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 909.880 1200.000 910.480 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 941.160 1200.000 941.760 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 88.440 1200.000 89.040 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 973.120 1200.000 973.720 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1004.400 1200.000 1005.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1036.360 1200.000 1036.960 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1067.640 1200.000 1068.240 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1099.600 1200.000 1100.200 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1130.880 1200.000 1131.480 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1162.840 1200.000 1163.440 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1194.120 1200.000 1194.720 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 120.400 1200.000 121.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 151.680 1200.000 152.280 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 183.640 1200.000 184.240 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 214.920 1200.000 215.520 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 246.880 1200.000 247.480 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 278.160 1200.000 278.760 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 309.440 1200.000 310.040 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1130.200 4.000 1130.800 ;
    END
  END la_data_in[0]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.160 4.000 1162.760 ;
    END
  END la_data_in[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.080 4.000 1141.680 ;
    END
  END la_data_out[0]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END la_data_out[1]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.120 4.000 1194.720 ;
    END
  END la_data_out[2]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1151.280 4.000 1151.880 ;
    END
  END la_oen[0]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.240 4.000 1183.840 ;
    END
  END la_oen[1]
  PIN one_e
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END one_e
  PIN one_n
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.730 1196.000 16.010 1200.000 ;
    END
  END one_n
  PIN ram_ce_e
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1194.250 0.000 1194.530 4.000 ;
    END
  END ram_ce_e
  PIN ram_ce_n
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1194.250 1196.000 1194.530 1200.000 ;
    END
  END ram_ce_n
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.000 4.000 780.600 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.960 4.000 812.560 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.200 4.000 875.800 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.160 4.000 907.760 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.120 4.000 939.720 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.080 4.000 971.680 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1035.000 4.000 1035.600 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.280 4.000 1066.880 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.240 4.000 1098.840 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.920 4.000 504.520 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.960 4.000 727.560 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.200 4.000 790.800 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.160 4.000 822.760 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.120 4.000 854.720 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.080 4.000 886.680 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.000 4.000 950.600 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 981.280 4.000 981.880 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.200 4.000 1045.800 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.160 4.000 1077.760 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.120 4.000 1109.720 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.080 4.000 376.680 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.880 4.000 451.480 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.160 4.000 482.760 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.080 4.000 546.680 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.000 4.000 610.600 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.920 4.000 674.520 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.200 4.000 705.800 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 4.000 737.760 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.120 4.000 769.720 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.080 4.000 801.680 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.960 4.000 897.560 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.200 4.000 960.800 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.160 4.000 992.760 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.120 4.000 1024.720 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.080 4.000 1056.680 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.000 4.000 1120.600 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wbs_we_i
  PIN zero_e
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END zero_e
  PIN zero_n
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.150 1196.000 5.430 1200.000 ;
    END
  END zero_n
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1188.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1194.935 1188.725 ;
      LAYER met1 ;
        RECT 4.670 4.460 1195.010 1192.000 ;
      LAYER met2 ;
        RECT 4.690 1195.720 4.870 1196.000 ;
        RECT 5.710 1195.720 15.450 1196.000 ;
        RECT 16.290 1195.720 26.490 1196.000 ;
        RECT 27.330 1195.720 37.530 1196.000 ;
        RECT 38.370 1195.720 48.570 1196.000 ;
        RECT 49.410 1195.720 59.610 1196.000 ;
        RECT 60.450 1195.720 70.650 1196.000 ;
        RECT 71.490 1195.720 81.690 1196.000 ;
        RECT 82.530 1195.720 92.730 1196.000 ;
        RECT 93.570 1195.720 103.770 1196.000 ;
        RECT 104.610 1195.720 114.810 1196.000 ;
        RECT 115.650 1195.720 125.850 1196.000 ;
        RECT 126.690 1195.720 136.890 1196.000 ;
        RECT 137.730 1195.720 147.930 1196.000 ;
        RECT 148.770 1195.720 158.970 1196.000 ;
        RECT 159.810 1195.720 170.010 1196.000 ;
        RECT 170.850 1195.720 180.590 1196.000 ;
        RECT 181.430 1195.720 191.630 1196.000 ;
        RECT 192.470 1195.720 202.670 1196.000 ;
        RECT 203.510 1195.720 213.710 1196.000 ;
        RECT 214.550 1195.720 224.750 1196.000 ;
        RECT 225.590 1195.720 235.790 1196.000 ;
        RECT 236.630 1195.720 246.830 1196.000 ;
        RECT 247.670 1195.720 257.870 1196.000 ;
        RECT 258.710 1195.720 268.910 1196.000 ;
        RECT 269.750 1195.720 279.950 1196.000 ;
        RECT 280.790 1195.720 290.990 1196.000 ;
        RECT 291.830 1195.720 302.030 1196.000 ;
        RECT 302.870 1195.720 313.070 1196.000 ;
        RECT 313.910 1195.720 324.110 1196.000 ;
        RECT 324.950 1195.720 335.150 1196.000 ;
        RECT 335.990 1195.720 346.190 1196.000 ;
        RECT 347.030 1195.720 356.770 1196.000 ;
        RECT 357.610 1195.720 367.810 1196.000 ;
        RECT 368.650 1195.720 378.850 1196.000 ;
        RECT 379.690 1195.720 389.890 1196.000 ;
        RECT 390.730 1195.720 400.930 1196.000 ;
        RECT 401.770 1195.720 411.970 1196.000 ;
        RECT 412.810 1195.720 423.010 1196.000 ;
        RECT 423.850 1195.720 434.050 1196.000 ;
        RECT 434.890 1195.720 445.090 1196.000 ;
        RECT 445.930 1195.720 456.130 1196.000 ;
        RECT 456.970 1195.720 467.170 1196.000 ;
        RECT 468.010 1195.720 478.210 1196.000 ;
        RECT 479.050 1195.720 489.250 1196.000 ;
        RECT 490.090 1195.720 500.290 1196.000 ;
        RECT 501.130 1195.720 511.330 1196.000 ;
        RECT 512.170 1195.720 521.910 1196.000 ;
        RECT 522.750 1195.720 532.950 1196.000 ;
        RECT 533.790 1195.720 543.990 1196.000 ;
        RECT 544.830 1195.720 555.030 1196.000 ;
        RECT 555.870 1195.720 566.070 1196.000 ;
        RECT 566.910 1195.720 577.110 1196.000 ;
        RECT 577.950 1195.720 588.150 1196.000 ;
        RECT 588.990 1195.720 599.190 1196.000 ;
        RECT 600.030 1195.720 610.230 1196.000 ;
        RECT 611.070 1195.720 621.270 1196.000 ;
        RECT 622.110 1195.720 632.310 1196.000 ;
        RECT 633.150 1195.720 643.350 1196.000 ;
        RECT 644.190 1195.720 654.390 1196.000 ;
        RECT 655.230 1195.720 665.430 1196.000 ;
        RECT 666.270 1195.720 676.470 1196.000 ;
        RECT 677.310 1195.720 687.510 1196.000 ;
        RECT 688.350 1195.720 698.090 1196.000 ;
        RECT 698.930 1195.720 709.130 1196.000 ;
        RECT 709.970 1195.720 720.170 1196.000 ;
        RECT 721.010 1195.720 731.210 1196.000 ;
        RECT 732.050 1195.720 742.250 1196.000 ;
        RECT 743.090 1195.720 753.290 1196.000 ;
        RECT 754.130 1195.720 764.330 1196.000 ;
        RECT 765.170 1195.720 775.370 1196.000 ;
        RECT 776.210 1195.720 786.410 1196.000 ;
        RECT 787.250 1195.720 797.450 1196.000 ;
        RECT 798.290 1195.720 808.490 1196.000 ;
        RECT 809.330 1195.720 819.530 1196.000 ;
        RECT 820.370 1195.720 830.570 1196.000 ;
        RECT 831.410 1195.720 841.610 1196.000 ;
        RECT 842.450 1195.720 852.650 1196.000 ;
        RECT 853.490 1195.720 863.230 1196.000 ;
        RECT 864.070 1195.720 874.270 1196.000 ;
        RECT 875.110 1195.720 885.310 1196.000 ;
        RECT 886.150 1195.720 896.350 1196.000 ;
        RECT 897.190 1195.720 907.390 1196.000 ;
        RECT 908.230 1195.720 918.430 1196.000 ;
        RECT 919.270 1195.720 929.470 1196.000 ;
        RECT 930.310 1195.720 940.510 1196.000 ;
        RECT 941.350 1195.720 951.550 1196.000 ;
        RECT 952.390 1195.720 962.590 1196.000 ;
        RECT 963.430 1195.720 973.630 1196.000 ;
        RECT 974.470 1195.720 984.670 1196.000 ;
        RECT 985.510 1195.720 995.710 1196.000 ;
        RECT 996.550 1195.720 1006.750 1196.000 ;
        RECT 1007.590 1195.720 1017.790 1196.000 ;
        RECT 1018.630 1195.720 1028.830 1196.000 ;
        RECT 1029.670 1195.720 1039.410 1196.000 ;
        RECT 1040.250 1195.720 1050.450 1196.000 ;
        RECT 1051.290 1195.720 1061.490 1196.000 ;
        RECT 1062.330 1195.720 1072.530 1196.000 ;
        RECT 1073.370 1195.720 1083.570 1196.000 ;
        RECT 1084.410 1195.720 1094.610 1196.000 ;
        RECT 1095.450 1195.720 1105.650 1196.000 ;
        RECT 1106.490 1195.720 1116.690 1196.000 ;
        RECT 1117.530 1195.720 1127.730 1196.000 ;
        RECT 1128.570 1195.720 1138.770 1196.000 ;
        RECT 1139.610 1195.720 1149.810 1196.000 ;
        RECT 1150.650 1195.720 1160.850 1196.000 ;
        RECT 1161.690 1195.720 1171.890 1196.000 ;
        RECT 1172.730 1195.720 1182.930 1196.000 ;
        RECT 1183.770 1195.720 1193.970 1196.000 ;
        RECT 1194.810 1195.720 1194.990 1196.000 ;
        RECT 4.690 4.280 1194.990 1195.720 ;
        RECT 4.690 4.000 4.870 4.280 ;
        RECT 5.710 4.000 15.450 4.280 ;
        RECT 16.290 4.000 26.490 4.280 ;
        RECT 27.330 4.000 37.530 4.280 ;
        RECT 38.370 4.000 48.570 4.280 ;
        RECT 49.410 4.000 59.610 4.280 ;
        RECT 60.450 4.000 70.650 4.280 ;
        RECT 71.490 4.000 81.690 4.280 ;
        RECT 82.530 4.000 92.730 4.280 ;
        RECT 93.570 4.000 103.770 4.280 ;
        RECT 104.610 4.000 114.810 4.280 ;
        RECT 115.650 4.000 125.850 4.280 ;
        RECT 126.690 4.000 136.890 4.280 ;
        RECT 137.730 4.000 147.930 4.280 ;
        RECT 148.770 4.000 158.970 4.280 ;
        RECT 159.810 4.000 170.010 4.280 ;
        RECT 170.850 4.000 180.590 4.280 ;
        RECT 181.430 4.000 191.630 4.280 ;
        RECT 192.470 4.000 202.670 4.280 ;
        RECT 203.510 4.000 213.710 4.280 ;
        RECT 214.550 4.000 224.750 4.280 ;
        RECT 225.590 4.000 235.790 4.280 ;
        RECT 236.630 4.000 246.830 4.280 ;
        RECT 247.670 4.000 257.870 4.280 ;
        RECT 258.710 4.000 268.910 4.280 ;
        RECT 269.750 4.000 279.950 4.280 ;
        RECT 280.790 4.000 290.990 4.280 ;
        RECT 291.830 4.000 302.030 4.280 ;
        RECT 302.870 4.000 313.070 4.280 ;
        RECT 313.910 4.000 324.110 4.280 ;
        RECT 324.950 4.000 335.150 4.280 ;
        RECT 335.990 4.000 346.190 4.280 ;
        RECT 347.030 4.000 356.770 4.280 ;
        RECT 357.610 4.000 367.810 4.280 ;
        RECT 368.650 4.000 378.850 4.280 ;
        RECT 379.690 4.000 389.890 4.280 ;
        RECT 390.730 4.000 400.930 4.280 ;
        RECT 401.770 4.000 411.970 4.280 ;
        RECT 412.810 4.000 423.010 4.280 ;
        RECT 423.850 4.000 434.050 4.280 ;
        RECT 434.890 4.000 445.090 4.280 ;
        RECT 445.930 4.000 456.130 4.280 ;
        RECT 456.970 4.000 467.170 4.280 ;
        RECT 468.010 4.000 478.210 4.280 ;
        RECT 479.050 4.000 489.250 4.280 ;
        RECT 490.090 4.000 500.290 4.280 ;
        RECT 501.130 4.000 511.330 4.280 ;
        RECT 512.170 4.000 521.910 4.280 ;
        RECT 522.750 4.000 532.950 4.280 ;
        RECT 533.790 4.000 543.990 4.280 ;
        RECT 544.830 4.000 555.030 4.280 ;
        RECT 555.870 4.000 566.070 4.280 ;
        RECT 566.910 4.000 577.110 4.280 ;
        RECT 577.950 4.000 588.150 4.280 ;
        RECT 588.990 4.000 599.190 4.280 ;
        RECT 600.030 4.000 610.230 4.280 ;
        RECT 611.070 4.000 621.270 4.280 ;
        RECT 622.110 4.000 632.310 4.280 ;
        RECT 633.150 4.000 643.350 4.280 ;
        RECT 644.190 4.000 654.390 4.280 ;
        RECT 655.230 4.000 665.430 4.280 ;
        RECT 666.270 4.000 676.470 4.280 ;
        RECT 677.310 4.000 687.510 4.280 ;
        RECT 688.350 4.000 698.090 4.280 ;
        RECT 698.930 4.000 709.130 4.280 ;
        RECT 709.970 4.000 720.170 4.280 ;
        RECT 721.010 4.000 731.210 4.280 ;
        RECT 732.050 4.000 742.250 4.280 ;
        RECT 743.090 4.000 753.290 4.280 ;
        RECT 754.130 4.000 764.330 4.280 ;
        RECT 765.170 4.000 775.370 4.280 ;
        RECT 776.210 4.000 786.410 4.280 ;
        RECT 787.250 4.000 797.450 4.280 ;
        RECT 798.290 4.000 808.490 4.280 ;
        RECT 809.330 4.000 819.530 4.280 ;
        RECT 820.370 4.000 830.570 4.280 ;
        RECT 831.410 4.000 841.610 4.280 ;
        RECT 842.450 4.000 852.650 4.280 ;
        RECT 853.490 4.000 863.230 4.280 ;
        RECT 864.070 4.000 874.270 4.280 ;
        RECT 875.110 4.000 885.310 4.280 ;
        RECT 886.150 4.000 896.350 4.280 ;
        RECT 897.190 4.000 907.390 4.280 ;
        RECT 908.230 4.000 918.430 4.280 ;
        RECT 919.270 4.000 929.470 4.280 ;
        RECT 930.310 4.000 940.510 4.280 ;
        RECT 941.350 4.000 951.550 4.280 ;
        RECT 952.390 4.000 962.590 4.280 ;
        RECT 963.430 4.000 973.630 4.280 ;
        RECT 974.470 4.000 984.670 4.280 ;
        RECT 985.510 4.000 995.710 4.280 ;
        RECT 996.550 4.000 1006.750 4.280 ;
        RECT 1007.590 4.000 1017.790 4.280 ;
        RECT 1018.630 4.000 1028.830 4.280 ;
        RECT 1029.670 4.000 1039.410 4.280 ;
        RECT 1040.250 4.000 1050.450 4.280 ;
        RECT 1051.290 4.000 1061.490 4.280 ;
        RECT 1062.330 4.000 1072.530 4.280 ;
        RECT 1073.370 4.000 1083.570 4.280 ;
        RECT 1084.410 4.000 1094.610 4.280 ;
        RECT 1095.450 4.000 1105.650 4.280 ;
        RECT 1106.490 4.000 1116.690 4.280 ;
        RECT 1117.530 4.000 1127.730 4.280 ;
        RECT 1128.570 4.000 1138.770 4.280 ;
        RECT 1139.610 4.000 1149.810 4.280 ;
        RECT 1150.650 4.000 1160.850 4.280 ;
        RECT 1161.690 4.000 1171.890 4.280 ;
        RECT 1172.730 4.000 1182.930 4.280 ;
        RECT 1183.770 4.000 1193.970 4.280 ;
        RECT 1194.810 4.000 1194.990 4.280 ;
      LAYER met3 ;
        RECT 3.990 1195.120 1196.000 1195.945 ;
        RECT 4.400 1193.720 1195.600 1195.120 ;
        RECT 3.990 1184.920 1196.000 1193.720 ;
        RECT 3.990 1184.240 1195.600 1184.920 ;
        RECT 4.400 1183.520 1195.600 1184.240 ;
        RECT 4.400 1182.840 1196.000 1183.520 ;
        RECT 3.990 1174.040 1196.000 1182.840 ;
        RECT 4.400 1172.640 1195.600 1174.040 ;
        RECT 3.990 1163.840 1196.000 1172.640 ;
        RECT 3.990 1163.160 1195.600 1163.840 ;
        RECT 4.400 1162.440 1195.600 1163.160 ;
        RECT 4.400 1161.760 1196.000 1162.440 ;
        RECT 3.990 1152.960 1196.000 1161.760 ;
        RECT 3.990 1152.280 1195.600 1152.960 ;
        RECT 4.400 1151.560 1195.600 1152.280 ;
        RECT 4.400 1150.880 1196.000 1151.560 ;
        RECT 3.990 1142.760 1196.000 1150.880 ;
        RECT 3.990 1142.080 1195.600 1142.760 ;
        RECT 4.400 1141.360 1195.600 1142.080 ;
        RECT 4.400 1140.680 1196.000 1141.360 ;
        RECT 3.990 1131.880 1196.000 1140.680 ;
        RECT 3.990 1131.200 1195.600 1131.880 ;
        RECT 4.400 1130.480 1195.600 1131.200 ;
        RECT 4.400 1129.800 1196.000 1130.480 ;
        RECT 3.990 1121.680 1196.000 1129.800 ;
        RECT 3.990 1121.000 1195.600 1121.680 ;
        RECT 4.400 1120.280 1195.600 1121.000 ;
        RECT 4.400 1119.600 1196.000 1120.280 ;
        RECT 3.990 1110.800 1196.000 1119.600 ;
        RECT 3.990 1110.120 1195.600 1110.800 ;
        RECT 4.400 1109.400 1195.600 1110.120 ;
        RECT 4.400 1108.720 1196.000 1109.400 ;
        RECT 3.990 1100.600 1196.000 1108.720 ;
        RECT 3.990 1099.240 1195.600 1100.600 ;
        RECT 4.400 1099.200 1195.600 1099.240 ;
        RECT 4.400 1097.840 1196.000 1099.200 ;
        RECT 3.990 1089.720 1196.000 1097.840 ;
        RECT 3.990 1089.040 1195.600 1089.720 ;
        RECT 4.400 1088.320 1195.600 1089.040 ;
        RECT 4.400 1087.640 1196.000 1088.320 ;
        RECT 3.990 1079.520 1196.000 1087.640 ;
        RECT 3.990 1078.160 1195.600 1079.520 ;
        RECT 4.400 1078.120 1195.600 1078.160 ;
        RECT 4.400 1076.760 1196.000 1078.120 ;
        RECT 3.990 1068.640 1196.000 1076.760 ;
        RECT 3.990 1067.280 1195.600 1068.640 ;
        RECT 4.400 1067.240 1195.600 1067.280 ;
        RECT 4.400 1065.880 1196.000 1067.240 ;
        RECT 3.990 1058.440 1196.000 1065.880 ;
        RECT 3.990 1057.080 1195.600 1058.440 ;
        RECT 4.400 1057.040 1195.600 1057.080 ;
        RECT 4.400 1055.680 1196.000 1057.040 ;
        RECT 3.990 1047.560 1196.000 1055.680 ;
        RECT 3.990 1046.200 1195.600 1047.560 ;
        RECT 4.400 1046.160 1195.600 1046.200 ;
        RECT 4.400 1044.800 1196.000 1046.160 ;
        RECT 3.990 1037.360 1196.000 1044.800 ;
        RECT 3.990 1036.000 1195.600 1037.360 ;
        RECT 4.400 1035.960 1195.600 1036.000 ;
        RECT 4.400 1034.600 1196.000 1035.960 ;
        RECT 3.990 1026.480 1196.000 1034.600 ;
        RECT 3.990 1025.120 1195.600 1026.480 ;
        RECT 4.400 1025.080 1195.600 1025.120 ;
        RECT 4.400 1023.720 1196.000 1025.080 ;
        RECT 3.990 1016.280 1196.000 1023.720 ;
        RECT 3.990 1014.880 1195.600 1016.280 ;
        RECT 3.990 1014.240 1196.000 1014.880 ;
        RECT 4.400 1012.840 1196.000 1014.240 ;
        RECT 3.990 1005.400 1196.000 1012.840 ;
        RECT 3.990 1004.040 1195.600 1005.400 ;
        RECT 4.400 1004.000 1195.600 1004.040 ;
        RECT 4.400 1002.640 1196.000 1004.000 ;
        RECT 3.990 995.200 1196.000 1002.640 ;
        RECT 3.990 993.800 1195.600 995.200 ;
        RECT 3.990 993.160 1196.000 993.800 ;
        RECT 4.400 991.760 1196.000 993.160 ;
        RECT 3.990 984.320 1196.000 991.760 ;
        RECT 3.990 982.920 1195.600 984.320 ;
        RECT 3.990 982.280 1196.000 982.920 ;
        RECT 4.400 980.880 1196.000 982.280 ;
        RECT 3.990 974.120 1196.000 980.880 ;
        RECT 3.990 972.720 1195.600 974.120 ;
        RECT 3.990 972.080 1196.000 972.720 ;
        RECT 4.400 970.680 1196.000 972.080 ;
        RECT 3.990 963.240 1196.000 970.680 ;
        RECT 3.990 961.840 1195.600 963.240 ;
        RECT 3.990 961.200 1196.000 961.840 ;
        RECT 4.400 959.800 1196.000 961.200 ;
        RECT 3.990 953.040 1196.000 959.800 ;
        RECT 3.990 951.640 1195.600 953.040 ;
        RECT 3.990 951.000 1196.000 951.640 ;
        RECT 4.400 949.600 1196.000 951.000 ;
        RECT 3.990 942.160 1196.000 949.600 ;
        RECT 3.990 940.760 1195.600 942.160 ;
        RECT 3.990 940.120 1196.000 940.760 ;
        RECT 4.400 938.720 1196.000 940.120 ;
        RECT 3.990 931.960 1196.000 938.720 ;
        RECT 3.990 930.560 1195.600 931.960 ;
        RECT 3.990 929.240 1196.000 930.560 ;
        RECT 4.400 927.840 1196.000 929.240 ;
        RECT 3.990 921.080 1196.000 927.840 ;
        RECT 3.990 919.680 1195.600 921.080 ;
        RECT 3.990 919.040 1196.000 919.680 ;
        RECT 4.400 917.640 1196.000 919.040 ;
        RECT 3.990 910.880 1196.000 917.640 ;
        RECT 3.990 909.480 1195.600 910.880 ;
        RECT 3.990 908.160 1196.000 909.480 ;
        RECT 4.400 906.760 1196.000 908.160 ;
        RECT 3.990 900.680 1196.000 906.760 ;
        RECT 3.990 899.280 1195.600 900.680 ;
        RECT 3.990 897.960 1196.000 899.280 ;
        RECT 4.400 896.560 1196.000 897.960 ;
        RECT 3.990 889.800 1196.000 896.560 ;
        RECT 3.990 888.400 1195.600 889.800 ;
        RECT 3.990 887.080 1196.000 888.400 ;
        RECT 4.400 885.680 1196.000 887.080 ;
        RECT 3.990 879.600 1196.000 885.680 ;
        RECT 3.990 878.200 1195.600 879.600 ;
        RECT 3.990 876.200 1196.000 878.200 ;
        RECT 4.400 874.800 1196.000 876.200 ;
        RECT 3.990 868.720 1196.000 874.800 ;
        RECT 3.990 867.320 1195.600 868.720 ;
        RECT 3.990 866.000 1196.000 867.320 ;
        RECT 4.400 864.600 1196.000 866.000 ;
        RECT 3.990 858.520 1196.000 864.600 ;
        RECT 3.990 857.120 1195.600 858.520 ;
        RECT 3.990 855.120 1196.000 857.120 ;
        RECT 4.400 853.720 1196.000 855.120 ;
        RECT 3.990 847.640 1196.000 853.720 ;
        RECT 3.990 846.240 1195.600 847.640 ;
        RECT 3.990 844.240 1196.000 846.240 ;
        RECT 4.400 842.840 1196.000 844.240 ;
        RECT 3.990 837.440 1196.000 842.840 ;
        RECT 3.990 836.040 1195.600 837.440 ;
        RECT 3.990 834.040 1196.000 836.040 ;
        RECT 4.400 832.640 1196.000 834.040 ;
        RECT 3.990 826.560 1196.000 832.640 ;
        RECT 3.990 825.160 1195.600 826.560 ;
        RECT 3.990 823.160 1196.000 825.160 ;
        RECT 4.400 821.760 1196.000 823.160 ;
        RECT 3.990 816.360 1196.000 821.760 ;
        RECT 3.990 814.960 1195.600 816.360 ;
        RECT 3.990 812.960 1196.000 814.960 ;
        RECT 4.400 811.560 1196.000 812.960 ;
        RECT 3.990 805.480 1196.000 811.560 ;
        RECT 3.990 804.080 1195.600 805.480 ;
        RECT 3.990 802.080 1196.000 804.080 ;
        RECT 4.400 800.680 1196.000 802.080 ;
        RECT 3.990 795.280 1196.000 800.680 ;
        RECT 3.990 793.880 1195.600 795.280 ;
        RECT 3.990 791.200 1196.000 793.880 ;
        RECT 4.400 789.800 1196.000 791.200 ;
        RECT 3.990 784.400 1196.000 789.800 ;
        RECT 3.990 783.000 1195.600 784.400 ;
        RECT 3.990 781.000 1196.000 783.000 ;
        RECT 4.400 779.600 1196.000 781.000 ;
        RECT 3.990 774.200 1196.000 779.600 ;
        RECT 3.990 772.800 1195.600 774.200 ;
        RECT 3.990 770.120 1196.000 772.800 ;
        RECT 4.400 768.720 1196.000 770.120 ;
        RECT 3.990 763.320 1196.000 768.720 ;
        RECT 3.990 761.920 1195.600 763.320 ;
        RECT 3.990 759.240 1196.000 761.920 ;
        RECT 4.400 757.840 1196.000 759.240 ;
        RECT 3.990 753.120 1196.000 757.840 ;
        RECT 3.990 751.720 1195.600 753.120 ;
        RECT 3.990 749.040 1196.000 751.720 ;
        RECT 4.400 747.640 1196.000 749.040 ;
        RECT 3.990 742.240 1196.000 747.640 ;
        RECT 3.990 740.840 1195.600 742.240 ;
        RECT 3.990 738.160 1196.000 740.840 ;
        RECT 4.400 736.760 1196.000 738.160 ;
        RECT 3.990 732.040 1196.000 736.760 ;
        RECT 3.990 730.640 1195.600 732.040 ;
        RECT 3.990 727.960 1196.000 730.640 ;
        RECT 4.400 726.560 1196.000 727.960 ;
        RECT 3.990 721.160 1196.000 726.560 ;
        RECT 3.990 719.760 1195.600 721.160 ;
        RECT 3.990 717.080 1196.000 719.760 ;
        RECT 4.400 715.680 1196.000 717.080 ;
        RECT 3.990 710.960 1196.000 715.680 ;
        RECT 3.990 709.560 1195.600 710.960 ;
        RECT 3.990 706.200 1196.000 709.560 ;
        RECT 4.400 704.800 1196.000 706.200 ;
        RECT 3.990 700.080 1196.000 704.800 ;
        RECT 3.990 698.680 1195.600 700.080 ;
        RECT 3.990 696.000 1196.000 698.680 ;
        RECT 4.400 694.600 1196.000 696.000 ;
        RECT 3.990 689.880 1196.000 694.600 ;
        RECT 3.990 688.480 1195.600 689.880 ;
        RECT 3.990 685.120 1196.000 688.480 ;
        RECT 4.400 683.720 1196.000 685.120 ;
        RECT 3.990 679.000 1196.000 683.720 ;
        RECT 3.990 677.600 1195.600 679.000 ;
        RECT 3.990 674.920 1196.000 677.600 ;
        RECT 4.400 673.520 1196.000 674.920 ;
        RECT 3.990 668.800 1196.000 673.520 ;
        RECT 3.990 667.400 1195.600 668.800 ;
        RECT 3.990 664.040 1196.000 667.400 ;
        RECT 4.400 662.640 1196.000 664.040 ;
        RECT 3.990 657.920 1196.000 662.640 ;
        RECT 3.990 656.520 1195.600 657.920 ;
        RECT 3.990 653.160 1196.000 656.520 ;
        RECT 4.400 651.760 1196.000 653.160 ;
        RECT 3.990 647.720 1196.000 651.760 ;
        RECT 3.990 646.320 1195.600 647.720 ;
        RECT 3.990 642.960 1196.000 646.320 ;
        RECT 4.400 641.560 1196.000 642.960 ;
        RECT 3.990 636.840 1196.000 641.560 ;
        RECT 3.990 635.440 1195.600 636.840 ;
        RECT 3.990 632.080 1196.000 635.440 ;
        RECT 4.400 630.680 1196.000 632.080 ;
        RECT 3.990 626.640 1196.000 630.680 ;
        RECT 3.990 625.240 1195.600 626.640 ;
        RECT 3.990 621.200 1196.000 625.240 ;
        RECT 4.400 619.800 1196.000 621.200 ;
        RECT 3.990 615.760 1196.000 619.800 ;
        RECT 3.990 614.360 1195.600 615.760 ;
        RECT 3.990 611.000 1196.000 614.360 ;
        RECT 4.400 609.600 1196.000 611.000 ;
        RECT 3.990 605.560 1196.000 609.600 ;
        RECT 3.990 604.160 1195.600 605.560 ;
        RECT 3.990 600.120 1196.000 604.160 ;
        RECT 4.400 598.720 1196.000 600.120 ;
        RECT 3.990 595.360 1196.000 598.720 ;
        RECT 3.990 593.960 1195.600 595.360 ;
        RECT 3.990 589.920 1196.000 593.960 ;
        RECT 4.400 588.520 1196.000 589.920 ;
        RECT 3.990 584.480 1196.000 588.520 ;
        RECT 3.990 583.080 1195.600 584.480 ;
        RECT 3.990 579.040 1196.000 583.080 ;
        RECT 4.400 577.640 1196.000 579.040 ;
        RECT 3.990 574.280 1196.000 577.640 ;
        RECT 3.990 572.880 1195.600 574.280 ;
        RECT 3.990 568.160 1196.000 572.880 ;
        RECT 4.400 566.760 1196.000 568.160 ;
        RECT 3.990 563.400 1196.000 566.760 ;
        RECT 3.990 562.000 1195.600 563.400 ;
        RECT 3.990 557.960 1196.000 562.000 ;
        RECT 4.400 556.560 1196.000 557.960 ;
        RECT 3.990 553.200 1196.000 556.560 ;
        RECT 3.990 551.800 1195.600 553.200 ;
        RECT 3.990 547.080 1196.000 551.800 ;
        RECT 4.400 545.680 1196.000 547.080 ;
        RECT 3.990 542.320 1196.000 545.680 ;
        RECT 3.990 540.920 1195.600 542.320 ;
        RECT 3.990 536.200 1196.000 540.920 ;
        RECT 4.400 534.800 1196.000 536.200 ;
        RECT 3.990 532.120 1196.000 534.800 ;
        RECT 3.990 530.720 1195.600 532.120 ;
        RECT 3.990 526.000 1196.000 530.720 ;
        RECT 4.400 524.600 1196.000 526.000 ;
        RECT 3.990 521.240 1196.000 524.600 ;
        RECT 3.990 519.840 1195.600 521.240 ;
        RECT 3.990 515.120 1196.000 519.840 ;
        RECT 4.400 513.720 1196.000 515.120 ;
        RECT 3.990 511.040 1196.000 513.720 ;
        RECT 3.990 509.640 1195.600 511.040 ;
        RECT 3.990 504.920 1196.000 509.640 ;
        RECT 4.400 503.520 1196.000 504.920 ;
        RECT 3.990 500.160 1196.000 503.520 ;
        RECT 3.990 498.760 1195.600 500.160 ;
        RECT 3.990 494.040 1196.000 498.760 ;
        RECT 4.400 492.640 1196.000 494.040 ;
        RECT 3.990 489.960 1196.000 492.640 ;
        RECT 3.990 488.560 1195.600 489.960 ;
        RECT 3.990 483.160 1196.000 488.560 ;
        RECT 4.400 481.760 1196.000 483.160 ;
        RECT 3.990 479.080 1196.000 481.760 ;
        RECT 3.990 477.680 1195.600 479.080 ;
        RECT 3.990 472.960 1196.000 477.680 ;
        RECT 4.400 471.560 1196.000 472.960 ;
        RECT 3.990 468.880 1196.000 471.560 ;
        RECT 3.990 467.480 1195.600 468.880 ;
        RECT 3.990 462.080 1196.000 467.480 ;
        RECT 4.400 460.680 1196.000 462.080 ;
        RECT 3.990 458.000 1196.000 460.680 ;
        RECT 3.990 456.600 1195.600 458.000 ;
        RECT 3.990 451.880 1196.000 456.600 ;
        RECT 4.400 450.480 1196.000 451.880 ;
        RECT 3.990 447.800 1196.000 450.480 ;
        RECT 3.990 446.400 1195.600 447.800 ;
        RECT 3.990 441.000 1196.000 446.400 ;
        RECT 4.400 439.600 1196.000 441.000 ;
        RECT 3.990 436.920 1196.000 439.600 ;
        RECT 3.990 435.520 1195.600 436.920 ;
        RECT 3.990 430.120 1196.000 435.520 ;
        RECT 4.400 428.720 1196.000 430.120 ;
        RECT 3.990 426.720 1196.000 428.720 ;
        RECT 3.990 425.320 1195.600 426.720 ;
        RECT 3.990 419.920 1196.000 425.320 ;
        RECT 4.400 418.520 1196.000 419.920 ;
        RECT 3.990 415.840 1196.000 418.520 ;
        RECT 3.990 414.440 1195.600 415.840 ;
        RECT 3.990 409.040 1196.000 414.440 ;
        RECT 4.400 407.640 1196.000 409.040 ;
        RECT 3.990 405.640 1196.000 407.640 ;
        RECT 3.990 404.240 1195.600 405.640 ;
        RECT 3.990 398.160 1196.000 404.240 ;
        RECT 4.400 396.760 1196.000 398.160 ;
        RECT 3.990 394.760 1196.000 396.760 ;
        RECT 3.990 393.360 1195.600 394.760 ;
        RECT 3.990 387.960 1196.000 393.360 ;
        RECT 4.400 386.560 1196.000 387.960 ;
        RECT 3.990 384.560 1196.000 386.560 ;
        RECT 3.990 383.160 1195.600 384.560 ;
        RECT 3.990 377.080 1196.000 383.160 ;
        RECT 4.400 375.680 1196.000 377.080 ;
        RECT 3.990 373.680 1196.000 375.680 ;
        RECT 3.990 372.280 1195.600 373.680 ;
        RECT 3.990 366.880 1196.000 372.280 ;
        RECT 4.400 365.480 1196.000 366.880 ;
        RECT 3.990 363.480 1196.000 365.480 ;
        RECT 3.990 362.080 1195.600 363.480 ;
        RECT 3.990 356.000 1196.000 362.080 ;
        RECT 4.400 354.600 1196.000 356.000 ;
        RECT 3.990 352.600 1196.000 354.600 ;
        RECT 3.990 351.200 1195.600 352.600 ;
        RECT 3.990 345.120 1196.000 351.200 ;
        RECT 4.400 343.720 1196.000 345.120 ;
        RECT 3.990 342.400 1196.000 343.720 ;
        RECT 3.990 341.000 1195.600 342.400 ;
        RECT 3.990 334.920 1196.000 341.000 ;
        RECT 4.400 333.520 1196.000 334.920 ;
        RECT 3.990 331.520 1196.000 333.520 ;
        RECT 3.990 330.120 1195.600 331.520 ;
        RECT 3.990 324.040 1196.000 330.120 ;
        RECT 4.400 322.640 1196.000 324.040 ;
        RECT 3.990 321.320 1196.000 322.640 ;
        RECT 3.990 319.920 1195.600 321.320 ;
        RECT 3.990 313.160 1196.000 319.920 ;
        RECT 4.400 311.760 1196.000 313.160 ;
        RECT 3.990 310.440 1196.000 311.760 ;
        RECT 3.990 309.040 1195.600 310.440 ;
        RECT 3.990 302.960 1196.000 309.040 ;
        RECT 4.400 301.560 1196.000 302.960 ;
        RECT 3.990 300.240 1196.000 301.560 ;
        RECT 3.990 298.840 1195.600 300.240 ;
        RECT 3.990 292.080 1196.000 298.840 ;
        RECT 4.400 290.680 1196.000 292.080 ;
        RECT 3.990 290.040 1196.000 290.680 ;
        RECT 3.990 288.640 1195.600 290.040 ;
        RECT 3.990 281.880 1196.000 288.640 ;
        RECT 4.400 280.480 1196.000 281.880 ;
        RECT 3.990 279.160 1196.000 280.480 ;
        RECT 3.990 277.760 1195.600 279.160 ;
        RECT 3.990 271.000 1196.000 277.760 ;
        RECT 4.400 269.600 1196.000 271.000 ;
        RECT 3.990 268.960 1196.000 269.600 ;
        RECT 3.990 267.560 1195.600 268.960 ;
        RECT 3.990 260.120 1196.000 267.560 ;
        RECT 4.400 258.720 1196.000 260.120 ;
        RECT 3.990 258.080 1196.000 258.720 ;
        RECT 3.990 256.680 1195.600 258.080 ;
        RECT 3.990 249.920 1196.000 256.680 ;
        RECT 4.400 248.520 1196.000 249.920 ;
        RECT 3.990 247.880 1196.000 248.520 ;
        RECT 3.990 246.480 1195.600 247.880 ;
        RECT 3.990 239.040 1196.000 246.480 ;
        RECT 4.400 237.640 1196.000 239.040 ;
        RECT 3.990 237.000 1196.000 237.640 ;
        RECT 3.990 235.600 1195.600 237.000 ;
        RECT 3.990 228.840 1196.000 235.600 ;
        RECT 4.400 227.440 1196.000 228.840 ;
        RECT 3.990 226.800 1196.000 227.440 ;
        RECT 3.990 225.400 1195.600 226.800 ;
        RECT 3.990 217.960 1196.000 225.400 ;
        RECT 4.400 216.560 1196.000 217.960 ;
        RECT 3.990 215.920 1196.000 216.560 ;
        RECT 3.990 214.520 1195.600 215.920 ;
        RECT 3.990 207.080 1196.000 214.520 ;
        RECT 4.400 205.720 1196.000 207.080 ;
        RECT 4.400 205.680 1195.600 205.720 ;
        RECT 3.990 204.320 1195.600 205.680 ;
        RECT 3.990 196.880 1196.000 204.320 ;
        RECT 4.400 195.480 1196.000 196.880 ;
        RECT 3.990 194.840 1196.000 195.480 ;
        RECT 3.990 193.440 1195.600 194.840 ;
        RECT 3.990 186.000 1196.000 193.440 ;
        RECT 4.400 184.640 1196.000 186.000 ;
        RECT 4.400 184.600 1195.600 184.640 ;
        RECT 3.990 183.240 1195.600 184.600 ;
        RECT 3.990 175.120 1196.000 183.240 ;
        RECT 4.400 173.760 1196.000 175.120 ;
        RECT 4.400 173.720 1195.600 173.760 ;
        RECT 3.990 172.360 1195.600 173.720 ;
        RECT 3.990 164.920 1196.000 172.360 ;
        RECT 4.400 163.560 1196.000 164.920 ;
        RECT 4.400 163.520 1195.600 163.560 ;
        RECT 3.990 162.160 1195.600 163.520 ;
        RECT 3.990 154.040 1196.000 162.160 ;
        RECT 4.400 152.680 1196.000 154.040 ;
        RECT 4.400 152.640 1195.600 152.680 ;
        RECT 3.990 151.280 1195.600 152.640 ;
        RECT 3.990 143.840 1196.000 151.280 ;
        RECT 4.400 142.480 1196.000 143.840 ;
        RECT 4.400 142.440 1195.600 142.480 ;
        RECT 3.990 141.080 1195.600 142.440 ;
        RECT 3.990 132.960 1196.000 141.080 ;
        RECT 4.400 131.600 1196.000 132.960 ;
        RECT 4.400 131.560 1195.600 131.600 ;
        RECT 3.990 130.200 1195.600 131.560 ;
        RECT 3.990 122.080 1196.000 130.200 ;
        RECT 4.400 121.400 1196.000 122.080 ;
        RECT 4.400 120.680 1195.600 121.400 ;
        RECT 3.990 120.000 1195.600 120.680 ;
        RECT 3.990 111.880 1196.000 120.000 ;
        RECT 4.400 110.520 1196.000 111.880 ;
        RECT 4.400 110.480 1195.600 110.520 ;
        RECT 3.990 109.120 1195.600 110.480 ;
        RECT 3.990 101.000 1196.000 109.120 ;
        RECT 4.400 100.320 1196.000 101.000 ;
        RECT 4.400 99.600 1195.600 100.320 ;
        RECT 3.990 98.920 1195.600 99.600 ;
        RECT 3.990 90.120 1196.000 98.920 ;
        RECT 4.400 89.440 1196.000 90.120 ;
        RECT 4.400 88.720 1195.600 89.440 ;
        RECT 3.990 88.040 1195.600 88.720 ;
        RECT 3.990 79.920 1196.000 88.040 ;
        RECT 4.400 79.240 1196.000 79.920 ;
        RECT 4.400 78.520 1195.600 79.240 ;
        RECT 3.990 77.840 1195.600 78.520 ;
        RECT 3.990 69.040 1196.000 77.840 ;
        RECT 4.400 68.360 1196.000 69.040 ;
        RECT 4.400 67.640 1195.600 68.360 ;
        RECT 3.990 66.960 1195.600 67.640 ;
        RECT 3.990 58.840 1196.000 66.960 ;
        RECT 4.400 58.160 1196.000 58.840 ;
        RECT 4.400 57.440 1195.600 58.160 ;
        RECT 3.990 56.760 1195.600 57.440 ;
        RECT 3.990 47.960 1196.000 56.760 ;
        RECT 4.400 47.280 1196.000 47.960 ;
        RECT 4.400 46.560 1195.600 47.280 ;
        RECT 3.990 45.880 1195.600 46.560 ;
        RECT 3.990 37.080 1196.000 45.880 ;
        RECT 4.400 35.680 1195.600 37.080 ;
        RECT 3.990 26.880 1196.000 35.680 ;
        RECT 4.400 26.200 1196.000 26.880 ;
        RECT 4.400 25.480 1195.600 26.200 ;
        RECT 3.990 24.800 1195.600 25.480 ;
        RECT 3.990 16.000 1196.000 24.800 ;
        RECT 4.400 14.600 1195.600 16.000 ;
        RECT 3.990 5.800 1196.000 14.600 ;
        RECT 4.400 4.935 1195.600 5.800 ;
      LAYER met4 ;
        RECT 15.935 1189.280 1188.345 1195.945 ;
        RECT 15.935 10.640 20.640 1189.280 ;
        RECT 23.040 10.640 97.440 1189.280 ;
        RECT 99.840 10.640 1188.345 1189.280 ;
  END
END hs32_core1
END LIBRARY

