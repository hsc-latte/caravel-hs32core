VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2433.460 2924.800 2434.660 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2903.340 2924.800 2904.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3410.620 2.400 3411.820 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 2.400 3124.860 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2836.020 2.400 2837.220 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 2.400 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 2.400 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1974.460 2.400 1975.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 2.400 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 2.400 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 2.400 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 2.400 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 2.400 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 2.400 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 2.400 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 2.400 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1964.260 2924.800 1965.460 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2198.860 2924.800 2200.060 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 2.400 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 2.400 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 2.400 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 2.400 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 2.400 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 2.400 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 2.400 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 2.400 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 2.400 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 2.400 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 2.400 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 2.400 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.220 2.400 3340.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 2.400 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 2.400 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2476.980 2.400 2478.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 2.400 2190.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 2.400 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 2.400 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 2.400 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 2.400 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 2.400 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 2.400 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 2.400 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 2.400 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 538.730 1590.420 539.050 1590.480 ;
        RECT 544.250 1590.420 544.570 1590.480 ;
        RECT 538.730 1590.280 544.570 1590.420 ;
        RECT 538.730 1590.220 539.050 1590.280 ;
        RECT 544.250 1590.220 544.570 1590.280 ;
        RECT 544.250 14.180 544.570 14.240 ;
        RECT 633.030 14.180 633.350 14.240 ;
        RECT 544.250 14.040 633.350 14.180 ;
        RECT 544.250 13.980 544.570 14.040 ;
        RECT 633.030 13.980 633.350 14.040 ;
      LAYER via ;
        RECT 538.760 1590.220 539.020 1590.480 ;
        RECT 544.280 1590.220 544.540 1590.480 ;
        RECT 544.280 13.980 544.540 14.240 ;
        RECT 633.060 13.980 633.320 14.240 ;
      LAYER met2 ;
        RECT 538.760 1600.000 539.040 1604.000 ;
        RECT 538.820 1590.510 538.960 1600.000 ;
        RECT 538.760 1590.190 539.020 1590.510 ;
        RECT 544.280 1590.190 544.540 1590.510 ;
        RECT 544.340 14.270 544.480 1590.190 ;
        RECT 544.280 13.950 544.540 14.270 ;
        RECT 633.060 13.950 633.320 14.270 ;
        RECT 633.120 2.400 633.260 13.950 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1212.630 79.120 1212.950 79.180 ;
        RECT 2415.070 79.120 2415.390 79.180 ;
        RECT 1212.630 78.980 2415.390 79.120 ;
        RECT 1212.630 78.920 1212.950 78.980 ;
        RECT 2415.070 78.920 2415.390 78.980 ;
      LAYER via ;
        RECT 1212.660 78.920 1212.920 79.180 ;
        RECT 2415.100 78.920 2415.360 79.180 ;
      LAYER met2 ;
        RECT 1212.200 1600.450 1212.480 1604.000 ;
        RECT 1212.200 1600.310 1212.860 1600.450 ;
        RECT 1212.200 1600.000 1212.480 1600.310 ;
        RECT 1212.720 79.210 1212.860 1600.310 ;
        RECT 1212.660 78.890 1212.920 79.210 ;
        RECT 2415.100 78.890 2415.360 79.210 ;
        RECT 2415.160 17.410 2415.300 78.890 ;
        RECT 2415.160 17.270 2417.600 17.410 ;
        RECT 2417.460 2.400 2417.600 17.270 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1219.990 82.860 1220.310 82.920 ;
        RECT 2428.870 82.860 2429.190 82.920 ;
        RECT 1219.990 82.720 2429.190 82.860 ;
        RECT 1219.990 82.660 1220.310 82.720 ;
        RECT 2428.870 82.660 2429.190 82.720 ;
        RECT 2428.870 17.920 2429.190 17.980 ;
        RECT 2434.850 17.920 2435.170 17.980 ;
        RECT 2428.870 17.780 2435.170 17.920 ;
        RECT 2428.870 17.720 2429.190 17.780 ;
        RECT 2434.850 17.720 2435.170 17.780 ;
      LAYER via ;
        RECT 1220.020 82.660 1220.280 82.920 ;
        RECT 2428.900 82.660 2429.160 82.920 ;
        RECT 2428.900 17.720 2429.160 17.980 ;
        RECT 2434.880 17.720 2435.140 17.980 ;
      LAYER met2 ;
        RECT 1218.640 1600.450 1218.920 1604.000 ;
        RECT 1218.640 1600.310 1220.220 1600.450 ;
        RECT 1218.640 1600.000 1218.920 1600.310 ;
        RECT 1220.080 82.950 1220.220 1600.310 ;
        RECT 1220.020 82.630 1220.280 82.950 ;
        RECT 2428.900 82.630 2429.160 82.950 ;
        RECT 2428.960 18.010 2429.100 82.630 ;
        RECT 2428.900 17.690 2429.160 18.010 ;
        RECT 2434.880 17.690 2435.140 18.010 ;
        RECT 2434.940 2.400 2435.080 17.690 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1226.890 82.520 1227.210 82.580 ;
        RECT 2449.570 82.520 2449.890 82.580 ;
        RECT 1226.890 82.380 2449.890 82.520 ;
        RECT 1226.890 82.320 1227.210 82.380 ;
        RECT 2449.570 82.320 2449.890 82.380 ;
        RECT 2449.570 2.960 2449.890 3.020 ;
        RECT 2452.790 2.960 2453.110 3.020 ;
        RECT 2449.570 2.820 2453.110 2.960 ;
        RECT 2449.570 2.760 2449.890 2.820 ;
        RECT 2452.790 2.760 2453.110 2.820 ;
      LAYER via ;
        RECT 1226.920 82.320 1227.180 82.580 ;
        RECT 2449.600 82.320 2449.860 82.580 ;
        RECT 2449.600 2.760 2449.860 3.020 ;
        RECT 2452.820 2.760 2453.080 3.020 ;
      LAYER met2 ;
        RECT 1225.540 1600.450 1225.820 1604.000 ;
        RECT 1225.540 1600.310 1227.120 1600.450 ;
        RECT 1225.540 1600.000 1225.820 1600.310 ;
        RECT 1226.980 82.610 1227.120 1600.310 ;
        RECT 1226.920 82.290 1227.180 82.610 ;
        RECT 2449.600 82.290 2449.860 82.610 ;
        RECT 2449.660 3.050 2449.800 82.290 ;
        RECT 2449.600 2.730 2449.860 3.050 ;
        RECT 2452.820 2.730 2453.080 3.050 ;
        RECT 2452.880 2.400 2453.020 2.730 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1233.790 81.840 1234.110 81.900 ;
        RECT 2470.730 81.840 2471.050 81.900 ;
        RECT 1233.790 81.700 2471.050 81.840 ;
        RECT 1233.790 81.640 1234.110 81.700 ;
        RECT 2470.730 81.640 2471.050 81.700 ;
      LAYER via ;
        RECT 1233.820 81.640 1234.080 81.900 ;
        RECT 2470.760 81.640 2471.020 81.900 ;
      LAYER met2 ;
        RECT 1232.440 1600.450 1232.720 1604.000 ;
        RECT 1232.440 1600.310 1234.020 1600.450 ;
        RECT 1232.440 1600.000 1232.720 1600.310 ;
        RECT 1233.880 81.930 1234.020 1600.310 ;
        RECT 1233.820 81.610 1234.080 81.930 ;
        RECT 2470.760 81.610 2471.020 81.930 ;
        RECT 2470.820 2.400 2470.960 81.610 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1240.690 81.500 1241.010 81.560 ;
        RECT 2484.070 81.500 2484.390 81.560 ;
        RECT 1240.690 81.360 2484.390 81.500 ;
        RECT 1240.690 81.300 1241.010 81.360 ;
        RECT 2484.070 81.300 2484.390 81.360 ;
        RECT 2484.070 2.960 2484.390 3.020 ;
        RECT 2488.670 2.960 2488.990 3.020 ;
        RECT 2484.070 2.820 2488.990 2.960 ;
        RECT 2484.070 2.760 2484.390 2.820 ;
        RECT 2488.670 2.760 2488.990 2.820 ;
      LAYER via ;
        RECT 1240.720 81.300 1240.980 81.560 ;
        RECT 2484.100 81.300 2484.360 81.560 ;
        RECT 2484.100 2.760 2484.360 3.020 ;
        RECT 2488.700 2.760 2488.960 3.020 ;
      LAYER met2 ;
        RECT 1238.880 1600.450 1239.160 1604.000 ;
        RECT 1238.880 1600.310 1240.920 1600.450 ;
        RECT 1238.880 1600.000 1239.160 1600.310 ;
        RECT 1240.780 81.590 1240.920 1600.310 ;
        RECT 1240.720 81.270 1240.980 81.590 ;
        RECT 2484.100 81.270 2484.360 81.590 ;
        RECT 2484.160 3.050 2484.300 81.270 ;
        RECT 2484.100 2.730 2484.360 3.050 ;
        RECT 2488.700 2.730 2488.960 3.050 ;
        RECT 2488.760 2.400 2488.900 2.730 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1247.590 81.160 1247.910 81.220 ;
        RECT 2504.770 81.160 2505.090 81.220 ;
        RECT 1247.590 81.020 2505.090 81.160 ;
        RECT 1247.590 80.960 1247.910 81.020 ;
        RECT 2504.770 80.960 2505.090 81.020 ;
        RECT 2504.770 2.960 2505.090 3.020 ;
        RECT 2506.150 2.960 2506.470 3.020 ;
        RECT 2504.770 2.820 2506.470 2.960 ;
        RECT 2504.770 2.760 2505.090 2.820 ;
        RECT 2506.150 2.760 2506.470 2.820 ;
      LAYER via ;
        RECT 1247.620 80.960 1247.880 81.220 ;
        RECT 2504.800 80.960 2505.060 81.220 ;
        RECT 2504.800 2.760 2505.060 3.020 ;
        RECT 2506.180 2.760 2506.440 3.020 ;
      LAYER met2 ;
        RECT 1245.780 1600.450 1246.060 1604.000 ;
        RECT 1245.780 1600.310 1247.820 1600.450 ;
        RECT 1245.780 1600.000 1246.060 1600.310 ;
        RECT 1247.680 81.250 1247.820 1600.310 ;
        RECT 1247.620 80.930 1247.880 81.250 ;
        RECT 2504.800 80.930 2505.060 81.250 ;
        RECT 2504.860 3.050 2505.000 80.930 ;
        RECT 2504.800 2.730 2505.060 3.050 ;
        RECT 2506.180 2.730 2506.440 3.050 ;
        RECT 2506.240 2.400 2506.380 2.730 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1254.490 80.820 1254.810 80.880 ;
        RECT 2518.570 80.820 2518.890 80.880 ;
        RECT 1254.490 80.680 2518.890 80.820 ;
        RECT 1254.490 80.620 1254.810 80.680 ;
        RECT 2518.570 80.620 2518.890 80.680 ;
        RECT 2518.570 2.960 2518.890 3.020 ;
        RECT 2524.090 2.960 2524.410 3.020 ;
        RECT 2518.570 2.820 2524.410 2.960 ;
        RECT 2518.570 2.760 2518.890 2.820 ;
        RECT 2524.090 2.760 2524.410 2.820 ;
      LAYER via ;
        RECT 1254.520 80.620 1254.780 80.880 ;
        RECT 2518.600 80.620 2518.860 80.880 ;
        RECT 2518.600 2.760 2518.860 3.020 ;
        RECT 2524.120 2.760 2524.380 3.020 ;
      LAYER met2 ;
        RECT 1252.220 1601.130 1252.500 1604.000 ;
        RECT 1252.220 1600.990 1254.260 1601.130 ;
        RECT 1252.220 1600.000 1252.500 1600.990 ;
        RECT 1254.120 1590.250 1254.260 1600.990 ;
        RECT 1254.120 1590.110 1254.720 1590.250 ;
        RECT 1254.580 80.910 1254.720 1590.110 ;
        RECT 1254.520 80.590 1254.780 80.910 ;
        RECT 2518.600 80.590 2518.860 80.910 ;
        RECT 2518.660 3.050 2518.800 80.590 ;
        RECT 2518.600 2.730 2518.860 3.050 ;
        RECT 2524.120 2.730 2524.380 3.050 ;
        RECT 2524.180 2.400 2524.320 2.730 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1261.390 80.480 1261.710 80.540 ;
        RECT 2539.270 80.480 2539.590 80.540 ;
        RECT 1261.390 80.340 2539.590 80.480 ;
        RECT 1261.390 80.280 1261.710 80.340 ;
        RECT 2539.270 80.280 2539.590 80.340 ;
        RECT 2539.270 2.960 2539.590 3.020 ;
        RECT 2542.030 2.960 2542.350 3.020 ;
        RECT 2539.270 2.820 2542.350 2.960 ;
        RECT 2539.270 2.760 2539.590 2.820 ;
        RECT 2542.030 2.760 2542.350 2.820 ;
      LAYER via ;
        RECT 1261.420 80.280 1261.680 80.540 ;
        RECT 2539.300 80.280 2539.560 80.540 ;
        RECT 2539.300 2.760 2539.560 3.020 ;
        RECT 2542.060 2.760 2542.320 3.020 ;
      LAYER met2 ;
        RECT 1259.120 1600.450 1259.400 1604.000 ;
        RECT 1259.120 1600.310 1260.700 1600.450 ;
        RECT 1259.120 1600.000 1259.400 1600.310 ;
        RECT 1260.560 1590.250 1260.700 1600.310 ;
        RECT 1260.560 1590.110 1261.620 1590.250 ;
        RECT 1261.480 80.570 1261.620 1590.110 ;
        RECT 1261.420 80.250 1261.680 80.570 ;
        RECT 2539.300 80.250 2539.560 80.570 ;
        RECT 2539.360 3.050 2539.500 80.250 ;
        RECT 2539.300 2.730 2539.560 3.050 ;
        RECT 2542.060 2.730 2542.320 3.050 ;
        RECT 2542.120 2.400 2542.260 2.730 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1265.990 1589.400 1266.310 1589.460 ;
        RECT 1269.210 1589.400 1269.530 1589.460 ;
        RECT 1265.990 1589.260 1269.530 1589.400 ;
        RECT 1265.990 1589.200 1266.310 1589.260 ;
        RECT 1269.210 1589.200 1269.530 1589.260 ;
        RECT 1269.210 22.000 1269.530 22.060 ;
        RECT 2559.970 22.000 2560.290 22.060 ;
        RECT 1269.210 21.860 2560.290 22.000 ;
        RECT 1269.210 21.800 1269.530 21.860 ;
        RECT 2559.970 21.800 2560.290 21.860 ;
      LAYER via ;
        RECT 1266.020 1589.200 1266.280 1589.460 ;
        RECT 1269.240 1589.200 1269.500 1589.460 ;
        RECT 1269.240 21.800 1269.500 22.060 ;
        RECT 2560.000 21.800 2560.260 22.060 ;
      LAYER met2 ;
        RECT 1266.020 1600.000 1266.300 1604.000 ;
        RECT 1266.080 1589.490 1266.220 1600.000 ;
        RECT 1266.020 1589.170 1266.280 1589.490 ;
        RECT 1269.240 1589.170 1269.500 1589.490 ;
        RECT 1269.300 22.090 1269.440 1589.170 ;
        RECT 1269.240 21.770 1269.500 22.090 ;
        RECT 2560.000 21.770 2560.260 22.090 ;
        RECT 2560.060 2.400 2560.200 21.770 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1272.430 1589.400 1272.750 1589.460 ;
        RECT 1276.110 1589.400 1276.430 1589.460 ;
        RECT 1272.430 1589.260 1276.430 1589.400 ;
        RECT 1272.430 1589.200 1272.750 1589.260 ;
        RECT 1276.110 1589.200 1276.430 1589.260 ;
        RECT 1276.110 22.340 1276.430 22.400 ;
        RECT 2577.910 22.340 2578.230 22.400 ;
        RECT 1276.110 22.200 2578.230 22.340 ;
        RECT 1276.110 22.140 1276.430 22.200 ;
        RECT 2577.910 22.140 2578.230 22.200 ;
      LAYER via ;
        RECT 1272.460 1589.200 1272.720 1589.460 ;
        RECT 1276.140 1589.200 1276.400 1589.460 ;
        RECT 1276.140 22.140 1276.400 22.400 ;
        RECT 2577.940 22.140 2578.200 22.400 ;
      LAYER met2 ;
        RECT 1272.460 1600.000 1272.740 1604.000 ;
        RECT 1272.520 1589.490 1272.660 1600.000 ;
        RECT 1272.460 1589.170 1272.720 1589.490 ;
        RECT 1276.140 1589.170 1276.400 1589.490 ;
        RECT 1276.200 22.430 1276.340 1589.170 ;
        RECT 1276.140 22.110 1276.400 22.430 ;
        RECT 2577.940 22.110 2578.200 22.430 ;
        RECT 2578.000 2.400 2578.140 22.110 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 605.920 1600.450 606.200 1604.000 ;
        RECT 605.920 1600.310 607.040 1600.450 ;
        RECT 605.920 1600.000 606.200 1600.310 ;
        RECT 606.900 18.205 607.040 1600.310 ;
        RECT 606.830 17.835 607.110 18.205 ;
        RECT 811.530 17.835 811.810 18.205 ;
        RECT 811.600 2.400 811.740 17.835 ;
        RECT 811.390 -4.800 811.950 2.400 ;
      LAYER via2 ;
        RECT 606.830 17.880 607.110 18.160 ;
        RECT 811.530 17.880 811.810 18.160 ;
      LAYER met3 ;
        RECT 606.805 18.170 607.135 18.185 ;
        RECT 811.505 18.170 811.835 18.185 ;
        RECT 606.805 17.870 811.835 18.170 ;
        RECT 606.805 17.855 607.135 17.870 ;
        RECT 811.505 17.855 811.835 17.870 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1279.330 1589.400 1279.650 1589.460 ;
        RECT 1283.010 1589.400 1283.330 1589.460 ;
        RECT 1279.330 1589.260 1283.330 1589.400 ;
        RECT 1279.330 1589.200 1279.650 1589.260 ;
        RECT 1283.010 1589.200 1283.330 1589.260 ;
        RECT 1283.010 22.680 1283.330 22.740 ;
        RECT 2595.390 22.680 2595.710 22.740 ;
        RECT 1283.010 22.540 2595.710 22.680 ;
        RECT 1283.010 22.480 1283.330 22.540 ;
        RECT 2595.390 22.480 2595.710 22.540 ;
      LAYER via ;
        RECT 1279.360 1589.200 1279.620 1589.460 ;
        RECT 1283.040 1589.200 1283.300 1589.460 ;
        RECT 1283.040 22.480 1283.300 22.740 ;
        RECT 2595.420 22.480 2595.680 22.740 ;
      LAYER met2 ;
        RECT 1279.360 1600.000 1279.640 1604.000 ;
        RECT 1279.420 1589.490 1279.560 1600.000 ;
        RECT 1279.360 1589.170 1279.620 1589.490 ;
        RECT 1283.040 1589.170 1283.300 1589.490 ;
        RECT 1283.100 22.770 1283.240 1589.170 ;
        RECT 1283.040 22.450 1283.300 22.770 ;
        RECT 2595.420 22.450 2595.680 22.770 ;
        RECT 2595.480 2.400 2595.620 22.450 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1286.230 1589.400 1286.550 1589.460 ;
        RECT 1289.910 1589.400 1290.230 1589.460 ;
        RECT 1286.230 1589.260 1290.230 1589.400 ;
        RECT 1286.230 1589.200 1286.550 1589.260 ;
        RECT 1289.910 1589.200 1290.230 1589.260 ;
        RECT 1289.910 23.020 1290.230 23.080 ;
        RECT 2613.330 23.020 2613.650 23.080 ;
        RECT 1289.910 22.880 2613.650 23.020 ;
        RECT 1289.910 22.820 1290.230 22.880 ;
        RECT 2613.330 22.820 2613.650 22.880 ;
      LAYER via ;
        RECT 1286.260 1589.200 1286.520 1589.460 ;
        RECT 1289.940 1589.200 1290.200 1589.460 ;
        RECT 1289.940 22.820 1290.200 23.080 ;
        RECT 2613.360 22.820 2613.620 23.080 ;
      LAYER met2 ;
        RECT 1286.260 1600.000 1286.540 1604.000 ;
        RECT 1286.320 1589.490 1286.460 1600.000 ;
        RECT 1286.260 1589.170 1286.520 1589.490 ;
        RECT 1289.940 1589.170 1290.200 1589.490 ;
        RECT 1290.000 23.110 1290.140 1589.170 ;
        RECT 1289.940 22.790 1290.200 23.110 ;
        RECT 2613.360 22.790 2613.620 23.110 ;
        RECT 2613.420 2.400 2613.560 22.790 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1292.670 1589.400 1292.990 1589.460 ;
        RECT 1296.810 1589.400 1297.130 1589.460 ;
        RECT 1292.670 1589.260 1297.130 1589.400 ;
        RECT 1292.670 1589.200 1292.990 1589.260 ;
        RECT 1296.810 1589.200 1297.130 1589.260 ;
        RECT 1296.810 23.360 1297.130 23.420 ;
        RECT 2631.270 23.360 2631.590 23.420 ;
        RECT 1296.810 23.220 2631.590 23.360 ;
        RECT 1296.810 23.160 1297.130 23.220 ;
        RECT 2631.270 23.160 2631.590 23.220 ;
      LAYER via ;
        RECT 1292.700 1589.200 1292.960 1589.460 ;
        RECT 1296.840 1589.200 1297.100 1589.460 ;
        RECT 1296.840 23.160 1297.100 23.420 ;
        RECT 2631.300 23.160 2631.560 23.420 ;
      LAYER met2 ;
        RECT 1292.700 1600.000 1292.980 1604.000 ;
        RECT 1292.760 1589.490 1292.900 1600.000 ;
        RECT 1292.700 1589.170 1292.960 1589.490 ;
        RECT 1296.840 1589.170 1297.100 1589.490 ;
        RECT 1296.900 23.450 1297.040 1589.170 ;
        RECT 1296.840 23.130 1297.100 23.450 ;
        RECT 2631.300 23.130 2631.560 23.450 ;
        RECT 2631.360 2.400 2631.500 23.130 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1299.570 1590.760 1299.890 1590.820 ;
        RECT 1303.710 1590.760 1304.030 1590.820 ;
        RECT 1299.570 1590.620 1304.030 1590.760 ;
        RECT 1299.570 1590.560 1299.890 1590.620 ;
        RECT 1303.710 1590.560 1304.030 1590.620 ;
        RECT 1303.710 23.700 1304.030 23.760 ;
        RECT 2649.210 23.700 2649.530 23.760 ;
        RECT 1303.710 23.560 2649.530 23.700 ;
        RECT 1303.710 23.500 1304.030 23.560 ;
        RECT 2649.210 23.500 2649.530 23.560 ;
      LAYER via ;
        RECT 1299.600 1590.560 1299.860 1590.820 ;
        RECT 1303.740 1590.560 1304.000 1590.820 ;
        RECT 1303.740 23.500 1304.000 23.760 ;
        RECT 2649.240 23.500 2649.500 23.760 ;
      LAYER met2 ;
        RECT 1299.600 1600.000 1299.880 1604.000 ;
        RECT 1299.660 1590.850 1299.800 1600.000 ;
        RECT 1299.600 1590.530 1299.860 1590.850 ;
        RECT 1303.740 1590.530 1304.000 1590.850 ;
        RECT 1303.800 23.790 1303.940 1590.530 ;
        RECT 1303.740 23.470 1304.000 23.790 ;
        RECT 2649.240 23.470 2649.500 23.790 ;
        RECT 2649.300 2.400 2649.440 23.470 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1306.470 1589.060 1306.790 1589.120 ;
        RECT 1310.610 1589.060 1310.930 1589.120 ;
        RECT 1306.470 1588.920 1310.930 1589.060 ;
        RECT 1306.470 1588.860 1306.790 1588.920 ;
        RECT 1310.610 1588.860 1310.930 1588.920 ;
        RECT 1310.610 27.440 1310.930 27.500 ;
        RECT 2667.150 27.440 2667.470 27.500 ;
        RECT 1310.610 27.300 2667.470 27.440 ;
        RECT 1310.610 27.240 1310.930 27.300 ;
        RECT 2667.150 27.240 2667.470 27.300 ;
      LAYER via ;
        RECT 1306.500 1588.860 1306.760 1589.120 ;
        RECT 1310.640 1588.860 1310.900 1589.120 ;
        RECT 1310.640 27.240 1310.900 27.500 ;
        RECT 2667.180 27.240 2667.440 27.500 ;
      LAYER met2 ;
        RECT 1306.500 1600.000 1306.780 1604.000 ;
        RECT 1306.560 1589.150 1306.700 1600.000 ;
        RECT 1306.500 1588.830 1306.760 1589.150 ;
        RECT 1310.640 1588.830 1310.900 1589.150 ;
        RECT 1310.700 27.530 1310.840 1588.830 ;
        RECT 1310.640 27.210 1310.900 27.530 ;
        RECT 2667.180 27.210 2667.440 27.530 ;
        RECT 2667.240 2.400 2667.380 27.210 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1312.910 1588.720 1313.230 1588.780 ;
        RECT 1317.510 1588.720 1317.830 1588.780 ;
        RECT 1312.910 1588.580 1317.830 1588.720 ;
        RECT 1312.910 1588.520 1313.230 1588.580 ;
        RECT 1317.510 1588.520 1317.830 1588.580 ;
        RECT 1317.510 27.100 1317.830 27.160 ;
        RECT 2684.630 27.100 2684.950 27.160 ;
        RECT 1317.510 26.960 2684.950 27.100 ;
        RECT 1317.510 26.900 1317.830 26.960 ;
        RECT 2684.630 26.900 2684.950 26.960 ;
      LAYER via ;
        RECT 1312.940 1588.520 1313.200 1588.780 ;
        RECT 1317.540 1588.520 1317.800 1588.780 ;
        RECT 1317.540 26.900 1317.800 27.160 ;
        RECT 2684.660 26.900 2684.920 27.160 ;
      LAYER met2 ;
        RECT 1312.940 1600.000 1313.220 1604.000 ;
        RECT 1313.000 1588.810 1313.140 1600.000 ;
        RECT 1312.940 1588.490 1313.200 1588.810 ;
        RECT 1317.540 1588.490 1317.800 1588.810 ;
        RECT 1317.600 27.190 1317.740 1588.490 ;
        RECT 1317.540 26.870 1317.800 27.190 ;
        RECT 2684.660 26.870 2684.920 27.190 ;
        RECT 2684.720 2.400 2684.860 26.870 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1319.810 1589.400 1320.130 1589.460 ;
        RECT 1324.410 1589.400 1324.730 1589.460 ;
        RECT 1319.810 1589.260 1324.730 1589.400 ;
        RECT 1319.810 1589.200 1320.130 1589.260 ;
        RECT 1324.410 1589.200 1324.730 1589.260 ;
        RECT 1324.410 26.760 1324.730 26.820 ;
        RECT 2702.570 26.760 2702.890 26.820 ;
        RECT 1324.410 26.620 2702.890 26.760 ;
        RECT 1324.410 26.560 1324.730 26.620 ;
        RECT 2702.570 26.560 2702.890 26.620 ;
      LAYER via ;
        RECT 1319.840 1589.200 1320.100 1589.460 ;
        RECT 1324.440 1589.200 1324.700 1589.460 ;
        RECT 1324.440 26.560 1324.700 26.820 ;
        RECT 2702.600 26.560 2702.860 26.820 ;
      LAYER met2 ;
        RECT 1319.840 1600.000 1320.120 1604.000 ;
        RECT 1319.900 1589.490 1320.040 1600.000 ;
        RECT 1319.840 1589.170 1320.100 1589.490 ;
        RECT 1324.440 1589.170 1324.700 1589.490 ;
        RECT 1324.500 26.850 1324.640 1589.170 ;
        RECT 1324.440 26.530 1324.700 26.850 ;
        RECT 2702.600 26.530 2702.860 26.850 ;
        RECT 2702.660 2.400 2702.800 26.530 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1326.250 1590.760 1326.570 1590.820 ;
        RECT 1331.310 1590.760 1331.630 1590.820 ;
        RECT 1326.250 1590.620 1331.630 1590.760 ;
        RECT 1326.250 1590.560 1326.570 1590.620 ;
        RECT 1331.310 1590.560 1331.630 1590.620 ;
        RECT 1331.310 26.420 1331.630 26.480 ;
        RECT 2720.510 26.420 2720.830 26.480 ;
        RECT 1331.310 26.280 2720.830 26.420 ;
        RECT 1331.310 26.220 1331.630 26.280 ;
        RECT 2720.510 26.220 2720.830 26.280 ;
      LAYER via ;
        RECT 1326.280 1590.560 1326.540 1590.820 ;
        RECT 1331.340 1590.560 1331.600 1590.820 ;
        RECT 1331.340 26.220 1331.600 26.480 ;
        RECT 2720.540 26.220 2720.800 26.480 ;
      LAYER met2 ;
        RECT 1326.280 1600.000 1326.560 1604.000 ;
        RECT 1326.340 1590.850 1326.480 1600.000 ;
        RECT 1326.280 1590.530 1326.540 1590.850 ;
        RECT 1331.340 1590.530 1331.600 1590.850 ;
        RECT 1331.400 26.510 1331.540 1590.530 ;
        RECT 1331.340 26.190 1331.600 26.510 ;
        RECT 2720.540 26.190 2720.800 26.510 ;
        RECT 2720.600 2.400 2720.740 26.190 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1333.150 1589.400 1333.470 1589.460 ;
        RECT 1338.210 1589.400 1338.530 1589.460 ;
        RECT 1333.150 1589.260 1338.530 1589.400 ;
        RECT 1333.150 1589.200 1333.470 1589.260 ;
        RECT 1338.210 1589.200 1338.530 1589.260 ;
        RECT 1338.210 26.080 1338.530 26.140 ;
        RECT 2738.450 26.080 2738.770 26.140 ;
        RECT 1338.210 25.940 2738.770 26.080 ;
        RECT 1338.210 25.880 1338.530 25.940 ;
        RECT 2738.450 25.880 2738.770 25.940 ;
      LAYER via ;
        RECT 1333.180 1589.200 1333.440 1589.460 ;
        RECT 1338.240 1589.200 1338.500 1589.460 ;
        RECT 1338.240 25.880 1338.500 26.140 ;
        RECT 2738.480 25.880 2738.740 26.140 ;
      LAYER met2 ;
        RECT 1333.180 1600.000 1333.460 1604.000 ;
        RECT 1333.240 1589.490 1333.380 1600.000 ;
        RECT 1333.180 1589.170 1333.440 1589.490 ;
        RECT 1338.240 1589.170 1338.500 1589.490 ;
        RECT 1338.300 26.170 1338.440 1589.170 ;
        RECT 1338.240 25.850 1338.500 26.170 ;
        RECT 2738.480 25.850 2738.740 26.170 ;
        RECT 2738.540 2.400 2738.680 25.850 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1340.050 1590.760 1340.370 1590.820 ;
        RECT 1345.110 1590.760 1345.430 1590.820 ;
        RECT 1340.050 1590.620 1345.430 1590.760 ;
        RECT 1340.050 1590.560 1340.370 1590.620 ;
        RECT 1345.110 1590.560 1345.430 1590.620 ;
        RECT 1345.110 25.740 1345.430 25.800 ;
        RECT 2755.930 25.740 2756.250 25.800 ;
        RECT 1345.110 25.600 2756.250 25.740 ;
        RECT 1345.110 25.540 1345.430 25.600 ;
        RECT 2755.930 25.540 2756.250 25.600 ;
      LAYER via ;
        RECT 1340.080 1590.560 1340.340 1590.820 ;
        RECT 1345.140 1590.560 1345.400 1590.820 ;
        RECT 1345.140 25.540 1345.400 25.800 ;
        RECT 2755.960 25.540 2756.220 25.800 ;
      LAYER met2 ;
        RECT 1340.080 1600.000 1340.360 1604.000 ;
        RECT 1340.140 1590.850 1340.280 1600.000 ;
        RECT 1340.080 1590.530 1340.340 1590.850 ;
        RECT 1345.140 1590.530 1345.400 1590.850 ;
        RECT 1345.200 25.830 1345.340 1590.530 ;
        RECT 1345.140 25.510 1345.400 25.830 ;
        RECT 2755.960 25.510 2756.220 25.830 ;
        RECT 2756.020 2.400 2756.160 25.510 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 796.865 14.365 797.035 19.295 ;
      LAYER mcon ;
        RECT 796.865 19.125 797.035 19.295 ;
      LAYER met1 ;
        RECT 613.710 19.280 614.030 19.340 ;
        RECT 796.805 19.280 797.095 19.325 ;
        RECT 613.710 19.140 797.095 19.280 ;
        RECT 613.710 19.080 614.030 19.140 ;
        RECT 796.805 19.095 797.095 19.140 ;
        RECT 796.805 14.520 797.095 14.565 ;
        RECT 829.450 14.520 829.770 14.580 ;
        RECT 796.805 14.380 829.770 14.520 ;
        RECT 796.805 14.335 797.095 14.380 ;
        RECT 829.450 14.320 829.770 14.380 ;
      LAYER via ;
        RECT 613.740 19.080 614.000 19.340 ;
        RECT 829.480 14.320 829.740 14.580 ;
      LAYER met2 ;
        RECT 612.820 1600.450 613.100 1604.000 ;
        RECT 612.820 1600.310 613.940 1600.450 ;
        RECT 612.820 1600.000 613.100 1600.310 ;
        RECT 613.800 19.370 613.940 1600.310 ;
        RECT 613.740 19.050 614.000 19.370 ;
        RECT 829.480 14.290 829.740 14.610 ;
        RECT 829.540 2.400 829.680 14.290 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.490 1590.760 1346.810 1590.820 ;
        RECT 1352.010 1590.760 1352.330 1590.820 ;
        RECT 1346.490 1590.620 1352.330 1590.760 ;
        RECT 1346.490 1590.560 1346.810 1590.620 ;
        RECT 1352.010 1590.560 1352.330 1590.620 ;
        RECT 1352.010 25.400 1352.330 25.460 ;
        RECT 2773.870 25.400 2774.190 25.460 ;
        RECT 1352.010 25.260 2774.190 25.400 ;
        RECT 1352.010 25.200 1352.330 25.260 ;
        RECT 2773.870 25.200 2774.190 25.260 ;
      LAYER via ;
        RECT 1346.520 1590.560 1346.780 1590.820 ;
        RECT 1352.040 1590.560 1352.300 1590.820 ;
        RECT 1352.040 25.200 1352.300 25.460 ;
        RECT 2773.900 25.200 2774.160 25.460 ;
      LAYER met2 ;
        RECT 1346.520 1600.000 1346.800 1604.000 ;
        RECT 1346.580 1590.850 1346.720 1600.000 ;
        RECT 1346.520 1590.530 1346.780 1590.850 ;
        RECT 1352.040 1590.530 1352.300 1590.850 ;
        RECT 1352.100 25.490 1352.240 1590.530 ;
        RECT 1352.040 25.170 1352.300 25.490 ;
        RECT 2773.900 25.170 2774.160 25.490 ;
        RECT 2773.960 2.400 2774.100 25.170 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1353.390 1590.760 1353.710 1590.820 ;
        RECT 1358.910 1590.760 1359.230 1590.820 ;
        RECT 1353.390 1590.620 1359.230 1590.760 ;
        RECT 1353.390 1590.560 1353.710 1590.620 ;
        RECT 1358.910 1590.560 1359.230 1590.620 ;
        RECT 1358.910 25.060 1359.230 25.120 ;
        RECT 2791.810 25.060 2792.130 25.120 ;
        RECT 1358.910 24.920 2792.130 25.060 ;
        RECT 1358.910 24.860 1359.230 24.920 ;
        RECT 2791.810 24.860 2792.130 24.920 ;
      LAYER via ;
        RECT 1353.420 1590.560 1353.680 1590.820 ;
        RECT 1358.940 1590.560 1359.200 1590.820 ;
        RECT 1358.940 24.860 1359.200 25.120 ;
        RECT 2791.840 24.860 2792.100 25.120 ;
      LAYER met2 ;
        RECT 1353.420 1600.000 1353.700 1604.000 ;
        RECT 1353.480 1590.850 1353.620 1600.000 ;
        RECT 1353.420 1590.530 1353.680 1590.850 ;
        RECT 1358.940 1590.530 1359.200 1590.850 ;
        RECT 1359.000 25.150 1359.140 1590.530 ;
        RECT 1358.940 24.830 1359.200 25.150 ;
        RECT 2791.840 24.830 2792.100 25.150 ;
        RECT 2791.900 2.400 2792.040 24.830 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1360.290 1590.420 1360.610 1590.480 ;
        RECT 1365.810 1590.420 1366.130 1590.480 ;
        RECT 1360.290 1590.280 1366.130 1590.420 ;
        RECT 1360.290 1590.220 1360.610 1590.280 ;
        RECT 1365.810 1590.220 1366.130 1590.280 ;
        RECT 1365.810 24.720 1366.130 24.780 ;
        RECT 2809.750 24.720 2810.070 24.780 ;
        RECT 1365.810 24.580 2810.070 24.720 ;
        RECT 1365.810 24.520 1366.130 24.580 ;
        RECT 2809.750 24.520 2810.070 24.580 ;
      LAYER via ;
        RECT 1360.320 1590.220 1360.580 1590.480 ;
        RECT 1365.840 1590.220 1366.100 1590.480 ;
        RECT 1365.840 24.520 1366.100 24.780 ;
        RECT 2809.780 24.520 2810.040 24.780 ;
      LAYER met2 ;
        RECT 1360.320 1600.000 1360.600 1604.000 ;
        RECT 1360.380 1590.510 1360.520 1600.000 ;
        RECT 1360.320 1590.190 1360.580 1590.510 ;
        RECT 1365.840 1590.190 1366.100 1590.510 ;
        RECT 1365.900 24.810 1366.040 1590.190 ;
        RECT 1365.840 24.490 1366.100 24.810 ;
        RECT 2809.780 24.490 2810.040 24.810 ;
        RECT 2809.840 2.400 2809.980 24.490 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1366.730 1590.760 1367.050 1590.820 ;
        RECT 1372.710 1590.760 1373.030 1590.820 ;
        RECT 1366.730 1590.620 1373.030 1590.760 ;
        RECT 1366.730 1590.560 1367.050 1590.620 ;
        RECT 1372.710 1590.560 1373.030 1590.620 ;
        RECT 1372.710 24.380 1373.030 24.440 ;
        RECT 2827.690 24.380 2828.010 24.440 ;
        RECT 1372.710 24.240 2828.010 24.380 ;
        RECT 1372.710 24.180 1373.030 24.240 ;
        RECT 2827.690 24.180 2828.010 24.240 ;
      LAYER via ;
        RECT 1366.760 1590.560 1367.020 1590.820 ;
        RECT 1372.740 1590.560 1373.000 1590.820 ;
        RECT 1372.740 24.180 1373.000 24.440 ;
        RECT 2827.720 24.180 2827.980 24.440 ;
      LAYER met2 ;
        RECT 1366.760 1600.000 1367.040 1604.000 ;
        RECT 1366.820 1590.850 1366.960 1600.000 ;
        RECT 1366.760 1590.530 1367.020 1590.850 ;
        RECT 1372.740 1590.530 1373.000 1590.850 ;
        RECT 1372.800 24.470 1372.940 1590.530 ;
        RECT 1372.740 24.150 1373.000 24.470 ;
        RECT 2827.720 24.150 2827.980 24.470 ;
        RECT 2827.780 2.400 2827.920 24.150 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1373.630 1590.420 1373.950 1590.480 ;
        RECT 1379.610 1590.420 1379.930 1590.480 ;
        RECT 1373.630 1590.280 1379.930 1590.420 ;
        RECT 1373.630 1590.220 1373.950 1590.280 ;
        RECT 1379.610 1590.220 1379.930 1590.280 ;
        RECT 1379.610 24.040 1379.930 24.100 ;
        RECT 2845.170 24.040 2845.490 24.100 ;
        RECT 1379.610 23.900 2845.490 24.040 ;
        RECT 1379.610 23.840 1379.930 23.900 ;
        RECT 2845.170 23.840 2845.490 23.900 ;
      LAYER via ;
        RECT 1373.660 1590.220 1373.920 1590.480 ;
        RECT 1379.640 1590.220 1379.900 1590.480 ;
        RECT 1379.640 23.840 1379.900 24.100 ;
        RECT 2845.200 23.840 2845.460 24.100 ;
      LAYER met2 ;
        RECT 1373.660 1600.000 1373.940 1604.000 ;
        RECT 1373.720 1590.510 1373.860 1600.000 ;
        RECT 1373.660 1590.190 1373.920 1590.510 ;
        RECT 1379.640 1590.190 1379.900 1590.510 ;
        RECT 1379.700 24.130 1379.840 1590.190 ;
        RECT 1379.640 23.810 1379.900 24.130 ;
        RECT 2845.200 23.810 2845.460 24.130 ;
        RECT 2845.260 2.400 2845.400 23.810 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.530 1589.400 1380.850 1589.460 ;
        RECT 1386.510 1589.400 1386.830 1589.460 ;
        RECT 1380.530 1589.260 1386.830 1589.400 ;
        RECT 1380.530 1589.200 1380.850 1589.260 ;
        RECT 1386.510 1589.200 1386.830 1589.260 ;
      LAYER via ;
        RECT 1380.560 1589.200 1380.820 1589.460 ;
        RECT 1386.540 1589.200 1386.800 1589.460 ;
      LAYER met2 ;
        RECT 1380.560 1600.000 1380.840 1604.000 ;
        RECT 1380.620 1589.490 1380.760 1600.000 ;
        RECT 1380.560 1589.170 1380.820 1589.490 ;
        RECT 1386.540 1589.170 1386.800 1589.490 ;
        RECT 1386.600 25.685 1386.740 1589.170 ;
        RECT 1386.530 25.315 1386.810 25.685 ;
        RECT 2863.130 25.315 2863.410 25.685 ;
        RECT 2863.200 2.400 2863.340 25.315 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
      LAYER via2 ;
        RECT 1386.530 25.360 1386.810 25.640 ;
        RECT 2863.130 25.360 2863.410 25.640 ;
      LAYER met3 ;
        RECT 1386.505 25.650 1386.835 25.665 ;
        RECT 2863.105 25.650 2863.435 25.665 ;
        RECT 1386.505 25.350 2863.435 25.650 ;
        RECT 1386.505 25.335 1386.835 25.350 ;
        RECT 2863.105 25.335 2863.435 25.350 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.970 1589.060 1387.290 1589.120 ;
        RECT 1393.410 1589.060 1393.730 1589.120 ;
        RECT 1386.970 1588.920 1393.730 1589.060 ;
        RECT 1386.970 1588.860 1387.290 1588.920 ;
        RECT 1393.410 1588.860 1393.730 1588.920 ;
      LAYER via ;
        RECT 1387.000 1588.860 1387.260 1589.120 ;
        RECT 1393.440 1588.860 1393.700 1589.120 ;
      LAYER met2 ;
        RECT 1387.000 1600.000 1387.280 1604.000 ;
        RECT 1387.060 1589.150 1387.200 1600.000 ;
        RECT 1387.000 1588.830 1387.260 1589.150 ;
        RECT 1393.440 1588.830 1393.700 1589.150 ;
        RECT 1393.500 25.005 1393.640 1588.830 ;
        RECT 1393.430 24.635 1393.710 25.005 ;
        RECT 2881.070 24.635 2881.350 25.005 ;
        RECT 2881.140 2.400 2881.280 24.635 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
      LAYER via2 ;
        RECT 1393.430 24.680 1393.710 24.960 ;
        RECT 2881.070 24.680 2881.350 24.960 ;
      LAYER met3 ;
        RECT 1393.405 24.970 1393.735 24.985 ;
        RECT 2881.045 24.970 2881.375 24.985 ;
        RECT 1393.405 24.670 2881.375 24.970 ;
        RECT 1393.405 24.655 1393.735 24.670 ;
        RECT 2881.045 24.655 2881.375 24.670 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1393.870 1589.400 1394.190 1589.460 ;
        RECT 1400.310 1589.400 1400.630 1589.460 ;
        RECT 1393.870 1589.260 1400.630 1589.400 ;
        RECT 1393.870 1589.200 1394.190 1589.260 ;
        RECT 1400.310 1589.200 1400.630 1589.260 ;
      LAYER via ;
        RECT 1393.900 1589.200 1394.160 1589.460 ;
        RECT 1400.340 1589.200 1400.600 1589.460 ;
      LAYER met2 ;
        RECT 1393.900 1600.000 1394.180 1604.000 ;
        RECT 1393.960 1589.490 1394.100 1600.000 ;
        RECT 1393.900 1589.170 1394.160 1589.490 ;
        RECT 1400.340 1589.170 1400.600 1589.490 ;
        RECT 1400.400 24.325 1400.540 1589.170 ;
        RECT 1400.330 23.955 1400.610 24.325 ;
        RECT 2899.010 23.955 2899.290 24.325 ;
        RECT 2899.080 2.400 2899.220 23.955 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
      LAYER via2 ;
        RECT 1400.330 24.000 1400.610 24.280 ;
        RECT 2899.010 24.000 2899.290 24.280 ;
      LAYER met3 ;
        RECT 1400.305 24.290 1400.635 24.305 ;
        RECT 2898.985 24.290 2899.315 24.305 ;
        RECT 1400.305 23.990 2899.315 24.290 ;
        RECT 1400.305 23.975 1400.635 23.990 ;
        RECT 2898.985 23.975 2899.315 23.990 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 619.260 1600.450 619.540 1604.000 ;
        RECT 619.260 1600.310 620.380 1600.450 ;
        RECT 619.260 1600.000 619.540 1600.310 ;
        RECT 620.240 16.165 620.380 1600.310 ;
        RECT 620.170 15.795 620.450 16.165 ;
        RECT 846.950 15.795 847.230 16.165 ;
        RECT 847.020 2.400 847.160 15.795 ;
        RECT 846.810 -4.800 847.370 2.400 ;
      LAYER via2 ;
        RECT 620.170 15.840 620.450 16.120 ;
        RECT 846.950 15.840 847.230 16.120 ;
      LAYER met3 ;
        RECT 620.145 16.130 620.475 16.145 ;
        RECT 846.925 16.130 847.255 16.145 ;
        RECT 620.145 15.830 847.255 16.130 ;
        RECT 620.145 15.815 620.475 15.830 ;
        RECT 846.925 15.815 847.255 15.830 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 665.765 18.785 665.935 19.635 ;
      LAYER mcon ;
        RECT 665.765 19.465 665.935 19.635 ;
      LAYER met1 ;
        RECT 627.510 19.620 627.830 19.680 ;
        RECT 665.705 19.620 665.995 19.665 ;
        RECT 627.510 19.480 665.995 19.620 ;
        RECT 627.510 19.420 627.830 19.480 ;
        RECT 665.705 19.435 665.995 19.480 ;
        RECT 849.690 19.620 850.010 19.680 ;
        RECT 864.870 19.620 865.190 19.680 ;
        RECT 849.690 19.480 865.190 19.620 ;
        RECT 849.690 19.420 850.010 19.480 ;
        RECT 864.870 19.420 865.190 19.480 ;
        RECT 665.705 18.940 665.995 18.985 ;
        RECT 849.690 18.940 850.010 19.000 ;
        RECT 665.705 18.800 850.010 18.940 ;
        RECT 665.705 18.755 665.995 18.800 ;
        RECT 849.690 18.740 850.010 18.800 ;
      LAYER via ;
        RECT 627.540 19.420 627.800 19.680 ;
        RECT 849.720 19.420 849.980 19.680 ;
        RECT 864.900 19.420 865.160 19.680 ;
        RECT 849.720 18.740 849.980 19.000 ;
      LAYER met2 ;
        RECT 626.160 1600.450 626.440 1604.000 ;
        RECT 626.160 1600.310 627.740 1600.450 ;
        RECT 626.160 1600.000 626.440 1600.310 ;
        RECT 627.600 19.710 627.740 1600.310 ;
        RECT 627.540 19.390 627.800 19.710 ;
        RECT 849.720 19.390 849.980 19.710 ;
        RECT 864.900 19.390 865.160 19.710 ;
        RECT 849.780 19.030 849.920 19.390 ;
        RECT 849.720 18.710 849.980 19.030 ;
        RECT 864.960 2.400 865.100 19.390 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 703.485 1588.225 704.575 1588.395 ;
        RECT 677.265 1586.525 677.435 1588.055 ;
        RECT 703.485 1587.545 703.655 1588.225 ;
        RECT 802.385 15.045 803.475 15.215 ;
      LAYER mcon ;
        RECT 704.405 1588.225 704.575 1588.395 ;
        RECT 677.265 1587.885 677.435 1588.055 ;
        RECT 803.305 15.045 803.475 15.215 ;
      LAYER met1 ;
        RECT 704.345 1588.380 704.635 1588.425 ;
        RECT 727.790 1588.380 728.110 1588.440 ;
        RECT 704.345 1588.240 728.110 1588.380 ;
        RECT 704.345 1588.195 704.635 1588.240 ;
        RECT 727.790 1588.180 728.110 1588.240 ;
        RECT 677.205 1588.040 677.495 1588.085 ;
        RECT 655.660 1587.900 677.495 1588.040 ;
        RECT 633.030 1587.020 633.350 1587.080 ;
        RECT 655.660 1587.020 655.800 1587.900 ;
        RECT 677.205 1587.855 677.495 1587.900 ;
        RECT 703.425 1587.700 703.715 1587.745 ;
        RECT 697.060 1587.560 703.715 1587.700 ;
        RECT 697.060 1587.360 697.200 1587.560 ;
        RECT 703.425 1587.515 703.715 1587.560 ;
        RECT 633.030 1586.880 655.800 1587.020 ;
        RECT 696.600 1587.220 697.200 1587.360 ;
        RECT 633.030 1586.820 633.350 1586.880 ;
        RECT 677.205 1586.680 677.495 1586.725 ;
        RECT 696.600 1586.680 696.740 1587.220 ;
        RECT 677.205 1586.540 696.740 1586.680 ;
        RECT 677.205 1586.495 677.495 1586.540 ;
        RECT 802.325 15.200 802.615 15.245 ;
        RECT 762.380 15.060 802.615 15.200 ;
        RECT 727.790 14.520 728.110 14.580 ;
        RECT 762.380 14.520 762.520 15.060 ;
        RECT 802.325 15.015 802.615 15.060 ;
        RECT 803.245 15.200 803.535 15.245 ;
        RECT 882.810 15.200 883.130 15.260 ;
        RECT 803.245 15.060 883.130 15.200 ;
        RECT 803.245 15.015 803.535 15.060 ;
        RECT 882.810 15.000 883.130 15.060 ;
        RECT 727.790 14.380 762.520 14.520 ;
        RECT 727.790 14.320 728.110 14.380 ;
      LAYER via ;
        RECT 727.820 1588.180 728.080 1588.440 ;
        RECT 633.060 1586.820 633.320 1587.080 ;
        RECT 727.820 14.320 728.080 14.580 ;
        RECT 882.840 15.000 883.100 15.260 ;
      LAYER met2 ;
        RECT 633.060 1600.000 633.340 1604.000 ;
        RECT 633.120 1587.110 633.260 1600.000 ;
        RECT 727.820 1588.150 728.080 1588.470 ;
        RECT 633.060 1586.790 633.320 1587.110 ;
        RECT 727.880 14.610 728.020 1588.150 ;
        RECT 882.840 14.970 883.100 15.290 ;
        RECT 727.820 14.290 728.080 14.610 ;
        RECT 882.900 2.400 883.040 14.970 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 789.965 14.705 790.135 15.895 ;
        RECT 865.865 13.685 866.035 15.895 ;
      LAYER mcon ;
        RECT 789.965 15.725 790.135 15.895 ;
        RECT 865.865 15.725 866.035 15.895 ;
      LAYER met1 ;
        RECT 639.470 1589.060 639.790 1589.120 ;
        RECT 742.050 1589.060 742.370 1589.120 ;
        RECT 639.470 1588.920 742.370 1589.060 ;
        RECT 639.470 1588.860 639.790 1588.920 ;
        RECT 742.050 1588.860 742.370 1588.920 ;
        RECT 789.905 15.880 790.195 15.925 ;
        RECT 865.805 15.880 866.095 15.925 ;
        RECT 789.905 15.740 866.095 15.880 ;
        RECT 789.905 15.695 790.195 15.740 ;
        RECT 865.805 15.695 866.095 15.740 ;
        RECT 789.905 14.860 790.195 14.905 ;
        RECT 762.840 14.720 790.195 14.860 ;
        RECT 742.050 14.180 742.370 14.240 ;
        RECT 762.840 14.180 762.980 14.720 ;
        RECT 789.905 14.675 790.195 14.720 ;
        RECT 742.050 14.040 762.980 14.180 ;
        RECT 742.050 13.980 742.370 14.040 ;
        RECT 865.805 13.840 866.095 13.885 ;
        RECT 900.750 13.840 901.070 13.900 ;
        RECT 865.805 13.700 901.070 13.840 ;
        RECT 865.805 13.655 866.095 13.700 ;
        RECT 900.750 13.640 901.070 13.700 ;
      LAYER via ;
        RECT 639.500 1588.860 639.760 1589.120 ;
        RECT 742.080 1588.860 742.340 1589.120 ;
        RECT 742.080 13.980 742.340 14.240 ;
        RECT 900.780 13.640 901.040 13.900 ;
      LAYER met2 ;
        RECT 639.500 1600.000 639.780 1604.000 ;
        RECT 639.560 1589.150 639.700 1600.000 ;
        RECT 639.500 1588.830 639.760 1589.150 ;
        RECT 742.080 1588.830 742.340 1589.150 ;
        RECT 742.140 14.270 742.280 1588.830 ;
        RECT 742.080 13.950 742.340 14.270 ;
        RECT 900.780 13.610 901.040 13.930 ;
        RECT 900.840 2.400 900.980 13.610 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 690.145 1589.245 690.315 1590.095 ;
        RECT 737.525 1589.925 738.155 1590.095 ;
        RECT 737.985 1587.205 738.155 1589.925 ;
        RECT 782.605 16.065 782.775 18.615 ;
      LAYER mcon ;
        RECT 690.145 1589.925 690.315 1590.095 ;
        RECT 782.605 18.445 782.775 18.615 ;
      LAYER met1 ;
        RECT 690.085 1590.080 690.375 1590.125 ;
        RECT 737.465 1590.080 737.755 1590.125 ;
        RECT 690.085 1589.940 737.755 1590.080 ;
        RECT 690.085 1589.895 690.375 1589.940 ;
        RECT 737.465 1589.895 737.755 1589.940 ;
        RECT 646.370 1589.400 646.690 1589.460 ;
        RECT 690.085 1589.400 690.375 1589.445 ;
        RECT 646.370 1589.260 690.375 1589.400 ;
        RECT 646.370 1589.200 646.690 1589.260 ;
        RECT 690.085 1589.215 690.375 1589.260 ;
        RECT 755.390 1587.700 755.710 1587.760 ;
        RECT 740.300 1587.560 755.710 1587.700 ;
        RECT 737.925 1587.360 738.215 1587.405 ;
        RECT 740.300 1587.360 740.440 1587.560 ;
        RECT 755.390 1587.500 755.710 1587.560 ;
        RECT 737.925 1587.220 740.440 1587.360 ;
        RECT 737.925 1587.175 738.215 1587.220 ;
        RECT 755.390 18.600 755.710 18.660 ;
        RECT 782.545 18.600 782.835 18.645 ;
        RECT 755.390 18.460 782.835 18.600 ;
        RECT 755.390 18.400 755.710 18.460 ;
        RECT 782.545 18.415 782.835 18.460 ;
        RECT 884.650 18.600 884.970 18.660 ;
        RECT 918.690 18.600 919.010 18.660 ;
        RECT 884.650 18.460 919.010 18.600 ;
        RECT 884.650 18.400 884.970 18.460 ;
        RECT 918.690 18.400 919.010 18.460 ;
        RECT 782.545 16.220 782.835 16.265 ;
        RECT 883.270 16.220 883.590 16.280 ;
        RECT 782.545 16.080 883.590 16.220 ;
        RECT 782.545 16.035 782.835 16.080 ;
        RECT 883.270 16.020 883.590 16.080 ;
      LAYER via ;
        RECT 646.400 1589.200 646.660 1589.460 ;
        RECT 755.420 1587.500 755.680 1587.760 ;
        RECT 755.420 18.400 755.680 18.660 ;
        RECT 884.680 18.400 884.940 18.660 ;
        RECT 918.720 18.400 918.980 18.660 ;
        RECT 883.300 16.020 883.560 16.280 ;
      LAYER met2 ;
        RECT 646.400 1600.000 646.680 1604.000 ;
        RECT 646.460 1589.490 646.600 1600.000 ;
        RECT 646.400 1589.170 646.660 1589.490 ;
        RECT 755.420 1587.470 755.680 1587.790 ;
        RECT 755.480 18.690 755.620 1587.470 ;
        RECT 755.420 18.370 755.680 18.690 ;
        RECT 884.680 18.370 884.940 18.690 ;
        RECT 918.720 18.370 918.980 18.690 ;
        RECT 884.740 18.090 884.880 18.370 ;
        RECT 883.360 17.950 884.880 18.090 ;
        RECT 883.360 16.310 883.500 17.950 ;
        RECT 883.300 15.990 883.560 16.310 ;
        RECT 918.780 2.400 918.920 18.370 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 737.065 1586.865 737.235 1588.055 ;
        RECT 739.365 1586.865 739.535 1588.395 ;
      LAYER mcon ;
        RECT 739.365 1588.225 739.535 1588.395 ;
        RECT 737.065 1587.885 737.235 1588.055 ;
      LAYER met1 ;
        RECT 653.270 1589.740 653.590 1589.800 ;
        RECT 673.050 1589.740 673.370 1589.800 ;
        RECT 653.270 1589.600 673.370 1589.740 ;
        RECT 653.270 1589.540 653.590 1589.600 ;
        RECT 673.050 1589.540 673.370 1589.600 ;
        RECT 739.305 1588.380 739.595 1588.425 ;
        RECT 762.750 1588.380 763.070 1588.440 ;
        RECT 739.305 1588.240 763.070 1588.380 ;
        RECT 739.305 1588.195 739.595 1588.240 ;
        RECT 762.750 1588.180 763.070 1588.240 ;
        RECT 689.610 1588.040 689.930 1588.100 ;
        RECT 737.005 1588.040 737.295 1588.085 ;
        RECT 689.610 1587.900 737.295 1588.040 ;
        RECT 689.610 1587.840 689.930 1587.900 ;
        RECT 737.005 1587.855 737.295 1587.900 ;
        RECT 737.005 1587.020 737.295 1587.065 ;
        RECT 739.305 1587.020 739.595 1587.065 ;
        RECT 737.005 1586.880 739.595 1587.020 ;
        RECT 737.005 1586.835 737.295 1586.880 ;
        RECT 739.305 1586.835 739.595 1586.880 ;
        RECT 932.030 17.920 932.350 17.980 ;
        RECT 936.170 17.920 936.490 17.980 ;
        RECT 932.030 17.780 936.490 17.920 ;
        RECT 932.030 17.720 932.350 17.780 ;
        RECT 936.170 17.720 936.490 17.780 ;
        RECT 931.570 16.560 931.890 16.620 ;
        RECT 782.160 16.420 931.890 16.560 ;
        RECT 762.750 16.220 763.070 16.280 ;
        RECT 782.160 16.220 782.300 16.420 ;
        RECT 931.570 16.360 931.890 16.420 ;
        RECT 762.750 16.080 782.300 16.220 ;
        RECT 762.750 16.020 763.070 16.080 ;
      LAYER via ;
        RECT 653.300 1589.540 653.560 1589.800 ;
        RECT 673.080 1589.540 673.340 1589.800 ;
        RECT 762.780 1588.180 763.040 1588.440 ;
        RECT 689.640 1587.840 689.900 1588.100 ;
        RECT 932.060 17.720 932.320 17.980 ;
        RECT 936.200 17.720 936.460 17.980 ;
        RECT 762.780 16.020 763.040 16.280 ;
        RECT 931.600 16.360 931.860 16.620 ;
      LAYER met2 ;
        RECT 653.300 1600.000 653.580 1604.000 ;
        RECT 653.360 1589.830 653.500 1600.000 ;
        RECT 653.300 1589.510 653.560 1589.830 ;
        RECT 673.080 1589.685 673.340 1589.830 ;
        RECT 673.070 1589.315 673.350 1589.685 ;
        RECT 689.630 1589.315 689.910 1589.685 ;
        RECT 689.700 1588.130 689.840 1589.315 ;
        RECT 762.780 1588.150 763.040 1588.470 ;
        RECT 689.640 1587.810 689.900 1588.130 ;
        RECT 762.840 16.310 762.980 1588.150 ;
        RECT 932.060 17.690 932.320 18.010 ;
        RECT 936.200 17.690 936.460 18.010 ;
        RECT 932.120 17.410 932.260 17.690 ;
        RECT 931.660 17.270 932.260 17.410 ;
        RECT 931.660 16.650 931.800 17.270 ;
        RECT 931.600 16.330 931.860 16.650 ;
        RECT 762.780 15.990 763.040 16.310 ;
        RECT 936.260 2.400 936.400 17.690 ;
        RECT 936.050 -4.800 936.610 2.400 ;
      LAYER via2 ;
        RECT 673.070 1589.360 673.350 1589.640 ;
        RECT 689.630 1589.360 689.910 1589.640 ;
      LAYER met3 ;
        RECT 673.045 1589.650 673.375 1589.665 ;
        RECT 689.605 1589.650 689.935 1589.665 ;
        RECT 673.045 1589.350 689.935 1589.650 ;
        RECT 673.045 1589.335 673.375 1589.350 ;
        RECT 689.605 1589.335 689.935 1589.350 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 749.025 1589.585 749.195 1593.495 ;
        RECT 763.745 1589.245 763.915 1590.435 ;
        RECT 809.285 20.485 810.375 20.655 ;
        RECT 809.285 20.145 809.455 20.485 ;
      LAYER mcon ;
        RECT 749.025 1593.325 749.195 1593.495 ;
        RECT 763.745 1590.265 763.915 1590.435 ;
        RECT 810.205 20.485 810.375 20.655 ;
      LAYER met1 ;
        RECT 690.530 1593.820 690.850 1593.880 ;
        RECT 690.530 1593.680 728.940 1593.820 ;
        RECT 690.530 1593.620 690.850 1593.680 ;
        RECT 728.800 1593.480 728.940 1593.680 ;
        RECT 748.965 1593.480 749.255 1593.525 ;
        RECT 728.800 1593.340 749.255 1593.480 ;
        RECT 748.965 1593.295 749.255 1593.340 ;
        RECT 763.685 1590.420 763.975 1590.465 ;
        RECT 769.190 1590.420 769.510 1590.480 ;
        RECT 763.685 1590.280 769.510 1590.420 ;
        RECT 763.685 1590.235 763.975 1590.280 ;
        RECT 769.190 1590.220 769.510 1590.280 ;
        RECT 748.965 1589.740 749.255 1589.785 ;
        RECT 748.965 1589.600 761.600 1589.740 ;
        RECT 748.965 1589.555 749.255 1589.600 ;
        RECT 761.460 1589.400 761.600 1589.600 ;
        RECT 763.685 1589.400 763.975 1589.445 ;
        RECT 761.460 1589.260 763.975 1589.400 ;
        RECT 763.685 1589.215 763.975 1589.260 ;
        RECT 659.710 1588.380 660.030 1588.440 ;
        RECT 690.070 1588.380 690.390 1588.440 ;
        RECT 659.710 1588.240 690.390 1588.380 ;
        RECT 659.710 1588.180 660.030 1588.240 ;
        RECT 690.070 1588.180 690.390 1588.240 ;
        RECT 810.145 20.640 810.435 20.685 ;
        RECT 810.145 20.500 935.020 20.640 ;
        RECT 810.145 20.455 810.435 20.500 ;
        RECT 769.190 20.300 769.510 20.360 ;
        RECT 809.225 20.300 809.515 20.345 ;
        RECT 769.190 20.160 809.515 20.300 ;
        RECT 769.190 20.100 769.510 20.160 ;
        RECT 809.225 20.115 809.515 20.160 ;
        RECT 934.880 19.960 935.020 20.500 ;
        RECT 954.110 19.960 954.430 20.020 ;
        RECT 934.880 19.820 954.430 19.960 ;
        RECT 954.110 19.760 954.430 19.820 ;
      LAYER via ;
        RECT 690.560 1593.620 690.820 1593.880 ;
        RECT 769.220 1590.220 769.480 1590.480 ;
        RECT 659.740 1588.180 660.000 1588.440 ;
        RECT 690.100 1588.180 690.360 1588.440 ;
        RECT 769.220 20.100 769.480 20.360 ;
        RECT 954.140 19.760 954.400 20.020 ;
      LAYER met2 ;
        RECT 659.740 1600.000 660.020 1604.000 ;
        RECT 659.800 1588.470 659.940 1600.000 ;
        RECT 690.560 1593.590 690.820 1593.910 ;
        RECT 690.620 1588.890 690.760 1593.590 ;
        RECT 769.220 1590.190 769.480 1590.510 ;
        RECT 690.160 1588.750 690.760 1588.890 ;
        RECT 690.160 1588.470 690.300 1588.750 ;
        RECT 659.740 1588.150 660.000 1588.470 ;
        RECT 690.100 1588.150 690.360 1588.470 ;
        RECT 769.280 20.390 769.420 1590.190 ;
        RECT 769.220 20.070 769.480 20.390 ;
        RECT 954.140 19.730 954.400 20.050 ;
        RECT 954.200 2.400 954.340 19.730 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 738.905 1588.735 739.075 1590.095 ;
        RECT 757.305 1588.905 757.475 1590.095 ;
        RECT 692.905 1587.205 693.075 1588.735 ;
        RECT 738.445 1588.565 739.075 1588.735 ;
        RECT 809.745 20.145 810.835 20.315 ;
        RECT 933.945 18.615 934.115 19.975 ;
        RECT 935.785 18.615 935.955 18.955 ;
        RECT 933.945 18.445 935.955 18.615 ;
        RECT 951.885 18.105 952.055 18.955 ;
      LAYER mcon ;
        RECT 738.905 1589.925 739.075 1590.095 ;
        RECT 757.305 1589.925 757.475 1590.095 ;
        RECT 692.905 1588.565 693.075 1588.735 ;
        RECT 810.665 20.145 810.835 20.315 ;
        RECT 933.945 19.805 934.115 19.975 ;
        RECT 935.785 18.785 935.955 18.955 ;
        RECT 951.885 18.785 952.055 18.955 ;
      LAYER met1 ;
        RECT 738.845 1590.080 739.135 1590.125 ;
        RECT 757.245 1590.080 757.535 1590.125 ;
        RECT 738.845 1589.940 757.535 1590.080 ;
        RECT 738.845 1589.895 739.135 1589.940 ;
        RECT 757.245 1589.895 757.535 1589.940 ;
        RECT 757.245 1589.060 757.535 1589.105 ;
        RECT 776.090 1589.060 776.410 1589.120 ;
        RECT 757.245 1588.920 776.410 1589.060 ;
        RECT 757.245 1588.875 757.535 1588.920 ;
        RECT 776.090 1588.860 776.410 1588.920 ;
        RECT 692.845 1588.720 693.135 1588.765 ;
        RECT 738.385 1588.720 738.675 1588.765 ;
        RECT 692.845 1588.580 738.675 1588.720 ;
        RECT 692.845 1588.535 693.135 1588.580 ;
        RECT 738.385 1588.535 738.675 1588.580 ;
        RECT 666.610 1587.700 666.930 1587.760 ;
        RECT 666.610 1587.560 688.920 1587.700 ;
        RECT 666.610 1587.500 666.930 1587.560 ;
        RECT 688.780 1587.360 688.920 1587.560 ;
        RECT 692.845 1587.360 693.135 1587.405 ;
        RECT 688.780 1587.220 693.135 1587.360 ;
        RECT 692.845 1587.175 693.135 1587.220 ;
        RECT 776.090 20.640 776.410 20.700 ;
        RECT 776.090 20.500 809.900 20.640 ;
        RECT 776.090 20.440 776.410 20.500 ;
        RECT 809.760 20.345 809.900 20.500 ;
        RECT 809.685 20.115 809.975 20.345 ;
        RECT 810.605 20.300 810.895 20.345 ;
        RECT 810.605 20.160 932.720 20.300 ;
        RECT 810.605 20.115 810.895 20.160 ;
        RECT 932.580 19.960 932.720 20.160 ;
        RECT 933.885 19.960 934.175 20.005 ;
        RECT 932.580 19.820 934.175 19.960 ;
        RECT 933.885 19.775 934.175 19.820 ;
        RECT 935.725 18.940 936.015 18.985 ;
        RECT 951.825 18.940 952.115 18.985 ;
        RECT 935.725 18.800 952.115 18.940 ;
        RECT 935.725 18.755 936.015 18.800 ;
        RECT 951.825 18.755 952.115 18.800 ;
        RECT 951.825 18.260 952.115 18.305 ;
        RECT 972.050 18.260 972.370 18.320 ;
        RECT 951.825 18.120 972.370 18.260 ;
        RECT 951.825 18.075 952.115 18.120 ;
        RECT 972.050 18.060 972.370 18.120 ;
      LAYER via ;
        RECT 776.120 1588.860 776.380 1589.120 ;
        RECT 666.640 1587.500 666.900 1587.760 ;
        RECT 776.120 20.440 776.380 20.700 ;
        RECT 972.080 18.060 972.340 18.320 ;
      LAYER met2 ;
        RECT 666.640 1600.000 666.920 1604.000 ;
        RECT 666.700 1587.790 666.840 1600.000 ;
        RECT 776.120 1588.830 776.380 1589.150 ;
        RECT 666.640 1587.470 666.900 1587.790 ;
        RECT 776.180 20.730 776.320 1588.830 ;
        RECT 776.120 20.410 776.380 20.730 ;
        RECT 972.080 18.030 972.340 18.350 ;
        RECT 972.140 2.400 972.280 18.030 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 545.170 1587.360 545.490 1587.420 ;
        RECT 551.610 1587.360 551.930 1587.420 ;
        RECT 545.170 1587.220 551.930 1587.360 ;
        RECT 545.170 1587.160 545.490 1587.220 ;
        RECT 551.610 1587.160 551.930 1587.220 ;
        RECT 551.610 15.540 551.930 15.600 ;
        RECT 650.970 15.540 651.290 15.600 ;
        RECT 551.610 15.400 651.290 15.540 ;
        RECT 551.610 15.340 551.930 15.400 ;
        RECT 650.970 15.340 651.290 15.400 ;
      LAYER via ;
        RECT 545.200 1587.160 545.460 1587.420 ;
        RECT 551.640 1587.160 551.900 1587.420 ;
        RECT 551.640 15.340 551.900 15.600 ;
        RECT 651.000 15.340 651.260 15.600 ;
      LAYER met2 ;
        RECT 545.200 1600.000 545.480 1604.000 ;
        RECT 545.260 1587.450 545.400 1600.000 ;
        RECT 545.200 1587.130 545.460 1587.450 ;
        RECT 551.640 1587.130 551.900 1587.450 ;
        RECT 551.700 15.630 551.840 1587.130 ;
        RECT 551.640 15.310 551.900 15.630 ;
        RECT 651.000 15.310 651.260 15.630 ;
        RECT 651.060 2.400 651.200 15.310 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 717.745 1587.545 717.915 1589.755 ;
        RECT 739.825 1587.885 742.295 1588.055 ;
        RECT 739.825 1587.545 739.995 1587.885 ;
      LAYER mcon ;
        RECT 717.745 1589.585 717.915 1589.755 ;
        RECT 742.125 1587.885 742.295 1588.055 ;
      LAYER met1 ;
        RECT 673.510 1589.740 673.830 1589.800 ;
        RECT 717.685 1589.740 717.975 1589.785 ;
        RECT 673.510 1589.600 717.975 1589.740 ;
        RECT 673.510 1589.540 673.830 1589.600 ;
        RECT 717.685 1589.555 717.975 1589.600 ;
        RECT 742.065 1588.040 742.355 1588.085 ;
        RECT 782.990 1588.040 783.310 1588.100 ;
        RECT 742.065 1587.900 783.310 1588.040 ;
        RECT 742.065 1587.855 742.355 1587.900 ;
        RECT 782.990 1587.840 783.310 1587.900 ;
        RECT 717.685 1587.700 717.975 1587.745 ;
        RECT 739.765 1587.700 740.055 1587.745 ;
        RECT 717.685 1587.560 740.055 1587.700 ;
        RECT 717.685 1587.515 717.975 1587.560 ;
        RECT 739.765 1587.515 740.055 1587.560 ;
        RECT 782.990 14.180 783.310 14.240 ;
        RECT 989.990 14.180 990.310 14.240 ;
        RECT 782.990 14.040 990.310 14.180 ;
        RECT 782.990 13.980 783.310 14.040 ;
        RECT 989.990 13.980 990.310 14.040 ;
      LAYER via ;
        RECT 673.540 1589.540 673.800 1589.800 ;
        RECT 783.020 1587.840 783.280 1588.100 ;
        RECT 783.020 13.980 783.280 14.240 ;
        RECT 990.020 13.980 990.280 14.240 ;
      LAYER met2 ;
        RECT 673.540 1600.000 673.820 1604.000 ;
        RECT 673.600 1589.830 673.740 1600.000 ;
        RECT 673.540 1589.510 673.800 1589.830 ;
        RECT 783.020 1587.810 783.280 1588.130 ;
        RECT 783.080 14.270 783.220 1587.810 ;
        RECT 783.020 13.950 783.280 14.270 ;
        RECT 990.020 13.950 990.280 14.270 ;
        RECT 990.080 2.400 990.220 13.950 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 679.950 1595.180 680.270 1595.240 ;
        RECT 682.710 1595.180 683.030 1595.240 ;
        RECT 679.950 1595.040 683.030 1595.180 ;
        RECT 679.950 1594.980 680.270 1595.040 ;
        RECT 682.710 1594.980 683.030 1595.040 ;
        RECT 682.710 20.980 683.030 21.040 ;
        RECT 1007.470 20.980 1007.790 21.040 ;
        RECT 682.710 20.840 1007.790 20.980 ;
        RECT 682.710 20.780 683.030 20.840 ;
        RECT 1007.470 20.780 1007.790 20.840 ;
      LAYER via ;
        RECT 679.980 1594.980 680.240 1595.240 ;
        RECT 682.740 1594.980 683.000 1595.240 ;
        RECT 682.740 20.780 683.000 21.040 ;
        RECT 1007.500 20.780 1007.760 21.040 ;
      LAYER met2 ;
        RECT 679.980 1600.000 680.260 1604.000 ;
        RECT 680.040 1595.270 680.180 1600.000 ;
        RECT 679.980 1594.950 680.240 1595.270 ;
        RECT 682.740 1594.950 683.000 1595.270 ;
        RECT 682.800 21.070 682.940 1594.950 ;
        RECT 682.740 20.750 683.000 21.070 ;
        RECT 1007.500 20.750 1007.760 21.070 ;
        RECT 1007.560 2.400 1007.700 20.750 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 689.150 21.320 689.470 21.380 ;
        RECT 1025.410 21.320 1025.730 21.380 ;
        RECT 689.150 21.180 1025.730 21.320 ;
        RECT 689.150 21.120 689.470 21.180 ;
        RECT 1025.410 21.120 1025.730 21.180 ;
      LAYER via ;
        RECT 689.180 21.120 689.440 21.380 ;
        RECT 1025.440 21.120 1025.700 21.380 ;
      LAYER met2 ;
        RECT 686.880 1600.450 687.160 1604.000 ;
        RECT 686.880 1600.310 688.000 1600.450 ;
        RECT 686.880 1600.000 687.160 1600.310 ;
        RECT 687.860 1580.050 688.000 1600.310 ;
        RECT 687.860 1579.910 689.380 1580.050 ;
        RECT 689.240 21.410 689.380 1579.910 ;
        RECT 689.180 21.090 689.440 21.410 ;
        RECT 1025.440 21.090 1025.700 21.410 ;
        RECT 1025.500 2.400 1025.640 21.090 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 693.290 1587.360 693.610 1587.420 ;
        RECT 696.050 1587.360 696.370 1587.420 ;
        RECT 693.290 1587.220 696.370 1587.360 ;
        RECT 693.290 1587.160 693.610 1587.220 ;
        RECT 696.050 1587.160 696.370 1587.220 ;
        RECT 696.050 21.660 696.370 21.720 ;
        RECT 1043.350 21.660 1043.670 21.720 ;
        RECT 696.050 21.520 1043.670 21.660 ;
        RECT 696.050 21.460 696.370 21.520 ;
        RECT 1043.350 21.460 1043.670 21.520 ;
      LAYER via ;
        RECT 693.320 1587.160 693.580 1587.420 ;
        RECT 696.080 1587.160 696.340 1587.420 ;
        RECT 696.080 21.460 696.340 21.720 ;
        RECT 1043.380 21.460 1043.640 21.720 ;
      LAYER met2 ;
        RECT 693.320 1600.000 693.600 1604.000 ;
        RECT 693.380 1587.450 693.520 1600.000 ;
        RECT 693.320 1587.130 693.580 1587.450 ;
        RECT 696.080 1587.130 696.340 1587.450 ;
        RECT 696.140 21.750 696.280 1587.130 ;
        RECT 696.080 21.430 696.340 21.750 ;
        RECT 1043.380 21.430 1043.640 21.750 ;
        RECT 1043.440 2.400 1043.580 21.430 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 700.190 1587.360 700.510 1587.420 ;
        RECT 702.950 1587.360 703.270 1587.420 ;
        RECT 700.190 1587.220 703.270 1587.360 ;
        RECT 700.190 1587.160 700.510 1587.220 ;
        RECT 702.950 1587.160 703.270 1587.220 ;
        RECT 702.950 22.000 703.270 22.060 ;
        RECT 1061.290 22.000 1061.610 22.060 ;
        RECT 702.950 21.860 1061.610 22.000 ;
        RECT 702.950 21.800 703.270 21.860 ;
        RECT 1061.290 21.800 1061.610 21.860 ;
      LAYER via ;
        RECT 700.220 1587.160 700.480 1587.420 ;
        RECT 702.980 1587.160 703.240 1587.420 ;
        RECT 702.980 21.800 703.240 22.060 ;
        RECT 1061.320 21.800 1061.580 22.060 ;
      LAYER met2 ;
        RECT 700.220 1600.000 700.500 1604.000 ;
        RECT 700.280 1587.450 700.420 1600.000 ;
        RECT 700.220 1587.130 700.480 1587.450 ;
        RECT 702.980 1587.130 703.240 1587.450 ;
        RECT 703.040 22.090 703.180 1587.130 ;
        RECT 702.980 21.770 703.240 22.090 ;
        RECT 1061.320 21.770 1061.580 22.090 ;
        RECT 1061.380 2.400 1061.520 21.770 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 707.090 1587.360 707.410 1587.420 ;
        RECT 709.850 1587.360 710.170 1587.420 ;
        RECT 707.090 1587.220 710.170 1587.360 ;
        RECT 707.090 1587.160 707.410 1587.220 ;
        RECT 709.850 1587.160 710.170 1587.220 ;
        RECT 709.850 22.340 710.170 22.400 ;
        RECT 1079.230 22.340 1079.550 22.400 ;
        RECT 709.850 22.200 1079.550 22.340 ;
        RECT 709.850 22.140 710.170 22.200 ;
        RECT 1079.230 22.140 1079.550 22.200 ;
      LAYER via ;
        RECT 707.120 1587.160 707.380 1587.420 ;
        RECT 709.880 1587.160 710.140 1587.420 ;
        RECT 709.880 22.140 710.140 22.400 ;
        RECT 1079.260 22.140 1079.520 22.400 ;
      LAYER met2 ;
        RECT 707.120 1600.000 707.400 1604.000 ;
        RECT 707.180 1587.450 707.320 1600.000 ;
        RECT 707.120 1587.130 707.380 1587.450 ;
        RECT 709.880 1587.130 710.140 1587.450 ;
        RECT 709.940 22.430 710.080 1587.130 ;
        RECT 709.880 22.110 710.140 22.430 ;
        RECT 1079.260 22.110 1079.520 22.430 ;
        RECT 1079.320 2.400 1079.460 22.110 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 713.530 1587.360 713.850 1587.420 ;
        RECT 716.750 1587.360 717.070 1587.420 ;
        RECT 713.530 1587.220 717.070 1587.360 ;
        RECT 713.530 1587.160 713.850 1587.220 ;
        RECT 716.750 1587.160 717.070 1587.220 ;
        RECT 716.750 22.680 717.070 22.740 ;
        RECT 1096.710 22.680 1097.030 22.740 ;
        RECT 716.750 22.540 1097.030 22.680 ;
        RECT 716.750 22.480 717.070 22.540 ;
        RECT 1096.710 22.480 1097.030 22.540 ;
      LAYER via ;
        RECT 713.560 1587.160 713.820 1587.420 ;
        RECT 716.780 1587.160 717.040 1587.420 ;
        RECT 716.780 22.480 717.040 22.740 ;
        RECT 1096.740 22.480 1097.000 22.740 ;
      LAYER met2 ;
        RECT 713.560 1600.000 713.840 1604.000 ;
        RECT 713.620 1587.450 713.760 1600.000 ;
        RECT 713.560 1587.130 713.820 1587.450 ;
        RECT 716.780 1587.130 717.040 1587.450 ;
        RECT 716.840 22.770 716.980 1587.130 ;
        RECT 716.780 22.450 717.040 22.770 ;
        RECT 1096.740 22.450 1097.000 22.770 ;
        RECT 1096.800 2.400 1096.940 22.450 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 720.430 1587.360 720.750 1587.420 ;
        RECT 723.650 1587.360 723.970 1587.420 ;
        RECT 720.430 1587.220 723.970 1587.360 ;
        RECT 720.430 1587.160 720.750 1587.220 ;
        RECT 723.650 1587.160 723.970 1587.220 ;
        RECT 723.650 23.020 723.970 23.080 ;
        RECT 1114.650 23.020 1114.970 23.080 ;
        RECT 723.650 22.880 1114.970 23.020 ;
        RECT 723.650 22.820 723.970 22.880 ;
        RECT 1114.650 22.820 1114.970 22.880 ;
      LAYER via ;
        RECT 720.460 1587.160 720.720 1587.420 ;
        RECT 723.680 1587.160 723.940 1587.420 ;
        RECT 723.680 22.820 723.940 23.080 ;
        RECT 1114.680 22.820 1114.940 23.080 ;
      LAYER met2 ;
        RECT 720.460 1600.000 720.740 1604.000 ;
        RECT 720.520 1587.450 720.660 1600.000 ;
        RECT 720.460 1587.130 720.720 1587.450 ;
        RECT 723.680 1587.130 723.940 1587.450 ;
        RECT 723.740 23.110 723.880 1587.130 ;
        RECT 723.680 22.790 723.940 23.110 ;
        RECT 1114.680 22.790 1114.940 23.110 ;
        RECT 1114.740 2.400 1114.880 22.790 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 727.330 1587.360 727.650 1587.420 ;
        RECT 731.010 1587.360 731.330 1587.420 ;
        RECT 727.330 1587.220 731.330 1587.360 ;
        RECT 727.330 1587.160 727.650 1587.220 ;
        RECT 731.010 1587.160 731.330 1587.220 ;
        RECT 731.010 23.360 731.330 23.420 ;
        RECT 1132.590 23.360 1132.910 23.420 ;
        RECT 731.010 23.220 1132.910 23.360 ;
        RECT 731.010 23.160 731.330 23.220 ;
        RECT 1132.590 23.160 1132.910 23.220 ;
      LAYER via ;
        RECT 727.360 1587.160 727.620 1587.420 ;
        RECT 731.040 1587.160 731.300 1587.420 ;
        RECT 731.040 23.160 731.300 23.420 ;
        RECT 1132.620 23.160 1132.880 23.420 ;
      LAYER met2 ;
        RECT 727.360 1600.000 727.640 1604.000 ;
        RECT 727.420 1587.450 727.560 1600.000 ;
        RECT 727.360 1587.130 727.620 1587.450 ;
        RECT 731.040 1587.130 731.300 1587.450 ;
        RECT 731.100 23.450 731.240 1587.130 ;
        RECT 731.040 23.130 731.300 23.450 ;
        RECT 1132.620 23.130 1132.880 23.450 ;
        RECT 1132.680 2.400 1132.820 23.130 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 733.770 1589.740 734.090 1589.800 ;
        RECT 737.910 1589.740 738.230 1589.800 ;
        RECT 733.770 1589.600 738.230 1589.740 ;
        RECT 733.770 1589.540 734.090 1589.600 ;
        RECT 737.910 1589.540 738.230 1589.600 ;
        RECT 737.910 23.700 738.230 23.760 ;
        RECT 1150.530 23.700 1150.850 23.760 ;
        RECT 737.910 23.560 1150.850 23.700 ;
        RECT 737.910 23.500 738.230 23.560 ;
        RECT 1150.530 23.500 1150.850 23.560 ;
      LAYER via ;
        RECT 733.800 1589.540 734.060 1589.800 ;
        RECT 737.940 1589.540 738.200 1589.800 ;
        RECT 737.940 23.500 738.200 23.760 ;
        RECT 1150.560 23.500 1150.820 23.760 ;
      LAYER met2 ;
        RECT 733.800 1600.000 734.080 1604.000 ;
        RECT 733.860 1589.830 734.000 1600.000 ;
        RECT 733.800 1589.510 734.060 1589.830 ;
        RECT 737.940 1589.510 738.200 1589.830 ;
        RECT 738.000 23.790 738.140 1589.510 ;
        RECT 737.940 23.470 738.200 23.790 ;
        RECT 1150.560 23.470 1150.820 23.790 ;
        RECT 1150.620 2.400 1150.760 23.470 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 656.565 18.445 658.115 18.615 ;
      LAYER mcon ;
        RECT 657.945 18.445 658.115 18.615 ;
      LAYER met1 ;
        RECT 552.070 1590.080 552.390 1590.140 ;
        RECT 638.090 1590.080 638.410 1590.140 ;
        RECT 552.070 1589.940 638.410 1590.080 ;
        RECT 552.070 1589.880 552.390 1589.940 ;
        RECT 638.090 1589.880 638.410 1589.940 ;
        RECT 638.090 18.600 638.410 18.660 ;
        RECT 656.505 18.600 656.795 18.645 ;
        RECT 638.090 18.460 656.795 18.600 ;
        RECT 638.090 18.400 638.410 18.460 ;
        RECT 656.505 18.415 656.795 18.460 ;
        RECT 657.885 18.600 658.175 18.645 ;
        RECT 668.910 18.600 669.230 18.660 ;
        RECT 657.885 18.460 669.230 18.600 ;
        RECT 657.885 18.415 658.175 18.460 ;
        RECT 668.910 18.400 669.230 18.460 ;
      LAYER via ;
        RECT 552.100 1589.880 552.360 1590.140 ;
        RECT 638.120 1589.880 638.380 1590.140 ;
        RECT 638.120 18.400 638.380 18.660 ;
        RECT 668.940 18.400 669.200 18.660 ;
      LAYER met2 ;
        RECT 552.100 1600.000 552.380 1604.000 ;
        RECT 552.160 1590.170 552.300 1600.000 ;
        RECT 552.100 1589.850 552.360 1590.170 ;
        RECT 638.120 1589.850 638.380 1590.170 ;
        RECT 638.180 18.690 638.320 1589.850 ;
        RECT 638.120 18.370 638.380 18.690 ;
        RECT 668.940 18.370 669.200 18.690 ;
        RECT 669.000 2.400 669.140 18.370 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 740.670 1587.360 740.990 1587.420 ;
        RECT 744.810 1587.360 745.130 1587.420 ;
        RECT 740.670 1587.220 745.130 1587.360 ;
        RECT 740.670 1587.160 740.990 1587.220 ;
        RECT 744.810 1587.160 745.130 1587.220 ;
        RECT 744.810 27.440 745.130 27.500 ;
        RECT 1168.470 27.440 1168.790 27.500 ;
        RECT 744.810 27.300 1168.790 27.440 ;
        RECT 744.810 27.240 745.130 27.300 ;
        RECT 1168.470 27.240 1168.790 27.300 ;
      LAYER via ;
        RECT 740.700 1587.160 740.960 1587.420 ;
        RECT 744.840 1587.160 745.100 1587.420 ;
        RECT 744.840 27.240 745.100 27.500 ;
        RECT 1168.500 27.240 1168.760 27.500 ;
      LAYER met2 ;
        RECT 740.700 1600.000 740.980 1604.000 ;
        RECT 740.760 1587.450 740.900 1600.000 ;
        RECT 740.700 1587.130 740.960 1587.450 ;
        RECT 744.840 1587.130 745.100 1587.450 ;
        RECT 744.900 27.530 745.040 1587.130 ;
        RECT 744.840 27.210 745.100 27.530 ;
        RECT 1168.500 27.210 1168.760 27.530 ;
        RECT 1168.560 2.400 1168.700 27.210 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 751.325 786.505 751.495 821.015 ;
        RECT 751.325 689.605 751.495 724.455 ;
        RECT 751.325 593.045 751.495 627.895 ;
        RECT 751.325 496.485 751.495 531.335 ;
        RECT 751.325 386.325 751.495 434.775 ;
        RECT 751.325 241.485 751.495 289.595 ;
        RECT 751.325 144.925 751.495 193.035 ;
      LAYER mcon ;
        RECT 751.325 820.845 751.495 821.015 ;
        RECT 751.325 724.285 751.495 724.455 ;
        RECT 751.325 627.725 751.495 627.895 ;
        RECT 751.325 531.165 751.495 531.335 ;
        RECT 751.325 434.605 751.495 434.775 ;
        RECT 751.325 289.425 751.495 289.595 ;
        RECT 751.325 192.865 751.495 193.035 ;
      LAYER met1 ;
        RECT 747.570 1587.360 747.890 1587.420 ;
        RECT 750.790 1587.360 751.110 1587.420 ;
        RECT 747.570 1587.220 751.110 1587.360 ;
        RECT 747.570 1587.160 747.890 1587.220 ;
        RECT 750.790 1587.160 751.110 1587.220 ;
        RECT 750.790 1414.640 751.110 1414.700 ;
        RECT 751.710 1414.640 752.030 1414.700 ;
        RECT 750.790 1414.500 752.030 1414.640 ;
        RECT 750.790 1414.440 751.110 1414.500 ;
        RECT 751.710 1414.440 752.030 1414.500 ;
        RECT 750.790 1318.080 751.110 1318.140 ;
        RECT 751.710 1318.080 752.030 1318.140 ;
        RECT 750.790 1317.940 752.030 1318.080 ;
        RECT 750.790 1317.880 751.110 1317.940 ;
        RECT 751.710 1317.880 752.030 1317.940 ;
        RECT 750.790 1221.520 751.110 1221.580 ;
        RECT 751.710 1221.520 752.030 1221.580 ;
        RECT 750.790 1221.380 752.030 1221.520 ;
        RECT 750.790 1221.320 751.110 1221.380 ;
        RECT 751.710 1221.320 752.030 1221.380 ;
        RECT 750.790 1124.960 751.110 1125.020 ;
        RECT 751.710 1124.960 752.030 1125.020 ;
        RECT 750.790 1124.820 752.030 1124.960 ;
        RECT 750.790 1124.760 751.110 1124.820 ;
        RECT 751.710 1124.760 752.030 1124.820 ;
        RECT 750.790 1028.400 751.110 1028.460 ;
        RECT 751.710 1028.400 752.030 1028.460 ;
        RECT 750.790 1028.260 752.030 1028.400 ;
        RECT 750.790 1028.200 751.110 1028.260 ;
        RECT 751.710 1028.200 752.030 1028.260 ;
        RECT 750.790 931.840 751.110 931.900 ;
        RECT 751.710 931.840 752.030 931.900 ;
        RECT 750.790 931.700 752.030 931.840 ;
        RECT 750.790 931.640 751.110 931.700 ;
        RECT 751.710 931.640 752.030 931.700 ;
        RECT 750.330 869.620 750.650 869.680 ;
        RECT 751.710 869.620 752.030 869.680 ;
        RECT 750.330 869.480 752.030 869.620 ;
        RECT 750.330 869.420 750.650 869.480 ;
        RECT 751.710 869.420 752.030 869.480 ;
        RECT 750.790 835.280 751.110 835.340 ;
        RECT 751.710 835.280 752.030 835.340 ;
        RECT 750.790 835.140 752.030 835.280 ;
        RECT 750.790 835.080 751.110 835.140 ;
        RECT 751.710 835.080 752.030 835.140 ;
        RECT 751.250 821.000 751.570 821.060 ;
        RECT 751.055 820.860 751.570 821.000 ;
        RECT 751.250 820.800 751.570 820.860 ;
        RECT 751.250 786.660 751.570 786.720 ;
        RECT 751.055 786.520 751.570 786.660 ;
        RECT 751.250 786.460 751.570 786.520 ;
        RECT 750.790 738.380 751.110 738.440 ;
        RECT 751.710 738.380 752.030 738.440 ;
        RECT 750.790 738.240 752.030 738.380 ;
        RECT 750.790 738.180 751.110 738.240 ;
        RECT 751.710 738.180 752.030 738.240 ;
        RECT 751.250 724.440 751.570 724.500 ;
        RECT 751.055 724.300 751.570 724.440 ;
        RECT 751.250 724.240 751.570 724.300 ;
        RECT 751.250 689.760 751.570 689.820 ;
        RECT 751.055 689.620 751.570 689.760 ;
        RECT 751.250 689.560 751.570 689.620 ;
        RECT 750.790 641.820 751.110 641.880 ;
        RECT 751.710 641.820 752.030 641.880 ;
        RECT 750.790 641.680 752.030 641.820 ;
        RECT 750.790 641.620 751.110 641.680 ;
        RECT 751.710 641.620 752.030 641.680 ;
        RECT 751.250 627.880 751.570 627.940 ;
        RECT 751.055 627.740 751.570 627.880 ;
        RECT 751.250 627.680 751.570 627.740 ;
        RECT 751.250 593.200 751.570 593.260 ;
        RECT 751.055 593.060 751.570 593.200 ;
        RECT 751.250 593.000 751.570 593.060 ;
        RECT 750.790 545.260 751.110 545.320 ;
        RECT 751.710 545.260 752.030 545.320 ;
        RECT 750.790 545.120 752.030 545.260 ;
        RECT 750.790 545.060 751.110 545.120 ;
        RECT 751.710 545.060 752.030 545.120 ;
        RECT 751.250 531.320 751.570 531.380 ;
        RECT 751.055 531.180 751.570 531.320 ;
        RECT 751.250 531.120 751.570 531.180 ;
        RECT 751.250 496.640 751.570 496.700 ;
        RECT 751.055 496.500 751.570 496.640 ;
        RECT 751.250 496.440 751.570 496.500 ;
        RECT 750.790 448.700 751.110 448.760 ;
        RECT 751.710 448.700 752.030 448.760 ;
        RECT 750.790 448.560 752.030 448.700 ;
        RECT 750.790 448.500 751.110 448.560 ;
        RECT 751.710 448.500 752.030 448.560 ;
        RECT 751.250 434.760 751.570 434.820 ;
        RECT 751.055 434.620 751.570 434.760 ;
        RECT 751.250 434.560 751.570 434.620 ;
        RECT 751.265 386.480 751.555 386.525 ;
        RECT 751.710 386.480 752.030 386.540 ;
        RECT 751.265 386.340 752.030 386.480 ;
        RECT 751.265 386.295 751.555 386.340 ;
        RECT 751.710 386.280 752.030 386.340 ;
        RECT 750.790 352.140 751.110 352.200 ;
        RECT 750.790 352.000 751.480 352.140 ;
        RECT 750.790 351.940 751.110 352.000 ;
        RECT 751.340 351.860 751.480 352.000 ;
        RECT 751.250 351.600 751.570 351.860 ;
        RECT 751.265 289.580 751.555 289.625 ;
        RECT 751.710 289.580 752.030 289.640 ;
        RECT 751.265 289.440 752.030 289.580 ;
        RECT 751.265 289.395 751.555 289.440 ;
        RECT 751.710 289.380 752.030 289.440 ;
        RECT 751.250 241.640 751.570 241.700 ;
        RECT 751.055 241.500 751.570 241.640 ;
        RECT 751.250 241.440 751.570 241.500 ;
        RECT 751.265 193.020 751.555 193.065 ;
        RECT 751.710 193.020 752.030 193.080 ;
        RECT 751.265 192.880 752.030 193.020 ;
        RECT 751.265 192.835 751.555 192.880 ;
        RECT 751.710 192.820 752.030 192.880 ;
        RECT 751.250 145.080 751.570 145.140 ;
        RECT 751.055 144.940 751.570 145.080 ;
        RECT 751.250 144.880 751.570 144.940 ;
        RECT 750.790 27.100 751.110 27.160 ;
        RECT 1185.950 27.100 1186.270 27.160 ;
        RECT 750.790 26.960 1186.270 27.100 ;
        RECT 750.790 26.900 751.110 26.960 ;
        RECT 1185.950 26.900 1186.270 26.960 ;
      LAYER via ;
        RECT 747.600 1587.160 747.860 1587.420 ;
        RECT 750.820 1587.160 751.080 1587.420 ;
        RECT 750.820 1414.440 751.080 1414.700 ;
        RECT 751.740 1414.440 752.000 1414.700 ;
        RECT 750.820 1317.880 751.080 1318.140 ;
        RECT 751.740 1317.880 752.000 1318.140 ;
        RECT 750.820 1221.320 751.080 1221.580 ;
        RECT 751.740 1221.320 752.000 1221.580 ;
        RECT 750.820 1124.760 751.080 1125.020 ;
        RECT 751.740 1124.760 752.000 1125.020 ;
        RECT 750.820 1028.200 751.080 1028.460 ;
        RECT 751.740 1028.200 752.000 1028.460 ;
        RECT 750.820 931.640 751.080 931.900 ;
        RECT 751.740 931.640 752.000 931.900 ;
        RECT 750.360 869.420 750.620 869.680 ;
        RECT 751.740 869.420 752.000 869.680 ;
        RECT 750.820 835.080 751.080 835.340 ;
        RECT 751.740 835.080 752.000 835.340 ;
        RECT 751.280 820.800 751.540 821.060 ;
        RECT 751.280 786.460 751.540 786.720 ;
        RECT 750.820 738.180 751.080 738.440 ;
        RECT 751.740 738.180 752.000 738.440 ;
        RECT 751.280 724.240 751.540 724.500 ;
        RECT 751.280 689.560 751.540 689.820 ;
        RECT 750.820 641.620 751.080 641.880 ;
        RECT 751.740 641.620 752.000 641.880 ;
        RECT 751.280 627.680 751.540 627.940 ;
        RECT 751.280 593.000 751.540 593.260 ;
        RECT 750.820 545.060 751.080 545.320 ;
        RECT 751.740 545.060 752.000 545.320 ;
        RECT 751.280 531.120 751.540 531.380 ;
        RECT 751.280 496.440 751.540 496.700 ;
        RECT 750.820 448.500 751.080 448.760 ;
        RECT 751.740 448.500 752.000 448.760 ;
        RECT 751.280 434.560 751.540 434.820 ;
        RECT 751.740 386.280 752.000 386.540 ;
        RECT 750.820 351.940 751.080 352.200 ;
        RECT 751.280 351.600 751.540 351.860 ;
        RECT 751.740 289.380 752.000 289.640 ;
        RECT 751.280 241.440 751.540 241.700 ;
        RECT 751.740 192.820 752.000 193.080 ;
        RECT 751.280 144.880 751.540 145.140 ;
        RECT 750.820 26.900 751.080 27.160 ;
        RECT 1185.980 26.900 1186.240 27.160 ;
      LAYER met2 ;
        RECT 747.600 1600.000 747.880 1604.000 ;
        RECT 747.660 1587.450 747.800 1600.000 ;
        RECT 747.600 1587.130 747.860 1587.450 ;
        RECT 750.820 1587.130 751.080 1587.450 ;
        RECT 750.880 1558.970 751.020 1587.130 ;
        RECT 750.880 1558.830 751.480 1558.970 ;
        RECT 751.340 1511.370 751.480 1558.830 ;
        RECT 751.340 1511.230 751.940 1511.370 ;
        RECT 751.800 1414.730 751.940 1511.230 ;
        RECT 750.820 1414.410 751.080 1414.730 ;
        RECT 751.740 1414.410 752.000 1414.730 ;
        RECT 750.880 1414.130 751.020 1414.410 ;
        RECT 750.880 1413.990 751.480 1414.130 ;
        RECT 751.340 1366.530 751.480 1413.990 ;
        RECT 751.340 1366.390 751.940 1366.530 ;
        RECT 751.800 1318.170 751.940 1366.390 ;
        RECT 750.820 1317.850 751.080 1318.170 ;
        RECT 751.740 1317.850 752.000 1318.170 ;
        RECT 750.880 1317.570 751.020 1317.850 ;
        RECT 750.880 1317.430 751.480 1317.570 ;
        RECT 751.340 1269.970 751.480 1317.430 ;
        RECT 751.340 1269.830 751.940 1269.970 ;
        RECT 751.800 1221.610 751.940 1269.830 ;
        RECT 750.820 1221.290 751.080 1221.610 ;
        RECT 751.740 1221.290 752.000 1221.610 ;
        RECT 750.880 1221.010 751.020 1221.290 ;
        RECT 750.880 1220.870 751.480 1221.010 ;
        RECT 751.340 1173.410 751.480 1220.870 ;
        RECT 751.340 1173.270 751.940 1173.410 ;
        RECT 751.800 1125.050 751.940 1173.270 ;
        RECT 750.820 1124.730 751.080 1125.050 ;
        RECT 751.740 1124.730 752.000 1125.050 ;
        RECT 750.880 1124.450 751.020 1124.730 ;
        RECT 750.880 1124.310 751.480 1124.450 ;
        RECT 751.340 1076.850 751.480 1124.310 ;
        RECT 751.340 1076.710 751.940 1076.850 ;
        RECT 751.800 1028.490 751.940 1076.710 ;
        RECT 750.820 1028.170 751.080 1028.490 ;
        RECT 751.740 1028.170 752.000 1028.490 ;
        RECT 750.880 1027.890 751.020 1028.170 ;
        RECT 750.880 1027.750 751.480 1027.890 ;
        RECT 751.340 980.290 751.480 1027.750 ;
        RECT 751.340 980.150 751.940 980.290 ;
        RECT 751.800 931.930 751.940 980.150 ;
        RECT 750.820 931.610 751.080 931.930 ;
        RECT 751.740 931.610 752.000 931.930 ;
        RECT 750.880 931.330 751.020 931.610 ;
        RECT 750.880 931.190 751.480 931.330 ;
        RECT 751.340 917.845 751.480 931.190 ;
        RECT 750.350 917.475 750.630 917.845 ;
        RECT 751.270 917.475 751.550 917.845 ;
        RECT 750.420 869.710 750.560 917.475 ;
        RECT 750.360 869.390 750.620 869.710 ;
        RECT 751.740 869.390 752.000 869.710 ;
        RECT 751.800 835.370 751.940 869.390 ;
        RECT 750.820 835.050 751.080 835.370 ;
        RECT 751.740 835.050 752.000 835.370 ;
        RECT 750.880 834.770 751.020 835.050 ;
        RECT 750.880 834.630 751.480 834.770 ;
        RECT 751.340 821.090 751.480 834.630 ;
        RECT 751.280 820.770 751.540 821.090 ;
        RECT 751.280 786.430 751.540 786.750 ;
        RECT 751.340 772.890 751.480 786.430 ;
        RECT 751.340 772.750 751.940 772.890 ;
        RECT 751.800 738.470 751.940 772.750 ;
        RECT 750.820 738.210 751.080 738.470 ;
        RECT 750.820 738.150 751.480 738.210 ;
        RECT 751.740 738.150 752.000 738.470 ;
        RECT 750.880 738.070 751.480 738.150 ;
        RECT 751.340 724.530 751.480 738.070 ;
        RECT 751.280 724.210 751.540 724.530 ;
        RECT 751.280 689.530 751.540 689.850 ;
        RECT 751.340 676.330 751.480 689.530 ;
        RECT 751.340 676.190 751.940 676.330 ;
        RECT 751.800 641.910 751.940 676.190 ;
        RECT 750.820 641.650 751.080 641.910 ;
        RECT 750.820 641.590 751.480 641.650 ;
        RECT 751.740 641.590 752.000 641.910 ;
        RECT 750.880 641.510 751.480 641.590 ;
        RECT 751.340 627.970 751.480 641.510 ;
        RECT 751.280 627.650 751.540 627.970 ;
        RECT 751.280 592.970 751.540 593.290 ;
        RECT 751.340 579.770 751.480 592.970 ;
        RECT 751.340 579.630 751.940 579.770 ;
        RECT 751.800 545.350 751.940 579.630 ;
        RECT 750.820 545.090 751.080 545.350 ;
        RECT 750.820 545.030 751.480 545.090 ;
        RECT 751.740 545.030 752.000 545.350 ;
        RECT 750.880 544.950 751.480 545.030 ;
        RECT 751.340 531.410 751.480 544.950 ;
        RECT 751.280 531.090 751.540 531.410 ;
        RECT 751.280 496.410 751.540 496.730 ;
        RECT 751.340 483.210 751.480 496.410 ;
        RECT 751.340 483.070 751.940 483.210 ;
        RECT 751.800 448.790 751.940 483.070 ;
        RECT 750.820 448.530 751.080 448.790 ;
        RECT 750.820 448.470 751.480 448.530 ;
        RECT 751.740 448.470 752.000 448.790 ;
        RECT 750.880 448.390 751.480 448.470 ;
        RECT 751.340 434.850 751.480 448.390 ;
        RECT 751.280 434.530 751.540 434.850 ;
        RECT 751.740 386.250 752.000 386.570 ;
        RECT 751.800 386.085 751.940 386.250 ;
        RECT 750.810 385.715 751.090 386.085 ;
        RECT 751.730 385.715 752.010 386.085 ;
        RECT 750.880 352.230 751.020 385.715 ;
        RECT 750.820 351.910 751.080 352.230 ;
        RECT 751.280 351.570 751.540 351.890 ;
        RECT 751.340 303.690 751.480 351.570 ;
        RECT 751.340 303.550 751.940 303.690 ;
        RECT 751.800 289.670 751.940 303.550 ;
        RECT 751.740 289.350 752.000 289.670 ;
        RECT 751.280 241.410 751.540 241.730 ;
        RECT 751.340 207.130 751.480 241.410 ;
        RECT 751.340 206.990 751.940 207.130 ;
        RECT 751.800 193.110 751.940 206.990 ;
        RECT 751.740 192.790 752.000 193.110 ;
        RECT 751.280 144.850 751.540 145.170 ;
        RECT 751.340 110.570 751.480 144.850 ;
        RECT 751.340 110.430 751.940 110.570 ;
        RECT 751.800 62.290 751.940 110.430 ;
        RECT 750.880 62.150 751.940 62.290 ;
        RECT 750.880 27.190 751.020 62.150 ;
        RECT 750.820 26.870 751.080 27.190 ;
        RECT 1185.980 26.870 1186.240 27.190 ;
        RECT 1186.040 2.400 1186.180 26.870 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
      LAYER via2 ;
        RECT 750.350 917.520 750.630 917.800 ;
        RECT 751.270 917.520 751.550 917.800 ;
        RECT 750.810 385.760 751.090 386.040 ;
        RECT 751.730 385.760 752.010 386.040 ;
      LAYER met3 ;
        RECT 750.325 917.810 750.655 917.825 ;
        RECT 751.245 917.810 751.575 917.825 ;
        RECT 750.325 917.510 751.575 917.810 ;
        RECT 750.325 917.495 750.655 917.510 ;
        RECT 751.245 917.495 751.575 917.510 ;
        RECT 750.785 386.050 751.115 386.065 ;
        RECT 751.705 386.050 752.035 386.065 ;
        RECT 750.785 385.750 752.035 386.050 ;
        RECT 750.785 385.735 751.115 385.750 ;
        RECT 751.705 385.735 752.035 385.750 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 754.010 1587.360 754.330 1587.420 ;
        RECT 758.610 1587.360 758.930 1587.420 ;
        RECT 754.010 1587.220 758.930 1587.360 ;
        RECT 754.010 1587.160 754.330 1587.220 ;
        RECT 758.610 1587.160 758.930 1587.220 ;
        RECT 758.610 26.760 758.930 26.820 ;
        RECT 1203.890 26.760 1204.210 26.820 ;
        RECT 758.610 26.620 1204.210 26.760 ;
        RECT 758.610 26.560 758.930 26.620 ;
        RECT 1203.890 26.560 1204.210 26.620 ;
      LAYER via ;
        RECT 754.040 1587.160 754.300 1587.420 ;
        RECT 758.640 1587.160 758.900 1587.420 ;
        RECT 758.640 26.560 758.900 26.820 ;
        RECT 1203.920 26.560 1204.180 26.820 ;
      LAYER met2 ;
        RECT 754.040 1600.000 754.320 1604.000 ;
        RECT 754.100 1587.450 754.240 1600.000 ;
        RECT 754.040 1587.130 754.300 1587.450 ;
        RECT 758.640 1587.130 758.900 1587.450 ;
        RECT 758.700 26.850 758.840 1587.130 ;
        RECT 758.640 26.530 758.900 26.850 ;
        RECT 1203.920 26.530 1204.180 26.850 ;
        RECT 1203.980 2.400 1204.120 26.530 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 760.910 1587.360 761.230 1587.420 ;
        RECT 765.510 1587.360 765.830 1587.420 ;
        RECT 760.910 1587.220 765.830 1587.360 ;
        RECT 760.910 1587.160 761.230 1587.220 ;
        RECT 765.510 1587.160 765.830 1587.220 ;
        RECT 765.510 26.420 765.830 26.480 ;
        RECT 1221.830 26.420 1222.150 26.480 ;
        RECT 765.510 26.280 1222.150 26.420 ;
        RECT 765.510 26.220 765.830 26.280 ;
        RECT 1221.830 26.220 1222.150 26.280 ;
      LAYER via ;
        RECT 760.940 1587.160 761.200 1587.420 ;
        RECT 765.540 1587.160 765.800 1587.420 ;
        RECT 765.540 26.220 765.800 26.480 ;
        RECT 1221.860 26.220 1222.120 26.480 ;
      LAYER met2 ;
        RECT 760.940 1600.000 761.220 1604.000 ;
        RECT 761.000 1587.450 761.140 1600.000 ;
        RECT 760.940 1587.130 761.200 1587.450 ;
        RECT 765.540 1587.130 765.800 1587.450 ;
        RECT 765.600 26.510 765.740 1587.130 ;
        RECT 765.540 26.190 765.800 26.510 ;
        RECT 1221.860 26.190 1222.120 26.510 ;
        RECT 1221.920 2.400 1222.060 26.190 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 767.350 1587.360 767.670 1587.420 ;
        RECT 772.410 1587.360 772.730 1587.420 ;
        RECT 767.350 1587.220 772.730 1587.360 ;
        RECT 767.350 1587.160 767.670 1587.220 ;
        RECT 772.410 1587.160 772.730 1587.220 ;
        RECT 772.410 26.080 772.730 26.140 ;
        RECT 1239.770 26.080 1240.090 26.140 ;
        RECT 772.410 25.940 1240.090 26.080 ;
        RECT 772.410 25.880 772.730 25.940 ;
        RECT 1239.770 25.880 1240.090 25.940 ;
      LAYER via ;
        RECT 767.380 1587.160 767.640 1587.420 ;
        RECT 772.440 1587.160 772.700 1587.420 ;
        RECT 772.440 25.880 772.700 26.140 ;
        RECT 1239.800 25.880 1240.060 26.140 ;
      LAYER met2 ;
        RECT 767.380 1600.000 767.660 1604.000 ;
        RECT 767.440 1587.450 767.580 1600.000 ;
        RECT 767.380 1587.130 767.640 1587.450 ;
        RECT 772.440 1587.130 772.700 1587.450 ;
        RECT 772.500 26.170 772.640 1587.130 ;
        RECT 772.440 25.850 772.700 26.170 ;
        RECT 1239.800 25.850 1240.060 26.170 ;
        RECT 1239.860 2.400 1240.000 25.850 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 774.250 1587.360 774.570 1587.420 ;
        RECT 779.310 1587.360 779.630 1587.420 ;
        RECT 774.250 1587.220 779.630 1587.360 ;
        RECT 774.250 1587.160 774.570 1587.220 ;
        RECT 779.310 1587.160 779.630 1587.220 ;
        RECT 779.310 25.740 779.630 25.800 ;
        RECT 1257.250 25.740 1257.570 25.800 ;
        RECT 779.310 25.600 1257.570 25.740 ;
        RECT 779.310 25.540 779.630 25.600 ;
        RECT 1257.250 25.540 1257.570 25.600 ;
      LAYER via ;
        RECT 774.280 1587.160 774.540 1587.420 ;
        RECT 779.340 1587.160 779.600 1587.420 ;
        RECT 779.340 25.540 779.600 25.800 ;
        RECT 1257.280 25.540 1257.540 25.800 ;
      LAYER met2 ;
        RECT 774.280 1600.000 774.560 1604.000 ;
        RECT 774.340 1587.450 774.480 1600.000 ;
        RECT 774.280 1587.130 774.540 1587.450 ;
        RECT 779.340 1587.130 779.600 1587.450 ;
        RECT 779.400 25.830 779.540 1587.130 ;
        RECT 779.340 25.510 779.600 25.830 ;
        RECT 1257.280 25.510 1257.540 25.830 ;
        RECT 1257.340 2.400 1257.480 25.510 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 781.150 1587.700 781.470 1587.760 ;
        RECT 786.210 1587.700 786.530 1587.760 ;
        RECT 781.150 1587.560 786.530 1587.700 ;
        RECT 781.150 1587.500 781.470 1587.560 ;
        RECT 786.210 1587.500 786.530 1587.560 ;
        RECT 786.210 25.400 786.530 25.460 ;
        RECT 1275.190 25.400 1275.510 25.460 ;
        RECT 786.210 25.260 1275.510 25.400 ;
        RECT 786.210 25.200 786.530 25.260 ;
        RECT 1275.190 25.200 1275.510 25.260 ;
      LAYER via ;
        RECT 781.180 1587.500 781.440 1587.760 ;
        RECT 786.240 1587.500 786.500 1587.760 ;
        RECT 786.240 25.200 786.500 25.460 ;
        RECT 1275.220 25.200 1275.480 25.460 ;
      LAYER met2 ;
        RECT 781.180 1600.000 781.460 1604.000 ;
        RECT 781.240 1587.790 781.380 1600.000 ;
        RECT 781.180 1587.470 781.440 1587.790 ;
        RECT 786.240 1587.470 786.500 1587.790 ;
        RECT 786.300 25.490 786.440 1587.470 ;
        RECT 786.240 25.170 786.500 25.490 ;
        RECT 1275.220 25.170 1275.480 25.490 ;
        RECT 1275.280 2.400 1275.420 25.170 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 787.590 1588.040 787.910 1588.100 ;
        RECT 793.110 1588.040 793.430 1588.100 ;
        RECT 787.590 1587.900 793.430 1588.040 ;
        RECT 787.590 1587.840 787.910 1587.900 ;
        RECT 793.110 1587.840 793.430 1587.900 ;
        RECT 793.110 25.060 793.430 25.120 ;
        RECT 1293.130 25.060 1293.450 25.120 ;
        RECT 793.110 24.920 1293.450 25.060 ;
        RECT 793.110 24.860 793.430 24.920 ;
        RECT 1293.130 24.860 1293.450 24.920 ;
      LAYER via ;
        RECT 787.620 1587.840 787.880 1588.100 ;
        RECT 793.140 1587.840 793.400 1588.100 ;
        RECT 793.140 24.860 793.400 25.120 ;
        RECT 1293.160 24.860 1293.420 25.120 ;
      LAYER met2 ;
        RECT 787.620 1600.000 787.900 1604.000 ;
        RECT 787.680 1588.130 787.820 1600.000 ;
        RECT 787.620 1587.810 787.880 1588.130 ;
        RECT 793.140 1587.810 793.400 1588.130 ;
        RECT 793.200 25.150 793.340 1587.810 ;
        RECT 793.140 24.830 793.400 25.150 ;
        RECT 1293.160 24.830 1293.420 25.150 ;
        RECT 1293.220 2.400 1293.360 24.830 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 794.490 1588.040 794.810 1588.100 ;
        RECT 800.010 1588.040 800.330 1588.100 ;
        RECT 794.490 1587.900 800.330 1588.040 ;
        RECT 794.490 1587.840 794.810 1587.900 ;
        RECT 800.010 1587.840 800.330 1587.900 ;
        RECT 800.010 24.720 800.330 24.780 ;
        RECT 1311.070 24.720 1311.390 24.780 ;
        RECT 800.010 24.580 1311.390 24.720 ;
        RECT 800.010 24.520 800.330 24.580 ;
        RECT 1311.070 24.520 1311.390 24.580 ;
      LAYER via ;
        RECT 794.520 1587.840 794.780 1588.100 ;
        RECT 800.040 1587.840 800.300 1588.100 ;
        RECT 800.040 24.520 800.300 24.780 ;
        RECT 1311.100 24.520 1311.360 24.780 ;
      LAYER met2 ;
        RECT 794.520 1600.000 794.800 1604.000 ;
        RECT 794.580 1588.130 794.720 1600.000 ;
        RECT 794.520 1587.810 794.780 1588.130 ;
        RECT 800.040 1587.810 800.300 1588.130 ;
        RECT 800.100 24.810 800.240 1587.810 ;
        RECT 800.040 24.490 800.300 24.810 ;
        RECT 1311.100 24.490 1311.360 24.810 ;
        RECT 1311.160 2.400 1311.300 24.490 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 801.390 1587.700 801.710 1587.760 ;
        RECT 806.910 1587.700 807.230 1587.760 ;
        RECT 801.390 1587.560 807.230 1587.700 ;
        RECT 801.390 1587.500 801.710 1587.560 ;
        RECT 806.910 1587.500 807.230 1587.560 ;
        RECT 806.910 24.380 807.230 24.440 ;
        RECT 1329.010 24.380 1329.330 24.440 ;
        RECT 806.910 24.240 1329.330 24.380 ;
        RECT 806.910 24.180 807.230 24.240 ;
        RECT 1329.010 24.180 1329.330 24.240 ;
      LAYER via ;
        RECT 801.420 1587.500 801.680 1587.760 ;
        RECT 806.940 1587.500 807.200 1587.760 ;
        RECT 806.940 24.180 807.200 24.440 ;
        RECT 1329.040 24.180 1329.300 24.440 ;
      LAYER met2 ;
        RECT 801.420 1600.000 801.700 1604.000 ;
        RECT 801.480 1587.790 801.620 1600.000 ;
        RECT 801.420 1587.470 801.680 1587.790 ;
        RECT 806.940 1587.470 807.200 1587.790 ;
        RECT 807.000 24.470 807.140 1587.470 ;
        RECT 806.940 24.150 807.200 24.470 ;
        RECT 1329.040 24.150 1329.300 24.470 ;
        RECT 1329.100 2.400 1329.240 24.150 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 558.970 1592.800 559.290 1592.860 ;
        RECT 665.690 1592.800 666.010 1592.860 ;
        RECT 558.970 1592.660 666.010 1592.800 ;
        RECT 558.970 1592.600 559.290 1592.660 ;
        RECT 665.690 1592.600 666.010 1592.660 ;
        RECT 665.690 18.260 666.010 18.320 ;
        RECT 686.390 18.260 686.710 18.320 ;
        RECT 665.690 18.120 686.710 18.260 ;
        RECT 665.690 18.060 666.010 18.120 ;
        RECT 686.390 18.060 686.710 18.120 ;
      LAYER via ;
        RECT 559.000 1592.600 559.260 1592.860 ;
        RECT 665.720 1592.600 665.980 1592.860 ;
        RECT 665.720 18.060 665.980 18.320 ;
        RECT 686.420 18.060 686.680 18.320 ;
      LAYER met2 ;
        RECT 559.000 1600.000 559.280 1604.000 ;
        RECT 559.060 1592.890 559.200 1600.000 ;
        RECT 559.000 1592.570 559.260 1592.890 ;
        RECT 665.720 1592.570 665.980 1592.890 ;
        RECT 665.780 18.350 665.920 1592.570 ;
        RECT 665.720 18.030 665.980 18.350 ;
        RECT 686.420 18.030 686.680 18.350 ;
        RECT 686.480 2.400 686.620 18.030 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 807.830 1587.360 808.150 1587.420 ;
        RECT 813.810 1587.360 814.130 1587.420 ;
        RECT 807.830 1587.220 814.130 1587.360 ;
        RECT 807.830 1587.160 808.150 1587.220 ;
        RECT 813.810 1587.160 814.130 1587.220 ;
        RECT 813.810 24.040 814.130 24.100 ;
        RECT 1346.490 24.040 1346.810 24.100 ;
        RECT 813.810 23.900 1346.810 24.040 ;
        RECT 813.810 23.840 814.130 23.900 ;
        RECT 1346.490 23.840 1346.810 23.900 ;
      LAYER via ;
        RECT 807.860 1587.160 808.120 1587.420 ;
        RECT 813.840 1587.160 814.100 1587.420 ;
        RECT 813.840 23.840 814.100 24.100 ;
        RECT 1346.520 23.840 1346.780 24.100 ;
      LAYER met2 ;
        RECT 807.860 1600.000 808.140 1604.000 ;
        RECT 807.920 1587.450 808.060 1600.000 ;
        RECT 807.860 1587.130 808.120 1587.450 ;
        RECT 813.840 1587.130 814.100 1587.450 ;
        RECT 813.900 24.130 814.040 1587.130 ;
        RECT 813.840 23.810 814.100 24.130 ;
        RECT 1346.520 23.810 1346.780 24.130 ;
        RECT 1346.580 2.400 1346.720 23.810 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 814.730 1587.360 815.050 1587.420 ;
        RECT 820.710 1587.360 821.030 1587.420 ;
        RECT 814.730 1587.220 821.030 1587.360 ;
        RECT 814.730 1587.160 815.050 1587.220 ;
        RECT 820.710 1587.160 821.030 1587.220 ;
      LAYER via ;
        RECT 814.760 1587.160 815.020 1587.420 ;
        RECT 820.740 1587.160 821.000 1587.420 ;
      LAYER met2 ;
        RECT 814.760 1600.000 815.040 1604.000 ;
        RECT 814.820 1587.450 814.960 1600.000 ;
        RECT 814.760 1587.130 815.020 1587.450 ;
        RECT 820.740 1587.130 821.000 1587.450 ;
        RECT 820.800 25.685 820.940 1587.130 ;
        RECT 820.730 25.315 821.010 25.685 ;
        RECT 1364.450 25.315 1364.730 25.685 ;
        RECT 1364.520 2.400 1364.660 25.315 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
      LAYER via2 ;
        RECT 820.730 25.360 821.010 25.640 ;
        RECT 1364.450 25.360 1364.730 25.640 ;
      LAYER met3 ;
        RECT 820.705 25.650 821.035 25.665 ;
        RECT 1364.425 25.650 1364.755 25.665 ;
        RECT 820.705 25.350 1364.755 25.650 ;
        RECT 820.705 25.335 821.035 25.350 ;
        RECT 1364.425 25.335 1364.755 25.350 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 821.630 1587.700 821.950 1587.760 ;
        RECT 827.610 1587.700 827.930 1587.760 ;
        RECT 821.630 1587.560 827.930 1587.700 ;
        RECT 821.630 1587.500 821.950 1587.560 ;
        RECT 827.610 1587.500 827.930 1587.560 ;
      LAYER via ;
        RECT 821.660 1587.500 821.920 1587.760 ;
        RECT 827.640 1587.500 827.900 1587.760 ;
      LAYER met2 ;
        RECT 821.660 1600.000 821.940 1604.000 ;
        RECT 821.720 1587.790 821.860 1600.000 ;
        RECT 821.660 1587.470 821.920 1587.790 ;
        RECT 827.640 1587.470 827.900 1587.790 ;
        RECT 827.700 25.005 827.840 1587.470 ;
        RECT 827.630 24.635 827.910 25.005 ;
        RECT 1382.390 24.635 1382.670 25.005 ;
        RECT 1382.460 2.400 1382.600 24.635 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
      LAYER via2 ;
        RECT 827.630 24.680 827.910 24.960 ;
        RECT 1382.390 24.680 1382.670 24.960 ;
      LAYER met3 ;
        RECT 827.605 24.970 827.935 24.985 ;
        RECT 1382.365 24.970 1382.695 24.985 ;
        RECT 827.605 24.670 1382.695 24.970 ;
        RECT 827.605 24.655 827.935 24.670 ;
        RECT 1382.365 24.655 1382.695 24.670 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 828.070 1587.360 828.390 1587.420 ;
        RECT 834.510 1587.360 834.830 1587.420 ;
        RECT 828.070 1587.220 834.830 1587.360 ;
        RECT 828.070 1587.160 828.390 1587.220 ;
        RECT 834.510 1587.160 834.830 1587.220 ;
        RECT 1367.190 11.800 1367.510 11.860 ;
        RECT 1400.310 11.800 1400.630 11.860 ;
        RECT 1367.190 11.660 1400.630 11.800 ;
        RECT 1367.190 11.600 1367.510 11.660 ;
        RECT 1400.310 11.600 1400.630 11.660 ;
      LAYER via ;
        RECT 828.100 1587.160 828.360 1587.420 ;
        RECT 834.540 1587.160 834.800 1587.420 ;
        RECT 1367.220 11.600 1367.480 11.860 ;
        RECT 1400.340 11.600 1400.600 11.860 ;
      LAYER met2 ;
        RECT 828.100 1600.000 828.380 1604.000 ;
        RECT 828.160 1587.450 828.300 1600.000 ;
        RECT 828.100 1587.130 828.360 1587.450 ;
        RECT 834.540 1587.130 834.800 1587.450 ;
        RECT 834.600 24.325 834.740 1587.130 ;
        RECT 834.530 23.955 834.810 24.325 ;
        RECT 861.670 24.210 861.950 24.325 ;
        RECT 862.590 24.210 862.870 24.325 ;
        RECT 861.670 24.070 862.870 24.210 ;
        RECT 861.670 23.955 861.950 24.070 ;
        RECT 862.590 23.955 862.870 24.070 ;
        RECT 903.530 23.955 903.810 24.325 ;
        RECT 910.430 23.955 910.710 24.325 ;
        RECT 1027.270 23.955 1027.550 24.325 ;
        RECT 1062.230 23.955 1062.510 24.325 ;
        RECT 903.600 22.965 903.740 23.955 ;
        RECT 910.500 22.965 910.640 23.955 ;
        RECT 1027.340 22.965 1027.480 23.955 ;
        RECT 1062.300 22.965 1062.440 23.955 ;
        RECT 903.530 22.595 903.810 22.965 ;
        RECT 910.430 22.595 910.710 22.965 ;
        RECT 1027.270 22.595 1027.550 22.965 ;
        RECT 1062.230 22.595 1062.510 22.965 ;
        RECT 1158.830 22.595 1159.110 22.965 ;
        RECT 1172.630 22.850 1172.910 22.965 ;
        RECT 1172.630 22.710 1173.760 22.850 ;
        RECT 1172.630 22.595 1172.910 22.710 ;
        RECT 1158.900 20.925 1159.040 22.595 ;
        RECT 1173.620 22.285 1173.760 22.710 ;
        RECT 1296.830 22.595 1297.110 22.965 ;
        RECT 1173.550 21.915 1173.830 22.285 ;
        RECT 1220.470 22.170 1220.750 22.285 ;
        RECT 1221.390 22.170 1221.670 22.285 ;
        RECT 1220.470 22.030 1221.670 22.170 ;
        RECT 1220.470 21.915 1220.750 22.030 ;
        RECT 1221.390 21.915 1221.670 22.030 ;
        RECT 1296.900 21.605 1297.040 22.595 ;
        RECT 1296.830 21.235 1297.110 21.605 ;
        RECT 1367.210 21.235 1367.490 21.605 ;
        RECT 1158.830 20.555 1159.110 20.925 ;
        RECT 1367.280 11.890 1367.420 21.235 ;
        RECT 1367.220 11.570 1367.480 11.890 ;
        RECT 1400.340 11.570 1400.600 11.890 ;
        RECT 1400.400 2.400 1400.540 11.570 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
      LAYER via2 ;
        RECT 834.530 24.000 834.810 24.280 ;
        RECT 861.670 24.000 861.950 24.280 ;
        RECT 862.590 24.000 862.870 24.280 ;
        RECT 903.530 24.000 903.810 24.280 ;
        RECT 910.430 24.000 910.710 24.280 ;
        RECT 1027.270 24.000 1027.550 24.280 ;
        RECT 1062.230 24.000 1062.510 24.280 ;
        RECT 903.530 22.640 903.810 22.920 ;
        RECT 910.430 22.640 910.710 22.920 ;
        RECT 1027.270 22.640 1027.550 22.920 ;
        RECT 1062.230 22.640 1062.510 22.920 ;
        RECT 1158.830 22.640 1159.110 22.920 ;
        RECT 1172.630 22.640 1172.910 22.920 ;
        RECT 1296.830 22.640 1297.110 22.920 ;
        RECT 1173.550 21.960 1173.830 22.240 ;
        RECT 1220.470 21.960 1220.750 22.240 ;
        RECT 1221.390 21.960 1221.670 22.240 ;
        RECT 1296.830 21.280 1297.110 21.560 ;
        RECT 1367.210 21.280 1367.490 21.560 ;
        RECT 1158.830 20.600 1159.110 20.880 ;
      LAYER met3 ;
        RECT 834.505 24.120 834.835 24.305 ;
        RECT 861.645 24.290 861.975 24.305 ;
        RECT 835.670 24.120 861.975 24.290 ;
        RECT 834.505 23.990 861.975 24.120 ;
        RECT 834.505 23.975 835.970 23.990 ;
        RECT 861.645 23.975 861.975 23.990 ;
        RECT 862.565 24.290 862.895 24.305 ;
        RECT 903.505 24.290 903.835 24.305 ;
        RECT 862.565 23.990 903.835 24.290 ;
        RECT 862.565 23.975 862.895 23.990 ;
        RECT 903.505 23.975 903.835 23.990 ;
        RECT 910.405 24.290 910.735 24.305 ;
        RECT 1027.245 24.290 1027.575 24.305 ;
        RECT 1062.205 24.290 1062.535 24.305 ;
        RECT 910.405 23.990 930.960 24.290 ;
        RECT 910.405 23.975 910.735 23.990 ;
        RECT 834.520 23.820 835.970 23.975 ;
        RECT 930.660 23.610 930.960 23.990 ;
        RECT 1027.245 23.990 1062.535 24.290 ;
        RECT 1027.245 23.975 1027.575 23.990 ;
        RECT 1062.205 23.975 1062.535 23.990 ;
        RECT 930.660 23.310 965.690 23.610 ;
        RECT 903.505 22.930 903.835 22.945 ;
        RECT 910.405 22.930 910.735 22.945 ;
        RECT 903.505 22.630 910.735 22.930 ;
        RECT 903.505 22.615 903.835 22.630 ;
        RECT 910.405 22.615 910.735 22.630 ;
        RECT 965.390 22.250 965.690 23.310 ;
        RECT 1027.245 22.930 1027.575 22.945 ;
        RECT 1014.150 22.630 1027.575 22.930 ;
        RECT 1014.150 22.250 1014.450 22.630 ;
        RECT 1027.245 22.615 1027.575 22.630 ;
        RECT 1062.205 22.930 1062.535 22.945 ;
        RECT 1158.805 22.930 1159.135 22.945 ;
        RECT 1172.605 22.930 1172.935 22.945 ;
        RECT 1248.710 22.930 1249.090 22.940 ;
        RECT 1062.205 22.630 1076.090 22.930 ;
        RECT 1062.205 22.615 1062.535 22.630 ;
        RECT 965.390 21.950 966.610 22.250 ;
        RECT 966.310 21.570 966.610 21.950 ;
        RECT 980.110 21.950 1014.450 22.250 ;
        RECT 1075.790 22.080 1076.090 22.630 ;
        RECT 1158.805 22.630 1172.935 22.930 ;
        RECT 1158.805 22.615 1159.135 22.630 ;
        RECT 1172.605 22.615 1172.935 22.630 ;
        RECT 1231.270 22.630 1249.090 22.930 ;
        RECT 1110.710 22.250 1111.090 22.260 ;
        RECT 1076.710 22.080 1111.090 22.250 ;
        RECT 1075.790 21.950 1111.090 22.080 ;
        RECT 980.110 21.570 980.410 21.950 ;
        RECT 1075.790 21.780 1077.010 21.950 ;
        RECT 1110.710 21.940 1111.090 21.950 ;
        RECT 1173.525 22.250 1173.855 22.265 ;
        RECT 1220.445 22.250 1220.775 22.265 ;
        RECT 1173.525 21.950 1220.775 22.250 ;
        RECT 1173.525 21.935 1173.855 21.950 ;
        RECT 1220.445 21.935 1220.775 21.950 ;
        RECT 1221.365 22.250 1221.695 22.265 ;
        RECT 1231.270 22.250 1231.570 22.630 ;
        RECT 1248.710 22.620 1249.090 22.630 ;
        RECT 1296.805 22.930 1297.135 22.945 ;
        RECT 1345.310 22.930 1345.690 22.940 ;
        RECT 1296.805 22.630 1345.690 22.930 ;
        RECT 1296.805 22.615 1297.135 22.630 ;
        RECT 1345.310 22.620 1345.690 22.630 ;
        RECT 1221.365 21.950 1231.570 22.250 ;
        RECT 1221.365 21.935 1221.695 21.950 ;
        RECT 966.310 21.270 980.410 21.570 ;
        RECT 1248.710 21.570 1249.090 21.580 ;
        RECT 1296.805 21.570 1297.135 21.585 ;
        RECT 1248.710 21.270 1297.135 21.570 ;
        RECT 1248.710 21.260 1249.090 21.270 ;
        RECT 1296.805 21.255 1297.135 21.270 ;
        RECT 1345.310 21.570 1345.690 21.580 ;
        RECT 1367.185 21.570 1367.515 21.585 ;
        RECT 1345.310 21.270 1367.515 21.570 ;
        RECT 1345.310 21.260 1345.690 21.270 ;
        RECT 1367.185 21.255 1367.515 21.270 ;
        RECT 1110.710 20.890 1111.090 20.900 ;
        RECT 1158.805 20.890 1159.135 20.905 ;
        RECT 1110.710 20.590 1159.135 20.890 ;
        RECT 1110.710 20.580 1111.090 20.590 ;
        RECT 1158.805 20.575 1159.135 20.590 ;
      LAYER via3 ;
        RECT 1110.740 21.940 1111.060 22.260 ;
        RECT 1248.740 22.620 1249.060 22.940 ;
        RECT 1345.340 22.620 1345.660 22.940 ;
        RECT 1248.740 21.260 1249.060 21.580 ;
        RECT 1345.340 21.260 1345.660 21.580 ;
        RECT 1110.740 20.580 1111.060 20.900 ;
      LAYER met4 ;
        RECT 1248.735 22.615 1249.065 22.945 ;
        RECT 1345.335 22.615 1345.665 22.945 ;
        RECT 1110.735 21.935 1111.065 22.265 ;
        RECT 1110.750 20.905 1111.050 21.935 ;
        RECT 1248.750 21.585 1249.050 22.615 ;
        RECT 1345.350 21.585 1345.650 22.615 ;
        RECT 1248.735 21.255 1249.065 21.585 ;
        RECT 1345.335 21.255 1345.665 21.585 ;
        RECT 1110.735 20.575 1111.065 20.905 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 834.970 1590.760 835.290 1590.820 ;
        RECT 841.410 1590.760 841.730 1590.820 ;
        RECT 834.970 1590.620 841.730 1590.760 ;
        RECT 834.970 1590.560 835.290 1590.620 ;
        RECT 841.410 1590.560 841.730 1590.620 ;
      LAYER via ;
        RECT 835.000 1590.560 835.260 1590.820 ;
        RECT 841.440 1590.560 841.700 1590.820 ;
      LAYER met2 ;
        RECT 835.000 1600.000 835.280 1604.000 ;
        RECT 835.060 1590.850 835.200 1600.000 ;
        RECT 835.000 1590.530 835.260 1590.850 ;
        RECT 841.440 1590.530 841.700 1590.850 ;
        RECT 841.500 27.725 841.640 1590.530 ;
        RECT 841.430 27.355 841.710 27.725 ;
        RECT 1418.270 27.355 1418.550 27.725 ;
        RECT 1418.340 2.400 1418.480 27.355 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
      LAYER via2 ;
        RECT 841.430 27.400 841.710 27.680 ;
        RECT 1418.270 27.400 1418.550 27.680 ;
      LAYER met3 ;
        RECT 841.405 27.690 841.735 27.705 ;
        RECT 1418.245 27.690 1418.575 27.705 ;
        RECT 841.405 27.390 1418.575 27.690 ;
        RECT 841.405 27.375 841.735 27.390 ;
        RECT 1418.245 27.375 1418.575 27.390 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.490 69.260 840.810 69.320 ;
        RECT 1435.270 69.260 1435.590 69.320 ;
        RECT 840.490 69.120 1435.590 69.260 ;
        RECT 840.490 69.060 840.810 69.120 ;
        RECT 1435.270 69.060 1435.590 69.120 ;
      LAYER via ;
        RECT 840.520 69.060 840.780 69.320 ;
        RECT 1435.300 69.060 1435.560 69.320 ;
      LAYER met2 ;
        RECT 841.440 1600.450 841.720 1604.000 ;
        RECT 840.580 1600.310 841.720 1600.450 ;
        RECT 840.580 69.350 840.720 1600.310 ;
        RECT 841.440 1600.000 841.720 1600.310 ;
        RECT 840.520 69.030 840.780 69.350 ;
        RECT 1435.300 69.030 1435.560 69.350 ;
        RECT 1435.360 3.130 1435.500 69.030 ;
        RECT 1435.360 2.990 1435.960 3.130 ;
        RECT 1435.820 2.400 1435.960 2.990 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 848.340 1600.000 848.620 1604.000 ;
        RECT 848.400 27.045 848.540 1600.000 ;
        RECT 848.330 26.675 848.610 27.045 ;
        RECT 1453.690 26.675 1453.970 27.045 ;
        RECT 1453.760 2.400 1453.900 26.675 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
      LAYER via2 ;
        RECT 848.330 26.720 848.610 27.000 ;
        RECT 1453.690 26.720 1453.970 27.000 ;
      LAYER met3 ;
        RECT 848.305 27.010 848.635 27.025 ;
        RECT 1453.665 27.010 1453.995 27.025 ;
        RECT 848.305 26.710 1453.995 27.010 ;
        RECT 848.305 26.695 848.635 26.710 ;
        RECT 1453.665 26.695 1453.995 26.710 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 854.750 69.940 855.070 70.000 ;
        RECT 1469.770 69.940 1470.090 70.000 ;
        RECT 854.750 69.800 1470.090 69.940 ;
        RECT 854.750 69.740 855.070 69.800 ;
        RECT 1469.770 69.740 1470.090 69.800 ;
      LAYER via ;
        RECT 854.780 69.740 855.040 70.000 ;
        RECT 1469.800 69.740 1470.060 70.000 ;
      LAYER met2 ;
        RECT 855.240 1600.450 855.520 1604.000 ;
        RECT 854.840 1600.310 855.520 1600.450 ;
        RECT 854.840 70.030 854.980 1600.310 ;
        RECT 855.240 1600.000 855.520 1600.310 ;
        RECT 854.780 69.710 855.040 70.030 ;
        RECT 1469.800 69.710 1470.060 70.030 ;
        RECT 1469.860 3.130 1470.000 69.710 ;
        RECT 1469.860 2.990 1471.840 3.130 ;
        RECT 1471.700 2.400 1471.840 2.990 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 862.110 27.780 862.430 27.840 ;
        RECT 1489.550 27.780 1489.870 27.840 ;
        RECT 862.110 27.640 1489.870 27.780 ;
        RECT 862.110 27.580 862.430 27.640 ;
        RECT 1489.550 27.580 1489.870 27.640 ;
      LAYER via ;
        RECT 862.140 27.580 862.400 27.840 ;
        RECT 1489.580 27.580 1489.840 27.840 ;
      LAYER met2 ;
        RECT 861.680 1600.450 861.960 1604.000 ;
        RECT 861.680 1600.310 862.340 1600.450 ;
        RECT 861.680 1600.000 861.960 1600.310 ;
        RECT 862.200 27.870 862.340 1600.310 ;
        RECT 862.140 27.550 862.400 27.870 ;
        RECT 1489.580 27.550 1489.840 27.870 ;
        RECT 1489.640 2.400 1489.780 27.550 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.010 28.120 869.330 28.180 ;
        RECT 1507.030 28.120 1507.350 28.180 ;
        RECT 869.010 27.980 1507.350 28.120 ;
        RECT 869.010 27.920 869.330 27.980 ;
        RECT 1507.030 27.920 1507.350 27.980 ;
      LAYER via ;
        RECT 869.040 27.920 869.300 28.180 ;
        RECT 1507.060 27.920 1507.320 28.180 ;
      LAYER met2 ;
        RECT 868.580 1600.450 868.860 1604.000 ;
        RECT 868.580 1600.310 869.240 1600.450 ;
        RECT 868.580 1600.000 868.860 1600.310 ;
        RECT 869.100 28.210 869.240 1600.310 ;
        RECT 869.040 27.890 869.300 28.210 ;
        RECT 1507.060 27.890 1507.320 28.210 ;
        RECT 1507.120 2.400 1507.260 27.890 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 579.745 1588.225 579.915 1589.075 ;
        RECT 628.045 1587.885 628.215 1588.735 ;
        RECT 704.405 786.505 704.575 821.015 ;
        RECT 704.405 689.605 704.575 724.455 ;
        RECT 704.405 593.045 704.575 627.895 ;
        RECT 704.405 496.485 704.575 531.335 ;
        RECT 704.405 386.325 704.575 434.775 ;
        RECT 704.405 338.045 704.575 385.815 ;
        RECT 704.405 255.085 704.575 289.595 ;
        RECT 704.405 158.525 704.575 193.035 ;
        RECT 704.405 2.805 704.575 48.195 ;
      LAYER mcon ;
        RECT 579.745 1588.905 579.915 1589.075 ;
        RECT 628.045 1588.565 628.215 1588.735 ;
        RECT 704.405 820.845 704.575 821.015 ;
        RECT 704.405 724.285 704.575 724.455 ;
        RECT 704.405 627.725 704.575 627.895 ;
        RECT 704.405 531.165 704.575 531.335 ;
        RECT 704.405 434.605 704.575 434.775 ;
        RECT 704.405 385.645 704.575 385.815 ;
        RECT 704.405 289.425 704.575 289.595 ;
        RECT 704.405 192.865 704.575 193.035 ;
        RECT 704.405 48.025 704.575 48.195 ;
      LAYER met1 ;
        RECT 565.410 1589.060 565.730 1589.120 ;
        RECT 579.685 1589.060 579.975 1589.105 ;
        RECT 565.410 1588.920 579.975 1589.060 ;
        RECT 565.410 1588.860 565.730 1588.920 ;
        RECT 579.685 1588.875 579.975 1588.920 ;
        RECT 627.985 1588.720 628.275 1588.765 ;
        RECT 594.480 1588.580 628.275 1588.720 ;
        RECT 579.685 1588.380 579.975 1588.425 ;
        RECT 594.480 1588.380 594.620 1588.580 ;
        RECT 627.985 1588.535 628.275 1588.580 ;
        RECT 641.860 1588.580 692.600 1588.720 ;
        RECT 641.860 1588.380 642.000 1588.580 ;
        RECT 579.685 1588.240 594.620 1588.380 ;
        RECT 635.420 1588.240 642.000 1588.380 ;
        RECT 692.460 1588.380 692.600 1588.580 ;
        RECT 703.870 1588.380 704.190 1588.440 ;
        RECT 692.460 1588.240 704.190 1588.380 ;
        RECT 579.685 1588.195 579.975 1588.240 ;
        RECT 627.985 1588.040 628.275 1588.085 ;
        RECT 635.420 1588.040 635.560 1588.240 ;
        RECT 703.870 1588.180 704.190 1588.240 ;
        RECT 627.985 1587.900 635.560 1588.040 ;
        RECT 627.985 1587.855 628.275 1587.900 ;
        RECT 703.870 1559.140 704.190 1559.200 ;
        RECT 704.790 1559.140 705.110 1559.200 ;
        RECT 703.870 1559.000 705.110 1559.140 ;
        RECT 703.870 1558.940 704.190 1559.000 ;
        RECT 704.790 1558.940 705.110 1559.000 ;
        RECT 703.870 1483.660 704.190 1483.720 ;
        RECT 704.790 1483.660 705.110 1483.720 ;
        RECT 703.870 1483.520 705.110 1483.660 ;
        RECT 703.870 1483.460 704.190 1483.520 ;
        RECT 704.790 1483.460 705.110 1483.520 ;
        RECT 703.870 1318.080 704.190 1318.140 ;
        RECT 704.790 1318.080 705.110 1318.140 ;
        RECT 703.870 1317.940 705.110 1318.080 ;
        RECT 703.870 1317.880 704.190 1317.940 ;
        RECT 704.790 1317.880 705.110 1317.940 ;
        RECT 703.870 1221.520 704.190 1221.580 ;
        RECT 704.790 1221.520 705.110 1221.580 ;
        RECT 703.870 1221.380 705.110 1221.520 ;
        RECT 703.870 1221.320 704.190 1221.380 ;
        RECT 704.790 1221.320 705.110 1221.380 ;
        RECT 703.870 1124.960 704.190 1125.020 ;
        RECT 704.790 1124.960 705.110 1125.020 ;
        RECT 703.870 1124.820 705.110 1124.960 ;
        RECT 703.870 1124.760 704.190 1124.820 ;
        RECT 704.790 1124.760 705.110 1124.820 ;
        RECT 703.870 1028.400 704.190 1028.460 ;
        RECT 704.790 1028.400 705.110 1028.460 ;
        RECT 703.870 1028.260 705.110 1028.400 ;
        RECT 703.870 1028.200 704.190 1028.260 ;
        RECT 704.790 1028.200 705.110 1028.260 ;
        RECT 703.870 931.840 704.190 931.900 ;
        RECT 704.790 931.840 705.110 931.900 ;
        RECT 703.870 931.700 705.110 931.840 ;
        RECT 703.870 931.640 704.190 931.700 ;
        RECT 704.790 931.640 705.110 931.700 ;
        RECT 704.790 869.620 705.110 869.680 ;
        RECT 705.710 869.620 706.030 869.680 ;
        RECT 704.790 869.480 706.030 869.620 ;
        RECT 704.790 869.420 705.110 869.480 ;
        RECT 705.710 869.420 706.030 869.480 ;
        RECT 703.870 835.280 704.190 835.340 ;
        RECT 704.790 835.280 705.110 835.340 ;
        RECT 703.870 835.140 705.110 835.280 ;
        RECT 703.870 835.080 704.190 835.140 ;
        RECT 704.790 835.080 705.110 835.140 ;
        RECT 704.330 821.000 704.650 821.060 ;
        RECT 704.135 820.860 704.650 821.000 ;
        RECT 704.330 820.800 704.650 820.860 ;
        RECT 704.330 786.660 704.650 786.720 ;
        RECT 704.135 786.520 704.650 786.660 ;
        RECT 704.330 786.460 704.650 786.520 ;
        RECT 703.870 738.380 704.190 738.440 ;
        RECT 704.790 738.380 705.110 738.440 ;
        RECT 703.870 738.240 705.110 738.380 ;
        RECT 703.870 738.180 704.190 738.240 ;
        RECT 704.790 738.180 705.110 738.240 ;
        RECT 704.330 724.440 704.650 724.500 ;
        RECT 704.135 724.300 704.650 724.440 ;
        RECT 704.330 724.240 704.650 724.300 ;
        RECT 704.330 689.760 704.650 689.820 ;
        RECT 704.135 689.620 704.650 689.760 ;
        RECT 704.330 689.560 704.650 689.620 ;
        RECT 703.870 641.820 704.190 641.880 ;
        RECT 704.790 641.820 705.110 641.880 ;
        RECT 703.870 641.680 705.110 641.820 ;
        RECT 703.870 641.620 704.190 641.680 ;
        RECT 704.790 641.620 705.110 641.680 ;
        RECT 704.330 627.880 704.650 627.940 ;
        RECT 704.135 627.740 704.650 627.880 ;
        RECT 704.330 627.680 704.650 627.740 ;
        RECT 704.330 593.200 704.650 593.260 ;
        RECT 704.135 593.060 704.650 593.200 ;
        RECT 704.330 593.000 704.650 593.060 ;
        RECT 703.870 545.260 704.190 545.320 ;
        RECT 704.790 545.260 705.110 545.320 ;
        RECT 703.870 545.120 705.110 545.260 ;
        RECT 703.870 545.060 704.190 545.120 ;
        RECT 704.790 545.060 705.110 545.120 ;
        RECT 704.330 531.320 704.650 531.380 ;
        RECT 704.135 531.180 704.650 531.320 ;
        RECT 704.330 531.120 704.650 531.180 ;
        RECT 704.330 496.640 704.650 496.700 ;
        RECT 704.135 496.500 704.650 496.640 ;
        RECT 704.330 496.440 704.650 496.500 ;
        RECT 703.870 448.700 704.190 448.760 ;
        RECT 704.790 448.700 705.110 448.760 ;
        RECT 703.870 448.560 705.110 448.700 ;
        RECT 703.870 448.500 704.190 448.560 ;
        RECT 704.790 448.500 705.110 448.560 ;
        RECT 704.330 434.760 704.650 434.820 ;
        RECT 704.135 434.620 704.650 434.760 ;
        RECT 704.330 434.560 704.650 434.620 ;
        RECT 704.345 386.480 704.635 386.525 ;
        RECT 704.790 386.480 705.110 386.540 ;
        RECT 704.345 386.340 705.110 386.480 ;
        RECT 704.345 386.295 704.635 386.340 ;
        RECT 704.790 386.280 705.110 386.340 ;
        RECT 704.345 385.800 704.635 385.845 ;
        RECT 704.790 385.800 705.110 385.860 ;
        RECT 704.345 385.660 705.110 385.800 ;
        RECT 704.345 385.615 704.635 385.660 ;
        RECT 704.790 385.600 705.110 385.660 ;
        RECT 704.330 338.200 704.650 338.260 ;
        RECT 704.135 338.060 704.650 338.200 ;
        RECT 704.330 338.000 704.650 338.060 ;
        RECT 704.345 289.580 704.635 289.625 ;
        RECT 704.790 289.580 705.110 289.640 ;
        RECT 704.345 289.440 705.110 289.580 ;
        RECT 704.345 289.395 704.635 289.440 ;
        RECT 704.790 289.380 705.110 289.440 ;
        RECT 704.330 255.240 704.650 255.300 ;
        RECT 704.135 255.100 704.650 255.240 ;
        RECT 704.330 255.040 704.650 255.100 ;
        RECT 704.345 193.020 704.635 193.065 ;
        RECT 704.790 193.020 705.110 193.080 ;
        RECT 704.345 192.880 705.110 193.020 ;
        RECT 704.345 192.835 704.635 192.880 ;
        RECT 704.790 192.820 705.110 192.880 ;
        RECT 704.330 158.680 704.650 158.740 ;
        RECT 704.135 158.540 704.650 158.680 ;
        RECT 704.330 158.480 704.650 158.540 ;
        RECT 703.870 48.180 704.190 48.240 ;
        RECT 704.345 48.180 704.635 48.225 ;
        RECT 703.870 48.040 704.635 48.180 ;
        RECT 703.870 47.980 704.190 48.040 ;
        RECT 704.345 47.995 704.635 48.040 ;
        RECT 704.330 2.960 704.650 3.020 ;
        RECT 704.135 2.820 704.650 2.960 ;
        RECT 704.330 2.760 704.650 2.820 ;
      LAYER via ;
        RECT 565.440 1588.860 565.700 1589.120 ;
        RECT 703.900 1588.180 704.160 1588.440 ;
        RECT 703.900 1558.940 704.160 1559.200 ;
        RECT 704.820 1558.940 705.080 1559.200 ;
        RECT 703.900 1483.460 704.160 1483.720 ;
        RECT 704.820 1483.460 705.080 1483.720 ;
        RECT 703.900 1317.880 704.160 1318.140 ;
        RECT 704.820 1317.880 705.080 1318.140 ;
        RECT 703.900 1221.320 704.160 1221.580 ;
        RECT 704.820 1221.320 705.080 1221.580 ;
        RECT 703.900 1124.760 704.160 1125.020 ;
        RECT 704.820 1124.760 705.080 1125.020 ;
        RECT 703.900 1028.200 704.160 1028.460 ;
        RECT 704.820 1028.200 705.080 1028.460 ;
        RECT 703.900 931.640 704.160 931.900 ;
        RECT 704.820 931.640 705.080 931.900 ;
        RECT 704.820 869.420 705.080 869.680 ;
        RECT 705.740 869.420 706.000 869.680 ;
        RECT 703.900 835.080 704.160 835.340 ;
        RECT 704.820 835.080 705.080 835.340 ;
        RECT 704.360 820.800 704.620 821.060 ;
        RECT 704.360 786.460 704.620 786.720 ;
        RECT 703.900 738.180 704.160 738.440 ;
        RECT 704.820 738.180 705.080 738.440 ;
        RECT 704.360 724.240 704.620 724.500 ;
        RECT 704.360 689.560 704.620 689.820 ;
        RECT 703.900 641.620 704.160 641.880 ;
        RECT 704.820 641.620 705.080 641.880 ;
        RECT 704.360 627.680 704.620 627.940 ;
        RECT 704.360 593.000 704.620 593.260 ;
        RECT 703.900 545.060 704.160 545.320 ;
        RECT 704.820 545.060 705.080 545.320 ;
        RECT 704.360 531.120 704.620 531.380 ;
        RECT 704.360 496.440 704.620 496.700 ;
        RECT 703.900 448.500 704.160 448.760 ;
        RECT 704.820 448.500 705.080 448.760 ;
        RECT 704.360 434.560 704.620 434.820 ;
        RECT 704.820 386.280 705.080 386.540 ;
        RECT 704.820 385.600 705.080 385.860 ;
        RECT 704.360 338.000 704.620 338.260 ;
        RECT 704.820 289.380 705.080 289.640 ;
        RECT 704.360 255.040 704.620 255.300 ;
        RECT 704.820 192.820 705.080 193.080 ;
        RECT 704.360 158.480 704.620 158.740 ;
        RECT 703.900 47.980 704.160 48.240 ;
        RECT 704.360 2.760 704.620 3.020 ;
      LAYER met2 ;
        RECT 565.440 1600.000 565.720 1604.000 ;
        RECT 565.500 1589.150 565.640 1600.000 ;
        RECT 565.440 1588.830 565.700 1589.150 ;
        RECT 703.900 1588.150 704.160 1588.470 ;
        RECT 703.960 1559.230 704.100 1588.150 ;
        RECT 703.900 1558.910 704.160 1559.230 ;
        RECT 704.820 1558.910 705.080 1559.230 ;
        RECT 704.880 1483.750 705.020 1558.910 ;
        RECT 703.900 1483.430 704.160 1483.750 ;
        RECT 704.820 1483.430 705.080 1483.750 ;
        RECT 703.960 1462.410 704.100 1483.430 ;
        RECT 703.960 1462.270 704.560 1462.410 ;
        RECT 704.420 1414.810 704.560 1462.270 ;
        RECT 704.420 1414.670 705.020 1414.810 ;
        RECT 704.880 1318.170 705.020 1414.670 ;
        RECT 703.900 1317.850 704.160 1318.170 ;
        RECT 704.820 1317.850 705.080 1318.170 ;
        RECT 703.960 1317.570 704.100 1317.850 ;
        RECT 703.960 1317.430 704.560 1317.570 ;
        RECT 704.420 1269.970 704.560 1317.430 ;
        RECT 704.420 1269.830 705.020 1269.970 ;
        RECT 704.880 1221.610 705.020 1269.830 ;
        RECT 703.900 1221.290 704.160 1221.610 ;
        RECT 704.820 1221.290 705.080 1221.610 ;
        RECT 703.960 1221.010 704.100 1221.290 ;
        RECT 703.960 1220.870 704.560 1221.010 ;
        RECT 704.420 1173.410 704.560 1220.870 ;
        RECT 704.420 1173.270 705.020 1173.410 ;
        RECT 704.880 1125.050 705.020 1173.270 ;
        RECT 703.900 1124.730 704.160 1125.050 ;
        RECT 704.820 1124.730 705.080 1125.050 ;
        RECT 703.960 1124.450 704.100 1124.730 ;
        RECT 703.960 1124.310 704.560 1124.450 ;
        RECT 704.420 1076.850 704.560 1124.310 ;
        RECT 704.420 1076.710 705.020 1076.850 ;
        RECT 704.880 1028.490 705.020 1076.710 ;
        RECT 703.900 1028.170 704.160 1028.490 ;
        RECT 704.820 1028.170 705.080 1028.490 ;
        RECT 703.960 1027.890 704.100 1028.170 ;
        RECT 703.960 1027.750 704.560 1027.890 ;
        RECT 704.420 980.290 704.560 1027.750 ;
        RECT 704.420 980.150 705.020 980.290 ;
        RECT 704.880 931.930 705.020 980.150 ;
        RECT 703.900 931.610 704.160 931.930 ;
        RECT 704.820 931.610 705.080 931.930 ;
        RECT 703.960 931.330 704.100 931.610 ;
        RECT 703.960 931.190 704.560 931.330 ;
        RECT 704.420 917.845 704.560 931.190 ;
        RECT 704.350 917.475 704.630 917.845 ;
        RECT 705.730 917.475 706.010 917.845 ;
        RECT 705.800 869.710 705.940 917.475 ;
        RECT 704.820 869.390 705.080 869.710 ;
        RECT 705.740 869.390 706.000 869.710 ;
        RECT 704.880 835.370 705.020 869.390 ;
        RECT 703.900 835.050 704.160 835.370 ;
        RECT 704.820 835.050 705.080 835.370 ;
        RECT 703.960 834.770 704.100 835.050 ;
        RECT 703.960 834.630 704.560 834.770 ;
        RECT 704.420 821.090 704.560 834.630 ;
        RECT 704.360 820.770 704.620 821.090 ;
        RECT 704.360 786.430 704.620 786.750 ;
        RECT 704.420 772.890 704.560 786.430 ;
        RECT 704.420 772.750 705.020 772.890 ;
        RECT 704.880 738.470 705.020 772.750 ;
        RECT 703.900 738.210 704.160 738.470 ;
        RECT 703.900 738.150 704.560 738.210 ;
        RECT 704.820 738.150 705.080 738.470 ;
        RECT 703.960 738.070 704.560 738.150 ;
        RECT 704.420 724.530 704.560 738.070 ;
        RECT 704.360 724.210 704.620 724.530 ;
        RECT 704.360 689.530 704.620 689.850 ;
        RECT 704.420 676.330 704.560 689.530 ;
        RECT 704.420 676.190 705.020 676.330 ;
        RECT 704.880 641.910 705.020 676.190 ;
        RECT 703.900 641.650 704.160 641.910 ;
        RECT 703.900 641.590 704.560 641.650 ;
        RECT 704.820 641.590 705.080 641.910 ;
        RECT 703.960 641.510 704.560 641.590 ;
        RECT 704.420 627.970 704.560 641.510 ;
        RECT 704.360 627.650 704.620 627.970 ;
        RECT 704.360 592.970 704.620 593.290 ;
        RECT 704.420 579.770 704.560 592.970 ;
        RECT 704.420 579.630 705.020 579.770 ;
        RECT 704.880 545.350 705.020 579.630 ;
        RECT 703.900 545.090 704.160 545.350 ;
        RECT 703.900 545.030 704.560 545.090 ;
        RECT 704.820 545.030 705.080 545.350 ;
        RECT 703.960 544.950 704.560 545.030 ;
        RECT 704.420 531.410 704.560 544.950 ;
        RECT 704.360 531.090 704.620 531.410 ;
        RECT 704.360 496.410 704.620 496.730 ;
        RECT 704.420 483.210 704.560 496.410 ;
        RECT 704.420 483.070 705.020 483.210 ;
        RECT 704.880 448.790 705.020 483.070 ;
        RECT 703.900 448.530 704.160 448.790 ;
        RECT 703.900 448.470 704.560 448.530 ;
        RECT 704.820 448.470 705.080 448.790 ;
        RECT 703.960 448.390 704.560 448.470 ;
        RECT 704.420 434.850 704.560 448.390 ;
        RECT 704.360 434.530 704.620 434.850 ;
        RECT 704.820 386.250 705.080 386.570 ;
        RECT 704.880 385.890 705.020 386.250 ;
        RECT 704.820 385.570 705.080 385.890 ;
        RECT 704.360 337.970 704.620 338.290 ;
        RECT 704.420 303.690 704.560 337.970 ;
        RECT 704.420 303.550 705.020 303.690 ;
        RECT 704.880 289.670 705.020 303.550 ;
        RECT 704.820 289.350 705.080 289.670 ;
        RECT 704.360 255.010 704.620 255.330 ;
        RECT 704.420 207.130 704.560 255.010 ;
        RECT 704.420 206.990 705.020 207.130 ;
        RECT 704.880 193.110 705.020 206.990 ;
        RECT 704.820 192.790 705.080 193.110 ;
        RECT 704.360 158.450 704.620 158.770 ;
        RECT 704.420 110.570 704.560 158.450 ;
        RECT 704.420 110.430 705.020 110.570 ;
        RECT 704.880 62.290 705.020 110.430 ;
        RECT 703.960 62.150 705.020 62.290 ;
        RECT 703.960 48.270 704.100 62.150 ;
        RECT 703.900 47.950 704.160 48.270 ;
        RECT 704.360 2.730 704.620 3.050 ;
        RECT 704.420 2.400 704.560 2.730 ;
        RECT 704.210 -4.800 704.770 2.400 ;
      LAYER via2 ;
        RECT 704.350 917.520 704.630 917.800 ;
        RECT 705.730 917.520 706.010 917.800 ;
      LAYER met3 ;
        RECT 704.325 917.810 704.655 917.825 ;
        RECT 705.705 917.810 706.035 917.825 ;
        RECT 704.325 917.510 706.035 917.810 ;
        RECT 704.325 917.495 704.655 917.510 ;
        RECT 705.705 917.495 706.035 917.510 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 875.910 28.460 876.230 28.520 ;
        RECT 1525.430 28.460 1525.750 28.520 ;
        RECT 875.910 28.320 1525.750 28.460 ;
        RECT 875.910 28.260 876.230 28.320 ;
        RECT 1525.430 28.260 1525.750 28.320 ;
      LAYER via ;
        RECT 875.940 28.260 876.200 28.520 ;
        RECT 1525.460 28.260 1525.720 28.520 ;
      LAYER met2 ;
        RECT 875.480 1600.450 875.760 1604.000 ;
        RECT 875.480 1600.310 876.140 1600.450 ;
        RECT 875.480 1600.000 875.760 1600.310 ;
        RECT 876.000 28.550 876.140 1600.310 ;
        RECT 875.940 28.230 876.200 28.550 ;
        RECT 1525.460 28.230 1525.720 28.550 ;
        RECT 1525.520 14.010 1525.660 28.230 ;
        RECT 1525.060 13.870 1525.660 14.010 ;
        RECT 1525.060 2.400 1525.200 13.870 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 28.800 883.130 28.860 ;
        RECT 1542.910 28.800 1543.230 28.860 ;
        RECT 882.810 28.660 1543.230 28.800 ;
        RECT 882.810 28.600 883.130 28.660 ;
        RECT 1542.910 28.600 1543.230 28.660 ;
      LAYER via ;
        RECT 882.840 28.600 883.100 28.860 ;
        RECT 1542.940 28.600 1543.200 28.860 ;
      LAYER met2 ;
        RECT 881.920 1600.450 882.200 1604.000 ;
        RECT 881.920 1600.310 883.040 1600.450 ;
        RECT 881.920 1600.000 882.200 1600.310 ;
        RECT 882.900 28.890 883.040 1600.310 ;
        RECT 882.840 28.570 883.100 28.890 ;
        RECT 1542.940 28.570 1543.200 28.890 ;
        RECT 1543.000 2.400 1543.140 28.570 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 889.710 29.140 890.030 29.200 ;
        RECT 1560.850 29.140 1561.170 29.200 ;
        RECT 889.710 29.000 1561.170 29.140 ;
        RECT 889.710 28.940 890.030 29.000 ;
        RECT 1560.850 28.940 1561.170 29.000 ;
      LAYER via ;
        RECT 889.740 28.940 890.000 29.200 ;
        RECT 1560.880 28.940 1561.140 29.200 ;
      LAYER met2 ;
        RECT 888.820 1600.450 889.100 1604.000 ;
        RECT 888.820 1600.310 889.940 1600.450 ;
        RECT 888.820 1600.000 889.100 1600.310 ;
        RECT 889.800 29.230 889.940 1600.310 ;
        RECT 889.740 28.910 890.000 29.230 ;
        RECT 1560.880 28.910 1561.140 29.230 ;
        RECT 1560.940 2.400 1561.080 28.910 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 896.610 29.480 896.930 29.540 ;
        RECT 1578.790 29.480 1579.110 29.540 ;
        RECT 896.610 29.340 1579.110 29.480 ;
        RECT 896.610 29.280 896.930 29.340 ;
        RECT 1578.790 29.280 1579.110 29.340 ;
      LAYER via ;
        RECT 896.640 29.280 896.900 29.540 ;
        RECT 1578.820 29.280 1579.080 29.540 ;
      LAYER met2 ;
        RECT 895.720 1600.450 896.000 1604.000 ;
        RECT 895.720 1600.310 896.840 1600.450 ;
        RECT 895.720 1600.000 896.000 1600.310 ;
        RECT 896.700 29.570 896.840 1600.310 ;
        RECT 896.640 29.250 896.900 29.570 ;
        RECT 1578.820 29.250 1579.080 29.570 ;
        RECT 1578.880 2.400 1579.020 29.250 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 903.510 29.820 903.830 29.880 ;
        RECT 1596.270 29.820 1596.590 29.880 ;
        RECT 903.510 29.680 1596.590 29.820 ;
        RECT 903.510 29.620 903.830 29.680 ;
        RECT 1596.270 29.620 1596.590 29.680 ;
      LAYER via ;
        RECT 903.540 29.620 903.800 29.880 ;
        RECT 1596.300 29.620 1596.560 29.880 ;
      LAYER met2 ;
        RECT 902.160 1600.450 902.440 1604.000 ;
        RECT 902.160 1600.310 903.740 1600.450 ;
        RECT 902.160 1600.000 902.440 1600.310 ;
        RECT 903.600 29.910 903.740 1600.310 ;
        RECT 903.540 29.590 903.800 29.910 ;
        RECT 1596.300 29.590 1596.560 29.910 ;
        RECT 1596.360 2.400 1596.500 29.590 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 910.410 30.160 910.730 30.220 ;
        RECT 1614.210 30.160 1614.530 30.220 ;
        RECT 910.410 30.020 1614.530 30.160 ;
        RECT 910.410 29.960 910.730 30.020 ;
        RECT 1614.210 29.960 1614.530 30.020 ;
      LAYER via ;
        RECT 910.440 29.960 910.700 30.220 ;
        RECT 1614.240 29.960 1614.500 30.220 ;
      LAYER met2 ;
        RECT 909.060 1600.450 909.340 1604.000 ;
        RECT 909.060 1600.310 910.640 1600.450 ;
        RECT 909.060 1600.000 909.340 1600.310 ;
        RECT 910.500 30.250 910.640 1600.310 ;
        RECT 910.440 29.930 910.700 30.250 ;
        RECT 1614.240 29.930 1614.500 30.250 ;
        RECT 1614.300 2.400 1614.440 29.930 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 917.310 30.500 917.630 30.560 ;
        RECT 1632.150 30.500 1632.470 30.560 ;
        RECT 917.310 30.360 1632.470 30.500 ;
        RECT 917.310 30.300 917.630 30.360 ;
        RECT 1632.150 30.300 1632.470 30.360 ;
      LAYER via ;
        RECT 917.340 30.300 917.600 30.560 ;
        RECT 1632.180 30.300 1632.440 30.560 ;
      LAYER met2 ;
        RECT 915.960 1600.450 916.240 1604.000 ;
        RECT 915.960 1600.310 917.540 1600.450 ;
        RECT 915.960 1600.000 916.240 1600.310 ;
        RECT 917.400 30.590 917.540 1600.310 ;
        RECT 917.340 30.270 917.600 30.590 ;
        RECT 1632.180 30.270 1632.440 30.590 ;
        RECT 1632.240 2.400 1632.380 30.270 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 924.210 34.240 924.530 34.300 ;
        RECT 1650.090 34.240 1650.410 34.300 ;
        RECT 924.210 34.100 1650.410 34.240 ;
        RECT 924.210 34.040 924.530 34.100 ;
        RECT 1650.090 34.040 1650.410 34.100 ;
      LAYER via ;
        RECT 924.240 34.040 924.500 34.300 ;
        RECT 1650.120 34.040 1650.380 34.300 ;
      LAYER met2 ;
        RECT 922.400 1600.450 922.680 1604.000 ;
        RECT 922.400 1600.310 924.440 1600.450 ;
        RECT 922.400 1600.000 922.680 1600.310 ;
        RECT 924.300 34.330 924.440 1600.310 ;
        RECT 924.240 34.010 924.500 34.330 ;
        RECT 1650.120 34.010 1650.380 34.330 ;
        RECT 1650.180 2.400 1650.320 34.010 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 931.110 33.900 931.430 33.960 ;
        RECT 1668.030 33.900 1668.350 33.960 ;
        RECT 931.110 33.760 1668.350 33.900 ;
        RECT 931.110 33.700 931.430 33.760 ;
        RECT 1668.030 33.700 1668.350 33.760 ;
      LAYER via ;
        RECT 931.140 33.700 931.400 33.960 ;
        RECT 1668.060 33.700 1668.320 33.960 ;
      LAYER met2 ;
        RECT 929.300 1600.450 929.580 1604.000 ;
        RECT 929.300 1600.310 931.340 1600.450 ;
        RECT 929.300 1600.000 929.580 1600.310 ;
        RECT 931.200 33.990 931.340 1600.310 ;
        RECT 931.140 33.670 931.400 33.990 ;
        RECT 1668.060 33.670 1668.320 33.990 ;
        RECT 1668.120 2.400 1668.260 33.670 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 935.710 1589.740 936.030 1589.800 ;
        RECT 938.010 1589.740 938.330 1589.800 ;
        RECT 935.710 1589.600 938.330 1589.740 ;
        RECT 935.710 1589.540 936.030 1589.600 ;
        RECT 938.010 1589.540 938.330 1589.600 ;
        RECT 938.010 33.560 938.330 33.620 ;
        RECT 1685.510 33.560 1685.830 33.620 ;
        RECT 938.010 33.420 1685.830 33.560 ;
        RECT 938.010 33.360 938.330 33.420 ;
        RECT 1685.510 33.360 1685.830 33.420 ;
      LAYER via ;
        RECT 935.740 1589.540 936.000 1589.800 ;
        RECT 938.040 1589.540 938.300 1589.800 ;
        RECT 938.040 33.360 938.300 33.620 ;
        RECT 1685.540 33.360 1685.800 33.620 ;
      LAYER met2 ;
        RECT 935.740 1600.000 936.020 1604.000 ;
        RECT 935.800 1589.830 935.940 1600.000 ;
        RECT 935.740 1589.510 936.000 1589.830 ;
        RECT 938.040 1589.510 938.300 1589.830 ;
        RECT 938.100 33.650 938.240 1589.510 ;
        RECT 938.040 33.330 938.300 33.650 ;
        RECT 1685.540 33.330 1685.800 33.650 ;
        RECT 1685.600 2.400 1685.740 33.330 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.340 1600.000 572.620 1604.000 ;
        RECT 572.400 16.845 572.540 1600.000 ;
        RECT 572.330 16.475 572.610 16.845 ;
        RECT 722.290 16.475 722.570 16.845 ;
        RECT 722.360 2.400 722.500 16.475 ;
        RECT 722.150 -4.800 722.710 2.400 ;
      LAYER via2 ;
        RECT 572.330 16.520 572.610 16.800 ;
        RECT 722.290 16.520 722.570 16.800 ;
      LAYER met3 ;
        RECT 572.305 16.810 572.635 16.825 ;
        RECT 722.265 16.810 722.595 16.825 ;
        RECT 572.305 16.510 722.595 16.810 ;
        RECT 572.305 16.495 572.635 16.510 ;
        RECT 722.265 16.495 722.595 16.510 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 942.610 1590.080 942.930 1590.140 ;
        RECT 944.910 1590.080 945.230 1590.140 ;
        RECT 942.610 1589.940 945.230 1590.080 ;
        RECT 942.610 1589.880 942.930 1589.940 ;
        RECT 944.910 1589.880 945.230 1589.940 ;
        RECT 944.910 33.220 945.230 33.280 ;
        RECT 1703.450 33.220 1703.770 33.280 ;
        RECT 944.910 33.080 1703.770 33.220 ;
        RECT 944.910 33.020 945.230 33.080 ;
        RECT 1703.450 33.020 1703.770 33.080 ;
      LAYER via ;
        RECT 942.640 1589.880 942.900 1590.140 ;
        RECT 944.940 1589.880 945.200 1590.140 ;
        RECT 944.940 33.020 945.200 33.280 ;
        RECT 1703.480 33.020 1703.740 33.280 ;
      LAYER met2 ;
        RECT 942.640 1600.000 942.920 1604.000 ;
        RECT 942.700 1590.170 942.840 1600.000 ;
        RECT 942.640 1589.850 942.900 1590.170 ;
        RECT 944.940 1589.850 945.200 1590.170 ;
        RECT 945.000 33.310 945.140 1589.850 ;
        RECT 944.940 32.990 945.200 33.310 ;
        RECT 1703.480 32.990 1703.740 33.310 ;
        RECT 1703.540 2.400 1703.680 32.990 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 949.510 1590.080 949.830 1590.140 ;
        RECT 951.810 1590.080 952.130 1590.140 ;
        RECT 949.510 1589.940 952.130 1590.080 ;
        RECT 949.510 1589.880 949.830 1589.940 ;
        RECT 951.810 1589.880 952.130 1589.940 ;
        RECT 951.810 32.880 952.130 32.940 ;
        RECT 1721.390 32.880 1721.710 32.940 ;
        RECT 951.810 32.740 1721.710 32.880 ;
        RECT 951.810 32.680 952.130 32.740 ;
        RECT 1721.390 32.680 1721.710 32.740 ;
      LAYER via ;
        RECT 949.540 1589.880 949.800 1590.140 ;
        RECT 951.840 1589.880 952.100 1590.140 ;
        RECT 951.840 32.680 952.100 32.940 ;
        RECT 1721.420 32.680 1721.680 32.940 ;
      LAYER met2 ;
        RECT 949.540 1600.000 949.820 1604.000 ;
        RECT 949.600 1590.170 949.740 1600.000 ;
        RECT 949.540 1589.850 949.800 1590.170 ;
        RECT 951.840 1589.850 952.100 1590.170 ;
        RECT 951.900 32.970 952.040 1589.850 ;
        RECT 951.840 32.650 952.100 32.970 ;
        RECT 1721.420 32.650 1721.680 32.970 ;
        RECT 1721.480 2.400 1721.620 32.650 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 955.950 1590.080 956.270 1590.140 ;
        RECT 958.250 1590.080 958.570 1590.140 ;
        RECT 955.950 1589.940 958.570 1590.080 ;
        RECT 955.950 1589.880 956.270 1589.940 ;
        RECT 958.250 1589.880 958.570 1589.940 ;
      LAYER via ;
        RECT 955.980 1589.880 956.240 1590.140 ;
        RECT 958.280 1589.880 958.540 1590.140 ;
      LAYER met2 ;
        RECT 955.980 1600.000 956.260 1604.000 ;
        RECT 956.040 1590.170 956.180 1600.000 ;
        RECT 955.980 1589.850 956.240 1590.170 ;
        RECT 958.280 1589.850 958.540 1590.170 ;
        RECT 958.340 26.365 958.480 1589.850 ;
        RECT 958.270 25.995 958.550 26.365 ;
        RECT 1739.350 25.995 1739.630 26.365 ;
        RECT 1739.420 2.400 1739.560 25.995 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
      LAYER via2 ;
        RECT 958.270 26.040 958.550 26.320 ;
        RECT 1739.350 26.040 1739.630 26.320 ;
      LAYER met3 ;
        RECT 958.245 26.330 958.575 26.345 ;
        RECT 1739.325 26.330 1739.655 26.345 ;
        RECT 958.245 26.030 1739.655 26.330 ;
        RECT 958.245 26.015 958.575 26.030 ;
        RECT 1739.325 26.015 1739.655 26.030 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 962.850 1589.740 963.170 1589.800 ;
        RECT 965.610 1589.740 965.930 1589.800 ;
        RECT 962.850 1589.600 965.930 1589.740 ;
        RECT 962.850 1589.540 963.170 1589.600 ;
        RECT 965.610 1589.540 965.930 1589.600 ;
        RECT 965.610 32.540 965.930 32.600 ;
        RECT 1756.810 32.540 1757.130 32.600 ;
        RECT 965.610 32.400 1757.130 32.540 ;
        RECT 965.610 32.340 965.930 32.400 ;
        RECT 1756.810 32.340 1757.130 32.400 ;
      LAYER via ;
        RECT 962.880 1589.540 963.140 1589.800 ;
        RECT 965.640 1589.540 965.900 1589.800 ;
        RECT 965.640 32.340 965.900 32.600 ;
        RECT 1756.840 32.340 1757.100 32.600 ;
      LAYER met2 ;
        RECT 962.880 1600.000 963.160 1604.000 ;
        RECT 962.940 1589.830 963.080 1600.000 ;
        RECT 962.880 1589.510 963.140 1589.830 ;
        RECT 965.640 1589.510 965.900 1589.830 ;
        RECT 965.700 32.630 965.840 1589.510 ;
        RECT 965.640 32.310 965.900 32.630 ;
        RECT 1756.840 32.310 1757.100 32.630 ;
        RECT 1756.900 2.400 1757.040 32.310 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 969.750 1590.080 970.070 1590.140 ;
        RECT 972.510 1590.080 972.830 1590.140 ;
        RECT 969.750 1589.940 972.830 1590.080 ;
        RECT 969.750 1589.880 970.070 1589.940 ;
        RECT 972.510 1589.880 972.830 1589.940 ;
        RECT 972.510 32.200 972.830 32.260 ;
        RECT 1774.750 32.200 1775.070 32.260 ;
        RECT 972.510 32.060 1775.070 32.200 ;
        RECT 972.510 32.000 972.830 32.060 ;
        RECT 1774.750 32.000 1775.070 32.060 ;
      LAYER via ;
        RECT 969.780 1589.880 970.040 1590.140 ;
        RECT 972.540 1589.880 972.800 1590.140 ;
        RECT 972.540 32.000 972.800 32.260 ;
        RECT 1774.780 32.000 1775.040 32.260 ;
      LAYER met2 ;
        RECT 969.780 1600.000 970.060 1604.000 ;
        RECT 969.840 1590.170 969.980 1600.000 ;
        RECT 969.780 1589.850 970.040 1590.170 ;
        RECT 972.540 1589.850 972.800 1590.170 ;
        RECT 972.600 32.290 972.740 1589.850 ;
        RECT 972.540 31.970 972.800 32.290 ;
        RECT 1774.780 31.970 1775.040 32.290 ;
        RECT 1774.840 2.400 1774.980 31.970 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 976.190 1589.740 976.510 1589.800 ;
        RECT 979.410 1589.740 979.730 1589.800 ;
        RECT 976.190 1589.600 979.730 1589.740 ;
        RECT 976.190 1589.540 976.510 1589.600 ;
        RECT 979.410 1589.540 979.730 1589.600 ;
        RECT 979.410 31.860 979.730 31.920 ;
        RECT 1792.690 31.860 1793.010 31.920 ;
        RECT 979.410 31.720 1793.010 31.860 ;
        RECT 979.410 31.660 979.730 31.720 ;
        RECT 1792.690 31.660 1793.010 31.720 ;
      LAYER via ;
        RECT 976.220 1589.540 976.480 1589.800 ;
        RECT 979.440 1589.540 979.700 1589.800 ;
        RECT 979.440 31.660 979.700 31.920 ;
        RECT 1792.720 31.660 1792.980 31.920 ;
      LAYER met2 ;
        RECT 976.220 1600.000 976.500 1604.000 ;
        RECT 976.280 1589.830 976.420 1600.000 ;
        RECT 976.220 1589.510 976.480 1589.830 ;
        RECT 979.440 1589.510 979.700 1589.830 ;
        RECT 979.500 31.950 979.640 1589.510 ;
        RECT 979.440 31.630 979.700 31.950 ;
        RECT 1792.720 31.630 1792.980 31.950 ;
        RECT 1792.780 2.400 1792.920 31.630 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 983.090 1590.080 983.410 1590.140 ;
        RECT 985.850 1590.080 986.170 1590.140 ;
        RECT 983.090 1589.940 986.170 1590.080 ;
        RECT 983.090 1589.880 983.410 1589.940 ;
        RECT 985.850 1589.880 986.170 1589.940 ;
      LAYER via ;
        RECT 983.120 1589.880 983.380 1590.140 ;
        RECT 985.880 1589.880 986.140 1590.140 ;
      LAYER met2 ;
        RECT 983.120 1600.000 983.400 1604.000 ;
        RECT 983.180 1590.170 983.320 1600.000 ;
        RECT 983.120 1589.850 983.380 1590.170 ;
        RECT 985.880 1589.850 986.140 1590.170 ;
        RECT 985.940 33.845 986.080 1589.850 ;
        RECT 985.870 33.475 986.150 33.845 ;
        RECT 1810.650 33.475 1810.930 33.845 ;
        RECT 1810.720 2.400 1810.860 33.475 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
      LAYER via2 ;
        RECT 985.870 33.520 986.150 33.800 ;
        RECT 1810.650 33.520 1810.930 33.800 ;
      LAYER met3 ;
        RECT 985.845 33.810 986.175 33.825 ;
        RECT 1810.625 33.810 1810.955 33.825 ;
        RECT 985.845 33.510 1810.955 33.810 ;
        RECT 985.845 33.495 986.175 33.510 ;
        RECT 1810.625 33.495 1810.955 33.510 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 989.990 1587.360 990.310 1587.420 ;
        RECT 993.210 1587.360 993.530 1587.420 ;
        RECT 989.990 1587.220 993.530 1587.360 ;
        RECT 989.990 1587.160 990.310 1587.220 ;
        RECT 993.210 1587.160 993.530 1587.220 ;
      LAYER via ;
        RECT 990.020 1587.160 990.280 1587.420 ;
        RECT 993.240 1587.160 993.500 1587.420 ;
      LAYER met2 ;
        RECT 990.020 1600.000 990.300 1604.000 ;
        RECT 990.080 1587.450 990.220 1600.000 ;
        RECT 990.020 1587.130 990.280 1587.450 ;
        RECT 993.240 1587.130 993.500 1587.450 ;
        RECT 993.300 33.165 993.440 1587.130 ;
        RECT 993.230 32.795 993.510 33.165 ;
        RECT 1829.050 32.795 1829.330 33.165 ;
        RECT 1829.120 3.130 1829.260 32.795 ;
        RECT 1828.660 2.990 1829.260 3.130 ;
        RECT 1828.660 2.400 1828.800 2.990 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
      LAYER via2 ;
        RECT 993.230 32.840 993.510 33.120 ;
        RECT 1829.050 32.840 1829.330 33.120 ;
      LAYER met3 ;
        RECT 993.205 33.130 993.535 33.145 ;
        RECT 1829.025 33.130 1829.355 33.145 ;
        RECT 993.205 32.830 1829.355 33.130 ;
        RECT 993.205 32.815 993.535 32.830 ;
        RECT 1829.025 32.815 1829.355 32.830 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 996.430 1590.080 996.750 1590.140 ;
        RECT 1000.110 1590.080 1000.430 1590.140 ;
        RECT 996.430 1589.940 1000.430 1590.080 ;
        RECT 996.430 1589.880 996.750 1589.940 ;
        RECT 1000.110 1589.880 1000.430 1589.940 ;
        RECT 1000.110 31.520 1000.430 31.580 ;
        RECT 1846.050 31.520 1846.370 31.580 ;
        RECT 1000.110 31.380 1846.370 31.520 ;
        RECT 1000.110 31.320 1000.430 31.380 ;
        RECT 1846.050 31.320 1846.370 31.380 ;
      LAYER via ;
        RECT 996.460 1589.880 996.720 1590.140 ;
        RECT 1000.140 1589.880 1000.400 1590.140 ;
        RECT 1000.140 31.320 1000.400 31.580 ;
        RECT 1846.080 31.320 1846.340 31.580 ;
      LAYER met2 ;
        RECT 996.460 1600.000 996.740 1604.000 ;
        RECT 996.520 1590.170 996.660 1600.000 ;
        RECT 996.460 1589.850 996.720 1590.170 ;
        RECT 1000.140 1589.850 1000.400 1590.170 ;
        RECT 1000.200 31.610 1000.340 1589.850 ;
        RECT 1000.140 31.290 1000.400 31.610 ;
        RECT 1846.080 31.290 1846.340 31.610 ;
        RECT 1846.140 2.400 1846.280 31.290 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1003.330 1589.740 1003.650 1589.800 ;
        RECT 1007.010 1589.740 1007.330 1589.800 ;
        RECT 1003.330 1589.600 1007.330 1589.740 ;
        RECT 1003.330 1589.540 1003.650 1589.600 ;
        RECT 1007.010 1589.540 1007.330 1589.600 ;
      LAYER via ;
        RECT 1003.360 1589.540 1003.620 1589.800 ;
        RECT 1007.040 1589.540 1007.300 1589.800 ;
      LAYER met2 ;
        RECT 1003.360 1600.000 1003.640 1604.000 ;
        RECT 1003.420 1589.830 1003.560 1600.000 ;
        RECT 1003.360 1589.510 1003.620 1589.830 ;
        RECT 1007.040 1589.510 1007.300 1589.830 ;
        RECT 1007.100 32.485 1007.240 1589.510 ;
        RECT 1007.030 32.115 1007.310 32.485 ;
        RECT 1864.010 32.115 1864.290 32.485 ;
        RECT 1864.080 2.400 1864.220 32.115 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
      LAYER via2 ;
        RECT 1007.030 32.160 1007.310 32.440 ;
        RECT 1864.010 32.160 1864.290 32.440 ;
      LAYER met3 ;
        RECT 1007.005 32.450 1007.335 32.465 ;
        RECT 1863.985 32.450 1864.315 32.465 ;
        RECT 1007.005 32.150 1864.315 32.450 ;
        RECT 1007.005 32.135 1007.335 32.150 ;
        RECT 1863.985 32.135 1864.315 32.150 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 728.250 1594.160 728.570 1594.220 ;
        RECT 690.160 1594.020 728.570 1594.160 ;
        RECT 579.210 1593.820 579.530 1593.880 ;
        RECT 690.160 1593.820 690.300 1594.020 ;
        RECT 728.250 1593.960 728.570 1594.020 ;
        RECT 579.210 1593.680 690.300 1593.820 ;
        RECT 579.210 1593.620 579.530 1593.680 ;
        RECT 729.170 16.560 729.490 16.620 ;
        RECT 740.210 16.560 740.530 16.620 ;
        RECT 729.170 16.420 740.530 16.560 ;
        RECT 729.170 16.360 729.490 16.420 ;
        RECT 740.210 16.360 740.530 16.420 ;
      LAYER via ;
        RECT 579.240 1593.620 579.500 1593.880 ;
        RECT 728.280 1593.960 728.540 1594.220 ;
        RECT 729.200 16.360 729.460 16.620 ;
        RECT 740.240 16.360 740.500 16.620 ;
      LAYER met2 ;
        RECT 579.240 1600.000 579.520 1604.000 ;
        RECT 579.300 1593.910 579.440 1600.000 ;
        RECT 728.280 1593.930 728.540 1594.250 ;
        RECT 579.240 1593.590 579.500 1593.910 ;
        RECT 728.340 39.170 728.480 1593.930 ;
        RECT 728.340 39.030 729.400 39.170 ;
        RECT 729.260 16.650 729.400 39.030 ;
        RECT 729.200 16.330 729.460 16.650 ;
        RECT 740.240 16.330 740.500 16.650 ;
        RECT 740.300 2.400 740.440 16.330 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1013.985 20.825 1014.155 34.595 ;
      LAYER mcon ;
        RECT 1013.985 34.425 1014.155 34.595 ;
      LAYER met1 ;
        RECT 1009.770 1587.360 1010.090 1587.420 ;
        RECT 1013.910 1587.360 1014.230 1587.420 ;
        RECT 1009.770 1587.220 1014.230 1587.360 ;
        RECT 1009.770 1587.160 1010.090 1587.220 ;
        RECT 1013.910 1587.160 1014.230 1587.220 ;
        RECT 1013.910 34.580 1014.230 34.640 ;
        RECT 1013.715 34.440 1014.230 34.580 ;
        RECT 1013.910 34.380 1014.230 34.440 ;
        RECT 1013.925 20.980 1014.215 21.025 ;
        RECT 1881.930 20.980 1882.250 21.040 ;
        RECT 1013.925 20.840 1882.250 20.980 ;
        RECT 1013.925 20.795 1014.215 20.840 ;
        RECT 1881.930 20.780 1882.250 20.840 ;
      LAYER via ;
        RECT 1009.800 1587.160 1010.060 1587.420 ;
        RECT 1013.940 1587.160 1014.200 1587.420 ;
        RECT 1013.940 34.380 1014.200 34.640 ;
        RECT 1881.960 20.780 1882.220 21.040 ;
      LAYER met2 ;
        RECT 1009.800 1600.000 1010.080 1604.000 ;
        RECT 1009.860 1587.450 1010.000 1600.000 ;
        RECT 1009.800 1587.130 1010.060 1587.450 ;
        RECT 1013.940 1587.130 1014.200 1587.450 ;
        RECT 1014.000 34.670 1014.140 1587.130 ;
        RECT 1013.940 34.350 1014.200 34.670 ;
        RECT 1881.960 20.750 1882.220 21.070 ;
        RECT 1882.020 2.400 1882.160 20.750 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1016.670 1589.740 1016.990 1589.800 ;
        RECT 1020.810 1589.740 1021.130 1589.800 ;
        RECT 1016.670 1589.600 1021.130 1589.740 ;
        RECT 1016.670 1589.540 1016.990 1589.600 ;
        RECT 1020.810 1589.540 1021.130 1589.600 ;
      LAYER via ;
        RECT 1016.700 1589.540 1016.960 1589.800 ;
        RECT 1020.840 1589.540 1021.100 1589.800 ;
      LAYER met2 ;
        RECT 1016.700 1600.000 1016.980 1604.000 ;
        RECT 1016.760 1589.830 1016.900 1600.000 ;
        RECT 1016.700 1589.510 1016.960 1589.830 ;
        RECT 1020.840 1589.510 1021.100 1589.830 ;
        RECT 1020.900 31.805 1021.040 1589.510 ;
        RECT 1020.830 31.435 1021.110 31.805 ;
        RECT 1899.890 31.435 1900.170 31.805 ;
        RECT 1899.960 2.400 1900.100 31.435 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
      LAYER via2 ;
        RECT 1020.830 31.480 1021.110 31.760 ;
        RECT 1899.890 31.480 1900.170 31.760 ;
      LAYER met3 ;
        RECT 1020.805 31.770 1021.135 31.785 ;
        RECT 1899.865 31.770 1900.195 31.785 ;
        RECT 1020.805 31.470 1900.195 31.770 ;
        RECT 1020.805 31.455 1021.135 31.470 ;
        RECT 1899.865 31.455 1900.195 31.470 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1023.570 1588.380 1023.890 1588.440 ;
        RECT 1027.710 1588.380 1028.030 1588.440 ;
        RECT 1023.570 1588.240 1028.030 1588.380 ;
        RECT 1023.570 1588.180 1023.890 1588.240 ;
        RECT 1027.710 1588.180 1028.030 1588.240 ;
        RECT 1027.710 21.320 1028.030 21.380 ;
        RECT 1917.810 21.320 1918.130 21.380 ;
        RECT 1027.710 21.180 1918.130 21.320 ;
        RECT 1027.710 21.120 1028.030 21.180 ;
        RECT 1917.810 21.120 1918.130 21.180 ;
      LAYER via ;
        RECT 1023.600 1588.180 1023.860 1588.440 ;
        RECT 1027.740 1588.180 1028.000 1588.440 ;
        RECT 1027.740 21.120 1028.000 21.380 ;
        RECT 1917.840 21.120 1918.100 21.380 ;
      LAYER met2 ;
        RECT 1023.600 1600.000 1023.880 1604.000 ;
        RECT 1023.660 1588.470 1023.800 1600.000 ;
        RECT 1023.600 1588.150 1023.860 1588.470 ;
        RECT 1027.740 1588.150 1028.000 1588.470 ;
        RECT 1027.800 21.410 1027.940 1588.150 ;
        RECT 1027.740 21.090 1028.000 21.410 ;
        RECT 1917.840 21.090 1918.100 21.410 ;
        RECT 1917.900 2.400 1918.040 21.090 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1030.010 1590.080 1030.330 1590.140 ;
        RECT 1034.150 1590.080 1034.470 1590.140 ;
        RECT 1030.010 1589.940 1034.470 1590.080 ;
        RECT 1030.010 1589.880 1030.330 1589.940 ;
        RECT 1034.150 1589.880 1034.470 1589.940 ;
      LAYER via ;
        RECT 1030.040 1589.880 1030.300 1590.140 ;
        RECT 1034.180 1589.880 1034.440 1590.140 ;
      LAYER met2 ;
        RECT 1030.040 1600.000 1030.320 1604.000 ;
        RECT 1030.100 1590.170 1030.240 1600.000 ;
        RECT 1030.040 1589.850 1030.300 1590.170 ;
        RECT 1034.180 1589.850 1034.440 1590.170 ;
        RECT 1034.240 31.125 1034.380 1589.850 ;
        RECT 1034.170 30.755 1034.450 31.125 ;
        RECT 1935.310 30.755 1935.590 31.125 ;
        RECT 1935.380 2.400 1935.520 30.755 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
      LAYER via2 ;
        RECT 1034.170 30.800 1034.450 31.080 ;
        RECT 1935.310 30.800 1935.590 31.080 ;
      LAYER met3 ;
        RECT 1034.145 31.090 1034.475 31.105 ;
        RECT 1935.285 31.090 1935.615 31.105 ;
        RECT 1034.145 30.790 1935.615 31.090 ;
        RECT 1034.145 30.775 1034.475 30.790 ;
        RECT 1935.285 30.775 1935.615 30.790 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1036.910 1590.080 1037.230 1590.140 ;
        RECT 1040.590 1590.080 1040.910 1590.140 ;
        RECT 1036.910 1589.940 1040.910 1590.080 ;
        RECT 1036.910 1589.880 1037.230 1589.940 ;
        RECT 1040.590 1589.880 1040.910 1589.940 ;
        RECT 1040.590 71.300 1040.910 71.360 ;
        RECT 1952.770 71.300 1953.090 71.360 ;
        RECT 1040.590 71.160 1953.090 71.300 ;
        RECT 1040.590 71.100 1040.910 71.160 ;
        RECT 1952.770 71.100 1953.090 71.160 ;
      LAYER via ;
        RECT 1036.940 1589.880 1037.200 1590.140 ;
        RECT 1040.620 1589.880 1040.880 1590.140 ;
        RECT 1040.620 71.100 1040.880 71.360 ;
        RECT 1952.800 71.100 1953.060 71.360 ;
      LAYER met2 ;
        RECT 1036.940 1600.000 1037.220 1604.000 ;
        RECT 1037.000 1590.170 1037.140 1600.000 ;
        RECT 1036.940 1589.850 1037.200 1590.170 ;
        RECT 1040.620 1589.850 1040.880 1590.170 ;
        RECT 1040.680 71.390 1040.820 1589.850 ;
        RECT 1040.620 71.070 1040.880 71.390 ;
        RECT 1952.800 71.070 1953.060 71.390 ;
        RECT 1952.860 7.890 1953.000 71.070 ;
        RECT 1952.860 7.750 1953.460 7.890 ;
        RECT 1953.320 2.400 1953.460 7.750 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1043.810 1590.080 1044.130 1590.140 ;
        RECT 1047.950 1590.080 1048.270 1590.140 ;
        RECT 1043.810 1589.940 1048.270 1590.080 ;
        RECT 1043.810 1589.880 1044.130 1589.940 ;
        RECT 1047.950 1589.880 1048.270 1589.940 ;
        RECT 1047.950 21.660 1048.270 21.720 ;
        RECT 1971.170 21.660 1971.490 21.720 ;
        RECT 1047.950 21.520 1971.490 21.660 ;
        RECT 1047.950 21.460 1048.270 21.520 ;
        RECT 1971.170 21.460 1971.490 21.520 ;
      LAYER via ;
        RECT 1043.840 1589.880 1044.100 1590.140 ;
        RECT 1047.980 1589.880 1048.240 1590.140 ;
        RECT 1047.980 21.460 1048.240 21.720 ;
        RECT 1971.200 21.460 1971.460 21.720 ;
      LAYER met2 ;
        RECT 1043.840 1600.000 1044.120 1604.000 ;
        RECT 1043.900 1590.170 1044.040 1600.000 ;
        RECT 1043.840 1589.850 1044.100 1590.170 ;
        RECT 1047.980 1589.850 1048.240 1590.170 ;
        RECT 1048.040 21.750 1048.180 1589.850 ;
        RECT 1047.980 21.430 1048.240 21.750 ;
        RECT 1971.200 21.430 1971.460 21.750 ;
        RECT 1971.260 2.400 1971.400 21.430 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1050.250 1590.080 1050.570 1590.140 ;
        RECT 1055.310 1590.080 1055.630 1590.140 ;
        RECT 1050.250 1589.940 1055.630 1590.080 ;
        RECT 1050.250 1589.880 1050.570 1589.940 ;
        RECT 1055.310 1589.880 1055.630 1589.940 ;
        RECT 1055.310 35.260 1055.630 35.320 ;
        RECT 1989.110 35.260 1989.430 35.320 ;
        RECT 1055.310 35.120 1989.430 35.260 ;
        RECT 1055.310 35.060 1055.630 35.120 ;
        RECT 1989.110 35.060 1989.430 35.120 ;
      LAYER via ;
        RECT 1050.280 1589.880 1050.540 1590.140 ;
        RECT 1055.340 1589.880 1055.600 1590.140 ;
        RECT 1055.340 35.060 1055.600 35.320 ;
        RECT 1989.140 35.060 1989.400 35.320 ;
      LAYER met2 ;
        RECT 1050.280 1600.000 1050.560 1604.000 ;
        RECT 1050.340 1590.170 1050.480 1600.000 ;
        RECT 1050.280 1589.850 1050.540 1590.170 ;
        RECT 1055.340 1589.850 1055.600 1590.170 ;
        RECT 1055.400 35.350 1055.540 1589.850 ;
        RECT 1055.340 35.030 1055.600 35.350 ;
        RECT 1989.140 35.030 1989.400 35.350 ;
        RECT 1989.200 2.400 1989.340 35.030 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1057.150 1590.080 1057.470 1590.140 ;
        RECT 1062.210 1590.080 1062.530 1590.140 ;
        RECT 1057.150 1589.940 1062.530 1590.080 ;
        RECT 1057.150 1589.880 1057.470 1589.940 ;
        RECT 1062.210 1589.880 1062.530 1589.940 ;
        RECT 1062.210 35.600 1062.530 35.660 ;
        RECT 2006.590 35.600 2006.910 35.660 ;
        RECT 1062.210 35.460 2006.910 35.600 ;
        RECT 1062.210 35.400 1062.530 35.460 ;
        RECT 2006.590 35.400 2006.910 35.460 ;
      LAYER via ;
        RECT 1057.180 1589.880 1057.440 1590.140 ;
        RECT 1062.240 1589.880 1062.500 1590.140 ;
        RECT 1062.240 35.400 1062.500 35.660 ;
        RECT 2006.620 35.400 2006.880 35.660 ;
      LAYER met2 ;
        RECT 1057.180 1600.000 1057.460 1604.000 ;
        RECT 1057.240 1590.170 1057.380 1600.000 ;
        RECT 1057.180 1589.850 1057.440 1590.170 ;
        RECT 1062.240 1589.850 1062.500 1590.170 ;
        RECT 1062.300 35.690 1062.440 1589.850 ;
        RECT 1062.240 35.370 1062.500 35.690 ;
        RECT 2006.620 35.370 2006.880 35.690 ;
        RECT 2006.680 2.400 2006.820 35.370 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1064.050 1589.740 1064.370 1589.800 ;
        RECT 1069.110 1589.740 1069.430 1589.800 ;
        RECT 1064.050 1589.600 1069.430 1589.740 ;
        RECT 1064.050 1589.540 1064.370 1589.600 ;
        RECT 1069.110 1589.540 1069.430 1589.600 ;
        RECT 1069.110 35.940 1069.430 36.000 ;
        RECT 2024.530 35.940 2024.850 36.000 ;
        RECT 1069.110 35.800 2024.850 35.940 ;
        RECT 1069.110 35.740 1069.430 35.800 ;
        RECT 2024.530 35.740 2024.850 35.800 ;
      LAYER via ;
        RECT 1064.080 1589.540 1064.340 1589.800 ;
        RECT 1069.140 1589.540 1069.400 1589.800 ;
        RECT 1069.140 35.740 1069.400 36.000 ;
        RECT 2024.560 35.740 2024.820 36.000 ;
      LAYER met2 ;
        RECT 1064.080 1600.000 1064.360 1604.000 ;
        RECT 1064.140 1589.830 1064.280 1600.000 ;
        RECT 1064.080 1589.510 1064.340 1589.830 ;
        RECT 1069.140 1589.510 1069.400 1589.830 ;
        RECT 1069.200 36.030 1069.340 1589.510 ;
        RECT 1069.140 35.710 1069.400 36.030 ;
        RECT 2024.560 35.710 2024.820 36.030 ;
        RECT 2024.620 2.400 2024.760 35.710 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1070.490 1590.080 1070.810 1590.140 ;
        RECT 1075.550 1590.080 1075.870 1590.140 ;
        RECT 1070.490 1589.940 1075.870 1590.080 ;
        RECT 1070.490 1589.880 1070.810 1589.940 ;
        RECT 1075.550 1589.880 1075.870 1589.940 ;
        RECT 1075.550 36.280 1075.870 36.340 ;
        RECT 2042.930 36.280 2043.250 36.340 ;
        RECT 1075.550 36.140 2043.250 36.280 ;
        RECT 1075.550 36.080 1075.870 36.140 ;
        RECT 2042.930 36.080 2043.250 36.140 ;
      LAYER via ;
        RECT 1070.520 1589.880 1070.780 1590.140 ;
        RECT 1075.580 1589.880 1075.840 1590.140 ;
        RECT 1075.580 36.080 1075.840 36.340 ;
        RECT 2042.960 36.080 2043.220 36.340 ;
      LAYER met2 ;
        RECT 1070.520 1600.000 1070.800 1604.000 ;
        RECT 1070.580 1590.170 1070.720 1600.000 ;
        RECT 1070.520 1589.850 1070.780 1590.170 ;
        RECT 1075.580 1589.850 1075.840 1590.170 ;
        RECT 1075.640 36.370 1075.780 1589.850 ;
        RECT 1075.580 36.050 1075.840 36.370 ;
        RECT 2042.960 36.050 2043.220 36.370 ;
        RECT 2043.020 17.410 2043.160 36.050 ;
        RECT 2042.560 17.270 2043.160 17.410 ;
        RECT 2042.560 2.400 2042.700 17.270 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 718.205 1589.585 718.375 1593.155 ;
        RECT 733.385 1588.395 733.555 1589.755 ;
        RECT 733.385 1588.225 737.695 1588.395 ;
        RECT 737.525 1587.885 737.695 1588.225 ;
      LAYER mcon ;
        RECT 718.205 1592.985 718.375 1593.155 ;
        RECT 733.385 1589.585 733.555 1589.755 ;
      LAYER met1 ;
        RECT 585.650 1593.480 585.970 1593.540 ;
        RECT 585.650 1593.340 714.680 1593.480 ;
        RECT 585.650 1593.280 585.970 1593.340 ;
        RECT 714.540 1593.140 714.680 1593.340 ;
        RECT 718.145 1593.140 718.435 1593.185 ;
        RECT 714.540 1593.000 718.435 1593.140 ;
        RECT 718.145 1592.955 718.435 1593.000 ;
        RECT 718.145 1589.740 718.435 1589.785 ;
        RECT 733.325 1589.740 733.615 1589.785 ;
        RECT 718.145 1589.600 733.615 1589.740 ;
        RECT 718.145 1589.555 718.435 1589.600 ;
        RECT 733.325 1589.555 733.615 1589.600 ;
        RECT 737.465 1588.040 737.755 1588.085 ;
        RECT 741.590 1588.040 741.910 1588.100 ;
        RECT 737.465 1587.900 741.910 1588.040 ;
        RECT 737.465 1587.855 737.755 1587.900 ;
        RECT 741.590 1587.840 741.910 1587.900 ;
        RECT 741.590 20.640 741.910 20.700 ;
        RECT 757.690 20.640 758.010 20.700 ;
        RECT 741.590 20.500 758.010 20.640 ;
        RECT 741.590 20.440 741.910 20.500 ;
        RECT 757.690 20.440 758.010 20.500 ;
      LAYER via ;
        RECT 585.680 1593.280 585.940 1593.540 ;
        RECT 741.620 1587.840 741.880 1588.100 ;
        RECT 741.620 20.440 741.880 20.700 ;
        RECT 757.720 20.440 757.980 20.700 ;
      LAYER met2 ;
        RECT 585.680 1600.000 585.960 1604.000 ;
        RECT 585.740 1593.570 585.880 1600.000 ;
        RECT 585.680 1593.250 585.940 1593.570 ;
        RECT 741.620 1587.810 741.880 1588.130 ;
        RECT 741.680 20.730 741.820 1587.810 ;
        RECT 741.620 20.410 741.880 20.730 ;
        RECT 757.720 20.410 757.980 20.730 ;
        RECT 757.780 2.400 757.920 20.410 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1077.390 1589.740 1077.710 1589.800 ;
        RECT 1082.910 1589.740 1083.230 1589.800 ;
        RECT 1077.390 1589.600 1083.230 1589.740 ;
        RECT 1077.390 1589.540 1077.710 1589.600 ;
        RECT 1082.910 1589.540 1083.230 1589.600 ;
        RECT 1082.910 36.620 1083.230 36.680 ;
        RECT 2060.410 36.620 2060.730 36.680 ;
        RECT 1082.910 36.480 2060.730 36.620 ;
        RECT 1082.910 36.420 1083.230 36.480 ;
        RECT 2060.410 36.420 2060.730 36.480 ;
      LAYER via ;
        RECT 1077.420 1589.540 1077.680 1589.800 ;
        RECT 1082.940 1589.540 1083.200 1589.800 ;
        RECT 1082.940 36.420 1083.200 36.680 ;
        RECT 2060.440 36.420 2060.700 36.680 ;
      LAYER met2 ;
        RECT 1077.420 1600.000 1077.700 1604.000 ;
        RECT 1077.480 1589.830 1077.620 1600.000 ;
        RECT 1077.420 1589.510 1077.680 1589.830 ;
        RECT 1082.940 1589.510 1083.200 1589.830 ;
        RECT 1083.000 36.710 1083.140 1589.510 ;
        RECT 1082.940 36.390 1083.200 36.710 ;
        RECT 2060.440 36.390 2060.700 36.710 ;
        RECT 2060.500 2.400 2060.640 36.390 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1083.830 1590.080 1084.150 1590.140 ;
        RECT 1089.810 1590.080 1090.130 1590.140 ;
        RECT 1083.830 1589.940 1090.130 1590.080 ;
        RECT 1083.830 1589.880 1084.150 1589.940 ;
        RECT 1089.810 1589.880 1090.130 1589.940 ;
        RECT 1089.810 36.960 1090.130 37.020 ;
        RECT 2078.350 36.960 2078.670 37.020 ;
        RECT 1089.810 36.820 2078.670 36.960 ;
        RECT 1089.810 36.760 1090.130 36.820 ;
        RECT 2078.350 36.760 2078.670 36.820 ;
      LAYER via ;
        RECT 1083.860 1589.880 1084.120 1590.140 ;
        RECT 1089.840 1589.880 1090.100 1590.140 ;
        RECT 1089.840 36.760 1090.100 37.020 ;
        RECT 2078.380 36.760 2078.640 37.020 ;
      LAYER met2 ;
        RECT 1083.860 1600.000 1084.140 1604.000 ;
        RECT 1083.920 1590.170 1084.060 1600.000 ;
        RECT 1083.860 1589.850 1084.120 1590.170 ;
        RECT 1089.840 1589.850 1090.100 1590.170 ;
        RECT 1089.900 37.050 1090.040 1589.850 ;
        RECT 1089.840 36.730 1090.100 37.050 ;
        RECT 2078.380 36.730 2078.640 37.050 ;
        RECT 2078.440 2.400 2078.580 36.730 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1090.730 1589.740 1091.050 1589.800 ;
        RECT 1096.710 1589.740 1097.030 1589.800 ;
        RECT 1090.730 1589.600 1097.030 1589.740 ;
        RECT 1090.730 1589.540 1091.050 1589.600 ;
        RECT 1096.710 1589.540 1097.030 1589.600 ;
        RECT 1096.710 37.300 1097.030 37.360 ;
        RECT 2095.830 37.300 2096.150 37.360 ;
        RECT 1096.710 37.160 2096.150 37.300 ;
        RECT 1096.710 37.100 1097.030 37.160 ;
        RECT 2095.830 37.100 2096.150 37.160 ;
      LAYER via ;
        RECT 1090.760 1589.540 1091.020 1589.800 ;
        RECT 1096.740 1589.540 1097.000 1589.800 ;
        RECT 1096.740 37.100 1097.000 37.360 ;
        RECT 2095.860 37.100 2096.120 37.360 ;
      LAYER met2 ;
        RECT 1090.760 1600.000 1091.040 1604.000 ;
        RECT 1090.820 1589.830 1090.960 1600.000 ;
        RECT 1090.760 1589.510 1091.020 1589.830 ;
        RECT 1096.740 1589.510 1097.000 1589.830 ;
        RECT 1096.800 37.390 1096.940 1589.510 ;
        RECT 1096.740 37.070 1097.000 37.390 ;
        RECT 2095.860 37.070 2096.120 37.390 ;
        RECT 2095.920 2.400 2096.060 37.070 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1097.630 1588.040 1097.950 1588.100 ;
        RECT 1103.610 1588.040 1103.930 1588.100 ;
        RECT 1097.630 1587.900 1103.930 1588.040 ;
        RECT 1097.630 1587.840 1097.950 1587.900 ;
        RECT 1103.610 1587.840 1103.930 1587.900 ;
        RECT 1103.610 37.640 1103.930 37.700 ;
        RECT 2113.770 37.640 2114.090 37.700 ;
        RECT 1103.610 37.500 2114.090 37.640 ;
        RECT 1103.610 37.440 1103.930 37.500 ;
        RECT 2113.770 37.440 2114.090 37.500 ;
      LAYER via ;
        RECT 1097.660 1587.840 1097.920 1588.100 ;
        RECT 1103.640 1587.840 1103.900 1588.100 ;
        RECT 1103.640 37.440 1103.900 37.700 ;
        RECT 2113.800 37.440 2114.060 37.700 ;
      LAYER met2 ;
        RECT 1097.660 1600.000 1097.940 1604.000 ;
        RECT 1097.720 1588.130 1097.860 1600.000 ;
        RECT 1097.660 1587.810 1097.920 1588.130 ;
        RECT 1103.640 1587.810 1103.900 1588.130 ;
        RECT 1103.700 37.730 1103.840 1587.810 ;
        RECT 1103.640 37.410 1103.900 37.730 ;
        RECT 2113.800 37.410 2114.060 37.730 ;
        RECT 2113.860 2.400 2114.000 37.410 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1104.070 1589.740 1104.390 1589.800 ;
        RECT 1110.050 1589.740 1110.370 1589.800 ;
        RECT 1104.070 1589.600 1110.370 1589.740 ;
        RECT 1104.070 1589.540 1104.390 1589.600 ;
        RECT 1110.050 1589.540 1110.370 1589.600 ;
        RECT 1110.050 41.380 1110.370 41.440 ;
        RECT 2131.710 41.380 2132.030 41.440 ;
        RECT 1110.050 41.240 2132.030 41.380 ;
        RECT 1110.050 41.180 1110.370 41.240 ;
        RECT 2131.710 41.180 2132.030 41.240 ;
      LAYER via ;
        RECT 1104.100 1589.540 1104.360 1589.800 ;
        RECT 1110.080 1589.540 1110.340 1589.800 ;
        RECT 1110.080 41.180 1110.340 41.440 ;
        RECT 2131.740 41.180 2132.000 41.440 ;
      LAYER met2 ;
        RECT 1104.100 1600.000 1104.380 1604.000 ;
        RECT 1104.160 1589.830 1104.300 1600.000 ;
        RECT 1104.100 1589.510 1104.360 1589.830 ;
        RECT 1110.080 1589.510 1110.340 1589.830 ;
        RECT 1110.140 41.470 1110.280 1589.510 ;
        RECT 1110.080 41.150 1110.340 41.470 ;
        RECT 2131.740 41.150 2132.000 41.470 ;
        RECT 2131.800 2.400 2131.940 41.150 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.970 1588.040 1111.290 1588.100 ;
        RECT 1117.410 1588.040 1117.730 1588.100 ;
        RECT 1110.970 1587.900 1117.730 1588.040 ;
        RECT 1110.970 1587.840 1111.290 1587.900 ;
        RECT 1117.410 1587.840 1117.730 1587.900 ;
        RECT 1117.410 41.040 1117.730 41.100 ;
        RECT 2149.650 41.040 2149.970 41.100 ;
        RECT 1117.410 40.900 2149.970 41.040 ;
        RECT 1117.410 40.840 1117.730 40.900 ;
        RECT 2149.650 40.840 2149.970 40.900 ;
      LAYER via ;
        RECT 1111.000 1587.840 1111.260 1588.100 ;
        RECT 1117.440 1587.840 1117.700 1588.100 ;
        RECT 1117.440 40.840 1117.700 41.100 ;
        RECT 2149.680 40.840 2149.940 41.100 ;
      LAYER met2 ;
        RECT 1111.000 1600.000 1111.280 1604.000 ;
        RECT 1111.060 1588.130 1111.200 1600.000 ;
        RECT 1111.000 1587.810 1111.260 1588.130 ;
        RECT 1117.440 1587.810 1117.700 1588.130 ;
        RECT 1117.500 41.130 1117.640 1587.810 ;
        RECT 1117.440 40.810 1117.700 41.130 ;
        RECT 2149.680 40.810 2149.940 41.130 ;
        RECT 2149.740 2.400 2149.880 40.810 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1117.870 1589.740 1118.190 1589.800 ;
        RECT 1124.310 1589.740 1124.630 1589.800 ;
        RECT 1117.870 1589.600 1124.630 1589.740 ;
        RECT 1117.870 1589.540 1118.190 1589.600 ;
        RECT 1124.310 1589.540 1124.630 1589.600 ;
        RECT 1124.310 40.700 1124.630 40.760 ;
        RECT 2167.590 40.700 2167.910 40.760 ;
        RECT 1124.310 40.560 2167.910 40.700 ;
        RECT 1124.310 40.500 1124.630 40.560 ;
        RECT 2167.590 40.500 2167.910 40.560 ;
      LAYER via ;
        RECT 1117.900 1589.540 1118.160 1589.800 ;
        RECT 1124.340 1589.540 1124.600 1589.800 ;
        RECT 1124.340 40.500 1124.600 40.760 ;
        RECT 2167.620 40.500 2167.880 40.760 ;
      LAYER met2 ;
        RECT 1117.900 1600.000 1118.180 1604.000 ;
        RECT 1117.960 1589.830 1118.100 1600.000 ;
        RECT 1117.900 1589.510 1118.160 1589.830 ;
        RECT 1124.340 1589.510 1124.600 1589.830 ;
        RECT 1124.400 40.790 1124.540 1589.510 ;
        RECT 1124.340 40.470 1124.600 40.790 ;
        RECT 2167.620 40.470 2167.880 40.790 ;
        RECT 2167.680 2.400 2167.820 40.470 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1123.850 40.360 1124.170 40.420 ;
        RECT 2185.070 40.360 2185.390 40.420 ;
        RECT 1123.850 40.220 2185.390 40.360 ;
        RECT 1123.850 40.160 1124.170 40.220 ;
        RECT 2185.070 40.160 2185.390 40.220 ;
      LAYER via ;
        RECT 1123.880 40.160 1124.140 40.420 ;
        RECT 2185.100 40.160 2185.360 40.420 ;
      LAYER met2 ;
        RECT 1124.340 1600.450 1124.620 1604.000 ;
        RECT 1123.940 1600.310 1124.620 1600.450 ;
        RECT 1123.940 40.450 1124.080 1600.310 ;
        RECT 1124.340 1600.000 1124.620 1600.310 ;
        RECT 1123.880 40.130 1124.140 40.450 ;
        RECT 2185.100 40.130 2185.360 40.450 ;
        RECT 2185.160 2.400 2185.300 40.130 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 40.020 1131.530 40.080 ;
        RECT 2203.010 40.020 2203.330 40.080 ;
        RECT 1131.210 39.880 2203.330 40.020 ;
        RECT 1131.210 39.820 1131.530 39.880 ;
        RECT 2203.010 39.820 2203.330 39.880 ;
      LAYER via ;
        RECT 1131.240 39.820 1131.500 40.080 ;
        RECT 2203.040 39.820 2203.300 40.080 ;
      LAYER met2 ;
        RECT 1131.240 1600.000 1131.520 1604.000 ;
        RECT 1131.300 40.110 1131.440 1600.000 ;
        RECT 1131.240 39.790 1131.500 40.110 ;
        RECT 2203.040 39.790 2203.300 40.110 ;
        RECT 2203.100 2.400 2203.240 39.790 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1138.110 39.680 1138.430 39.740 ;
        RECT 2220.950 39.680 2221.270 39.740 ;
        RECT 1138.110 39.540 2221.270 39.680 ;
        RECT 1138.110 39.480 1138.430 39.540 ;
        RECT 2220.950 39.480 2221.270 39.540 ;
      LAYER via ;
        RECT 1138.140 39.480 1138.400 39.740 ;
        RECT 2220.980 39.480 2221.240 39.740 ;
      LAYER met2 ;
        RECT 1138.140 1600.000 1138.420 1604.000 ;
        RECT 1138.200 39.770 1138.340 1600.000 ;
        RECT 1138.140 39.450 1138.400 39.770 ;
        RECT 2220.980 39.450 2221.240 39.770 ;
        RECT 2221.040 2.400 2221.180 39.450 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 714.065 1593.325 715.155 1593.495 ;
        RECT 714.065 1592.985 714.235 1593.325 ;
        RECT 728.325 1588.225 728.495 1593.495 ;
      LAYER mcon ;
        RECT 714.985 1593.325 715.155 1593.495 ;
        RECT 728.325 1593.325 728.495 1593.495 ;
      LAYER met1 ;
        RECT 714.925 1593.480 715.215 1593.525 ;
        RECT 728.265 1593.480 728.555 1593.525 ;
        RECT 714.925 1593.340 728.555 1593.480 ;
        RECT 714.925 1593.295 715.215 1593.340 ;
        RECT 728.265 1593.295 728.555 1593.340 ;
        RECT 592.550 1593.140 592.870 1593.200 ;
        RECT 714.005 1593.140 714.295 1593.185 ;
        RECT 592.550 1593.000 714.295 1593.140 ;
        RECT 592.550 1592.940 592.870 1593.000 ;
        RECT 714.005 1592.955 714.295 1593.000 ;
        RECT 761.370 1588.720 761.690 1588.780 ;
        RECT 738.920 1588.580 761.690 1588.720 ;
        RECT 728.265 1588.380 728.555 1588.425 ;
        RECT 738.920 1588.380 739.060 1588.580 ;
        RECT 761.370 1588.520 761.690 1588.580 ;
        RECT 728.265 1588.240 739.060 1588.380 ;
        RECT 728.265 1588.195 728.555 1588.240 ;
        RECT 762.290 20.640 762.610 20.700 ;
        RECT 775.630 20.640 775.950 20.700 ;
        RECT 762.290 20.500 775.950 20.640 ;
        RECT 762.290 20.440 762.610 20.500 ;
        RECT 775.630 20.440 775.950 20.500 ;
      LAYER via ;
        RECT 592.580 1592.940 592.840 1593.200 ;
        RECT 761.400 1588.520 761.660 1588.780 ;
        RECT 762.320 20.440 762.580 20.700 ;
        RECT 775.660 20.440 775.920 20.700 ;
      LAYER met2 ;
        RECT 592.580 1600.000 592.860 1604.000 ;
        RECT 592.640 1593.230 592.780 1600.000 ;
        RECT 592.580 1592.910 592.840 1593.230 ;
        RECT 761.460 1588.810 762.520 1588.890 ;
        RECT 761.400 1588.750 762.520 1588.810 ;
        RECT 761.400 1588.490 761.660 1588.750 ;
        RECT 762.380 20.730 762.520 1588.750 ;
        RECT 762.320 20.410 762.580 20.730 ;
        RECT 775.660 20.410 775.920 20.730 ;
        RECT 775.720 2.400 775.860 20.410 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.010 39.340 1145.330 39.400 ;
        RECT 2238.890 39.340 2239.210 39.400 ;
        RECT 1145.010 39.200 2239.210 39.340 ;
        RECT 1145.010 39.140 1145.330 39.200 ;
        RECT 2238.890 39.140 2239.210 39.200 ;
      LAYER via ;
        RECT 1145.040 39.140 1145.300 39.400 ;
        RECT 2238.920 39.140 2239.180 39.400 ;
      LAYER met2 ;
        RECT 1144.580 1600.450 1144.860 1604.000 ;
        RECT 1144.580 1600.310 1145.240 1600.450 ;
        RECT 1144.580 1600.000 1144.860 1600.310 ;
        RECT 1145.100 39.430 1145.240 1600.310 ;
        RECT 1145.040 39.110 1145.300 39.430 ;
        RECT 2238.920 39.110 2239.180 39.430 ;
        RECT 2238.980 2.400 2239.120 39.110 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1151.450 39.000 1151.770 39.060 ;
        RECT 2256.830 39.000 2257.150 39.060 ;
        RECT 1151.450 38.860 2257.150 39.000 ;
        RECT 1151.450 38.800 1151.770 38.860 ;
        RECT 2256.830 38.800 2257.150 38.860 ;
      LAYER via ;
        RECT 1151.480 38.800 1151.740 39.060 ;
        RECT 2256.860 38.800 2257.120 39.060 ;
      LAYER met2 ;
        RECT 1151.480 1600.000 1151.760 1604.000 ;
        RECT 1151.540 39.090 1151.680 1600.000 ;
        RECT 1151.480 38.770 1151.740 39.090 ;
        RECT 2256.860 38.770 2257.120 39.090 ;
        RECT 2256.920 7.210 2257.060 38.770 ;
        RECT 2256.460 7.070 2257.060 7.210 ;
        RECT 2256.460 2.400 2256.600 7.070 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1158.810 38.660 1159.130 38.720 ;
        RECT 2274.310 38.660 2274.630 38.720 ;
        RECT 1158.810 38.520 2274.630 38.660 ;
        RECT 1158.810 38.460 1159.130 38.520 ;
        RECT 2274.310 38.460 2274.630 38.520 ;
      LAYER via ;
        RECT 1158.840 38.460 1159.100 38.720 ;
        RECT 2274.340 38.460 2274.600 38.720 ;
      LAYER met2 ;
        RECT 1158.380 1600.450 1158.660 1604.000 ;
        RECT 1158.380 1600.310 1159.040 1600.450 ;
        RECT 1158.380 1600.000 1158.660 1600.310 ;
        RECT 1158.900 38.750 1159.040 1600.310 ;
        RECT 1158.840 38.430 1159.100 38.750 ;
        RECT 2274.340 38.430 2274.600 38.750 ;
        RECT 2274.400 2.400 2274.540 38.430 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1165.250 38.320 1165.570 38.380 ;
        RECT 2292.250 38.320 2292.570 38.380 ;
        RECT 1165.250 38.180 2292.570 38.320 ;
        RECT 1165.250 38.120 1165.570 38.180 ;
        RECT 2292.250 38.120 2292.570 38.180 ;
      LAYER via ;
        RECT 1165.280 38.120 1165.540 38.380 ;
        RECT 2292.280 38.120 2292.540 38.380 ;
      LAYER met2 ;
        RECT 1164.820 1600.450 1165.100 1604.000 ;
        RECT 1164.820 1600.310 1165.480 1600.450 ;
        RECT 1164.820 1600.000 1165.100 1600.310 ;
        RECT 1165.340 38.410 1165.480 1600.310 ;
        RECT 1165.280 38.090 1165.540 38.410 ;
        RECT 2292.280 38.090 2292.540 38.410 ;
        RECT 2292.340 2.400 2292.480 38.090 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1172.610 37.980 1172.930 38.040 ;
        RECT 2310.190 37.980 2310.510 38.040 ;
        RECT 1172.610 37.840 2310.510 37.980 ;
        RECT 1172.610 37.780 1172.930 37.840 ;
        RECT 2310.190 37.780 2310.510 37.840 ;
      LAYER via ;
        RECT 1172.640 37.780 1172.900 38.040 ;
        RECT 2310.220 37.780 2310.480 38.040 ;
      LAYER met2 ;
        RECT 1171.720 1600.450 1172.000 1604.000 ;
        RECT 1171.720 1600.310 1172.840 1600.450 ;
        RECT 1171.720 1600.000 1172.000 1600.310 ;
        RECT 1172.700 38.070 1172.840 1600.310 ;
        RECT 1172.640 37.750 1172.900 38.070 ;
        RECT 2310.220 37.750 2310.480 38.070 ;
        RECT 2310.280 2.400 2310.420 37.750 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1178.160 1600.450 1178.440 1604.000 ;
        RECT 1178.160 1600.310 1179.280 1600.450 ;
        RECT 1178.160 1600.000 1178.440 1600.310 ;
        RECT 1179.140 41.325 1179.280 1600.310 ;
        RECT 1179.070 40.955 1179.350 41.325 ;
        RECT 2328.150 40.955 2328.430 41.325 ;
        RECT 2328.220 2.400 2328.360 40.955 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
      LAYER via2 ;
        RECT 1179.070 41.000 1179.350 41.280 ;
        RECT 2328.150 41.000 2328.430 41.280 ;
      LAYER met3 ;
        RECT 1179.045 41.290 1179.375 41.305 ;
        RECT 2328.125 41.290 2328.455 41.305 ;
        RECT 1179.045 40.990 2328.455 41.290 ;
        RECT 1179.045 40.975 1179.375 40.990 ;
        RECT 2328.125 40.975 2328.455 40.990 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.060 1600.450 1185.340 1604.000 ;
        RECT 1185.060 1600.310 1186.640 1600.450 ;
        RECT 1185.060 1600.000 1185.340 1600.310 ;
        RECT 1186.500 40.645 1186.640 1600.310 ;
        RECT 1186.430 40.275 1186.710 40.645 ;
        RECT 2345.630 40.275 2345.910 40.645 ;
        RECT 2345.700 2.400 2345.840 40.275 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
      LAYER via2 ;
        RECT 1186.430 40.320 1186.710 40.600 ;
        RECT 2345.630 40.320 2345.910 40.600 ;
      LAYER met3 ;
        RECT 1186.405 40.610 1186.735 40.625 ;
        RECT 2345.605 40.610 2345.935 40.625 ;
        RECT 1186.405 40.310 2345.935 40.610 ;
        RECT 1186.405 40.295 1186.735 40.310 ;
        RECT 2345.605 40.295 2345.935 40.310 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1191.960 1600.450 1192.240 1604.000 ;
        RECT 1191.960 1600.310 1193.080 1600.450 ;
        RECT 1191.960 1600.000 1192.240 1600.310 ;
        RECT 1192.940 39.965 1193.080 1600.310 ;
        RECT 1192.870 39.595 1193.150 39.965 ;
        RECT 2363.570 39.595 2363.850 39.965 ;
        RECT 2363.640 2.400 2363.780 39.595 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
      LAYER via2 ;
        RECT 1192.870 39.640 1193.150 39.920 ;
        RECT 2363.570 39.640 2363.850 39.920 ;
      LAYER met3 ;
        RECT 1192.845 39.930 1193.175 39.945 ;
        RECT 2363.545 39.930 2363.875 39.945 ;
        RECT 1192.845 39.630 2363.875 39.930 ;
        RECT 1192.845 39.615 1193.175 39.630 ;
        RECT 2363.545 39.615 2363.875 39.630 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1198.400 1600.450 1198.680 1604.000 ;
        RECT 1198.400 1600.310 1200.440 1600.450 ;
        RECT 1198.400 1600.000 1198.680 1600.310 ;
        RECT 1200.300 39.285 1200.440 1600.310 ;
        RECT 1200.230 38.915 1200.510 39.285 ;
        RECT 2381.510 38.915 2381.790 39.285 ;
        RECT 2381.580 2.400 2381.720 38.915 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
      LAYER via2 ;
        RECT 1200.230 38.960 1200.510 39.240 ;
        RECT 2381.510 38.960 2381.790 39.240 ;
      LAYER met3 ;
        RECT 1200.205 39.250 1200.535 39.265 ;
        RECT 2381.485 39.250 2381.815 39.265 ;
        RECT 1200.205 38.950 2381.815 39.250 ;
        RECT 1200.205 38.935 1200.535 38.950 ;
        RECT 2381.485 38.935 2381.815 38.950 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1205.300 1600.450 1205.580 1604.000 ;
        RECT 1205.300 1600.310 1206.880 1600.450 ;
        RECT 1205.300 1600.000 1205.580 1600.310 ;
        RECT 1206.740 38.605 1206.880 1600.310 ;
        RECT 1206.670 38.235 1206.950 38.605 ;
        RECT 2399.450 38.235 2399.730 38.605 ;
        RECT 2399.520 2.400 2399.660 38.235 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
      LAYER via2 ;
        RECT 1206.670 38.280 1206.950 38.560 ;
        RECT 2399.450 38.280 2399.730 38.560 ;
      LAYER met3 ;
        RECT 1206.645 38.570 1206.975 38.585 ;
        RECT 2399.425 38.570 2399.755 38.585 ;
        RECT 1206.645 38.270 2399.755 38.570 ;
        RECT 1206.645 38.255 1206.975 38.270 ;
        RECT 2399.425 38.255 2399.755 38.270 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 599.020 1600.450 599.300 1604.000 ;
        RECT 599.020 1600.310 600.140 1600.450 ;
        RECT 599.020 1600.000 599.300 1600.310 ;
        RECT 600.000 17.525 600.140 1600.310 ;
        RECT 599.930 17.155 600.210 17.525 ;
        RECT 793.590 17.155 793.870 17.525 ;
        RECT 793.660 2.400 793.800 17.155 ;
        RECT 793.450 -4.800 794.010 2.400 ;
      LAYER via2 ;
        RECT 599.930 17.200 600.210 17.480 ;
        RECT 793.590 17.200 793.870 17.480 ;
      LAYER met3 ;
        RECT 599.905 17.490 600.235 17.505 ;
        RECT 793.565 17.490 793.895 17.505 ;
        RECT 599.905 17.190 793.895 17.490 ;
        RECT 599.905 17.175 600.235 17.190 ;
        RECT 793.565 17.175 793.895 17.190 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 603.665 16.745 603.835 18.615 ;
      LAYER mcon ;
        RECT 603.665 18.445 603.835 18.615 ;
      LAYER met1 ;
        RECT 541.030 1588.720 541.350 1588.780 ;
        RECT 544.710 1588.720 545.030 1588.780 ;
        RECT 541.030 1588.580 545.030 1588.720 ;
        RECT 541.030 1588.520 541.350 1588.580 ;
        RECT 544.710 1588.520 545.030 1588.580 ;
        RECT 544.710 18.600 545.030 18.660 ;
        RECT 603.605 18.600 603.895 18.645 ;
        RECT 544.710 18.460 603.895 18.600 ;
        RECT 544.710 18.400 545.030 18.460 ;
        RECT 603.605 18.415 603.895 18.460 ;
        RECT 603.605 16.900 603.895 16.945 ;
        RECT 639.010 16.900 639.330 16.960 ;
        RECT 603.605 16.760 639.330 16.900 ;
        RECT 603.605 16.715 603.895 16.760 ;
        RECT 639.010 16.700 639.330 16.760 ;
      LAYER via ;
        RECT 541.060 1588.520 541.320 1588.780 ;
        RECT 544.740 1588.520 545.000 1588.780 ;
        RECT 544.740 18.400 545.000 18.660 ;
        RECT 639.040 16.700 639.300 16.960 ;
      LAYER met2 ;
        RECT 541.060 1600.000 541.340 1604.000 ;
        RECT 541.120 1588.810 541.260 1600.000 ;
        RECT 541.060 1588.490 541.320 1588.810 ;
        RECT 544.740 1588.490 545.000 1588.810 ;
        RECT 544.800 18.690 544.940 1588.490 ;
        RECT 544.740 18.370 545.000 18.690 ;
        RECT 639.040 16.670 639.300 16.990 ;
        RECT 639.100 2.400 639.240 16.670 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1214.040 1600.000 1214.320 1604.000 ;
        RECT 1214.100 37.925 1214.240 1600.000 ;
        RECT 1214.030 37.555 1214.310 37.925 ;
        RECT 2422.910 37.555 2423.190 37.925 ;
        RECT 2422.980 2.400 2423.120 37.555 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
      LAYER via2 ;
        RECT 1214.030 37.600 1214.310 37.880 ;
        RECT 2422.910 37.600 2423.190 37.880 ;
      LAYER met3 ;
        RECT 1214.005 37.890 1214.335 37.905 ;
        RECT 2422.885 37.890 2423.215 37.905 ;
        RECT 1214.005 37.590 2423.215 37.890 ;
        RECT 1214.005 37.575 1214.335 37.590 ;
        RECT 2422.885 37.575 2423.215 37.590 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1220.450 72.660 1220.770 72.720 ;
        RECT 2435.770 72.660 2436.090 72.720 ;
        RECT 1220.450 72.520 2436.090 72.660 ;
        RECT 1220.450 72.460 1220.770 72.520 ;
        RECT 2435.770 72.460 2436.090 72.520 ;
      LAYER via ;
        RECT 1220.480 72.460 1220.740 72.720 ;
        RECT 2435.800 72.460 2436.060 72.720 ;
      LAYER met2 ;
        RECT 1220.940 1600.450 1221.220 1604.000 ;
        RECT 1220.540 1600.310 1221.220 1600.450 ;
        RECT 1220.540 72.750 1220.680 1600.310 ;
        RECT 1220.940 1600.000 1221.220 1600.310 ;
        RECT 1220.480 72.430 1220.740 72.750 ;
        RECT 2435.800 72.430 2436.060 72.750 ;
        RECT 2435.860 17.410 2436.000 72.430 ;
        RECT 2435.860 17.270 2441.060 17.410 ;
        RECT 2440.920 2.400 2441.060 17.270 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.350 72.320 1227.670 72.380 ;
        RECT 2456.470 72.320 2456.790 72.380 ;
        RECT 1227.350 72.180 2456.790 72.320 ;
        RECT 1227.350 72.120 1227.670 72.180 ;
        RECT 2456.470 72.120 2456.790 72.180 ;
      LAYER via ;
        RECT 1227.380 72.120 1227.640 72.380 ;
        RECT 2456.500 72.120 2456.760 72.380 ;
      LAYER met2 ;
        RECT 1227.840 1600.450 1228.120 1604.000 ;
        RECT 1227.440 1600.310 1228.120 1600.450 ;
        RECT 1227.440 72.410 1227.580 1600.310 ;
        RECT 1227.840 1600.000 1228.120 1600.310 ;
        RECT 1227.380 72.090 1227.640 72.410 ;
        RECT 2456.500 72.090 2456.760 72.410 ;
        RECT 2456.560 3.130 2456.700 72.090 ;
        RECT 2456.560 2.990 2458.540 3.130 ;
        RECT 2458.400 2.960 2458.540 2.990 ;
        RECT 2458.400 2.820 2459.000 2.960 ;
        RECT 2458.860 2.400 2459.000 2.820 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1234.250 82.180 1234.570 82.240 ;
        RECT 2470.270 82.180 2470.590 82.240 ;
        RECT 1234.250 82.040 2470.590 82.180 ;
        RECT 1234.250 81.980 1234.570 82.040 ;
        RECT 2470.270 81.980 2470.590 82.040 ;
        RECT 2470.270 17.240 2470.590 17.300 ;
        RECT 2476.710 17.240 2477.030 17.300 ;
        RECT 2470.270 17.100 2477.030 17.240 ;
        RECT 2470.270 17.040 2470.590 17.100 ;
        RECT 2476.710 17.040 2477.030 17.100 ;
      LAYER via ;
        RECT 1234.280 81.980 1234.540 82.240 ;
        RECT 2470.300 81.980 2470.560 82.240 ;
        RECT 2470.300 17.040 2470.560 17.300 ;
        RECT 2476.740 17.040 2477.000 17.300 ;
      LAYER met2 ;
        RECT 1234.280 1600.000 1234.560 1604.000 ;
        RECT 1234.340 82.270 1234.480 1600.000 ;
        RECT 1234.280 81.950 1234.540 82.270 ;
        RECT 2470.300 81.950 2470.560 82.270 ;
        RECT 2470.360 17.330 2470.500 81.950 ;
        RECT 2470.300 17.010 2470.560 17.330 ;
        RECT 2476.740 17.010 2477.000 17.330 ;
        RECT 2476.800 2.400 2476.940 17.010 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1241.610 43.420 1241.930 43.480 ;
        RECT 2494.650 43.420 2494.970 43.480 ;
        RECT 1241.610 43.280 2494.970 43.420 ;
        RECT 1241.610 43.220 1241.930 43.280 ;
        RECT 2494.650 43.220 2494.970 43.280 ;
      LAYER via ;
        RECT 1241.640 43.220 1241.900 43.480 ;
        RECT 2494.680 43.220 2494.940 43.480 ;
      LAYER met2 ;
        RECT 1241.180 1600.450 1241.460 1604.000 ;
        RECT 1241.180 1600.310 1241.840 1600.450 ;
        RECT 1241.180 1600.000 1241.460 1600.310 ;
        RECT 1241.700 43.510 1241.840 1600.310 ;
        RECT 1241.640 43.190 1241.900 43.510 ;
        RECT 2494.680 43.190 2494.940 43.510 ;
        RECT 2494.740 2.400 2494.880 43.190 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.510 43.760 1248.830 43.820 ;
        RECT 2512.130 43.760 2512.450 43.820 ;
        RECT 1248.510 43.620 2512.450 43.760 ;
        RECT 1248.510 43.560 1248.830 43.620 ;
        RECT 2512.130 43.560 2512.450 43.620 ;
      LAYER via ;
        RECT 1248.540 43.560 1248.800 43.820 ;
        RECT 2512.160 43.560 2512.420 43.820 ;
      LAYER met2 ;
        RECT 1248.080 1600.450 1248.360 1604.000 ;
        RECT 1248.080 1600.310 1248.740 1600.450 ;
        RECT 1248.080 1600.000 1248.360 1600.310 ;
        RECT 1248.600 43.850 1248.740 1600.310 ;
        RECT 1248.540 43.530 1248.800 43.850 ;
        RECT 2512.160 43.530 2512.420 43.850 ;
        RECT 2512.220 2.400 2512.360 43.530 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1255.410 44.100 1255.730 44.160 ;
        RECT 2530.070 44.100 2530.390 44.160 ;
        RECT 1255.410 43.960 2530.390 44.100 ;
        RECT 1255.410 43.900 1255.730 43.960 ;
        RECT 2530.070 43.900 2530.390 43.960 ;
      LAYER via ;
        RECT 1255.440 43.900 1255.700 44.160 ;
        RECT 2530.100 43.900 2530.360 44.160 ;
      LAYER met2 ;
        RECT 1254.520 1600.450 1254.800 1604.000 ;
        RECT 1254.520 1600.310 1255.640 1600.450 ;
        RECT 1254.520 1600.000 1254.800 1600.310 ;
        RECT 1255.500 44.190 1255.640 1600.310 ;
        RECT 1255.440 43.870 1255.700 44.190 ;
        RECT 2530.100 43.870 2530.360 44.190 ;
        RECT 2530.160 2.400 2530.300 43.870 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1262.310 44.440 1262.630 44.500 ;
        RECT 2548.010 44.440 2548.330 44.500 ;
        RECT 1262.310 44.300 2548.330 44.440 ;
        RECT 1262.310 44.240 1262.630 44.300 ;
        RECT 2548.010 44.240 2548.330 44.300 ;
      LAYER via ;
        RECT 1262.340 44.240 1262.600 44.500 ;
        RECT 2548.040 44.240 2548.300 44.500 ;
      LAYER met2 ;
        RECT 1261.420 1600.450 1261.700 1604.000 ;
        RECT 1261.420 1600.310 1262.540 1600.450 ;
        RECT 1261.420 1600.000 1261.700 1600.310 ;
        RECT 1262.400 44.530 1262.540 1600.310 ;
        RECT 1262.340 44.210 1262.600 44.530 ;
        RECT 2548.040 44.210 2548.300 44.530 ;
        RECT 2548.100 2.400 2548.240 44.210 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1268.750 48.180 1269.070 48.240 ;
        RECT 2565.950 48.180 2566.270 48.240 ;
        RECT 1268.750 48.040 2566.270 48.180 ;
        RECT 1268.750 47.980 1269.070 48.040 ;
        RECT 2565.950 47.980 2566.270 48.040 ;
      LAYER via ;
        RECT 1268.780 47.980 1269.040 48.240 ;
        RECT 2565.980 47.980 2566.240 48.240 ;
      LAYER met2 ;
        RECT 1268.320 1600.450 1268.600 1604.000 ;
        RECT 1268.320 1600.310 1268.980 1600.450 ;
        RECT 1268.320 1600.000 1268.600 1600.310 ;
        RECT 1268.840 48.270 1268.980 1600.310 ;
        RECT 1268.780 47.950 1269.040 48.270 ;
        RECT 2565.980 47.950 2566.240 48.270 ;
        RECT 2566.040 2.400 2566.180 47.950 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1275.650 47.840 1275.970 47.900 ;
        RECT 2583.890 47.840 2584.210 47.900 ;
        RECT 1275.650 47.700 2584.210 47.840 ;
        RECT 1275.650 47.640 1275.970 47.700 ;
        RECT 2583.890 47.640 2584.210 47.700 ;
      LAYER via ;
        RECT 1275.680 47.640 1275.940 47.900 ;
        RECT 2583.920 47.640 2584.180 47.900 ;
      LAYER met2 ;
        RECT 1274.760 1600.450 1275.040 1604.000 ;
        RECT 1274.760 1600.310 1275.880 1600.450 ;
        RECT 1274.760 1600.000 1275.040 1600.310 ;
        RECT 1275.740 47.930 1275.880 1600.310 ;
        RECT 1275.680 47.610 1275.940 47.930 ;
        RECT 2583.920 47.610 2584.180 47.930 ;
        RECT 2583.980 2.400 2584.120 47.610 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 608.190 1587.360 608.510 1587.420 ;
        RECT 613.250 1587.360 613.570 1587.420 ;
        RECT 608.190 1587.220 613.570 1587.360 ;
        RECT 608.190 1587.160 608.510 1587.220 ;
        RECT 613.250 1587.160 613.570 1587.220 ;
        RECT 613.250 30.160 613.570 30.220 ;
        RECT 817.490 30.160 817.810 30.220 ;
        RECT 613.250 30.020 817.810 30.160 ;
        RECT 613.250 29.960 613.570 30.020 ;
        RECT 817.490 29.960 817.810 30.020 ;
      LAYER via ;
        RECT 608.220 1587.160 608.480 1587.420 ;
        RECT 613.280 1587.160 613.540 1587.420 ;
        RECT 613.280 29.960 613.540 30.220 ;
        RECT 817.520 29.960 817.780 30.220 ;
      LAYER met2 ;
        RECT 608.220 1600.000 608.500 1604.000 ;
        RECT 608.280 1587.450 608.420 1600.000 ;
        RECT 608.220 1587.130 608.480 1587.450 ;
        RECT 613.280 1587.130 613.540 1587.450 ;
        RECT 613.340 30.250 613.480 1587.130 ;
        RECT 613.280 29.930 613.540 30.250 ;
        RECT 817.520 29.930 817.780 30.250 ;
        RECT 817.580 2.400 817.720 29.930 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1282.550 47.500 1282.870 47.560 ;
        RECT 2601.830 47.500 2602.150 47.560 ;
        RECT 1282.550 47.360 2602.150 47.500 ;
        RECT 1282.550 47.300 1282.870 47.360 ;
        RECT 2601.830 47.300 2602.150 47.360 ;
      LAYER via ;
        RECT 1282.580 47.300 1282.840 47.560 ;
        RECT 2601.860 47.300 2602.120 47.560 ;
      LAYER met2 ;
        RECT 1281.660 1600.450 1281.940 1604.000 ;
        RECT 1281.660 1600.310 1282.780 1600.450 ;
        RECT 1281.660 1600.000 1281.940 1600.310 ;
        RECT 1282.640 47.590 1282.780 1600.310 ;
        RECT 1282.580 47.270 1282.840 47.590 ;
        RECT 2601.860 47.270 2602.120 47.590 ;
        RECT 2601.920 7.210 2602.060 47.270 ;
        RECT 2601.460 7.070 2602.060 7.210 ;
        RECT 2601.460 2.400 2601.600 7.070 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1289.450 47.160 1289.770 47.220 ;
        RECT 2619.310 47.160 2619.630 47.220 ;
        RECT 1289.450 47.020 2619.630 47.160 ;
        RECT 1289.450 46.960 1289.770 47.020 ;
        RECT 2619.310 46.960 2619.630 47.020 ;
      LAYER via ;
        RECT 1289.480 46.960 1289.740 47.220 ;
        RECT 2619.340 46.960 2619.600 47.220 ;
      LAYER met2 ;
        RECT 1288.560 1600.450 1288.840 1604.000 ;
        RECT 1288.560 1600.310 1289.680 1600.450 ;
        RECT 1288.560 1600.000 1288.840 1600.310 ;
        RECT 1289.540 47.250 1289.680 1600.310 ;
        RECT 1289.480 46.930 1289.740 47.250 ;
        RECT 2619.340 46.930 2619.600 47.250 ;
        RECT 2619.400 2.400 2619.540 46.930 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1296.350 46.820 1296.670 46.880 ;
        RECT 2637.250 46.820 2637.570 46.880 ;
        RECT 1296.350 46.680 2637.570 46.820 ;
        RECT 1296.350 46.620 1296.670 46.680 ;
        RECT 2637.250 46.620 2637.570 46.680 ;
      LAYER via ;
        RECT 1296.380 46.620 1296.640 46.880 ;
        RECT 2637.280 46.620 2637.540 46.880 ;
      LAYER met2 ;
        RECT 1295.000 1600.450 1295.280 1604.000 ;
        RECT 1295.000 1600.310 1296.580 1600.450 ;
        RECT 1295.000 1600.000 1295.280 1600.310 ;
        RECT 1296.440 46.910 1296.580 1600.310 ;
        RECT 1296.380 46.590 1296.640 46.910 ;
        RECT 2637.280 46.590 2637.540 46.910 ;
        RECT 2637.340 2.400 2637.480 46.590 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1301.900 1600.450 1302.180 1604.000 ;
        RECT 1301.900 1600.310 1303.480 1600.450 ;
        RECT 1301.900 1600.000 1302.180 1600.310 ;
        RECT 1303.340 48.125 1303.480 1600.310 ;
        RECT 1303.270 47.755 1303.550 48.125 ;
        RECT 2655.210 47.755 2655.490 48.125 ;
        RECT 2655.280 2.400 2655.420 47.755 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
      LAYER via2 ;
        RECT 1303.270 47.800 1303.550 48.080 ;
        RECT 2655.210 47.800 2655.490 48.080 ;
      LAYER met3 ;
        RECT 1303.245 48.090 1303.575 48.105 ;
        RECT 2655.185 48.090 2655.515 48.105 ;
        RECT 1303.245 47.790 2655.515 48.090 ;
        RECT 1303.245 47.775 1303.575 47.790 ;
        RECT 2655.185 47.775 2655.515 47.790 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1310.150 46.480 1310.470 46.540 ;
        RECT 2672.670 46.480 2672.990 46.540 ;
        RECT 1310.150 46.340 2672.990 46.480 ;
        RECT 1310.150 46.280 1310.470 46.340 ;
        RECT 2672.670 46.280 2672.990 46.340 ;
      LAYER via ;
        RECT 1310.180 46.280 1310.440 46.540 ;
        RECT 2672.700 46.280 2672.960 46.540 ;
      LAYER met2 ;
        RECT 1308.340 1600.450 1308.620 1604.000 ;
        RECT 1308.340 1600.310 1310.380 1600.450 ;
        RECT 1308.340 1600.000 1308.620 1600.310 ;
        RECT 1310.240 46.570 1310.380 1600.310 ;
        RECT 1310.180 46.250 1310.440 46.570 ;
        RECT 2672.700 46.250 2672.960 46.570 ;
        RECT 2672.760 2.400 2672.900 46.250 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1315.240 1600.450 1315.520 1604.000 ;
        RECT 1315.240 1600.310 1317.280 1600.450 ;
        RECT 1315.240 1600.000 1315.520 1600.310 ;
        RECT 1317.140 47.445 1317.280 1600.310 ;
        RECT 1317.070 47.075 1317.350 47.445 ;
        RECT 2690.630 47.075 2690.910 47.445 ;
        RECT 2690.700 2.400 2690.840 47.075 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
      LAYER via2 ;
        RECT 1317.070 47.120 1317.350 47.400 ;
        RECT 2690.630 47.120 2690.910 47.400 ;
      LAYER met3 ;
        RECT 1317.045 47.410 1317.375 47.425 ;
        RECT 2690.605 47.410 2690.935 47.425 ;
        RECT 1317.045 47.110 2690.935 47.410 ;
        RECT 1317.045 47.095 1317.375 47.110 ;
        RECT 2690.605 47.095 2690.935 47.110 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1323.950 46.140 1324.270 46.200 ;
        RECT 2708.550 46.140 2708.870 46.200 ;
        RECT 1323.950 46.000 2708.870 46.140 ;
        RECT 1323.950 45.940 1324.270 46.000 ;
        RECT 2708.550 45.940 2708.870 46.000 ;
      LAYER via ;
        RECT 1323.980 45.940 1324.240 46.200 ;
        RECT 2708.580 45.940 2708.840 46.200 ;
      LAYER met2 ;
        RECT 1322.140 1600.450 1322.420 1604.000 ;
        RECT 1322.140 1600.310 1324.180 1600.450 ;
        RECT 1322.140 1600.000 1322.420 1600.310 ;
        RECT 1324.040 46.230 1324.180 1600.310 ;
        RECT 1323.980 45.910 1324.240 46.230 ;
        RECT 2708.580 45.910 2708.840 46.230 ;
        RECT 2708.640 2.400 2708.780 45.910 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1328.580 1600.450 1328.860 1604.000 ;
        RECT 1328.580 1600.310 1330.620 1600.450 ;
        RECT 1328.580 1600.000 1328.860 1600.310 ;
        RECT 1330.480 72.605 1330.620 1600.310 ;
        RECT 1330.410 72.235 1330.690 72.605 ;
        RECT 2725.590 72.235 2725.870 72.605 ;
        RECT 2725.660 3.130 2725.800 72.235 ;
        RECT 2725.660 2.990 2726.720 3.130 ;
        RECT 2726.580 2.400 2726.720 2.990 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
      LAYER via2 ;
        RECT 1330.410 72.280 1330.690 72.560 ;
        RECT 2725.590 72.280 2725.870 72.560 ;
      LAYER met3 ;
        RECT 1330.385 72.570 1330.715 72.585 ;
        RECT 2725.565 72.570 2725.895 72.585 ;
        RECT 1330.385 72.270 2725.895 72.570 ;
        RECT 1330.385 72.255 1330.715 72.270 ;
        RECT 2725.565 72.255 2725.895 72.270 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1335.450 1590.760 1335.770 1590.820 ;
        RECT 1337.750 1590.760 1338.070 1590.820 ;
        RECT 1335.450 1590.620 1338.070 1590.760 ;
        RECT 1335.450 1590.560 1335.770 1590.620 ;
        RECT 1337.750 1590.560 1338.070 1590.620 ;
      LAYER via ;
        RECT 1335.480 1590.560 1335.740 1590.820 ;
        RECT 1337.780 1590.560 1338.040 1590.820 ;
      LAYER met2 ;
        RECT 1335.480 1600.000 1335.760 1604.000 ;
        RECT 1335.540 1590.850 1335.680 1600.000 ;
        RECT 1335.480 1590.530 1335.740 1590.850 ;
        RECT 1337.780 1590.530 1338.040 1590.850 ;
        RECT 1337.840 46.765 1337.980 1590.530 ;
        RECT 1337.770 46.395 1338.050 46.765 ;
        RECT 2744.450 46.395 2744.730 46.765 ;
        RECT 2744.520 2.400 2744.660 46.395 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
      LAYER via2 ;
        RECT 1337.770 46.440 1338.050 46.720 ;
        RECT 2744.450 46.440 2744.730 46.720 ;
      LAYER met3 ;
        RECT 1337.745 46.730 1338.075 46.745 ;
        RECT 2744.425 46.730 2744.755 46.745 ;
        RECT 1337.745 46.430 2744.755 46.730 ;
        RECT 1337.745 46.415 1338.075 46.430 ;
        RECT 2744.425 46.415 2744.755 46.430 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1342.350 1590.420 1342.670 1590.480 ;
        RECT 1344.650 1590.420 1344.970 1590.480 ;
        RECT 1342.350 1590.280 1344.970 1590.420 ;
        RECT 1342.350 1590.220 1342.670 1590.280 ;
        RECT 1344.650 1590.220 1344.970 1590.280 ;
        RECT 1344.650 45.800 1344.970 45.860 ;
        RECT 2761.910 45.800 2762.230 45.860 ;
        RECT 1344.650 45.660 2762.230 45.800 ;
        RECT 1344.650 45.600 1344.970 45.660 ;
        RECT 2761.910 45.600 2762.230 45.660 ;
      LAYER via ;
        RECT 1342.380 1590.220 1342.640 1590.480 ;
        RECT 1344.680 1590.220 1344.940 1590.480 ;
        RECT 1344.680 45.600 1344.940 45.860 ;
        RECT 2761.940 45.600 2762.200 45.860 ;
      LAYER met2 ;
        RECT 1342.380 1600.000 1342.660 1604.000 ;
        RECT 1342.440 1590.510 1342.580 1600.000 ;
        RECT 1342.380 1590.190 1342.640 1590.510 ;
        RECT 1344.680 1590.190 1344.940 1590.510 ;
        RECT 1344.740 45.890 1344.880 1590.190 ;
        RECT 1344.680 45.570 1344.940 45.890 ;
        RECT 2761.940 45.570 2762.200 45.890 ;
        RECT 2762.000 2.400 2762.140 45.570 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 615.090 1587.360 615.410 1587.420 ;
        RECT 619.690 1587.360 620.010 1587.420 ;
        RECT 615.090 1587.220 620.010 1587.360 ;
        RECT 615.090 1587.160 615.410 1587.220 ;
        RECT 619.690 1587.160 620.010 1587.220 ;
        RECT 619.690 30.500 620.010 30.560 ;
        RECT 835.430 30.500 835.750 30.560 ;
        RECT 619.690 30.360 835.750 30.500 ;
        RECT 619.690 30.300 620.010 30.360 ;
        RECT 835.430 30.300 835.750 30.360 ;
      LAYER via ;
        RECT 615.120 1587.160 615.380 1587.420 ;
        RECT 619.720 1587.160 619.980 1587.420 ;
        RECT 619.720 30.300 619.980 30.560 ;
        RECT 835.460 30.300 835.720 30.560 ;
      LAYER met2 ;
        RECT 615.120 1600.000 615.400 1604.000 ;
        RECT 615.180 1587.450 615.320 1600.000 ;
        RECT 615.120 1587.130 615.380 1587.450 ;
        RECT 619.720 1587.130 619.980 1587.450 ;
        RECT 619.780 30.590 619.920 1587.130 ;
        RECT 619.720 30.270 619.980 30.590 ;
        RECT 835.460 30.270 835.720 30.590 ;
        RECT 835.520 2.400 835.660 30.270 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1348.790 1590.420 1349.110 1590.480 ;
        RECT 1351.550 1590.420 1351.870 1590.480 ;
        RECT 1348.790 1590.280 1351.870 1590.420 ;
        RECT 1348.790 1590.220 1349.110 1590.280 ;
        RECT 1351.550 1590.220 1351.870 1590.280 ;
      LAYER via ;
        RECT 1348.820 1590.220 1349.080 1590.480 ;
        RECT 1351.580 1590.220 1351.840 1590.480 ;
      LAYER met2 ;
        RECT 1348.820 1600.000 1349.100 1604.000 ;
        RECT 1348.880 1590.510 1349.020 1600.000 ;
        RECT 1348.820 1590.190 1349.080 1590.510 ;
        RECT 1351.580 1590.190 1351.840 1590.510 ;
        RECT 1351.640 46.085 1351.780 1590.190 ;
        RECT 1351.570 45.715 1351.850 46.085 ;
        RECT 2779.870 45.715 2780.150 46.085 ;
        RECT 2779.940 2.400 2780.080 45.715 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
      LAYER via2 ;
        RECT 1351.570 45.760 1351.850 46.040 ;
        RECT 2779.870 45.760 2780.150 46.040 ;
      LAYER met3 ;
        RECT 1351.545 46.050 1351.875 46.065 ;
        RECT 2779.845 46.050 2780.175 46.065 ;
        RECT 1351.545 45.750 2780.175 46.050 ;
        RECT 1351.545 45.735 1351.875 45.750 ;
        RECT 2779.845 45.735 2780.175 45.750 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1355.690 1590.420 1356.010 1590.480 ;
        RECT 1358.450 1590.420 1358.770 1590.480 ;
        RECT 1355.690 1590.280 1358.770 1590.420 ;
        RECT 1355.690 1590.220 1356.010 1590.280 ;
        RECT 1358.450 1590.220 1358.770 1590.280 ;
        RECT 1358.450 45.460 1358.770 45.520 ;
        RECT 2797.790 45.460 2798.110 45.520 ;
        RECT 1358.450 45.320 2798.110 45.460 ;
        RECT 1358.450 45.260 1358.770 45.320 ;
        RECT 2797.790 45.260 2798.110 45.320 ;
      LAYER via ;
        RECT 1355.720 1590.220 1355.980 1590.480 ;
        RECT 1358.480 1590.220 1358.740 1590.480 ;
        RECT 1358.480 45.260 1358.740 45.520 ;
        RECT 2797.820 45.260 2798.080 45.520 ;
      LAYER met2 ;
        RECT 1355.720 1600.000 1356.000 1604.000 ;
        RECT 1355.780 1590.510 1355.920 1600.000 ;
        RECT 1355.720 1590.190 1355.980 1590.510 ;
        RECT 1358.480 1590.190 1358.740 1590.510 ;
        RECT 1358.540 45.550 1358.680 1590.190 ;
        RECT 1358.480 45.230 1358.740 45.550 ;
        RECT 2797.820 45.230 2798.080 45.550 ;
        RECT 2797.880 2.400 2798.020 45.230 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1362.590 1590.760 1362.910 1590.820 ;
        RECT 1365.350 1590.760 1365.670 1590.820 ;
        RECT 1362.590 1590.620 1365.670 1590.760 ;
        RECT 1362.590 1590.560 1362.910 1590.620 ;
        RECT 1365.350 1590.560 1365.670 1590.620 ;
        RECT 1365.350 31.180 1365.670 31.240 ;
        RECT 2815.730 31.180 2816.050 31.240 ;
        RECT 1365.350 31.040 2816.050 31.180 ;
        RECT 1365.350 30.980 1365.670 31.040 ;
        RECT 2815.730 30.980 2816.050 31.040 ;
      LAYER via ;
        RECT 1362.620 1590.560 1362.880 1590.820 ;
        RECT 1365.380 1590.560 1365.640 1590.820 ;
        RECT 1365.380 30.980 1365.640 31.240 ;
        RECT 2815.760 30.980 2816.020 31.240 ;
      LAYER met2 ;
        RECT 1362.620 1600.000 1362.900 1604.000 ;
        RECT 1362.680 1590.850 1362.820 1600.000 ;
        RECT 1362.620 1590.530 1362.880 1590.850 ;
        RECT 1365.380 1590.530 1365.640 1590.850 ;
        RECT 1365.440 31.270 1365.580 1590.530 ;
        RECT 1365.380 30.950 1365.640 31.270 ;
        RECT 2815.760 30.950 2816.020 31.270 ;
        RECT 2815.820 2.400 2815.960 30.950 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1369.030 1590.420 1369.350 1590.480 ;
        RECT 1372.250 1590.420 1372.570 1590.480 ;
        RECT 1369.030 1590.280 1372.570 1590.420 ;
        RECT 1369.030 1590.220 1369.350 1590.280 ;
        RECT 1372.250 1590.220 1372.570 1590.280 ;
        RECT 1372.250 45.120 1372.570 45.180 ;
        RECT 2833.670 45.120 2833.990 45.180 ;
        RECT 1372.250 44.980 2833.990 45.120 ;
        RECT 1372.250 44.920 1372.570 44.980 ;
        RECT 2833.670 44.920 2833.990 44.980 ;
      LAYER via ;
        RECT 1369.060 1590.220 1369.320 1590.480 ;
        RECT 1372.280 1590.220 1372.540 1590.480 ;
        RECT 1372.280 44.920 1372.540 45.180 ;
        RECT 2833.700 44.920 2833.960 45.180 ;
      LAYER met2 ;
        RECT 1369.060 1600.000 1369.340 1604.000 ;
        RECT 1369.120 1590.510 1369.260 1600.000 ;
        RECT 1369.060 1590.190 1369.320 1590.510 ;
        RECT 1372.280 1590.190 1372.540 1590.510 ;
        RECT 1372.340 45.210 1372.480 1590.190 ;
        RECT 1372.280 44.890 1372.540 45.210 ;
        RECT 2833.700 44.890 2833.960 45.210 ;
        RECT 2833.760 2.400 2833.900 44.890 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1375.930 1589.060 1376.250 1589.120 ;
        RECT 1379.150 1589.060 1379.470 1589.120 ;
        RECT 1375.930 1588.920 1379.470 1589.060 ;
        RECT 1375.930 1588.860 1376.250 1588.920 ;
        RECT 1379.150 1588.860 1379.470 1588.920 ;
      LAYER via ;
        RECT 1375.960 1588.860 1376.220 1589.120 ;
        RECT 1379.180 1588.860 1379.440 1589.120 ;
      LAYER met2 ;
        RECT 1375.960 1600.000 1376.240 1604.000 ;
        RECT 1376.020 1589.150 1376.160 1600.000 ;
        RECT 1375.960 1588.830 1376.220 1589.150 ;
        RECT 1379.180 1588.830 1379.440 1589.150 ;
        RECT 1379.240 45.405 1379.380 1588.830 ;
        RECT 1379.170 45.035 1379.450 45.405 ;
        RECT 2851.170 45.035 2851.450 45.405 ;
        RECT 2851.240 2.400 2851.380 45.035 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
      LAYER via2 ;
        RECT 1379.170 45.080 1379.450 45.360 ;
        RECT 2851.170 45.080 2851.450 45.360 ;
      LAYER met3 ;
        RECT 1379.145 45.370 1379.475 45.385 ;
        RECT 2851.145 45.370 2851.475 45.385 ;
        RECT 1379.145 45.070 2851.475 45.370 ;
        RECT 1379.145 45.055 1379.475 45.070 ;
        RECT 2851.145 45.055 2851.475 45.070 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1382.370 1590.420 1382.690 1590.480 ;
        RECT 1386.050 1590.420 1386.370 1590.480 ;
        RECT 1382.370 1590.280 1386.370 1590.420 ;
        RECT 1382.370 1590.220 1382.690 1590.280 ;
        RECT 1386.050 1590.220 1386.370 1590.280 ;
        RECT 1386.050 30.840 1386.370 30.900 ;
        RECT 2869.090 30.840 2869.410 30.900 ;
        RECT 1386.050 30.700 2869.410 30.840 ;
        RECT 1386.050 30.640 1386.370 30.700 ;
        RECT 2869.090 30.640 2869.410 30.700 ;
      LAYER via ;
        RECT 1382.400 1590.220 1382.660 1590.480 ;
        RECT 1386.080 1590.220 1386.340 1590.480 ;
        RECT 1386.080 30.640 1386.340 30.900 ;
        RECT 2869.120 30.640 2869.380 30.900 ;
      LAYER met2 ;
        RECT 1382.400 1600.000 1382.680 1604.000 ;
        RECT 1382.460 1590.510 1382.600 1600.000 ;
        RECT 1382.400 1590.190 1382.660 1590.510 ;
        RECT 1386.080 1590.190 1386.340 1590.510 ;
        RECT 1386.140 30.930 1386.280 1590.190 ;
        RECT 1386.080 30.610 1386.340 30.930 ;
        RECT 2869.120 30.610 2869.380 30.930 ;
        RECT 2869.180 2.400 2869.320 30.610 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1389.270 1589.400 1389.590 1589.460 ;
        RECT 1392.950 1589.400 1393.270 1589.460 ;
        RECT 1389.270 1589.260 1393.270 1589.400 ;
        RECT 1389.270 1589.200 1389.590 1589.260 ;
        RECT 1392.950 1589.200 1393.270 1589.260 ;
        RECT 1392.950 44.780 1393.270 44.840 ;
        RECT 2887.030 44.780 2887.350 44.840 ;
        RECT 1392.950 44.640 2887.350 44.780 ;
        RECT 1392.950 44.580 1393.270 44.640 ;
        RECT 2887.030 44.580 2887.350 44.640 ;
      LAYER via ;
        RECT 1389.300 1589.200 1389.560 1589.460 ;
        RECT 1392.980 1589.200 1393.240 1589.460 ;
        RECT 1392.980 44.580 1393.240 44.840 ;
        RECT 2887.060 44.580 2887.320 44.840 ;
      LAYER met2 ;
        RECT 1389.300 1600.000 1389.580 1604.000 ;
        RECT 1389.360 1589.490 1389.500 1600.000 ;
        RECT 1389.300 1589.170 1389.560 1589.490 ;
        RECT 1392.980 1589.170 1393.240 1589.490 ;
        RECT 1393.040 44.870 1393.180 1589.170 ;
        RECT 1392.980 44.550 1393.240 44.870 ;
        RECT 2887.060 44.550 2887.320 44.870 ;
        RECT 2887.120 2.400 2887.260 44.550 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1396.200 1600.450 1396.480 1604.000 ;
        RECT 1396.200 1600.310 1398.240 1600.450 ;
        RECT 1396.200 1600.000 1396.480 1600.310 ;
        RECT 1398.100 1590.250 1398.240 1600.310 ;
        RECT 1398.100 1590.110 1400.080 1590.250 ;
        RECT 1399.940 44.725 1400.080 1590.110 ;
        RECT 1399.870 44.355 1400.150 44.725 ;
        RECT 2904.990 44.355 2905.270 44.725 ;
        RECT 2905.060 2.400 2905.200 44.355 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 1399.870 44.400 1400.150 44.680 ;
        RECT 2904.990 44.400 2905.270 44.680 ;
      LAYER met3 ;
        RECT 1399.845 44.690 1400.175 44.705 ;
        RECT 2904.965 44.690 2905.295 44.705 ;
        RECT 1399.845 44.390 2905.295 44.690 ;
        RECT 1399.845 44.375 1400.175 44.390 ;
        RECT 2904.965 44.375 2905.295 44.390 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 621.530 1587.360 621.850 1587.420 ;
        RECT 627.050 1587.360 627.370 1587.420 ;
        RECT 621.530 1587.220 627.370 1587.360 ;
        RECT 621.530 1587.160 621.850 1587.220 ;
        RECT 627.050 1587.160 627.370 1587.220 ;
        RECT 627.050 34.240 627.370 34.300 ;
        RECT 852.910 34.240 853.230 34.300 ;
        RECT 627.050 34.100 853.230 34.240 ;
        RECT 627.050 34.040 627.370 34.100 ;
        RECT 852.910 34.040 853.230 34.100 ;
      LAYER via ;
        RECT 621.560 1587.160 621.820 1587.420 ;
        RECT 627.080 1587.160 627.340 1587.420 ;
        RECT 627.080 34.040 627.340 34.300 ;
        RECT 852.940 34.040 853.200 34.300 ;
      LAYER met2 ;
        RECT 621.560 1600.000 621.840 1604.000 ;
        RECT 621.620 1587.450 621.760 1600.000 ;
        RECT 621.560 1587.130 621.820 1587.450 ;
        RECT 627.080 1587.130 627.340 1587.450 ;
        RECT 627.140 34.330 627.280 1587.130 ;
        RECT 627.080 34.010 627.340 34.330 ;
        RECT 852.940 34.010 853.200 34.330 ;
        RECT 853.000 2.400 853.140 34.010 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 628.430 1587.360 628.750 1587.420 ;
        RECT 634.410 1587.360 634.730 1587.420 ;
        RECT 628.430 1587.220 634.730 1587.360 ;
        RECT 628.430 1587.160 628.750 1587.220 ;
        RECT 634.410 1587.160 634.730 1587.220 ;
        RECT 634.410 33.900 634.730 33.960 ;
        RECT 870.850 33.900 871.170 33.960 ;
        RECT 634.410 33.760 871.170 33.900 ;
        RECT 634.410 33.700 634.730 33.760 ;
        RECT 870.850 33.700 871.170 33.760 ;
      LAYER via ;
        RECT 628.460 1587.160 628.720 1587.420 ;
        RECT 634.440 1587.160 634.700 1587.420 ;
        RECT 634.440 33.700 634.700 33.960 ;
        RECT 870.880 33.700 871.140 33.960 ;
      LAYER met2 ;
        RECT 628.460 1600.000 628.740 1604.000 ;
        RECT 628.520 1587.450 628.660 1600.000 ;
        RECT 628.460 1587.130 628.720 1587.450 ;
        RECT 634.440 1587.130 634.700 1587.450 ;
        RECT 634.500 33.990 634.640 1587.130 ;
        RECT 634.440 33.670 634.700 33.990 ;
        RECT 870.880 33.670 871.140 33.990 ;
        RECT 870.940 2.400 871.080 33.670 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 635.330 1589.400 635.650 1589.460 ;
        RECT 641.310 1589.400 641.630 1589.460 ;
        RECT 635.330 1589.260 641.630 1589.400 ;
        RECT 635.330 1589.200 635.650 1589.260 ;
        RECT 641.310 1589.200 641.630 1589.260 ;
        RECT 641.310 33.560 641.630 33.620 ;
        RECT 888.790 33.560 889.110 33.620 ;
        RECT 641.310 33.420 889.110 33.560 ;
        RECT 641.310 33.360 641.630 33.420 ;
        RECT 888.790 33.360 889.110 33.420 ;
      LAYER via ;
        RECT 635.360 1589.200 635.620 1589.460 ;
        RECT 641.340 1589.200 641.600 1589.460 ;
        RECT 641.340 33.360 641.600 33.620 ;
        RECT 888.820 33.360 889.080 33.620 ;
      LAYER met2 ;
        RECT 635.360 1600.000 635.640 1604.000 ;
        RECT 635.420 1589.490 635.560 1600.000 ;
        RECT 635.360 1589.170 635.620 1589.490 ;
        RECT 641.340 1589.170 641.600 1589.490 ;
        RECT 641.400 33.650 641.540 1589.170 ;
        RECT 641.340 33.330 641.600 33.650 ;
        RECT 888.820 33.330 889.080 33.650 ;
        RECT 888.880 2.400 889.020 33.330 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 641.770 1577.160 642.090 1577.220 ;
        RECT 647.750 1577.160 648.070 1577.220 ;
        RECT 641.770 1577.020 648.070 1577.160 ;
        RECT 641.770 1576.960 642.090 1577.020 ;
        RECT 647.750 1576.960 648.070 1577.020 ;
        RECT 647.750 33.220 648.070 33.280 ;
        RECT 906.730 33.220 907.050 33.280 ;
        RECT 647.750 33.080 907.050 33.220 ;
        RECT 647.750 33.020 648.070 33.080 ;
        RECT 906.730 33.020 907.050 33.080 ;
      LAYER via ;
        RECT 641.800 1576.960 642.060 1577.220 ;
        RECT 647.780 1576.960 648.040 1577.220 ;
        RECT 647.780 33.020 648.040 33.280 ;
        RECT 906.760 33.020 907.020 33.280 ;
      LAYER met2 ;
        RECT 641.800 1600.000 642.080 1604.000 ;
        RECT 641.860 1577.250 642.000 1600.000 ;
        RECT 641.800 1576.930 642.060 1577.250 ;
        RECT 647.780 1576.930 648.040 1577.250 ;
        RECT 647.840 33.310 647.980 1576.930 ;
        RECT 647.780 32.990 648.040 33.310 ;
        RECT 906.760 32.990 907.020 33.310 ;
        RECT 906.820 2.400 906.960 32.990 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 648.670 1587.360 648.990 1587.420 ;
        RECT 655.110 1587.360 655.430 1587.420 ;
        RECT 648.670 1587.220 655.430 1587.360 ;
        RECT 648.670 1587.160 648.990 1587.220 ;
        RECT 655.110 1587.160 655.430 1587.220 ;
        RECT 655.110 32.880 655.430 32.940 ;
        RECT 924.210 32.880 924.530 32.940 ;
        RECT 655.110 32.740 924.530 32.880 ;
        RECT 655.110 32.680 655.430 32.740 ;
        RECT 924.210 32.680 924.530 32.740 ;
      LAYER via ;
        RECT 648.700 1587.160 648.960 1587.420 ;
        RECT 655.140 1587.160 655.400 1587.420 ;
        RECT 655.140 32.680 655.400 32.940 ;
        RECT 924.240 32.680 924.500 32.940 ;
      LAYER met2 ;
        RECT 648.700 1600.000 648.980 1604.000 ;
        RECT 648.760 1587.450 648.900 1600.000 ;
        RECT 648.700 1587.130 648.960 1587.450 ;
        RECT 655.140 1587.130 655.400 1587.450 ;
        RECT 655.200 32.970 655.340 1587.130 ;
        RECT 655.140 32.650 655.400 32.970 ;
        RECT 924.240 32.650 924.500 32.970 ;
        RECT 924.300 2.400 924.440 32.650 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 654.650 32.540 654.970 32.600 ;
        RECT 942.150 32.540 942.470 32.600 ;
        RECT 654.650 32.400 942.470 32.540 ;
        RECT 654.650 32.340 654.970 32.400 ;
        RECT 942.150 32.340 942.470 32.400 ;
      LAYER via ;
        RECT 654.680 32.340 654.940 32.600 ;
        RECT 942.180 32.340 942.440 32.600 ;
      LAYER met2 ;
        RECT 655.140 1600.450 655.420 1604.000 ;
        RECT 654.740 1600.310 655.420 1600.450 ;
        RECT 654.740 32.630 654.880 1600.310 ;
        RECT 655.140 1600.000 655.420 1600.310 ;
        RECT 654.680 32.310 654.940 32.630 ;
        RECT 942.180 32.310 942.440 32.630 ;
        RECT 942.240 2.400 942.380 32.310 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 661.550 32.200 661.870 32.260 ;
        RECT 960.090 32.200 960.410 32.260 ;
        RECT 661.550 32.060 960.410 32.200 ;
        RECT 661.550 32.000 661.870 32.060 ;
        RECT 960.090 32.000 960.410 32.060 ;
      LAYER via ;
        RECT 661.580 32.000 661.840 32.260 ;
        RECT 960.120 32.000 960.380 32.260 ;
      LAYER met2 ;
        RECT 662.040 1600.450 662.320 1604.000 ;
        RECT 661.640 1600.310 662.320 1600.450 ;
        RECT 661.640 32.290 661.780 1600.310 ;
        RECT 662.040 1600.000 662.320 1600.310 ;
        RECT 661.580 31.970 661.840 32.290 ;
        RECT 960.120 31.970 960.380 32.290 ;
        RECT 960.180 2.400 960.320 31.970 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 668.450 31.860 668.770 31.920 ;
        RECT 978.030 31.860 978.350 31.920 ;
        RECT 668.450 31.720 978.350 31.860 ;
        RECT 668.450 31.660 668.770 31.720 ;
        RECT 978.030 31.660 978.350 31.720 ;
      LAYER via ;
        RECT 668.480 31.660 668.740 31.920 ;
        RECT 978.060 31.660 978.320 31.920 ;
      LAYER met2 ;
        RECT 668.940 1600.450 669.220 1604.000 ;
        RECT 668.540 1600.310 669.220 1600.450 ;
        RECT 668.540 31.950 668.680 1600.310 ;
        RECT 668.940 1600.000 669.220 1600.310 ;
        RECT 668.480 31.630 668.740 31.950 ;
        RECT 978.060 31.630 978.320 31.950 ;
        RECT 978.120 2.400 978.260 31.630 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 547.470 1587.700 547.790 1587.760 ;
        RECT 550.690 1587.700 551.010 1587.760 ;
        RECT 547.470 1587.560 551.010 1587.700 ;
        RECT 547.470 1587.500 547.790 1587.560 ;
        RECT 550.690 1587.500 551.010 1587.560 ;
        RECT 656.950 18.940 657.270 19.000 ;
        RECT 617.020 18.800 657.270 18.940 ;
        RECT 550.690 18.260 551.010 18.320 ;
        RECT 617.020 18.260 617.160 18.800 ;
        RECT 656.950 18.740 657.270 18.800 ;
        RECT 550.690 18.120 617.160 18.260 ;
        RECT 550.690 18.060 551.010 18.120 ;
      LAYER via ;
        RECT 547.500 1587.500 547.760 1587.760 ;
        RECT 550.720 1587.500 550.980 1587.760 ;
        RECT 550.720 18.060 550.980 18.320 ;
        RECT 656.980 18.740 657.240 19.000 ;
      LAYER met2 ;
        RECT 547.500 1600.000 547.780 1604.000 ;
        RECT 547.560 1587.790 547.700 1600.000 ;
        RECT 547.500 1587.470 547.760 1587.790 ;
        RECT 550.720 1587.470 550.980 1587.790 ;
        RECT 550.780 18.350 550.920 1587.470 ;
        RECT 656.980 18.710 657.240 19.030 ;
        RECT 550.720 18.030 550.980 18.350 ;
        RECT 657.040 2.400 657.180 18.710 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 675.425 1545.725 675.595 1559.835 ;
        RECT 674.965 1497.445 675.135 1511.215 ;
        RECT 674.505 1400.885 674.675 1448.995 ;
        RECT 674.505 1304.325 674.675 1352.435 ;
        RECT 674.505 1207.425 674.675 1255.875 ;
        RECT 674.505 1110.865 674.675 1124.975 ;
        RECT 674.505 1014.305 674.675 1028.415 ;
        RECT 675.425 772.905 675.595 787.355 ;
        RECT 675.425 724.625 675.595 738.395 ;
        RECT 674.965 572.645 675.135 620.755 ;
        RECT 674.965 448.205 675.135 524.195 ;
        RECT 674.505 89.845 674.675 137.955 ;
      LAYER mcon ;
        RECT 675.425 1559.665 675.595 1559.835 ;
        RECT 674.965 1511.045 675.135 1511.215 ;
        RECT 674.505 1448.825 674.675 1448.995 ;
        RECT 674.505 1352.265 674.675 1352.435 ;
        RECT 674.505 1255.705 674.675 1255.875 ;
        RECT 674.505 1124.805 674.675 1124.975 ;
        RECT 674.505 1028.245 674.675 1028.415 ;
        RECT 675.425 787.185 675.595 787.355 ;
        RECT 675.425 738.225 675.595 738.395 ;
        RECT 674.965 620.585 675.135 620.755 ;
        RECT 674.965 524.025 675.135 524.195 ;
        RECT 674.505 137.785 674.675 137.955 ;
      LAYER met1 ;
        RECT 675.365 1559.820 675.655 1559.865 ;
        RECT 675.810 1559.820 676.130 1559.880 ;
        RECT 675.365 1559.680 676.130 1559.820 ;
        RECT 675.365 1559.635 675.655 1559.680 ;
        RECT 675.810 1559.620 676.130 1559.680 ;
        RECT 675.350 1545.880 675.670 1545.940 ;
        RECT 675.155 1545.740 675.670 1545.880 ;
        RECT 675.350 1545.680 675.670 1545.740 ;
        RECT 674.890 1511.200 675.210 1511.260 ;
        RECT 674.695 1511.060 675.210 1511.200 ;
        RECT 674.890 1511.000 675.210 1511.060 ;
        RECT 674.890 1497.600 675.210 1497.660 ;
        RECT 674.695 1497.460 675.210 1497.600 ;
        RECT 674.890 1497.400 675.210 1497.460 ;
        RECT 674.445 1448.980 674.735 1449.025 ;
        RECT 675.810 1448.980 676.130 1449.040 ;
        RECT 674.445 1448.840 676.130 1448.980 ;
        RECT 674.445 1448.795 674.735 1448.840 ;
        RECT 675.810 1448.780 676.130 1448.840 ;
        RECT 674.430 1401.040 674.750 1401.100 ;
        RECT 674.235 1400.900 674.750 1401.040 ;
        RECT 674.430 1400.840 674.750 1400.900 ;
        RECT 674.445 1352.420 674.735 1352.465 ;
        RECT 674.890 1352.420 675.210 1352.480 ;
        RECT 674.445 1352.280 675.210 1352.420 ;
        RECT 674.445 1352.235 674.735 1352.280 ;
        RECT 674.890 1352.220 675.210 1352.280 ;
        RECT 674.430 1304.480 674.750 1304.540 ;
        RECT 674.235 1304.340 674.750 1304.480 ;
        RECT 674.430 1304.280 674.750 1304.340 ;
        RECT 674.445 1255.860 674.735 1255.905 ;
        RECT 674.890 1255.860 675.210 1255.920 ;
        RECT 674.445 1255.720 675.210 1255.860 ;
        RECT 674.445 1255.675 674.735 1255.720 ;
        RECT 674.890 1255.660 675.210 1255.720 ;
        RECT 674.430 1207.580 674.750 1207.640 ;
        RECT 674.235 1207.440 674.750 1207.580 ;
        RECT 674.430 1207.380 674.750 1207.440 ;
        RECT 674.430 1173.040 674.750 1173.300 ;
        RECT 674.520 1172.560 674.660 1173.040 ;
        RECT 674.890 1172.560 675.210 1172.620 ;
        RECT 674.520 1172.420 675.210 1172.560 ;
        RECT 674.890 1172.360 675.210 1172.420 ;
        RECT 674.430 1124.960 674.750 1125.020 ;
        RECT 674.235 1124.820 674.750 1124.960 ;
        RECT 674.430 1124.760 674.750 1124.820 ;
        RECT 674.430 1111.020 674.750 1111.080 ;
        RECT 674.235 1110.880 674.750 1111.020 ;
        RECT 674.430 1110.820 674.750 1110.880 ;
        RECT 674.430 1076.480 674.750 1076.740 ;
        RECT 674.520 1076.000 674.660 1076.480 ;
        RECT 674.890 1076.000 675.210 1076.060 ;
        RECT 674.520 1075.860 675.210 1076.000 ;
        RECT 674.890 1075.800 675.210 1075.860 ;
        RECT 674.430 1028.400 674.750 1028.460 ;
        RECT 674.235 1028.260 674.750 1028.400 ;
        RECT 674.430 1028.200 674.750 1028.260 ;
        RECT 674.430 1014.460 674.750 1014.520 ;
        RECT 674.235 1014.320 674.750 1014.460 ;
        RECT 674.430 1014.260 674.750 1014.320 ;
        RECT 674.430 979.920 674.750 980.180 ;
        RECT 674.520 979.440 674.660 979.920 ;
        RECT 674.890 979.440 675.210 979.500 ;
        RECT 674.520 979.300 675.210 979.440 ;
        RECT 674.890 979.240 675.210 979.300 ;
        RECT 673.970 917.900 674.290 917.960 ;
        RECT 675.350 917.900 675.670 917.960 ;
        RECT 673.970 917.760 675.670 917.900 ;
        RECT 673.970 917.700 674.290 917.760 ;
        RECT 675.350 917.700 675.670 917.760 ;
        RECT 675.350 883.700 675.670 883.960 ;
        RECT 674.890 882.880 675.210 882.940 ;
        RECT 675.440 882.880 675.580 883.700 ;
        RECT 674.890 882.740 675.580 882.880 ;
        RECT 674.890 882.680 675.210 882.740 ;
        RECT 673.970 834.940 674.290 835.000 ;
        RECT 674.890 834.940 675.210 835.000 ;
        RECT 673.970 834.800 675.210 834.940 ;
        RECT 673.970 834.740 674.290 834.800 ;
        RECT 674.890 834.740 675.210 834.800 ;
        RECT 675.350 787.340 675.670 787.400 ;
        RECT 675.155 787.200 675.670 787.340 ;
        RECT 675.350 787.140 675.670 787.200 ;
        RECT 675.350 773.060 675.670 773.120 ;
        RECT 675.155 772.920 675.670 773.060 ;
        RECT 675.350 772.860 675.670 772.920 ;
        RECT 675.350 738.380 675.670 738.440 ;
        RECT 675.155 738.240 675.670 738.380 ;
        RECT 675.350 738.180 675.670 738.240 ;
        RECT 675.350 724.780 675.670 724.840 ;
        RECT 675.155 724.640 675.670 724.780 ;
        RECT 675.350 724.580 675.670 724.640 ;
        RECT 675.350 690.440 675.670 690.500 ;
        RECT 674.980 690.300 675.670 690.440 ;
        RECT 674.980 689.820 675.120 690.300 ;
        RECT 675.350 690.240 675.670 690.300 ;
        RECT 674.890 689.560 675.210 689.820 ;
        RECT 674.890 641.620 675.210 641.880 ;
        RECT 674.980 641.480 675.120 641.620 ;
        RECT 675.350 641.480 675.670 641.540 ;
        RECT 674.980 641.340 675.670 641.480 ;
        RECT 675.350 641.280 675.670 641.340 ;
        RECT 674.905 620.740 675.195 620.785 ;
        RECT 675.350 620.740 675.670 620.800 ;
        RECT 674.905 620.600 675.670 620.740 ;
        RECT 674.905 620.555 675.195 620.600 ;
        RECT 675.350 620.540 675.670 620.600 ;
        RECT 674.890 572.800 675.210 572.860 ;
        RECT 674.695 572.660 675.210 572.800 ;
        RECT 674.890 572.600 675.210 572.660 ;
        RECT 674.890 545.060 675.210 545.320 ;
        RECT 674.980 544.920 675.120 545.060 ;
        RECT 675.350 544.920 675.670 544.980 ;
        RECT 674.980 544.780 675.670 544.920 ;
        RECT 675.350 544.720 675.670 544.780 ;
        RECT 674.905 524.180 675.195 524.225 ;
        RECT 675.350 524.180 675.670 524.240 ;
        RECT 674.905 524.040 675.670 524.180 ;
        RECT 674.905 523.995 675.195 524.040 ;
        RECT 675.350 523.980 675.670 524.040 ;
        RECT 674.890 448.360 675.210 448.420 ;
        RECT 674.695 448.220 675.210 448.360 ;
        RECT 674.890 448.160 675.210 448.220 ;
        RECT 673.510 410.620 673.830 410.680 ;
        RECT 675.350 410.620 675.670 410.680 ;
        RECT 673.510 410.480 675.670 410.620 ;
        RECT 673.510 410.420 673.830 410.480 ;
        RECT 675.350 410.420 675.670 410.480 ;
        RECT 674.890 352.480 675.210 352.540 ;
        RECT 674.520 352.340 675.210 352.480 ;
        RECT 674.520 351.860 674.660 352.340 ;
        RECT 674.890 352.280 675.210 352.340 ;
        RECT 674.430 351.600 674.750 351.860 ;
        RECT 674.430 331.060 674.750 331.120 ;
        RECT 675.350 331.060 675.670 331.120 ;
        RECT 674.430 330.920 675.670 331.060 ;
        RECT 674.430 330.860 674.750 330.920 ;
        RECT 675.350 330.860 675.670 330.920 ;
        RECT 674.430 234.500 674.750 234.560 ;
        RECT 675.350 234.500 675.670 234.560 ;
        RECT 674.430 234.360 675.670 234.500 ;
        RECT 674.430 234.300 674.750 234.360 ;
        RECT 675.350 234.300 675.670 234.360 ;
        RECT 674.430 137.940 674.750 138.000 ;
        RECT 674.235 137.800 674.750 137.940 ;
        RECT 674.430 137.740 674.750 137.800 ;
        RECT 674.445 90.000 674.735 90.045 ;
        RECT 674.890 90.000 675.210 90.060 ;
        RECT 674.445 89.860 675.210 90.000 ;
        RECT 674.445 89.815 674.735 89.860 ;
        RECT 674.890 89.800 675.210 89.860 ;
        RECT 674.890 62.460 675.210 62.520 ;
        RECT 674.520 62.320 675.210 62.460 ;
        RECT 674.520 62.180 674.660 62.320 ;
        RECT 674.890 62.260 675.210 62.320 ;
        RECT 674.430 61.920 674.750 62.180 ;
        RECT 674.430 31.520 674.750 31.580 ;
        RECT 995.970 31.520 996.290 31.580 ;
        RECT 674.430 31.380 996.290 31.520 ;
        RECT 674.430 31.320 674.750 31.380 ;
        RECT 995.970 31.320 996.290 31.380 ;
      LAYER via ;
        RECT 675.840 1559.620 676.100 1559.880 ;
        RECT 675.380 1545.680 675.640 1545.940 ;
        RECT 674.920 1511.000 675.180 1511.260 ;
        RECT 674.920 1497.400 675.180 1497.660 ;
        RECT 675.840 1448.780 676.100 1449.040 ;
        RECT 674.460 1400.840 674.720 1401.100 ;
        RECT 674.920 1352.220 675.180 1352.480 ;
        RECT 674.460 1304.280 674.720 1304.540 ;
        RECT 674.920 1255.660 675.180 1255.920 ;
        RECT 674.460 1207.380 674.720 1207.640 ;
        RECT 674.460 1173.040 674.720 1173.300 ;
        RECT 674.920 1172.360 675.180 1172.620 ;
        RECT 674.460 1124.760 674.720 1125.020 ;
        RECT 674.460 1110.820 674.720 1111.080 ;
        RECT 674.460 1076.480 674.720 1076.740 ;
        RECT 674.920 1075.800 675.180 1076.060 ;
        RECT 674.460 1028.200 674.720 1028.460 ;
        RECT 674.460 1014.260 674.720 1014.520 ;
        RECT 674.460 979.920 674.720 980.180 ;
        RECT 674.920 979.240 675.180 979.500 ;
        RECT 674.000 917.700 674.260 917.960 ;
        RECT 675.380 917.700 675.640 917.960 ;
        RECT 675.380 883.700 675.640 883.960 ;
        RECT 674.920 882.680 675.180 882.940 ;
        RECT 674.000 834.740 674.260 835.000 ;
        RECT 674.920 834.740 675.180 835.000 ;
        RECT 675.380 787.140 675.640 787.400 ;
        RECT 675.380 772.860 675.640 773.120 ;
        RECT 675.380 738.180 675.640 738.440 ;
        RECT 675.380 724.580 675.640 724.840 ;
        RECT 675.380 690.240 675.640 690.500 ;
        RECT 674.920 689.560 675.180 689.820 ;
        RECT 674.920 641.620 675.180 641.880 ;
        RECT 675.380 641.280 675.640 641.540 ;
        RECT 675.380 620.540 675.640 620.800 ;
        RECT 674.920 572.600 675.180 572.860 ;
        RECT 674.920 545.060 675.180 545.320 ;
        RECT 675.380 544.720 675.640 544.980 ;
        RECT 675.380 523.980 675.640 524.240 ;
        RECT 674.920 448.160 675.180 448.420 ;
        RECT 673.540 410.420 673.800 410.680 ;
        RECT 675.380 410.420 675.640 410.680 ;
        RECT 674.920 352.280 675.180 352.540 ;
        RECT 674.460 351.600 674.720 351.860 ;
        RECT 674.460 330.860 674.720 331.120 ;
        RECT 675.380 330.860 675.640 331.120 ;
        RECT 674.460 234.300 674.720 234.560 ;
        RECT 675.380 234.300 675.640 234.560 ;
        RECT 674.460 137.740 674.720 138.000 ;
        RECT 674.920 89.800 675.180 90.060 ;
        RECT 674.920 62.260 675.180 62.520 ;
        RECT 674.460 61.920 674.720 62.180 ;
        RECT 674.460 31.320 674.720 31.580 ;
        RECT 996.000 31.320 996.260 31.580 ;
      LAYER met2 ;
        RECT 675.380 1600.450 675.660 1604.000 ;
        RECT 675.380 1600.310 676.040 1600.450 ;
        RECT 675.380 1600.000 675.660 1600.310 ;
        RECT 675.900 1559.910 676.040 1600.310 ;
        RECT 675.840 1559.590 676.100 1559.910 ;
        RECT 675.380 1545.650 675.640 1545.970 ;
        RECT 675.440 1545.370 675.580 1545.650 ;
        RECT 674.980 1545.230 675.580 1545.370 ;
        RECT 674.980 1511.290 675.120 1545.230 ;
        RECT 674.920 1510.970 675.180 1511.290 ;
        RECT 674.920 1497.370 675.180 1497.690 ;
        RECT 674.980 1463.090 675.120 1497.370 ;
        RECT 674.980 1462.950 676.040 1463.090 ;
        RECT 675.900 1449.070 676.040 1462.950 ;
        RECT 675.840 1448.750 676.100 1449.070 ;
        RECT 674.460 1400.810 674.720 1401.130 ;
        RECT 674.520 1400.530 674.660 1400.810 ;
        RECT 674.910 1400.530 675.190 1400.645 ;
        RECT 674.520 1400.390 675.190 1400.530 ;
        RECT 674.910 1400.275 675.190 1400.390 ;
        RECT 674.910 1352.675 675.190 1353.045 ;
        RECT 674.980 1352.510 675.120 1352.675 ;
        RECT 674.920 1352.190 675.180 1352.510 ;
        RECT 674.460 1304.250 674.720 1304.570 ;
        RECT 674.520 1303.970 674.660 1304.250 ;
        RECT 674.910 1303.970 675.190 1304.085 ;
        RECT 674.520 1303.830 675.190 1303.970 ;
        RECT 674.910 1303.715 675.190 1303.830 ;
        RECT 674.910 1256.115 675.190 1256.485 ;
        RECT 674.980 1255.950 675.120 1256.115 ;
        RECT 674.920 1255.630 675.180 1255.950 ;
        RECT 674.460 1207.350 674.720 1207.670 ;
        RECT 674.520 1173.330 674.660 1207.350 ;
        RECT 674.460 1173.010 674.720 1173.330 ;
        RECT 674.920 1172.330 675.180 1172.650 ;
        RECT 674.980 1159.130 675.120 1172.330 ;
        RECT 674.520 1158.990 675.120 1159.130 ;
        RECT 674.520 1125.050 674.660 1158.990 ;
        RECT 674.460 1124.730 674.720 1125.050 ;
        RECT 674.460 1110.790 674.720 1111.110 ;
        RECT 674.520 1076.770 674.660 1110.790 ;
        RECT 674.460 1076.450 674.720 1076.770 ;
        RECT 674.920 1075.770 675.180 1076.090 ;
        RECT 674.980 1062.570 675.120 1075.770 ;
        RECT 674.520 1062.430 675.120 1062.570 ;
        RECT 674.520 1028.490 674.660 1062.430 ;
        RECT 674.460 1028.170 674.720 1028.490 ;
        RECT 674.460 1014.230 674.720 1014.550 ;
        RECT 674.520 980.210 674.660 1014.230 ;
        RECT 674.460 979.890 674.720 980.210 ;
        RECT 674.920 979.210 675.180 979.530 ;
        RECT 674.980 966.125 675.120 979.210 ;
        RECT 673.990 965.755 674.270 966.125 ;
        RECT 674.910 965.755 675.190 966.125 ;
        RECT 674.060 917.990 674.200 965.755 ;
        RECT 674.000 917.670 674.260 917.990 ;
        RECT 675.380 917.670 675.640 917.990 ;
        RECT 675.440 883.990 675.580 917.670 ;
        RECT 675.380 883.670 675.640 883.990 ;
        RECT 674.920 882.650 675.180 882.970 ;
        RECT 674.980 869.565 675.120 882.650 ;
        RECT 673.990 869.195 674.270 869.565 ;
        RECT 674.910 869.195 675.190 869.565 ;
        RECT 674.060 835.030 674.200 869.195 ;
        RECT 674.000 834.710 674.260 835.030 ;
        RECT 674.920 834.710 675.180 835.030 ;
        RECT 674.980 821.170 675.120 834.710 ;
        RECT 674.980 821.030 675.580 821.170 ;
        RECT 675.440 787.430 675.580 821.030 ;
        RECT 675.380 787.110 675.640 787.430 ;
        RECT 675.380 772.830 675.640 773.150 ;
        RECT 675.440 738.470 675.580 772.830 ;
        RECT 675.380 738.150 675.640 738.470 ;
        RECT 675.380 724.550 675.640 724.870 ;
        RECT 675.440 690.530 675.580 724.550 ;
        RECT 675.380 690.210 675.640 690.530 ;
        RECT 674.920 689.530 675.180 689.850 ;
        RECT 674.980 641.910 675.120 689.530 ;
        RECT 674.920 641.590 675.180 641.910 ;
        RECT 675.380 641.250 675.640 641.570 ;
        RECT 675.440 620.830 675.580 641.250 ;
        RECT 675.380 620.510 675.640 620.830 ;
        RECT 674.920 572.570 675.180 572.890 ;
        RECT 674.980 545.350 675.120 572.570 ;
        RECT 674.920 545.030 675.180 545.350 ;
        RECT 675.380 544.690 675.640 545.010 ;
        RECT 675.440 524.270 675.580 544.690 ;
        RECT 675.380 523.950 675.640 524.270 ;
        RECT 674.920 448.130 675.180 448.450 ;
        RECT 674.980 434.930 675.120 448.130 ;
        RECT 674.980 434.790 675.580 434.930 ;
        RECT 675.440 410.710 675.580 434.790 ;
        RECT 673.540 410.390 673.800 410.710 ;
        RECT 675.380 410.390 675.640 410.710 ;
        RECT 673.600 386.765 673.740 410.390 ;
        RECT 673.530 386.395 673.810 386.765 ;
        RECT 674.450 386.650 674.730 386.765 ;
        RECT 674.450 386.510 675.120 386.650 ;
        RECT 674.450 386.395 674.730 386.510 ;
        RECT 674.980 352.570 675.120 386.510 ;
        RECT 674.920 352.250 675.180 352.570 ;
        RECT 674.460 351.570 674.720 351.890 ;
        RECT 674.520 339.165 674.660 351.570 ;
        RECT 674.450 338.795 674.730 339.165 ;
        RECT 674.450 338.115 674.730 338.485 ;
        RECT 674.520 331.150 674.660 338.115 ;
        RECT 674.460 330.830 674.720 331.150 ;
        RECT 675.380 330.830 675.640 331.150 ;
        RECT 675.440 307.205 675.580 330.830 ;
        RECT 675.370 306.835 675.650 307.205 ;
        RECT 674.910 241.810 675.190 241.925 ;
        RECT 674.520 241.670 675.190 241.810 ;
        RECT 674.520 234.590 674.660 241.670 ;
        RECT 674.910 241.555 675.190 241.670 ;
        RECT 674.460 234.270 674.720 234.590 ;
        RECT 675.380 234.270 675.640 234.590 ;
        RECT 675.440 210.645 675.580 234.270 ;
        RECT 675.370 210.275 675.650 210.645 ;
        RECT 674.910 145.250 675.190 145.365 ;
        RECT 674.520 145.110 675.190 145.250 ;
        RECT 674.520 138.030 674.660 145.110 ;
        RECT 674.910 144.995 675.190 145.110 ;
        RECT 674.460 137.710 674.720 138.030 ;
        RECT 674.920 89.770 675.180 90.090 ;
        RECT 674.980 62.550 675.120 89.770 ;
        RECT 674.920 62.230 675.180 62.550 ;
        RECT 674.460 61.890 674.720 62.210 ;
        RECT 674.520 31.610 674.660 61.890 ;
        RECT 674.460 31.290 674.720 31.610 ;
        RECT 996.000 31.290 996.260 31.610 ;
        RECT 996.060 2.400 996.200 31.290 ;
        RECT 995.850 -4.800 996.410 2.400 ;
      LAYER via2 ;
        RECT 674.910 1400.320 675.190 1400.600 ;
        RECT 674.910 1352.720 675.190 1353.000 ;
        RECT 674.910 1303.760 675.190 1304.040 ;
        RECT 674.910 1256.160 675.190 1256.440 ;
        RECT 673.990 965.800 674.270 966.080 ;
        RECT 674.910 965.800 675.190 966.080 ;
        RECT 673.990 869.240 674.270 869.520 ;
        RECT 674.910 869.240 675.190 869.520 ;
        RECT 673.530 386.440 673.810 386.720 ;
        RECT 674.450 386.440 674.730 386.720 ;
        RECT 674.450 338.840 674.730 339.120 ;
        RECT 674.450 338.160 674.730 338.440 ;
        RECT 675.370 306.880 675.650 307.160 ;
        RECT 674.910 241.600 675.190 241.880 ;
        RECT 675.370 210.320 675.650 210.600 ;
        RECT 674.910 145.040 675.190 145.320 ;
      LAYER met3 ;
        RECT 674.885 1400.610 675.215 1400.625 ;
        RECT 675.550 1400.610 675.930 1400.620 ;
        RECT 674.885 1400.310 675.930 1400.610 ;
        RECT 674.885 1400.295 675.215 1400.310 ;
        RECT 675.550 1400.300 675.930 1400.310 ;
        RECT 674.885 1353.010 675.215 1353.025 ;
        RECT 675.550 1353.010 675.930 1353.020 ;
        RECT 674.885 1352.710 675.930 1353.010 ;
        RECT 674.885 1352.695 675.215 1352.710 ;
        RECT 675.550 1352.700 675.930 1352.710 ;
        RECT 674.885 1304.050 675.215 1304.065 ;
        RECT 675.550 1304.050 675.930 1304.060 ;
        RECT 674.885 1303.750 675.930 1304.050 ;
        RECT 674.885 1303.735 675.215 1303.750 ;
        RECT 675.550 1303.740 675.930 1303.750 ;
        RECT 674.885 1256.450 675.215 1256.465 ;
        RECT 675.550 1256.450 675.930 1256.460 ;
        RECT 674.885 1256.150 675.930 1256.450 ;
        RECT 674.885 1256.135 675.215 1256.150 ;
        RECT 675.550 1256.140 675.930 1256.150 ;
        RECT 673.965 966.090 674.295 966.105 ;
        RECT 674.885 966.090 675.215 966.105 ;
        RECT 673.965 965.790 675.215 966.090 ;
        RECT 673.965 965.775 674.295 965.790 ;
        RECT 674.885 965.775 675.215 965.790 ;
        RECT 673.965 869.530 674.295 869.545 ;
        RECT 674.885 869.530 675.215 869.545 ;
        RECT 673.965 869.230 675.215 869.530 ;
        RECT 673.965 869.215 674.295 869.230 ;
        RECT 674.885 869.215 675.215 869.230 ;
        RECT 673.505 386.730 673.835 386.745 ;
        RECT 674.425 386.730 674.755 386.745 ;
        RECT 673.505 386.430 674.755 386.730 ;
        RECT 673.505 386.415 673.835 386.430 ;
        RECT 674.425 386.415 674.755 386.430 ;
        RECT 674.425 338.815 674.755 339.145 ;
        RECT 674.440 338.465 674.740 338.815 ;
        RECT 674.425 338.135 674.755 338.465 ;
        RECT 675.345 307.180 675.675 307.185 ;
        RECT 675.345 307.170 675.930 307.180 ;
        RECT 675.120 306.870 675.930 307.170 ;
        RECT 675.345 306.860 675.930 306.870 ;
        RECT 675.345 306.855 675.675 306.860 ;
        RECT 674.885 241.890 675.215 241.905 ;
        RECT 675.550 241.890 675.930 241.900 ;
        RECT 674.885 241.590 675.930 241.890 ;
        RECT 674.885 241.575 675.215 241.590 ;
        RECT 675.550 241.580 675.930 241.590 ;
        RECT 675.345 210.620 675.675 210.625 ;
        RECT 675.345 210.610 675.930 210.620 ;
        RECT 675.120 210.310 675.930 210.610 ;
        RECT 675.345 210.300 675.930 210.310 ;
        RECT 675.345 210.295 675.675 210.300 ;
        RECT 674.885 145.330 675.215 145.345 ;
        RECT 675.550 145.330 675.930 145.340 ;
        RECT 674.885 145.030 675.930 145.330 ;
        RECT 674.885 145.015 675.215 145.030 ;
        RECT 675.550 145.020 675.930 145.030 ;
      LAYER via3 ;
        RECT 675.580 1400.300 675.900 1400.620 ;
        RECT 675.580 1352.700 675.900 1353.020 ;
        RECT 675.580 1303.740 675.900 1304.060 ;
        RECT 675.580 1256.140 675.900 1256.460 ;
        RECT 675.580 306.860 675.900 307.180 ;
        RECT 675.580 241.580 675.900 241.900 ;
        RECT 675.580 210.300 675.900 210.620 ;
        RECT 675.580 145.020 675.900 145.340 ;
      LAYER met4 ;
        RECT 675.575 1400.295 675.905 1400.625 ;
        RECT 675.590 1353.025 675.890 1400.295 ;
        RECT 675.575 1352.695 675.905 1353.025 ;
        RECT 675.575 1303.735 675.905 1304.065 ;
        RECT 675.590 1256.465 675.890 1303.735 ;
        RECT 675.575 1256.135 675.905 1256.465 ;
        RECT 675.575 306.855 675.905 307.185 ;
        RECT 675.590 241.905 675.890 306.855 ;
        RECT 675.575 241.575 675.905 241.905 ;
        RECT 675.575 210.295 675.905 210.625 ;
        RECT 675.590 145.345 675.890 210.295 ;
        RECT 675.575 145.015 675.905 145.345 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 810.205 18.785 811.295 18.955 ;
        RECT 810.205 18.445 810.375 18.785 ;
        RECT 811.125 16.745 811.295 18.785 ;
        RECT 829.985 14.365 830.155 16.915 ;
      LAYER mcon ;
        RECT 829.985 16.745 830.155 16.915 ;
      LAYER met1 ;
        RECT 789.890 18.600 790.210 18.660 ;
        RECT 810.145 18.600 810.435 18.645 ;
        RECT 789.890 18.460 810.435 18.600 ;
        RECT 789.890 18.400 790.210 18.460 ;
        RECT 810.145 18.415 810.435 18.460 ;
        RECT 811.065 16.900 811.355 16.945 ;
        RECT 829.925 16.900 830.215 16.945 ;
        RECT 811.065 16.760 830.215 16.900 ;
        RECT 811.065 16.715 811.355 16.760 ;
        RECT 829.925 16.715 830.215 16.760 ;
        RECT 829.925 14.520 830.215 14.565 ;
        RECT 1013.450 14.520 1013.770 14.580 ;
        RECT 829.925 14.380 1013.770 14.520 ;
        RECT 829.925 14.335 830.215 14.380 ;
        RECT 1013.450 14.320 1013.770 14.380 ;
      LAYER via ;
        RECT 789.920 18.400 790.180 18.660 ;
        RECT 1013.480 14.320 1013.740 14.580 ;
      LAYER met2 ;
        RECT 682.280 1600.000 682.560 1604.000 ;
        RECT 682.340 1591.045 682.480 1600.000 ;
        RECT 748.510 1592.035 748.790 1592.405 ;
        RECT 748.580 1591.045 748.720 1592.035 ;
        RECT 682.270 1590.675 682.550 1591.045 ;
        RECT 748.510 1590.675 748.790 1591.045 ;
        RECT 789.450 1590.675 789.730 1591.045 ;
        RECT 789.520 1558.970 789.660 1590.675 ;
        RECT 789.520 1558.830 790.120 1558.970 ;
        RECT 789.980 18.690 790.120 1558.830 ;
        RECT 789.920 18.370 790.180 18.690 ;
        RECT 1013.480 14.290 1013.740 14.610 ;
        RECT 1013.540 2.400 1013.680 14.290 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
      LAYER via2 ;
        RECT 748.510 1592.080 748.790 1592.360 ;
        RECT 682.270 1590.720 682.550 1591.000 ;
        RECT 748.510 1590.720 748.790 1591.000 ;
        RECT 789.450 1590.720 789.730 1591.000 ;
      LAYER met3 ;
        RECT 724.310 1592.370 724.690 1592.380 ;
        RECT 748.485 1592.370 748.815 1592.385 ;
        RECT 724.310 1592.070 748.815 1592.370 ;
        RECT 724.310 1592.060 724.690 1592.070 ;
        RECT 748.485 1592.055 748.815 1592.070 ;
        RECT 682.245 1591.010 682.575 1591.025 ;
        RECT 724.310 1591.010 724.690 1591.020 ;
        RECT 682.245 1590.710 724.690 1591.010 ;
        RECT 682.245 1590.695 682.575 1590.710 ;
        RECT 724.310 1590.700 724.690 1590.710 ;
        RECT 748.485 1591.010 748.815 1591.025 ;
        RECT 789.425 1591.010 789.755 1591.025 ;
        RECT 748.485 1590.710 772.490 1591.010 ;
        RECT 748.485 1590.695 748.815 1590.710 ;
        RECT 772.190 1590.500 772.490 1590.710 ;
        RECT 773.110 1590.710 789.755 1591.010 ;
        RECT 773.110 1590.500 773.410 1590.710 ;
        RECT 789.425 1590.695 789.755 1590.710 ;
        RECT 772.190 1590.200 773.410 1590.500 ;
      LAYER via3 ;
        RECT 724.340 1592.060 724.660 1592.380 ;
        RECT 724.340 1590.700 724.660 1591.020 ;
      LAYER met4 ;
        RECT 724.335 1592.055 724.665 1592.385 ;
        RECT 724.350 1591.025 724.650 1592.055 ;
        RECT 724.335 1590.695 724.665 1591.025 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 688.690 1559.480 689.010 1559.540 ;
        RECT 689.610 1559.480 689.930 1559.540 ;
        RECT 688.690 1559.340 689.930 1559.480 ;
        RECT 688.690 1559.280 689.010 1559.340 ;
        RECT 689.610 1559.280 689.930 1559.340 ;
        RECT 688.690 41.040 689.010 41.100 ;
        RECT 1031.390 41.040 1031.710 41.100 ;
        RECT 688.690 40.900 1031.710 41.040 ;
        RECT 688.690 40.840 689.010 40.900 ;
        RECT 1031.390 40.840 1031.710 40.900 ;
      LAYER via ;
        RECT 688.720 1559.280 688.980 1559.540 ;
        RECT 689.640 1559.280 689.900 1559.540 ;
        RECT 688.720 40.840 688.980 41.100 ;
        RECT 1031.420 40.840 1031.680 41.100 ;
      LAYER met2 ;
        RECT 689.180 1600.000 689.460 1604.000 ;
        RECT 689.240 1580.730 689.380 1600.000 ;
        RECT 689.240 1580.590 689.840 1580.730 ;
        RECT 689.700 1559.570 689.840 1580.590 ;
        RECT 688.720 1559.250 688.980 1559.570 ;
        RECT 689.640 1559.250 689.900 1559.570 ;
        RECT 688.780 41.130 688.920 1559.250 ;
        RECT 688.720 40.810 688.980 41.130 ;
        RECT 1031.420 40.810 1031.680 41.130 ;
        RECT 1031.480 2.400 1031.620 40.810 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 695.590 40.700 695.910 40.760 ;
        RECT 1049.330 40.700 1049.650 40.760 ;
        RECT 695.590 40.560 1049.650 40.700 ;
        RECT 695.590 40.500 695.910 40.560 ;
        RECT 1049.330 40.500 1049.650 40.560 ;
      LAYER via ;
        RECT 695.620 40.500 695.880 40.760 ;
        RECT 1049.360 40.500 1049.620 40.760 ;
      LAYER met2 ;
        RECT 695.620 1600.000 695.900 1604.000 ;
        RECT 695.680 40.790 695.820 1600.000 ;
        RECT 695.620 40.470 695.880 40.790 ;
        RECT 1049.360 40.470 1049.620 40.790 ;
        RECT 1049.420 2.400 1049.560 40.470 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 702.490 40.360 702.810 40.420 ;
        RECT 1067.270 40.360 1067.590 40.420 ;
        RECT 702.490 40.220 1067.590 40.360 ;
        RECT 702.490 40.160 702.810 40.220 ;
        RECT 1067.270 40.160 1067.590 40.220 ;
      LAYER via ;
        RECT 702.520 40.160 702.780 40.420 ;
        RECT 1067.300 40.160 1067.560 40.420 ;
      LAYER met2 ;
        RECT 702.520 1600.000 702.800 1604.000 ;
        RECT 702.580 40.450 702.720 1600.000 ;
        RECT 702.520 40.130 702.780 40.450 ;
        RECT 1067.300 40.130 1067.560 40.450 ;
        RECT 1067.360 2.400 1067.500 40.130 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 709.390 40.020 709.710 40.080 ;
        RECT 1085.210 40.020 1085.530 40.080 ;
        RECT 709.390 39.880 1085.530 40.020 ;
        RECT 709.390 39.820 709.710 39.880 ;
        RECT 1085.210 39.820 1085.530 39.880 ;
      LAYER via ;
        RECT 709.420 39.820 709.680 40.080 ;
        RECT 1085.240 39.820 1085.500 40.080 ;
      LAYER met2 ;
        RECT 709.420 1600.000 709.700 1604.000 ;
        RECT 709.480 40.110 709.620 1600.000 ;
        RECT 709.420 39.790 709.680 40.110 ;
        RECT 1085.240 39.790 1085.500 40.110 ;
        RECT 1085.300 2.400 1085.440 39.790 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 716.290 39.680 716.610 39.740 ;
        RECT 1102.690 39.680 1103.010 39.740 ;
        RECT 716.290 39.540 1103.010 39.680 ;
        RECT 716.290 39.480 716.610 39.540 ;
        RECT 1102.690 39.480 1103.010 39.540 ;
      LAYER via ;
        RECT 716.320 39.480 716.580 39.740 ;
        RECT 1102.720 39.480 1102.980 39.740 ;
      LAYER met2 ;
        RECT 715.860 1600.450 716.140 1604.000 ;
        RECT 715.860 1600.310 716.520 1600.450 ;
        RECT 715.860 1600.000 716.140 1600.310 ;
        RECT 716.380 39.770 716.520 1600.310 ;
        RECT 716.320 39.450 716.580 39.770 ;
        RECT 1102.720 39.450 1102.980 39.770 ;
        RECT 1102.780 2.400 1102.920 39.450 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 723.190 39.340 723.510 39.400 ;
        RECT 1120.630 39.340 1120.950 39.400 ;
        RECT 723.190 39.200 1120.950 39.340 ;
        RECT 723.190 39.140 723.510 39.200 ;
        RECT 1120.630 39.140 1120.950 39.200 ;
      LAYER via ;
        RECT 723.220 39.140 723.480 39.400 ;
        RECT 1120.660 39.140 1120.920 39.400 ;
      LAYER met2 ;
        RECT 722.760 1600.450 723.040 1604.000 ;
        RECT 722.760 1600.310 723.420 1600.450 ;
        RECT 722.760 1600.000 723.040 1600.310 ;
        RECT 723.280 39.430 723.420 1600.310 ;
        RECT 723.220 39.110 723.480 39.430 ;
        RECT 1120.660 39.110 1120.920 39.430 ;
        RECT 1120.720 2.400 1120.860 39.110 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 730.550 38.660 730.870 38.720 ;
        RECT 1138.570 38.660 1138.890 38.720 ;
        RECT 730.550 38.520 1138.890 38.660 ;
        RECT 730.550 38.460 730.870 38.520 ;
        RECT 1138.570 38.460 1138.890 38.520 ;
      LAYER via ;
        RECT 730.580 38.460 730.840 38.720 ;
        RECT 1138.600 38.460 1138.860 38.720 ;
      LAYER met2 ;
        RECT 729.660 1600.450 729.940 1604.000 ;
        RECT 729.660 1600.310 730.780 1600.450 ;
        RECT 729.660 1600.000 729.940 1600.310 ;
        RECT 730.640 38.750 730.780 1600.310 ;
        RECT 730.580 38.430 730.840 38.750 ;
        RECT 1138.600 38.430 1138.860 38.750 ;
        RECT 1138.660 2.400 1138.800 38.430 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 736.990 37.980 737.310 38.040 ;
        RECT 1156.510 37.980 1156.830 38.040 ;
        RECT 736.990 37.840 1156.830 37.980 ;
        RECT 736.990 37.780 737.310 37.840 ;
        RECT 1156.510 37.780 1156.830 37.840 ;
      LAYER via ;
        RECT 737.020 37.780 737.280 38.040 ;
        RECT 1156.540 37.780 1156.800 38.040 ;
      LAYER met2 ;
        RECT 736.100 1600.450 736.380 1604.000 ;
        RECT 736.100 1600.310 737.220 1600.450 ;
        RECT 736.100 1600.000 736.380 1600.310 ;
        RECT 737.080 38.070 737.220 1600.310 ;
        RECT 737.020 37.750 737.280 38.070 ;
        RECT 1156.540 37.750 1156.800 38.070 ;
        RECT 1156.600 2.400 1156.740 37.750 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 554.370 1587.360 554.690 1587.420 ;
        RECT 558.050 1587.360 558.370 1587.420 ;
        RECT 554.370 1587.220 558.370 1587.360 ;
        RECT 554.370 1587.160 554.690 1587.220 ;
        RECT 558.050 1587.160 558.370 1587.220 ;
        RECT 558.050 14.520 558.370 14.580 ;
        RECT 674.430 14.520 674.750 14.580 ;
        RECT 558.050 14.380 674.750 14.520 ;
        RECT 558.050 14.320 558.370 14.380 ;
        RECT 674.430 14.320 674.750 14.380 ;
      LAYER via ;
        RECT 554.400 1587.160 554.660 1587.420 ;
        RECT 558.080 1587.160 558.340 1587.420 ;
        RECT 558.080 14.320 558.340 14.580 ;
        RECT 674.460 14.320 674.720 14.580 ;
      LAYER met2 ;
        RECT 554.400 1600.000 554.680 1604.000 ;
        RECT 554.460 1587.450 554.600 1600.000 ;
        RECT 554.400 1587.130 554.660 1587.450 ;
        RECT 558.080 1587.130 558.340 1587.450 ;
        RECT 558.140 14.610 558.280 1587.130 ;
        RECT 558.080 14.290 558.340 14.610 ;
        RECT 674.460 14.290 674.720 14.610 ;
        RECT 674.520 2.400 674.660 14.290 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 762.365 1592.985 762.535 1594.175 ;
        RECT 777.085 1587.545 777.255 1593.155 ;
      LAYER mcon ;
        RECT 762.365 1594.005 762.535 1594.175 ;
        RECT 777.085 1592.985 777.255 1593.155 ;
      LAYER met1 ;
        RECT 762.305 1594.160 762.595 1594.205 ;
        RECT 751.340 1594.020 762.595 1594.160 ;
        RECT 742.970 1593.820 743.290 1593.880 ;
        RECT 751.340 1593.820 751.480 1594.020 ;
        RECT 762.305 1593.975 762.595 1594.020 ;
        RECT 742.970 1593.680 751.480 1593.820 ;
        RECT 742.970 1593.620 743.290 1593.680 ;
        RECT 762.305 1593.140 762.595 1593.185 ;
        RECT 777.025 1593.140 777.315 1593.185 ;
        RECT 762.305 1593.000 777.315 1593.140 ;
        RECT 762.305 1592.955 762.595 1593.000 ;
        RECT 777.025 1592.955 777.315 1593.000 ;
        RECT 777.025 1587.700 777.315 1587.745 ;
        RECT 777.025 1587.560 780.000 1587.700 ;
        RECT 777.025 1587.515 777.315 1587.560 ;
        RECT 779.860 1587.360 780.000 1587.560 ;
        RECT 789.520 1587.560 796.560 1587.700 ;
        RECT 789.520 1587.360 789.660 1587.560 ;
        RECT 779.860 1587.220 789.660 1587.360 ;
        RECT 796.420 1587.020 796.560 1587.560 ;
        RECT 796.420 1586.880 797.020 1587.020 ;
        RECT 796.880 1586.740 797.020 1586.880 ;
        RECT 796.790 1586.480 797.110 1586.740 ;
      LAYER via ;
        RECT 743.000 1593.620 743.260 1593.880 ;
        RECT 796.820 1586.480 797.080 1586.740 ;
      LAYER met2 ;
        RECT 743.000 1600.000 743.280 1604.000 ;
        RECT 743.060 1593.910 743.200 1600.000 ;
        RECT 743.000 1593.590 743.260 1593.910 ;
        RECT 796.820 1586.450 797.080 1586.770 ;
        RECT 796.880 15.485 797.020 1586.450 ;
        RECT 813.830 17.155 814.110 17.525 ;
        RECT 1174.010 17.155 1174.290 17.525 ;
        RECT 813.900 15.485 814.040 17.155 ;
        RECT 796.810 15.115 797.090 15.485 ;
        RECT 813.830 15.115 814.110 15.485 ;
        RECT 1174.080 2.400 1174.220 17.155 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
      LAYER via2 ;
        RECT 813.830 17.200 814.110 17.480 ;
        RECT 1174.010 17.200 1174.290 17.480 ;
        RECT 796.810 15.160 797.090 15.440 ;
        RECT 813.830 15.160 814.110 15.440 ;
      LAYER met3 ;
        RECT 813.805 17.490 814.135 17.505 ;
        RECT 1173.985 17.490 1174.315 17.505 ;
        RECT 813.805 17.190 1174.315 17.490 ;
        RECT 813.805 17.175 814.135 17.190 ;
        RECT 1173.985 17.175 1174.315 17.190 ;
        RECT 796.785 15.450 797.115 15.465 ;
        RECT 813.805 15.450 814.135 15.465 ;
        RECT 796.785 15.150 814.135 15.450 ;
        RECT 796.785 15.135 797.115 15.150 ;
        RECT 813.805 15.135 814.135 15.150 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 749.410 1593.480 749.730 1593.540 ;
        RECT 810.590 1593.480 810.910 1593.540 ;
        RECT 749.410 1593.340 810.910 1593.480 ;
        RECT 749.410 1593.280 749.730 1593.340 ;
        RECT 810.590 1593.280 810.910 1593.340 ;
      LAYER via ;
        RECT 749.440 1593.280 749.700 1593.540 ;
        RECT 810.620 1593.280 810.880 1593.540 ;
      LAYER met2 ;
        RECT 749.440 1600.000 749.720 1604.000 ;
        RECT 749.500 1593.570 749.640 1600.000 ;
        RECT 749.440 1593.250 749.700 1593.570 ;
        RECT 810.620 1593.250 810.880 1593.570 ;
        RECT 810.680 17.525 810.820 1593.250 ;
        RECT 1191.950 17.835 1192.230 18.205 ;
        RECT 810.610 17.155 810.890 17.525 ;
        RECT 1192.020 2.400 1192.160 17.835 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
      LAYER via2 ;
        RECT 1191.950 17.880 1192.230 18.160 ;
        RECT 810.610 17.200 810.890 17.480 ;
      LAYER met3 ;
        RECT 1191.925 18.170 1192.255 18.185 ;
        RECT 812.670 17.870 1192.255 18.170 ;
        RECT 810.585 17.490 810.915 17.505 ;
        RECT 812.670 17.490 812.970 17.870 ;
        RECT 1191.925 17.855 1192.255 17.870 ;
        RECT 810.585 17.190 812.970 17.490 ;
        RECT 810.585 17.175 810.915 17.190 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 757.690 43.760 758.010 43.820 ;
        RECT 1209.870 43.760 1210.190 43.820 ;
        RECT 757.690 43.620 1210.190 43.760 ;
        RECT 757.690 43.560 758.010 43.620 ;
        RECT 1209.870 43.560 1210.190 43.620 ;
      LAYER via ;
        RECT 757.720 43.560 757.980 43.820 ;
        RECT 1209.900 43.560 1210.160 43.820 ;
      LAYER met2 ;
        RECT 756.340 1600.450 756.620 1604.000 ;
        RECT 756.340 1600.310 757.920 1600.450 ;
        RECT 756.340 1600.000 756.620 1600.310 ;
        RECT 757.780 43.850 757.920 1600.310 ;
        RECT 757.720 43.530 757.980 43.850 ;
        RECT 1209.900 43.530 1210.160 43.850 ;
        RECT 1209.960 2.400 1210.100 43.530 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 765.050 44.100 765.370 44.160 ;
        RECT 1227.810 44.100 1228.130 44.160 ;
        RECT 765.050 43.960 1228.130 44.100 ;
        RECT 765.050 43.900 765.370 43.960 ;
        RECT 1227.810 43.900 1228.130 43.960 ;
      LAYER via ;
        RECT 765.080 43.900 765.340 44.160 ;
        RECT 1227.840 43.900 1228.100 44.160 ;
      LAYER met2 ;
        RECT 763.240 1600.450 763.520 1604.000 ;
        RECT 763.240 1600.310 765.280 1600.450 ;
        RECT 763.240 1600.000 763.520 1600.310 ;
        RECT 765.140 44.190 765.280 1600.310 ;
        RECT 765.080 43.870 765.340 44.190 ;
        RECT 1227.840 43.870 1228.100 44.190 ;
        RECT 1227.900 2.400 1228.040 43.870 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 771.490 48.180 771.810 48.240 ;
        RECT 1245.750 48.180 1246.070 48.240 ;
        RECT 771.490 48.040 1246.070 48.180 ;
        RECT 771.490 47.980 771.810 48.040 ;
        RECT 1245.750 47.980 1246.070 48.040 ;
      LAYER via ;
        RECT 771.520 47.980 771.780 48.240 ;
        RECT 1245.780 47.980 1246.040 48.240 ;
      LAYER met2 ;
        RECT 769.680 1600.450 769.960 1604.000 ;
        RECT 769.680 1600.310 771.720 1600.450 ;
        RECT 769.680 1600.000 769.960 1600.310 ;
        RECT 771.580 48.270 771.720 1600.310 ;
        RECT 771.520 47.950 771.780 48.270 ;
        RECT 1245.780 47.950 1246.040 48.270 ;
        RECT 1245.840 2.400 1245.980 47.950 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 776.550 1590.420 776.870 1590.480 ;
        RECT 778.850 1590.420 779.170 1590.480 ;
        RECT 776.550 1590.280 779.170 1590.420 ;
        RECT 776.550 1590.220 776.870 1590.280 ;
        RECT 778.850 1590.220 779.170 1590.280 ;
        RECT 778.850 47.500 779.170 47.560 ;
        RECT 1263.230 47.500 1263.550 47.560 ;
        RECT 778.850 47.360 1263.550 47.500 ;
        RECT 778.850 47.300 779.170 47.360 ;
        RECT 1263.230 47.300 1263.550 47.360 ;
      LAYER via ;
        RECT 776.580 1590.220 776.840 1590.480 ;
        RECT 778.880 1590.220 779.140 1590.480 ;
        RECT 778.880 47.300 779.140 47.560 ;
        RECT 1263.260 47.300 1263.520 47.560 ;
      LAYER met2 ;
        RECT 776.580 1600.000 776.860 1604.000 ;
        RECT 776.640 1590.510 776.780 1600.000 ;
        RECT 776.580 1590.190 776.840 1590.510 ;
        RECT 778.880 1590.190 779.140 1590.510 ;
        RECT 778.940 47.590 779.080 1590.190 ;
        RECT 778.880 47.270 779.140 47.590 ;
        RECT 1263.260 47.270 1263.520 47.590 ;
        RECT 1263.320 2.400 1263.460 47.270 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 783.450 1588.040 783.770 1588.100 ;
        RECT 785.290 1588.040 785.610 1588.100 ;
        RECT 783.450 1587.900 785.610 1588.040 ;
        RECT 783.450 1587.840 783.770 1587.900 ;
        RECT 785.290 1587.840 785.610 1587.900 ;
        RECT 785.290 47.160 785.610 47.220 ;
        RECT 1281.170 47.160 1281.490 47.220 ;
        RECT 785.290 47.020 1281.490 47.160 ;
        RECT 785.290 46.960 785.610 47.020 ;
        RECT 1281.170 46.960 1281.490 47.020 ;
      LAYER via ;
        RECT 783.480 1587.840 783.740 1588.100 ;
        RECT 785.320 1587.840 785.580 1588.100 ;
        RECT 785.320 46.960 785.580 47.220 ;
        RECT 1281.200 46.960 1281.460 47.220 ;
      LAYER met2 ;
        RECT 783.480 1600.000 783.760 1604.000 ;
        RECT 783.540 1588.130 783.680 1600.000 ;
        RECT 783.480 1587.810 783.740 1588.130 ;
        RECT 785.320 1587.810 785.580 1588.130 ;
        RECT 785.380 47.250 785.520 1587.810 ;
        RECT 785.320 46.930 785.580 47.250 ;
        RECT 1281.200 46.930 1281.460 47.250 ;
        RECT 1281.260 2.400 1281.400 46.930 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 789.890 1587.360 790.210 1587.420 ;
        RECT 792.650 1587.360 792.970 1587.420 ;
        RECT 789.890 1587.220 792.970 1587.360 ;
        RECT 789.890 1587.160 790.210 1587.220 ;
        RECT 792.650 1587.160 792.970 1587.220 ;
        RECT 792.650 31.180 792.970 31.240 ;
        RECT 1299.110 31.180 1299.430 31.240 ;
        RECT 792.650 31.040 1299.430 31.180 ;
        RECT 792.650 30.980 792.970 31.040 ;
        RECT 1299.110 30.980 1299.430 31.040 ;
      LAYER via ;
        RECT 789.920 1587.160 790.180 1587.420 ;
        RECT 792.680 1587.160 792.940 1587.420 ;
        RECT 792.680 30.980 792.940 31.240 ;
        RECT 1299.140 30.980 1299.400 31.240 ;
      LAYER met2 ;
        RECT 789.920 1600.000 790.200 1604.000 ;
        RECT 789.980 1587.450 790.120 1600.000 ;
        RECT 789.920 1587.130 790.180 1587.450 ;
        RECT 792.680 1587.130 792.940 1587.450 ;
        RECT 792.740 31.270 792.880 1587.130 ;
        RECT 792.680 30.950 792.940 31.270 ;
        RECT 1299.140 30.950 1299.400 31.270 ;
        RECT 1299.200 2.400 1299.340 30.950 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 796.790 1587.360 797.110 1587.420 ;
        RECT 799.550 1587.360 799.870 1587.420 ;
        RECT 796.790 1587.220 799.870 1587.360 ;
        RECT 796.790 1587.160 797.110 1587.220 ;
        RECT 799.550 1587.160 799.870 1587.220 ;
        RECT 799.550 30.840 799.870 30.900 ;
        RECT 1317.050 30.840 1317.370 30.900 ;
        RECT 799.550 30.700 1317.370 30.840 ;
        RECT 799.550 30.640 799.870 30.700 ;
        RECT 1317.050 30.640 1317.370 30.700 ;
      LAYER via ;
        RECT 796.820 1587.160 797.080 1587.420 ;
        RECT 799.580 1587.160 799.840 1587.420 ;
        RECT 799.580 30.640 799.840 30.900 ;
        RECT 1317.080 30.640 1317.340 30.900 ;
      LAYER met2 ;
        RECT 796.820 1600.000 797.100 1604.000 ;
        RECT 796.880 1587.450 797.020 1600.000 ;
        RECT 796.820 1587.130 797.080 1587.450 ;
        RECT 799.580 1587.130 799.840 1587.450 ;
        RECT 799.640 30.930 799.780 1587.130 ;
        RECT 799.580 30.610 799.840 30.930 ;
        RECT 1317.080 30.610 1317.340 30.930 ;
        RECT 1317.140 2.400 1317.280 30.610 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 803.690 1587.360 804.010 1587.420 ;
        RECT 806.450 1587.360 806.770 1587.420 ;
        RECT 803.690 1587.220 806.770 1587.360 ;
        RECT 803.690 1587.160 804.010 1587.220 ;
        RECT 806.450 1587.160 806.770 1587.220 ;
        RECT 806.450 34.920 806.770 34.980 ;
        RECT 1334.990 34.920 1335.310 34.980 ;
        RECT 806.450 34.780 1335.310 34.920 ;
        RECT 806.450 34.720 806.770 34.780 ;
        RECT 1334.990 34.720 1335.310 34.780 ;
      LAYER via ;
        RECT 803.720 1587.160 803.980 1587.420 ;
        RECT 806.480 1587.160 806.740 1587.420 ;
        RECT 806.480 34.720 806.740 34.980 ;
        RECT 1335.020 34.720 1335.280 34.980 ;
      LAYER met2 ;
        RECT 803.720 1600.000 804.000 1604.000 ;
        RECT 803.780 1587.450 803.920 1600.000 ;
        RECT 803.720 1587.130 803.980 1587.450 ;
        RECT 806.480 1587.130 806.740 1587.450 ;
        RECT 806.540 35.010 806.680 1587.130 ;
        RECT 806.480 34.690 806.740 35.010 ;
        RECT 1335.020 34.690 1335.280 35.010 ;
        RECT 1335.080 2.400 1335.220 34.690 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 665.765 15.385 665.935 17.255 ;
      LAYER mcon ;
        RECT 665.765 17.085 665.935 17.255 ;
      LAYER met1 ;
        RECT 561.270 1587.360 561.590 1587.420 ;
        RECT 564.950 1587.360 565.270 1587.420 ;
        RECT 561.270 1587.220 565.270 1587.360 ;
        RECT 561.270 1587.160 561.590 1587.220 ;
        RECT 564.950 1587.160 565.270 1587.220 ;
        RECT 564.950 17.240 565.270 17.300 ;
        RECT 665.705 17.240 665.995 17.285 ;
        RECT 564.950 17.100 665.995 17.240 ;
        RECT 564.950 17.040 565.270 17.100 ;
        RECT 665.705 17.055 665.995 17.100 ;
        RECT 665.705 15.540 665.995 15.585 ;
        RECT 692.370 15.540 692.690 15.600 ;
        RECT 665.705 15.400 692.690 15.540 ;
        RECT 665.705 15.355 665.995 15.400 ;
        RECT 692.370 15.340 692.690 15.400 ;
      LAYER via ;
        RECT 561.300 1587.160 561.560 1587.420 ;
        RECT 564.980 1587.160 565.240 1587.420 ;
        RECT 564.980 17.040 565.240 17.300 ;
        RECT 692.400 15.340 692.660 15.600 ;
      LAYER met2 ;
        RECT 561.300 1600.000 561.580 1604.000 ;
        RECT 561.360 1587.450 561.500 1600.000 ;
        RECT 561.300 1587.130 561.560 1587.450 ;
        RECT 564.980 1587.130 565.240 1587.450 ;
        RECT 565.040 17.330 565.180 1587.130 ;
        RECT 564.980 17.010 565.240 17.330 ;
        RECT 692.400 15.310 692.660 15.630 ;
        RECT 692.460 2.400 692.600 15.310 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 810.130 1587.700 810.450 1587.760 ;
        RECT 813.350 1587.700 813.670 1587.760 ;
        RECT 810.130 1587.560 813.670 1587.700 ;
        RECT 810.130 1587.500 810.450 1587.560 ;
        RECT 813.350 1587.500 813.670 1587.560 ;
        RECT 813.350 45.460 813.670 45.520 ;
        RECT 1352.470 45.460 1352.790 45.520 ;
        RECT 813.350 45.320 1352.790 45.460 ;
        RECT 813.350 45.260 813.670 45.320 ;
        RECT 1352.470 45.260 1352.790 45.320 ;
      LAYER via ;
        RECT 810.160 1587.500 810.420 1587.760 ;
        RECT 813.380 1587.500 813.640 1587.760 ;
        RECT 813.380 45.260 813.640 45.520 ;
        RECT 1352.500 45.260 1352.760 45.520 ;
      LAYER met2 ;
        RECT 810.160 1600.000 810.440 1604.000 ;
        RECT 810.220 1587.790 810.360 1600.000 ;
        RECT 810.160 1587.470 810.420 1587.790 ;
        RECT 813.380 1587.470 813.640 1587.790 ;
        RECT 813.440 45.550 813.580 1587.470 ;
        RECT 813.380 45.230 813.640 45.550 ;
        RECT 1352.500 45.230 1352.760 45.550 ;
        RECT 1352.560 2.400 1352.700 45.230 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 817.030 1587.700 817.350 1587.760 ;
        RECT 820.250 1587.700 820.570 1587.760 ;
        RECT 817.030 1587.560 820.570 1587.700 ;
        RECT 817.030 1587.500 817.350 1587.560 ;
        RECT 820.250 1587.500 820.570 1587.560 ;
        RECT 820.250 45.120 820.570 45.180 ;
        RECT 1370.410 45.120 1370.730 45.180 ;
        RECT 820.250 44.980 1370.730 45.120 ;
        RECT 820.250 44.920 820.570 44.980 ;
        RECT 1370.410 44.920 1370.730 44.980 ;
      LAYER via ;
        RECT 817.060 1587.500 817.320 1587.760 ;
        RECT 820.280 1587.500 820.540 1587.760 ;
        RECT 820.280 44.920 820.540 45.180 ;
        RECT 1370.440 44.920 1370.700 45.180 ;
      LAYER met2 ;
        RECT 817.060 1600.000 817.340 1604.000 ;
        RECT 817.120 1587.790 817.260 1600.000 ;
        RECT 817.060 1587.470 817.320 1587.790 ;
        RECT 820.280 1587.470 820.540 1587.790 ;
        RECT 820.340 45.210 820.480 1587.470 ;
        RECT 820.280 44.890 820.540 45.210 ;
        RECT 1370.440 44.890 1370.700 45.210 ;
        RECT 1370.500 2.400 1370.640 44.890 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 823.470 1587.360 823.790 1587.420 ;
        RECT 827.150 1587.360 827.470 1587.420 ;
        RECT 823.470 1587.220 827.470 1587.360 ;
        RECT 823.470 1587.160 823.790 1587.220 ;
        RECT 827.150 1587.160 827.470 1587.220 ;
        RECT 827.150 44.780 827.470 44.840 ;
        RECT 1388.350 44.780 1388.670 44.840 ;
        RECT 827.150 44.640 1388.670 44.780 ;
        RECT 827.150 44.580 827.470 44.640 ;
        RECT 1388.350 44.580 1388.670 44.640 ;
      LAYER via ;
        RECT 823.500 1587.160 823.760 1587.420 ;
        RECT 827.180 1587.160 827.440 1587.420 ;
        RECT 827.180 44.580 827.440 44.840 ;
        RECT 1388.380 44.580 1388.640 44.840 ;
      LAYER met2 ;
        RECT 823.500 1600.000 823.780 1604.000 ;
        RECT 823.560 1587.450 823.700 1600.000 ;
        RECT 823.500 1587.130 823.760 1587.450 ;
        RECT 827.180 1587.130 827.440 1587.450 ;
        RECT 827.240 44.870 827.380 1587.130 ;
        RECT 827.180 44.550 827.440 44.870 ;
        RECT 1388.380 44.550 1388.640 44.870 ;
        RECT 1388.440 2.400 1388.580 44.550 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 830.370 1588.040 830.690 1588.100 ;
        RECT 834.050 1588.040 834.370 1588.100 ;
        RECT 830.370 1587.900 834.370 1588.040 ;
        RECT 830.370 1587.840 830.690 1587.900 ;
        RECT 834.050 1587.840 834.370 1587.900 ;
        RECT 834.050 41.720 834.370 41.780 ;
        RECT 1406.290 41.720 1406.610 41.780 ;
        RECT 834.050 41.580 1406.610 41.720 ;
        RECT 834.050 41.520 834.370 41.580 ;
        RECT 1406.290 41.520 1406.610 41.580 ;
      LAYER via ;
        RECT 830.400 1587.840 830.660 1588.100 ;
        RECT 834.080 1587.840 834.340 1588.100 ;
        RECT 834.080 41.520 834.340 41.780 ;
        RECT 1406.320 41.520 1406.580 41.780 ;
      LAYER met2 ;
        RECT 830.400 1600.000 830.680 1604.000 ;
        RECT 830.460 1588.130 830.600 1600.000 ;
        RECT 830.400 1587.810 830.660 1588.130 ;
        RECT 834.080 1587.810 834.340 1588.130 ;
        RECT 834.140 41.810 834.280 1587.810 ;
        RECT 834.080 41.490 834.340 41.810 ;
        RECT 1406.320 41.490 1406.580 41.810 ;
        RECT 1406.380 2.400 1406.520 41.490 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 837.270 1590.420 837.590 1590.480 ;
        RECT 840.950 1590.420 841.270 1590.480 ;
        RECT 837.270 1590.280 841.270 1590.420 ;
        RECT 837.270 1590.220 837.590 1590.280 ;
        RECT 840.950 1590.220 841.270 1590.280 ;
        RECT 840.950 42.060 841.270 42.120 ;
        RECT 1423.770 42.060 1424.090 42.120 ;
        RECT 840.950 41.920 1424.090 42.060 ;
        RECT 840.950 41.860 841.270 41.920 ;
        RECT 1423.770 41.860 1424.090 41.920 ;
      LAYER via ;
        RECT 837.300 1590.220 837.560 1590.480 ;
        RECT 840.980 1590.220 841.240 1590.480 ;
        RECT 840.980 41.860 841.240 42.120 ;
        RECT 1423.800 41.860 1424.060 42.120 ;
      LAYER met2 ;
        RECT 837.300 1600.000 837.580 1604.000 ;
        RECT 837.360 1590.510 837.500 1600.000 ;
        RECT 837.300 1590.190 837.560 1590.510 ;
        RECT 840.980 1590.190 841.240 1590.510 ;
        RECT 841.040 42.150 841.180 1590.190 ;
        RECT 840.980 41.830 841.240 42.150 ;
        RECT 1423.800 41.830 1424.060 42.150 ;
        RECT 1423.860 2.400 1424.000 41.830 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 843.710 1590.420 844.030 1590.480 ;
        RECT 847.850 1590.420 848.170 1590.480 ;
        RECT 843.710 1590.280 848.170 1590.420 ;
        RECT 843.710 1590.220 844.030 1590.280 ;
        RECT 847.850 1590.220 848.170 1590.280 ;
        RECT 847.850 42.400 848.170 42.460 ;
        RECT 1441.710 42.400 1442.030 42.460 ;
        RECT 847.850 42.260 1442.030 42.400 ;
        RECT 847.850 42.200 848.170 42.260 ;
        RECT 1441.710 42.200 1442.030 42.260 ;
      LAYER via ;
        RECT 843.740 1590.220 844.000 1590.480 ;
        RECT 847.880 1590.220 848.140 1590.480 ;
        RECT 847.880 42.200 848.140 42.460 ;
        RECT 1441.740 42.200 1442.000 42.460 ;
      LAYER met2 ;
        RECT 843.740 1600.000 844.020 1604.000 ;
        RECT 843.800 1590.510 843.940 1600.000 ;
        RECT 843.740 1590.190 844.000 1590.510 ;
        RECT 847.880 1590.190 848.140 1590.510 ;
        RECT 847.940 42.490 848.080 1590.190 ;
        RECT 847.880 42.170 848.140 42.490 ;
        RECT 1441.740 42.170 1442.000 42.490 ;
        RECT 1441.800 2.400 1441.940 42.170 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 850.610 1589.740 850.930 1589.800 ;
        RECT 855.210 1589.740 855.530 1589.800 ;
        RECT 850.610 1589.600 855.530 1589.740 ;
        RECT 850.610 1589.540 850.930 1589.600 ;
        RECT 855.210 1589.540 855.530 1589.600 ;
        RECT 855.210 42.740 855.530 42.800 ;
        RECT 1459.650 42.740 1459.970 42.800 ;
        RECT 855.210 42.600 1459.970 42.740 ;
        RECT 855.210 42.540 855.530 42.600 ;
        RECT 1459.650 42.540 1459.970 42.600 ;
      LAYER via ;
        RECT 850.640 1589.540 850.900 1589.800 ;
        RECT 855.240 1589.540 855.500 1589.800 ;
        RECT 855.240 42.540 855.500 42.800 ;
        RECT 1459.680 42.540 1459.940 42.800 ;
      LAYER met2 ;
        RECT 850.640 1600.000 850.920 1604.000 ;
        RECT 850.700 1589.830 850.840 1600.000 ;
        RECT 850.640 1589.510 850.900 1589.830 ;
        RECT 855.240 1589.510 855.500 1589.830 ;
        RECT 855.300 42.830 855.440 1589.510 ;
        RECT 855.240 42.510 855.500 42.830 ;
        RECT 1459.680 42.510 1459.940 42.830 ;
        RECT 1459.740 2.400 1459.880 42.510 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 857.510 1587.360 857.830 1587.420 ;
        RECT 861.650 1587.360 861.970 1587.420 ;
        RECT 857.510 1587.220 861.970 1587.360 ;
        RECT 857.510 1587.160 857.830 1587.220 ;
        RECT 861.650 1587.160 861.970 1587.220 ;
        RECT 861.650 69.600 861.970 69.660 ;
        RECT 1476.670 69.600 1476.990 69.660 ;
        RECT 861.650 69.460 1476.990 69.600 ;
        RECT 861.650 69.400 861.970 69.460 ;
        RECT 1476.670 69.400 1476.990 69.460 ;
        RECT 1476.670 2.960 1476.990 3.020 ;
        RECT 1477.590 2.960 1477.910 3.020 ;
        RECT 1476.670 2.820 1477.910 2.960 ;
        RECT 1476.670 2.760 1476.990 2.820 ;
        RECT 1477.590 2.760 1477.910 2.820 ;
      LAYER via ;
        RECT 857.540 1587.160 857.800 1587.420 ;
        RECT 861.680 1587.160 861.940 1587.420 ;
        RECT 861.680 69.400 861.940 69.660 ;
        RECT 1476.700 69.400 1476.960 69.660 ;
        RECT 1476.700 2.760 1476.960 3.020 ;
        RECT 1477.620 2.760 1477.880 3.020 ;
      LAYER met2 ;
        RECT 857.540 1600.000 857.820 1604.000 ;
        RECT 857.600 1587.450 857.740 1600.000 ;
        RECT 857.540 1587.130 857.800 1587.450 ;
        RECT 861.680 1587.130 861.940 1587.450 ;
        RECT 861.740 69.690 861.880 1587.130 ;
        RECT 861.680 69.370 861.940 69.690 ;
        RECT 1476.700 69.370 1476.960 69.690 ;
        RECT 1476.760 3.050 1476.900 69.370 ;
        RECT 1476.700 2.730 1476.960 3.050 ;
        RECT 1477.620 2.730 1477.880 3.050 ;
        RECT 1477.680 2.400 1477.820 2.730 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 863.950 1589.740 864.270 1589.800 ;
        RECT 868.550 1589.740 868.870 1589.800 ;
        RECT 863.950 1589.600 868.870 1589.740 ;
        RECT 863.950 1589.540 864.270 1589.600 ;
        RECT 868.550 1589.540 868.870 1589.600 ;
        RECT 868.550 70.280 868.870 70.340 ;
        RECT 1490.470 70.280 1490.790 70.340 ;
        RECT 868.550 70.140 1490.790 70.280 ;
        RECT 868.550 70.080 868.870 70.140 ;
        RECT 1490.470 70.080 1490.790 70.140 ;
        RECT 1490.470 2.960 1490.790 3.020 ;
        RECT 1495.530 2.960 1495.850 3.020 ;
        RECT 1490.470 2.820 1495.850 2.960 ;
        RECT 1490.470 2.760 1490.790 2.820 ;
        RECT 1495.530 2.760 1495.850 2.820 ;
      LAYER via ;
        RECT 863.980 1589.540 864.240 1589.800 ;
        RECT 868.580 1589.540 868.840 1589.800 ;
        RECT 868.580 70.080 868.840 70.340 ;
        RECT 1490.500 70.080 1490.760 70.340 ;
        RECT 1490.500 2.760 1490.760 3.020 ;
        RECT 1495.560 2.760 1495.820 3.020 ;
      LAYER met2 ;
        RECT 863.980 1600.000 864.260 1604.000 ;
        RECT 864.040 1589.830 864.180 1600.000 ;
        RECT 863.980 1589.510 864.240 1589.830 ;
        RECT 868.580 1589.510 868.840 1589.830 ;
        RECT 868.640 70.370 868.780 1589.510 ;
        RECT 868.580 70.050 868.840 70.370 ;
        RECT 1490.500 70.050 1490.760 70.370 ;
        RECT 1490.560 3.050 1490.700 70.050 ;
        RECT 1490.500 2.730 1490.760 3.050 ;
        RECT 1495.560 2.730 1495.820 3.050 ;
        RECT 1495.620 2.400 1495.760 2.730 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 870.850 1589.740 871.170 1589.800 ;
        RECT 875.450 1589.740 875.770 1589.800 ;
        RECT 870.850 1589.600 875.770 1589.740 ;
        RECT 870.850 1589.540 871.170 1589.600 ;
        RECT 875.450 1589.540 875.770 1589.600 ;
        RECT 875.450 70.620 875.770 70.680 ;
        RECT 1511.170 70.620 1511.490 70.680 ;
        RECT 875.450 70.480 1511.490 70.620 ;
        RECT 875.450 70.420 875.770 70.480 ;
        RECT 1511.170 70.420 1511.490 70.480 ;
      LAYER via ;
        RECT 870.880 1589.540 871.140 1589.800 ;
        RECT 875.480 1589.540 875.740 1589.800 ;
        RECT 875.480 70.420 875.740 70.680 ;
        RECT 1511.200 70.420 1511.460 70.680 ;
      LAYER met2 ;
        RECT 870.880 1600.000 871.160 1604.000 ;
        RECT 870.940 1589.830 871.080 1600.000 ;
        RECT 870.880 1589.510 871.140 1589.830 ;
        RECT 875.480 1589.510 875.740 1589.830 ;
        RECT 875.540 70.710 875.680 1589.510 ;
        RECT 875.480 70.390 875.740 70.710 ;
        RECT 1511.200 70.390 1511.460 70.710 ;
        RECT 1511.260 3.130 1511.400 70.390 ;
        RECT 1511.260 2.990 1513.240 3.130 ;
        RECT 1513.100 2.400 1513.240 2.990 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 567.710 1587.360 568.030 1587.420 ;
        RECT 571.850 1587.360 572.170 1587.420 ;
        RECT 567.710 1587.220 572.170 1587.360 ;
        RECT 567.710 1587.160 568.030 1587.220 ;
        RECT 571.850 1587.160 572.170 1587.220 ;
        RECT 571.850 15.200 572.170 15.260 ;
        RECT 710.310 15.200 710.630 15.260 ;
        RECT 571.850 15.060 710.630 15.200 ;
        RECT 571.850 15.000 572.170 15.060 ;
        RECT 710.310 15.000 710.630 15.060 ;
      LAYER via ;
        RECT 567.740 1587.160 568.000 1587.420 ;
        RECT 571.880 1587.160 572.140 1587.420 ;
        RECT 571.880 15.000 572.140 15.260 ;
        RECT 710.340 15.000 710.600 15.260 ;
      LAYER met2 ;
        RECT 567.740 1600.000 568.020 1604.000 ;
        RECT 567.800 1587.450 567.940 1600.000 ;
        RECT 567.740 1587.130 568.000 1587.450 ;
        RECT 571.880 1587.130 572.140 1587.450 ;
        RECT 571.940 15.290 572.080 1587.130 ;
        RECT 571.880 14.970 572.140 15.290 ;
        RECT 710.340 14.970 710.600 15.290 ;
        RECT 710.400 2.400 710.540 14.970 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 877.750 1587.360 878.070 1587.420 ;
        RECT 882.350 1587.360 882.670 1587.420 ;
        RECT 877.750 1587.220 882.670 1587.360 ;
        RECT 877.750 1587.160 878.070 1587.220 ;
        RECT 882.350 1587.160 882.670 1587.220 ;
        RECT 882.350 70.960 882.670 71.020 ;
        RECT 1524.970 70.960 1525.290 71.020 ;
        RECT 882.350 70.820 1525.290 70.960 ;
        RECT 882.350 70.760 882.670 70.820 ;
        RECT 1524.970 70.760 1525.290 70.820 ;
        RECT 1524.970 14.520 1525.290 14.580 ;
        RECT 1530.950 14.520 1531.270 14.580 ;
        RECT 1524.970 14.380 1531.270 14.520 ;
        RECT 1524.970 14.320 1525.290 14.380 ;
        RECT 1530.950 14.320 1531.270 14.380 ;
      LAYER via ;
        RECT 877.780 1587.160 878.040 1587.420 ;
        RECT 882.380 1587.160 882.640 1587.420 ;
        RECT 882.380 70.760 882.640 71.020 ;
        RECT 1525.000 70.760 1525.260 71.020 ;
        RECT 1525.000 14.320 1525.260 14.580 ;
        RECT 1530.980 14.320 1531.240 14.580 ;
      LAYER met2 ;
        RECT 877.780 1600.000 878.060 1604.000 ;
        RECT 877.840 1587.450 877.980 1600.000 ;
        RECT 877.780 1587.130 878.040 1587.450 ;
        RECT 882.380 1587.130 882.640 1587.450 ;
        RECT 882.440 71.050 882.580 1587.130 ;
        RECT 882.380 70.730 882.640 71.050 ;
        RECT 1525.000 70.730 1525.260 71.050 ;
        RECT 1525.060 14.610 1525.200 70.730 ;
        RECT 1525.000 14.290 1525.260 14.610 ;
        RECT 1530.980 14.290 1531.240 14.610 ;
        RECT 1531.040 2.400 1531.180 14.290 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 884.190 1589.740 884.510 1589.800 ;
        RECT 889.250 1589.740 889.570 1589.800 ;
        RECT 884.190 1589.600 889.570 1589.740 ;
        RECT 884.190 1589.540 884.510 1589.600 ;
        RECT 889.250 1589.540 889.570 1589.600 ;
        RECT 889.250 48.520 889.570 48.580 ;
        RECT 1545.670 48.520 1545.990 48.580 ;
        RECT 889.250 48.380 1545.990 48.520 ;
        RECT 889.250 48.320 889.570 48.380 ;
        RECT 1545.670 48.320 1545.990 48.380 ;
        RECT 1545.670 2.960 1545.990 3.020 ;
        RECT 1548.890 2.960 1549.210 3.020 ;
        RECT 1545.670 2.820 1549.210 2.960 ;
        RECT 1545.670 2.760 1545.990 2.820 ;
        RECT 1548.890 2.760 1549.210 2.820 ;
      LAYER via ;
        RECT 884.220 1589.540 884.480 1589.800 ;
        RECT 889.280 1589.540 889.540 1589.800 ;
        RECT 889.280 48.320 889.540 48.580 ;
        RECT 1545.700 48.320 1545.960 48.580 ;
        RECT 1545.700 2.760 1545.960 3.020 ;
        RECT 1548.920 2.760 1549.180 3.020 ;
      LAYER met2 ;
        RECT 884.220 1600.000 884.500 1604.000 ;
        RECT 884.280 1589.830 884.420 1600.000 ;
        RECT 884.220 1589.510 884.480 1589.830 ;
        RECT 889.280 1589.510 889.540 1589.830 ;
        RECT 889.340 48.610 889.480 1589.510 ;
        RECT 889.280 48.290 889.540 48.610 ;
        RECT 1545.700 48.290 1545.960 48.610 ;
        RECT 1545.760 3.050 1545.900 48.290 ;
        RECT 1545.700 2.730 1545.960 3.050 ;
        RECT 1548.920 2.730 1549.180 3.050 ;
        RECT 1548.980 2.400 1549.120 2.730 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 891.090 1589.740 891.410 1589.800 ;
        RECT 896.150 1589.740 896.470 1589.800 ;
        RECT 891.090 1589.600 896.470 1589.740 ;
        RECT 891.090 1589.540 891.410 1589.600 ;
        RECT 896.150 1589.540 896.470 1589.600 ;
        RECT 896.150 48.860 896.470 48.920 ;
        RECT 1566.370 48.860 1566.690 48.920 ;
        RECT 896.150 48.720 1566.690 48.860 ;
        RECT 896.150 48.660 896.470 48.720 ;
        RECT 1566.370 48.660 1566.690 48.720 ;
      LAYER via ;
        RECT 891.120 1589.540 891.380 1589.800 ;
        RECT 896.180 1589.540 896.440 1589.800 ;
        RECT 896.180 48.660 896.440 48.920 ;
        RECT 1566.400 48.660 1566.660 48.920 ;
      LAYER met2 ;
        RECT 891.120 1600.000 891.400 1604.000 ;
        RECT 891.180 1589.830 891.320 1600.000 ;
        RECT 891.120 1589.510 891.380 1589.830 ;
        RECT 896.180 1589.510 896.440 1589.830 ;
        RECT 896.240 48.950 896.380 1589.510 ;
        RECT 896.180 48.630 896.440 48.950 ;
        RECT 1566.400 48.630 1566.660 48.950 ;
        RECT 1566.460 3.130 1566.600 48.630 ;
        RECT 1566.460 2.990 1567.060 3.130 ;
        RECT 1566.920 2.400 1567.060 2.990 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 897.530 1589.740 897.850 1589.800 ;
        RECT 903.050 1589.740 903.370 1589.800 ;
        RECT 897.530 1589.600 903.370 1589.740 ;
        RECT 897.530 1589.540 897.850 1589.600 ;
        RECT 903.050 1589.540 903.370 1589.600 ;
        RECT 903.050 49.200 903.370 49.260 ;
        RECT 1580.170 49.200 1580.490 49.260 ;
        RECT 903.050 49.060 1580.490 49.200 ;
        RECT 903.050 49.000 903.370 49.060 ;
        RECT 1580.170 49.000 1580.490 49.060 ;
        RECT 1580.170 2.960 1580.490 3.020 ;
        RECT 1584.770 2.960 1585.090 3.020 ;
        RECT 1580.170 2.820 1585.090 2.960 ;
        RECT 1580.170 2.760 1580.490 2.820 ;
        RECT 1584.770 2.760 1585.090 2.820 ;
      LAYER via ;
        RECT 897.560 1589.540 897.820 1589.800 ;
        RECT 903.080 1589.540 903.340 1589.800 ;
        RECT 903.080 49.000 903.340 49.260 ;
        RECT 1580.200 49.000 1580.460 49.260 ;
        RECT 1580.200 2.760 1580.460 3.020 ;
        RECT 1584.800 2.760 1585.060 3.020 ;
      LAYER met2 ;
        RECT 897.560 1600.000 897.840 1604.000 ;
        RECT 897.620 1589.830 897.760 1600.000 ;
        RECT 897.560 1589.510 897.820 1589.830 ;
        RECT 903.080 1589.510 903.340 1589.830 ;
        RECT 903.140 49.290 903.280 1589.510 ;
        RECT 903.080 48.970 903.340 49.290 ;
        RECT 1580.200 48.970 1580.460 49.290 ;
        RECT 1580.260 3.050 1580.400 48.970 ;
        RECT 1580.200 2.730 1580.460 3.050 ;
        RECT 1584.800 2.730 1585.060 3.050 ;
        RECT 1584.860 2.400 1585.000 2.730 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 904.430 1589.060 904.750 1589.120 ;
        RECT 909.950 1589.060 910.270 1589.120 ;
        RECT 904.430 1588.920 910.270 1589.060 ;
        RECT 904.430 1588.860 904.750 1588.920 ;
        RECT 909.950 1588.860 910.270 1588.920 ;
        RECT 909.950 49.540 910.270 49.600 ;
        RECT 1600.870 49.540 1601.190 49.600 ;
        RECT 909.950 49.400 1601.190 49.540 ;
        RECT 909.950 49.340 910.270 49.400 ;
        RECT 1600.870 49.340 1601.190 49.400 ;
      LAYER via ;
        RECT 904.460 1588.860 904.720 1589.120 ;
        RECT 909.980 1588.860 910.240 1589.120 ;
        RECT 909.980 49.340 910.240 49.600 ;
        RECT 1600.900 49.340 1601.160 49.600 ;
      LAYER met2 ;
        RECT 904.460 1600.000 904.740 1604.000 ;
        RECT 904.520 1589.150 904.660 1600.000 ;
        RECT 904.460 1588.830 904.720 1589.150 ;
        RECT 909.980 1588.830 910.240 1589.150 ;
        RECT 910.040 49.630 910.180 1588.830 ;
        RECT 909.980 49.310 910.240 49.630 ;
        RECT 1600.900 49.310 1601.160 49.630 ;
        RECT 1600.960 3.130 1601.100 49.310 ;
        RECT 1600.960 2.990 1602.480 3.130 ;
        RECT 1602.340 2.400 1602.480 2.990 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 911.330 1590.080 911.650 1590.140 ;
        RECT 916.850 1590.080 917.170 1590.140 ;
        RECT 911.330 1589.940 917.170 1590.080 ;
        RECT 911.330 1589.880 911.650 1589.940 ;
        RECT 916.850 1589.880 917.170 1589.940 ;
        RECT 916.850 49.880 917.170 49.940 ;
        RECT 1614.670 49.880 1614.990 49.940 ;
        RECT 916.850 49.740 1614.990 49.880 ;
        RECT 916.850 49.680 917.170 49.740 ;
        RECT 1614.670 49.680 1614.990 49.740 ;
        RECT 1614.670 2.960 1614.990 3.020 ;
        RECT 1620.190 2.960 1620.510 3.020 ;
        RECT 1614.670 2.820 1620.510 2.960 ;
        RECT 1614.670 2.760 1614.990 2.820 ;
        RECT 1620.190 2.760 1620.510 2.820 ;
      LAYER via ;
        RECT 911.360 1589.880 911.620 1590.140 ;
        RECT 916.880 1589.880 917.140 1590.140 ;
        RECT 916.880 49.680 917.140 49.940 ;
        RECT 1614.700 49.680 1614.960 49.940 ;
        RECT 1614.700 2.760 1614.960 3.020 ;
        RECT 1620.220 2.760 1620.480 3.020 ;
      LAYER met2 ;
        RECT 911.360 1600.000 911.640 1604.000 ;
        RECT 911.420 1590.170 911.560 1600.000 ;
        RECT 911.360 1589.850 911.620 1590.170 ;
        RECT 916.880 1589.850 917.140 1590.170 ;
        RECT 916.940 49.970 917.080 1589.850 ;
        RECT 916.880 49.650 917.140 49.970 ;
        RECT 1614.700 49.650 1614.960 49.970 ;
        RECT 1614.760 3.050 1614.900 49.650 ;
        RECT 1614.700 2.730 1614.960 3.050 ;
        RECT 1620.220 2.730 1620.480 3.050 ;
        RECT 1620.280 2.400 1620.420 2.730 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 917.770 1590.080 918.090 1590.140 ;
        RECT 923.750 1590.080 924.070 1590.140 ;
        RECT 917.770 1589.940 924.070 1590.080 ;
        RECT 917.770 1589.880 918.090 1589.940 ;
        RECT 923.750 1589.880 924.070 1589.940 ;
        RECT 923.750 50.220 924.070 50.280 ;
        RECT 1635.370 50.220 1635.690 50.280 ;
        RECT 923.750 50.080 1635.690 50.220 ;
        RECT 923.750 50.020 924.070 50.080 ;
        RECT 1635.370 50.020 1635.690 50.080 ;
        RECT 1635.370 2.960 1635.690 3.020 ;
        RECT 1638.130 2.960 1638.450 3.020 ;
        RECT 1635.370 2.820 1638.450 2.960 ;
        RECT 1635.370 2.760 1635.690 2.820 ;
        RECT 1638.130 2.760 1638.450 2.820 ;
      LAYER via ;
        RECT 917.800 1589.880 918.060 1590.140 ;
        RECT 923.780 1589.880 924.040 1590.140 ;
        RECT 923.780 50.020 924.040 50.280 ;
        RECT 1635.400 50.020 1635.660 50.280 ;
        RECT 1635.400 2.760 1635.660 3.020 ;
        RECT 1638.160 2.760 1638.420 3.020 ;
      LAYER met2 ;
        RECT 917.800 1600.000 918.080 1604.000 ;
        RECT 917.860 1590.170 918.000 1600.000 ;
        RECT 917.800 1589.850 918.060 1590.170 ;
        RECT 923.780 1589.850 924.040 1590.170 ;
        RECT 923.840 50.310 923.980 1589.850 ;
        RECT 923.780 49.990 924.040 50.310 ;
        RECT 1635.400 49.990 1635.660 50.310 ;
        RECT 1635.460 3.050 1635.600 49.990 ;
        RECT 1635.400 2.730 1635.660 3.050 ;
        RECT 1638.160 2.730 1638.420 3.050 ;
        RECT 1638.220 2.400 1638.360 2.730 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.670 1590.080 924.990 1590.140 ;
        RECT 930.650 1590.080 930.970 1590.140 ;
        RECT 924.670 1589.940 930.970 1590.080 ;
        RECT 924.670 1589.880 924.990 1589.940 ;
        RECT 930.650 1589.880 930.970 1589.940 ;
        RECT 930.650 50.560 930.970 50.620 ;
        RECT 1656.530 50.560 1656.850 50.620 ;
        RECT 930.650 50.420 1656.850 50.560 ;
        RECT 930.650 50.360 930.970 50.420 ;
        RECT 1656.530 50.360 1656.850 50.420 ;
      LAYER via ;
        RECT 924.700 1589.880 924.960 1590.140 ;
        RECT 930.680 1589.880 930.940 1590.140 ;
        RECT 930.680 50.360 930.940 50.620 ;
        RECT 1656.560 50.360 1656.820 50.620 ;
      LAYER met2 ;
        RECT 924.700 1600.000 924.980 1604.000 ;
        RECT 924.760 1590.170 924.900 1600.000 ;
        RECT 924.700 1589.850 924.960 1590.170 ;
        RECT 930.680 1589.850 930.940 1590.170 ;
        RECT 930.740 50.650 930.880 1589.850 ;
        RECT 930.680 50.330 930.940 50.650 ;
        RECT 1656.560 50.330 1656.820 50.650 ;
        RECT 1656.620 3.130 1656.760 50.330 ;
        RECT 1656.160 2.990 1656.760 3.130 ;
        RECT 1656.160 2.400 1656.300 2.990 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 931.570 1590.080 931.890 1590.140 ;
        RECT 937.090 1590.080 937.410 1590.140 ;
        RECT 931.570 1589.940 937.410 1590.080 ;
        RECT 931.570 1589.880 931.890 1589.940 ;
        RECT 937.090 1589.880 937.410 1589.940 ;
        RECT 937.090 50.900 937.410 50.960 ;
        RECT 1669.870 50.900 1670.190 50.960 ;
        RECT 937.090 50.760 1670.190 50.900 ;
        RECT 937.090 50.700 937.410 50.760 ;
        RECT 1669.870 50.700 1670.190 50.760 ;
        RECT 1669.870 2.960 1670.190 3.020 ;
        RECT 1673.550 2.960 1673.870 3.020 ;
        RECT 1669.870 2.820 1673.870 2.960 ;
        RECT 1669.870 2.760 1670.190 2.820 ;
        RECT 1673.550 2.760 1673.870 2.820 ;
      LAYER via ;
        RECT 931.600 1589.880 931.860 1590.140 ;
        RECT 937.120 1589.880 937.380 1590.140 ;
        RECT 937.120 50.700 937.380 50.960 ;
        RECT 1669.900 50.700 1670.160 50.960 ;
        RECT 1669.900 2.760 1670.160 3.020 ;
        RECT 1673.580 2.760 1673.840 3.020 ;
      LAYER met2 ;
        RECT 931.600 1600.000 931.880 1604.000 ;
        RECT 931.660 1590.170 931.800 1600.000 ;
        RECT 931.600 1589.850 931.860 1590.170 ;
        RECT 937.120 1589.850 937.380 1590.170 ;
        RECT 937.180 50.990 937.320 1589.850 ;
        RECT 937.120 50.670 937.380 50.990 ;
        RECT 1669.900 50.670 1670.160 50.990 ;
        RECT 1669.960 3.050 1670.100 50.670 ;
        RECT 1669.900 2.730 1670.160 3.050 ;
        RECT 1673.580 2.730 1673.840 3.050 ;
        RECT 1673.640 2.400 1673.780 2.730 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 937.550 51.240 937.870 51.300 ;
        RECT 1690.570 51.240 1690.890 51.300 ;
        RECT 937.550 51.100 1690.890 51.240 ;
        RECT 937.550 51.040 937.870 51.100 ;
        RECT 1690.570 51.040 1690.890 51.100 ;
      LAYER via ;
        RECT 937.580 51.040 937.840 51.300 ;
        RECT 1690.600 51.040 1690.860 51.300 ;
      LAYER met2 ;
        RECT 938.040 1600.450 938.320 1604.000 ;
        RECT 937.640 1600.310 938.320 1600.450 ;
        RECT 937.640 51.330 937.780 1600.310 ;
        RECT 938.040 1600.000 938.320 1600.310 ;
        RECT 937.580 51.010 937.840 51.330 ;
        RECT 1690.600 51.010 1690.860 51.330 ;
        RECT 1690.660 3.130 1690.800 51.010 ;
        RECT 1690.660 2.990 1691.720 3.130 ;
        RECT 1691.580 2.400 1691.720 2.990 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 574.610 1587.360 574.930 1587.420 ;
        RECT 579.210 1587.360 579.530 1587.420 ;
        RECT 574.610 1587.220 579.530 1587.360 ;
        RECT 574.610 1587.160 574.930 1587.220 ;
        RECT 579.210 1587.160 579.530 1587.220 ;
        RECT 579.210 16.220 579.530 16.280 ;
        RECT 728.250 16.220 728.570 16.280 ;
        RECT 579.210 16.080 728.570 16.220 ;
        RECT 579.210 16.020 579.530 16.080 ;
        RECT 728.250 16.020 728.570 16.080 ;
      LAYER via ;
        RECT 574.640 1587.160 574.900 1587.420 ;
        RECT 579.240 1587.160 579.500 1587.420 ;
        RECT 579.240 16.020 579.500 16.280 ;
        RECT 728.280 16.020 728.540 16.280 ;
      LAYER met2 ;
        RECT 574.640 1600.000 574.920 1604.000 ;
        RECT 574.700 1587.450 574.840 1600.000 ;
        RECT 574.640 1587.130 574.900 1587.450 ;
        RECT 579.240 1587.130 579.500 1587.450 ;
        RECT 579.300 16.310 579.440 1587.130 ;
        RECT 579.240 15.990 579.500 16.310 ;
        RECT 728.280 15.990 728.540 16.310 ;
        RECT 728.340 2.400 728.480 15.990 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 944.450 54.980 944.770 55.040 ;
        RECT 1704.370 54.980 1704.690 55.040 ;
        RECT 944.450 54.840 1704.690 54.980 ;
        RECT 944.450 54.780 944.770 54.840 ;
        RECT 1704.370 54.780 1704.690 54.840 ;
        RECT 1704.370 2.960 1704.690 3.020 ;
        RECT 1709.430 2.960 1709.750 3.020 ;
        RECT 1704.370 2.820 1709.750 2.960 ;
        RECT 1704.370 2.760 1704.690 2.820 ;
        RECT 1709.430 2.760 1709.750 2.820 ;
      LAYER via ;
        RECT 944.480 54.780 944.740 55.040 ;
        RECT 1704.400 54.780 1704.660 55.040 ;
        RECT 1704.400 2.760 1704.660 3.020 ;
        RECT 1709.460 2.760 1709.720 3.020 ;
      LAYER met2 ;
        RECT 944.940 1600.450 945.220 1604.000 ;
        RECT 944.540 1600.310 945.220 1600.450 ;
        RECT 944.540 55.070 944.680 1600.310 ;
        RECT 944.940 1600.000 945.220 1600.310 ;
        RECT 944.480 54.750 944.740 55.070 ;
        RECT 1704.400 54.750 1704.660 55.070 ;
        RECT 1704.460 3.050 1704.600 54.750 ;
        RECT 1704.400 2.730 1704.660 3.050 ;
        RECT 1709.460 2.730 1709.720 3.050 ;
        RECT 1709.520 2.400 1709.660 2.730 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 951.350 54.640 951.670 54.700 ;
        RECT 1725.070 54.640 1725.390 54.700 ;
        RECT 951.350 54.500 1725.390 54.640 ;
        RECT 951.350 54.440 951.670 54.500 ;
        RECT 1725.070 54.440 1725.390 54.500 ;
      LAYER via ;
        RECT 951.380 54.440 951.640 54.700 ;
        RECT 1725.100 54.440 1725.360 54.700 ;
      LAYER met2 ;
        RECT 951.840 1600.450 952.120 1604.000 ;
        RECT 951.440 1600.310 952.120 1600.450 ;
        RECT 951.440 54.730 951.580 1600.310 ;
        RECT 951.840 1600.000 952.120 1600.310 ;
        RECT 951.380 54.410 951.640 54.730 ;
        RECT 1725.100 54.410 1725.360 54.730 ;
        RECT 1725.160 16.730 1725.300 54.410 ;
        RECT 1725.160 16.590 1727.600 16.730 ;
        RECT 1727.460 2.400 1727.600 16.590 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 957.790 54.300 958.110 54.360 ;
        RECT 1738.870 54.300 1739.190 54.360 ;
        RECT 957.790 54.160 1739.190 54.300 ;
        RECT 957.790 54.100 958.110 54.160 ;
        RECT 1738.870 54.100 1739.190 54.160 ;
        RECT 1738.870 16.220 1739.190 16.280 ;
        RECT 1745.310 16.220 1745.630 16.280 ;
        RECT 1738.870 16.080 1745.630 16.220 ;
        RECT 1738.870 16.020 1739.190 16.080 ;
        RECT 1745.310 16.020 1745.630 16.080 ;
      LAYER via ;
        RECT 957.820 54.100 958.080 54.360 ;
        RECT 1738.900 54.100 1739.160 54.360 ;
        RECT 1738.900 16.020 1739.160 16.280 ;
        RECT 1745.340 16.020 1745.600 16.280 ;
      LAYER met2 ;
        RECT 958.280 1600.450 958.560 1604.000 ;
        RECT 957.880 1600.310 958.560 1600.450 ;
        RECT 957.880 54.390 958.020 1600.310 ;
        RECT 958.280 1600.000 958.560 1600.310 ;
        RECT 957.820 54.070 958.080 54.390 ;
        RECT 1738.900 54.070 1739.160 54.390 ;
        RECT 1738.960 16.310 1739.100 54.070 ;
        RECT 1738.900 15.990 1739.160 16.310 ;
        RECT 1745.340 15.990 1745.600 16.310 ;
        RECT 1745.400 2.400 1745.540 15.990 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 965.150 53.960 965.470 54.020 ;
        RECT 1759.570 53.960 1759.890 54.020 ;
        RECT 965.150 53.820 1759.890 53.960 ;
        RECT 965.150 53.760 965.470 53.820 ;
        RECT 1759.570 53.760 1759.890 53.820 ;
      LAYER via ;
        RECT 965.180 53.760 965.440 54.020 ;
        RECT 1759.600 53.760 1759.860 54.020 ;
      LAYER met2 ;
        RECT 965.180 1600.000 965.460 1604.000 ;
        RECT 965.240 54.050 965.380 1600.000 ;
        RECT 965.180 53.730 965.440 54.050 ;
        RECT 1759.600 53.730 1759.860 54.050 ;
        RECT 1759.660 16.730 1759.800 53.730 ;
        RECT 1759.660 16.590 1763.020 16.730 ;
        RECT 1762.880 2.400 1763.020 16.590 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 972.050 53.620 972.370 53.680 ;
        RECT 1780.730 53.620 1781.050 53.680 ;
        RECT 972.050 53.480 1781.050 53.620 ;
        RECT 972.050 53.420 972.370 53.480 ;
        RECT 1780.730 53.420 1781.050 53.480 ;
      LAYER via ;
        RECT 972.080 53.420 972.340 53.680 ;
        RECT 1780.760 53.420 1781.020 53.680 ;
      LAYER met2 ;
        RECT 971.620 1600.450 971.900 1604.000 ;
        RECT 971.620 1600.310 972.280 1600.450 ;
        RECT 971.620 1600.000 971.900 1600.310 ;
        RECT 972.140 53.710 972.280 1600.310 ;
        RECT 972.080 53.390 972.340 53.710 ;
        RECT 1780.760 53.390 1781.020 53.710 ;
        RECT 1780.820 2.400 1780.960 53.390 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 978.950 53.280 979.270 53.340 ;
        RECT 1794.070 53.280 1794.390 53.340 ;
        RECT 978.950 53.140 1794.390 53.280 ;
        RECT 978.950 53.080 979.270 53.140 ;
        RECT 1794.070 53.080 1794.390 53.140 ;
      LAYER via ;
        RECT 978.980 53.080 979.240 53.340 ;
        RECT 1794.100 53.080 1794.360 53.340 ;
      LAYER met2 ;
        RECT 978.520 1600.450 978.800 1604.000 ;
        RECT 978.520 1600.310 979.180 1600.450 ;
        RECT 978.520 1600.000 978.800 1600.310 ;
        RECT 979.040 53.370 979.180 1600.310 ;
        RECT 978.980 53.050 979.240 53.370 ;
        RECT 1794.100 53.050 1794.360 53.370 ;
        RECT 1794.160 16.730 1794.300 53.050 ;
        RECT 1794.160 16.590 1798.900 16.730 ;
        RECT 1798.760 2.400 1798.900 16.590 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 985.390 52.940 985.710 53.000 ;
        RECT 1814.770 52.940 1815.090 53.000 ;
        RECT 985.390 52.800 1815.090 52.940 ;
        RECT 985.390 52.740 985.710 52.800 ;
        RECT 1814.770 52.740 1815.090 52.800 ;
      LAYER via ;
        RECT 985.420 52.740 985.680 53.000 ;
        RECT 1814.800 52.740 1815.060 53.000 ;
      LAYER met2 ;
        RECT 985.420 1600.000 985.700 1604.000 ;
        RECT 985.480 53.030 985.620 1600.000 ;
        RECT 985.420 52.710 985.680 53.030 ;
        RECT 1814.800 52.710 1815.060 53.030 ;
        RECT 1814.860 16.730 1815.000 52.710 ;
        RECT 1814.860 16.590 1816.840 16.730 ;
        RECT 1816.700 2.400 1816.840 16.590 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 992.750 52.600 993.070 52.660 ;
        RECT 1828.570 52.600 1828.890 52.660 ;
        RECT 992.750 52.460 1828.890 52.600 ;
        RECT 992.750 52.400 993.070 52.460 ;
        RECT 1828.570 52.400 1828.890 52.460 ;
        RECT 1828.570 7.040 1828.890 7.100 ;
        RECT 1834.550 7.040 1834.870 7.100 ;
        RECT 1828.570 6.900 1834.870 7.040 ;
        RECT 1828.570 6.840 1828.890 6.900 ;
        RECT 1834.550 6.840 1834.870 6.900 ;
      LAYER via ;
        RECT 992.780 52.400 993.040 52.660 ;
        RECT 1828.600 52.400 1828.860 52.660 ;
        RECT 1828.600 6.840 1828.860 7.100 ;
        RECT 1834.580 6.840 1834.840 7.100 ;
      LAYER met2 ;
        RECT 991.860 1600.450 992.140 1604.000 ;
        RECT 991.860 1600.310 992.980 1600.450 ;
        RECT 991.860 1600.000 992.140 1600.310 ;
        RECT 992.840 52.690 992.980 1600.310 ;
        RECT 992.780 52.370 993.040 52.690 ;
        RECT 1828.600 52.370 1828.860 52.690 ;
        RECT 1828.660 7.130 1828.800 52.370 ;
        RECT 1828.600 6.810 1828.860 7.130 ;
        RECT 1834.580 6.810 1834.840 7.130 ;
        RECT 1834.640 2.400 1834.780 6.810 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 999.650 52.260 999.970 52.320 ;
        RECT 1849.270 52.260 1849.590 52.320 ;
        RECT 999.650 52.120 1849.590 52.260 ;
        RECT 999.650 52.060 999.970 52.120 ;
        RECT 1849.270 52.060 1849.590 52.120 ;
        RECT 1849.270 2.960 1849.590 3.020 ;
        RECT 1852.030 2.960 1852.350 3.020 ;
        RECT 1849.270 2.820 1852.350 2.960 ;
        RECT 1849.270 2.760 1849.590 2.820 ;
        RECT 1852.030 2.760 1852.350 2.820 ;
      LAYER via ;
        RECT 999.680 52.060 999.940 52.320 ;
        RECT 1849.300 52.060 1849.560 52.320 ;
        RECT 1849.300 2.760 1849.560 3.020 ;
        RECT 1852.060 2.760 1852.320 3.020 ;
      LAYER met2 ;
        RECT 998.760 1600.450 999.040 1604.000 ;
        RECT 998.760 1600.310 999.880 1600.450 ;
        RECT 998.760 1600.000 999.040 1600.310 ;
        RECT 999.740 52.350 999.880 1600.310 ;
        RECT 999.680 52.030 999.940 52.350 ;
        RECT 1849.300 52.030 1849.560 52.350 ;
        RECT 1849.360 3.050 1849.500 52.030 ;
        RECT 1849.300 2.730 1849.560 3.050 ;
        RECT 1852.060 2.730 1852.320 3.050 ;
        RECT 1852.120 2.400 1852.260 2.730 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1006.550 51.920 1006.870 51.980 ;
        RECT 1870.430 51.920 1870.750 51.980 ;
        RECT 1006.550 51.780 1870.750 51.920 ;
        RECT 1006.550 51.720 1006.870 51.780 ;
        RECT 1870.430 51.720 1870.750 51.780 ;
      LAYER via ;
        RECT 1006.580 51.720 1006.840 51.980 ;
        RECT 1870.460 51.720 1870.720 51.980 ;
      LAYER met2 ;
        RECT 1005.660 1600.450 1005.940 1604.000 ;
        RECT 1005.660 1600.310 1006.780 1600.450 ;
        RECT 1005.660 1600.000 1005.940 1600.310 ;
        RECT 1006.640 52.010 1006.780 1600.310 ;
        RECT 1006.580 51.690 1006.840 52.010 ;
        RECT 1870.460 51.690 1870.720 52.010 ;
        RECT 1870.520 7.210 1870.660 51.690 ;
        RECT 1870.060 7.070 1870.660 7.210 ;
        RECT 1870.060 2.400 1870.200 7.070 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 714.065 15.045 714.235 16.575 ;
      LAYER mcon ;
        RECT 714.065 16.405 714.235 16.575 ;
      LAYER met1 ;
        RECT 581.050 1587.360 581.370 1587.420 ;
        RECT 584.730 1587.360 585.050 1587.420 ;
        RECT 581.050 1587.220 585.050 1587.360 ;
        RECT 581.050 1587.160 581.370 1587.220 ;
        RECT 584.730 1587.160 585.050 1587.220 ;
        RECT 584.730 16.560 585.050 16.620 ;
        RECT 714.005 16.560 714.295 16.605 ;
        RECT 584.730 16.420 714.295 16.560 ;
        RECT 584.730 16.360 585.050 16.420 ;
        RECT 714.005 16.375 714.295 16.420 ;
        RECT 714.005 15.200 714.295 15.245 ;
        RECT 746.190 15.200 746.510 15.260 ;
        RECT 714.005 15.060 746.510 15.200 ;
        RECT 714.005 15.015 714.295 15.060 ;
        RECT 746.190 15.000 746.510 15.060 ;
      LAYER via ;
        RECT 581.080 1587.160 581.340 1587.420 ;
        RECT 584.760 1587.160 585.020 1587.420 ;
        RECT 584.760 16.360 585.020 16.620 ;
        RECT 746.220 15.000 746.480 15.260 ;
      LAYER met2 ;
        RECT 581.080 1600.000 581.360 1604.000 ;
        RECT 581.140 1587.450 581.280 1600.000 ;
        RECT 581.080 1587.130 581.340 1587.450 ;
        RECT 584.760 1587.130 585.020 1587.450 ;
        RECT 584.820 1579.370 584.960 1587.130 ;
        RECT 584.820 1579.230 585.880 1579.370 ;
        RECT 585.740 34.410 585.880 1579.230 ;
        RECT 584.820 34.270 585.880 34.410 ;
        RECT 584.820 16.650 584.960 34.270 ;
        RECT 584.760 16.330 585.020 16.650 ;
        RECT 746.220 14.970 746.480 15.290 ;
        RECT 746.280 2.400 746.420 14.970 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.450 51.580 1013.770 51.640 ;
        RECT 1883.770 51.580 1884.090 51.640 ;
        RECT 1013.450 51.440 1884.090 51.580 ;
        RECT 1013.450 51.380 1013.770 51.440 ;
        RECT 1883.770 51.380 1884.090 51.440 ;
        RECT 1883.770 2.960 1884.090 3.020 ;
        RECT 1887.910 2.960 1888.230 3.020 ;
        RECT 1883.770 2.820 1888.230 2.960 ;
        RECT 1883.770 2.760 1884.090 2.820 ;
        RECT 1887.910 2.760 1888.230 2.820 ;
      LAYER via ;
        RECT 1013.480 51.380 1013.740 51.640 ;
        RECT 1883.800 51.380 1884.060 51.640 ;
        RECT 1883.800 2.760 1884.060 3.020 ;
        RECT 1887.940 2.760 1888.200 3.020 ;
      LAYER met2 ;
        RECT 1012.100 1600.450 1012.380 1604.000 ;
        RECT 1012.100 1600.310 1013.680 1600.450 ;
        RECT 1012.100 1600.000 1012.380 1600.310 ;
        RECT 1013.540 51.670 1013.680 1600.310 ;
        RECT 1013.480 51.350 1013.740 51.670 ;
        RECT 1883.800 51.350 1884.060 51.670 ;
        RECT 1883.860 3.050 1884.000 51.350 ;
        RECT 1883.800 2.730 1884.060 3.050 ;
        RECT 1887.940 2.730 1888.200 3.050 ;
        RECT 1888.000 2.400 1888.140 2.730 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1019.000 1600.450 1019.280 1604.000 ;
        RECT 1019.000 1600.310 1020.580 1600.450 ;
        RECT 1019.000 1600.000 1019.280 1600.310 ;
        RECT 1020.440 54.245 1020.580 1600.310 ;
        RECT 1020.370 53.875 1020.650 54.245 ;
        RECT 1904.490 53.875 1904.770 54.245 ;
        RECT 1904.560 3.130 1904.700 53.875 ;
        RECT 1904.560 2.990 1906.080 3.130 ;
        RECT 1905.940 2.400 1906.080 2.990 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
      LAYER via2 ;
        RECT 1020.370 53.920 1020.650 54.200 ;
        RECT 1904.490 53.920 1904.770 54.200 ;
      LAYER met3 ;
        RECT 1020.345 54.210 1020.675 54.225 ;
        RECT 1904.465 54.210 1904.795 54.225 ;
        RECT 1020.345 53.910 1904.795 54.210 ;
        RECT 1020.345 53.895 1020.675 53.910 ;
        RECT 1904.465 53.895 1904.795 53.910 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1025.900 1600.450 1026.180 1604.000 ;
        RECT 1025.900 1600.310 1027.480 1600.450 ;
        RECT 1025.900 1600.000 1026.180 1600.310 ;
        RECT 1027.340 53.565 1027.480 1600.310 ;
        RECT 1027.270 53.195 1027.550 53.565 ;
        RECT 1918.290 53.195 1918.570 53.565 ;
        RECT 1918.360 16.730 1918.500 53.195 ;
        RECT 1918.360 16.590 1923.560 16.730 ;
        RECT 1923.420 2.400 1923.560 16.590 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
      LAYER via2 ;
        RECT 1027.270 53.240 1027.550 53.520 ;
        RECT 1918.290 53.240 1918.570 53.520 ;
      LAYER met3 ;
        RECT 1027.245 53.530 1027.575 53.545 ;
        RECT 1918.265 53.530 1918.595 53.545 ;
        RECT 1027.245 53.230 1918.595 53.530 ;
        RECT 1027.245 53.215 1027.575 53.230 ;
        RECT 1918.265 53.215 1918.595 53.230 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1033.690 43.080 1034.010 43.140 ;
        RECT 1941.270 43.080 1941.590 43.140 ;
        RECT 1033.690 42.940 1941.590 43.080 ;
        RECT 1033.690 42.880 1034.010 42.940 ;
        RECT 1941.270 42.880 1941.590 42.940 ;
      LAYER via ;
        RECT 1033.720 42.880 1033.980 43.140 ;
        RECT 1941.300 42.880 1941.560 43.140 ;
      LAYER met2 ;
        RECT 1032.340 1600.450 1032.620 1604.000 ;
        RECT 1032.340 1600.310 1033.920 1600.450 ;
        RECT 1032.340 1600.000 1032.620 1600.310 ;
        RECT 1033.780 43.170 1033.920 1600.310 ;
        RECT 1033.720 42.850 1033.980 43.170 ;
        RECT 1941.300 42.850 1941.560 43.170 ;
        RECT 1941.360 2.400 1941.500 42.850 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1039.210 1589.740 1039.530 1589.800 ;
        RECT 1041.510 1589.740 1041.830 1589.800 ;
        RECT 1039.210 1589.600 1041.830 1589.740 ;
        RECT 1039.210 1589.540 1039.530 1589.600 ;
        RECT 1041.510 1589.540 1041.830 1589.600 ;
        RECT 1953.230 16.900 1953.550 16.960 ;
        RECT 1959.210 16.900 1959.530 16.960 ;
        RECT 1953.230 16.760 1959.530 16.900 ;
        RECT 1953.230 16.700 1953.550 16.760 ;
        RECT 1959.210 16.700 1959.530 16.760 ;
      LAYER via ;
        RECT 1039.240 1589.540 1039.500 1589.800 ;
        RECT 1041.540 1589.540 1041.800 1589.800 ;
        RECT 1953.260 16.700 1953.520 16.960 ;
        RECT 1959.240 16.700 1959.500 16.960 ;
      LAYER met2 ;
        RECT 1039.240 1600.000 1039.520 1604.000 ;
        RECT 1039.300 1589.830 1039.440 1600.000 ;
        RECT 1039.240 1589.510 1039.500 1589.830 ;
        RECT 1041.540 1589.510 1041.800 1589.830 ;
        RECT 1041.600 52.885 1041.740 1589.510 ;
        RECT 1041.530 52.515 1041.810 52.885 ;
        RECT 1953.250 52.515 1953.530 52.885 ;
        RECT 1953.320 16.990 1953.460 52.515 ;
        RECT 1953.260 16.670 1953.520 16.990 ;
        RECT 1959.240 16.670 1959.500 16.990 ;
        RECT 1959.300 2.400 1959.440 16.670 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
      LAYER via2 ;
        RECT 1041.530 52.560 1041.810 52.840 ;
        RECT 1953.250 52.560 1953.530 52.840 ;
      LAYER met3 ;
        RECT 1041.505 52.850 1041.835 52.865 ;
        RECT 1953.225 52.850 1953.555 52.865 ;
        RECT 1041.505 52.550 1953.555 52.850 ;
        RECT 1041.505 52.535 1041.835 52.550 ;
        RECT 1953.225 52.535 1953.555 52.550 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1046.140 1600.450 1046.420 1604.000 ;
        RECT 1046.140 1600.310 1047.720 1600.450 ;
        RECT 1046.140 1600.000 1046.420 1600.310 ;
        RECT 1047.580 52.205 1047.720 1600.310 ;
        RECT 1047.510 51.835 1047.790 52.205 ;
        RECT 1973.490 51.835 1973.770 52.205 ;
        RECT 1973.560 16.730 1973.700 51.835 ;
        RECT 1973.560 16.590 1977.380 16.730 ;
        RECT 1977.240 2.400 1977.380 16.590 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
      LAYER via2 ;
        RECT 1047.510 51.880 1047.790 52.160 ;
        RECT 1973.490 51.880 1973.770 52.160 ;
      LAYER met3 ;
        RECT 1047.485 52.170 1047.815 52.185 ;
        RECT 1973.465 52.170 1973.795 52.185 ;
        RECT 1047.485 51.870 1973.795 52.170 ;
        RECT 1047.485 51.855 1047.815 51.870 ;
        RECT 1973.465 51.855 1973.795 51.870 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1052.580 1601.130 1052.860 1604.000 ;
        RECT 1052.580 1600.990 1054.620 1601.130 ;
        RECT 1052.580 1600.000 1052.860 1600.990 ;
        RECT 1054.480 1590.250 1054.620 1600.990 ;
        RECT 1054.480 1590.110 1055.080 1590.250 ;
        RECT 1054.940 51.525 1055.080 1590.110 ;
        RECT 1054.870 51.155 1055.150 51.525 ;
        RECT 1994.190 51.155 1994.470 51.525 ;
        RECT 1994.260 16.730 1994.400 51.155 ;
        RECT 1994.260 16.590 1995.320 16.730 ;
        RECT 1995.180 2.400 1995.320 16.590 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
      LAYER via2 ;
        RECT 1054.870 51.200 1055.150 51.480 ;
        RECT 1994.190 51.200 1994.470 51.480 ;
      LAYER met3 ;
        RECT 1054.845 51.490 1055.175 51.505 ;
        RECT 1994.165 51.490 1994.495 51.505 ;
        RECT 1054.845 51.190 1994.495 51.490 ;
        RECT 1054.845 51.175 1055.175 51.190 ;
        RECT 1994.165 51.175 1994.495 51.190 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1061.290 71.640 1061.610 71.700 ;
        RECT 2007.970 71.640 2008.290 71.700 ;
        RECT 1061.290 71.500 2008.290 71.640 ;
        RECT 1061.290 71.440 1061.610 71.500 ;
        RECT 2007.970 71.440 2008.290 71.500 ;
      LAYER via ;
        RECT 1061.320 71.440 1061.580 71.700 ;
        RECT 2008.000 71.440 2008.260 71.700 ;
      LAYER met2 ;
        RECT 1059.480 1600.450 1059.760 1604.000 ;
        RECT 1059.480 1600.310 1061.520 1600.450 ;
        RECT 1059.480 1600.000 1059.760 1600.310 ;
        RECT 1061.380 71.730 1061.520 1600.310 ;
        RECT 1061.320 71.410 1061.580 71.730 ;
        RECT 2008.000 71.410 2008.260 71.730 ;
        RECT 2008.060 16.730 2008.200 71.410 ;
        RECT 2008.060 16.590 2012.800 16.730 ;
        RECT 2012.660 2.400 2012.800 16.590 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1065.890 1590.080 1066.210 1590.140 ;
        RECT 1068.650 1590.080 1068.970 1590.140 ;
        RECT 1065.890 1589.940 1068.970 1590.080 ;
        RECT 1065.890 1589.880 1066.210 1589.940 ;
        RECT 1068.650 1589.880 1068.970 1589.940 ;
        RECT 1068.650 71.980 1068.970 72.040 ;
        RECT 2028.670 71.980 2028.990 72.040 ;
        RECT 1068.650 71.840 2028.990 71.980 ;
        RECT 1068.650 71.780 1068.970 71.840 ;
        RECT 2028.670 71.780 2028.990 71.840 ;
      LAYER via ;
        RECT 1065.920 1589.880 1066.180 1590.140 ;
        RECT 1068.680 1589.880 1068.940 1590.140 ;
        RECT 1068.680 71.780 1068.940 72.040 ;
        RECT 2028.700 71.780 2028.960 72.040 ;
      LAYER met2 ;
        RECT 1065.920 1600.000 1066.200 1604.000 ;
        RECT 1065.980 1590.170 1066.120 1600.000 ;
        RECT 1065.920 1589.850 1066.180 1590.170 ;
        RECT 1068.680 1589.850 1068.940 1590.170 ;
        RECT 1068.740 72.070 1068.880 1589.850 ;
        RECT 1068.680 71.750 1068.940 72.070 ;
        RECT 2028.700 71.750 2028.960 72.070 ;
        RECT 2028.760 17.410 2028.900 71.750 ;
        RECT 2028.760 17.270 2030.740 17.410 ;
        RECT 2030.600 2.400 2030.740 17.270 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1075.090 75.720 1075.410 75.780 ;
        RECT 2042.470 75.720 2042.790 75.780 ;
        RECT 1075.090 75.580 2042.790 75.720 ;
        RECT 1075.090 75.520 1075.410 75.580 ;
        RECT 2042.470 75.520 2042.790 75.580 ;
        RECT 2042.470 17.920 2042.790 17.980 ;
        RECT 2048.450 17.920 2048.770 17.980 ;
        RECT 2042.470 17.780 2048.770 17.920 ;
        RECT 2042.470 17.720 2042.790 17.780 ;
        RECT 2048.450 17.720 2048.770 17.780 ;
      LAYER via ;
        RECT 1075.120 75.520 1075.380 75.780 ;
        RECT 2042.500 75.520 2042.760 75.780 ;
        RECT 2042.500 17.720 2042.760 17.980 ;
        RECT 2048.480 17.720 2048.740 17.980 ;
      LAYER met2 ;
        RECT 1072.820 1601.130 1073.100 1604.000 ;
        RECT 1072.820 1600.990 1074.860 1601.130 ;
        RECT 1072.820 1600.000 1073.100 1600.990 ;
        RECT 1074.720 1590.250 1074.860 1600.990 ;
        RECT 1074.720 1590.110 1075.320 1590.250 ;
        RECT 1075.180 75.810 1075.320 1590.110 ;
        RECT 1075.120 75.490 1075.380 75.810 ;
        RECT 2042.500 75.490 2042.760 75.810 ;
        RECT 2042.560 18.010 2042.700 75.490 ;
        RECT 2042.500 17.690 2042.760 18.010 ;
        RECT 2048.480 17.690 2048.740 18.010 ;
        RECT 2048.540 2.400 2048.680 17.690 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 717.285 15.725 717.455 20.315 ;
      LAYER mcon ;
        RECT 717.285 20.145 717.455 20.315 ;
      LAYER met1 ;
        RECT 589.330 1579.540 589.650 1579.600 ;
        RECT 592.550 1579.540 592.870 1579.600 ;
        RECT 589.330 1579.400 592.870 1579.540 ;
        RECT 589.330 1579.340 589.650 1579.400 ;
        RECT 592.550 1579.340 592.870 1579.400 ;
        RECT 592.550 20.300 592.870 20.360 ;
        RECT 717.225 20.300 717.515 20.345 ;
        RECT 592.550 20.160 717.515 20.300 ;
        RECT 592.550 20.100 592.870 20.160 ;
        RECT 717.225 20.115 717.515 20.160 ;
        RECT 717.225 15.880 717.515 15.925 ;
        RECT 763.670 15.880 763.990 15.940 ;
        RECT 717.225 15.740 763.990 15.880 ;
        RECT 717.225 15.695 717.515 15.740 ;
        RECT 763.670 15.680 763.990 15.740 ;
      LAYER via ;
        RECT 589.360 1579.340 589.620 1579.600 ;
        RECT 592.580 1579.340 592.840 1579.600 ;
        RECT 592.580 20.100 592.840 20.360 ;
        RECT 763.700 15.680 763.960 15.940 ;
      LAYER met2 ;
        RECT 587.980 1600.450 588.260 1604.000 ;
        RECT 587.980 1600.310 589.560 1600.450 ;
        RECT 587.980 1600.000 588.260 1600.310 ;
        RECT 589.420 1579.630 589.560 1600.310 ;
        RECT 589.360 1579.310 589.620 1579.630 ;
        RECT 592.580 1579.310 592.840 1579.630 ;
        RECT 592.640 20.390 592.780 1579.310 ;
        RECT 592.580 20.070 592.840 20.390 ;
        RECT 763.700 15.650 763.960 15.970 ;
        RECT 763.760 2.400 763.900 15.650 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1079.690 1590.080 1080.010 1590.140 ;
        RECT 1082.450 1590.080 1082.770 1590.140 ;
        RECT 1079.690 1589.940 1082.770 1590.080 ;
        RECT 1079.690 1589.880 1080.010 1589.940 ;
        RECT 1082.450 1589.880 1082.770 1589.940 ;
        RECT 1082.450 55.660 1082.770 55.720 ;
        RECT 2063.170 55.660 2063.490 55.720 ;
        RECT 1082.450 55.520 2063.490 55.660 ;
        RECT 1082.450 55.460 1082.770 55.520 ;
        RECT 2063.170 55.460 2063.490 55.520 ;
        RECT 2063.170 2.960 2063.490 3.020 ;
        RECT 2066.390 2.960 2066.710 3.020 ;
        RECT 2063.170 2.820 2066.710 2.960 ;
        RECT 2063.170 2.760 2063.490 2.820 ;
        RECT 2066.390 2.760 2066.710 2.820 ;
      LAYER via ;
        RECT 1079.720 1589.880 1079.980 1590.140 ;
        RECT 1082.480 1589.880 1082.740 1590.140 ;
        RECT 1082.480 55.460 1082.740 55.720 ;
        RECT 2063.200 55.460 2063.460 55.720 ;
        RECT 2063.200 2.760 2063.460 3.020 ;
        RECT 2066.420 2.760 2066.680 3.020 ;
      LAYER met2 ;
        RECT 1079.720 1600.000 1080.000 1604.000 ;
        RECT 1079.780 1590.170 1079.920 1600.000 ;
        RECT 1079.720 1589.850 1079.980 1590.170 ;
        RECT 1082.480 1589.850 1082.740 1590.170 ;
        RECT 1082.540 55.750 1082.680 1589.850 ;
        RECT 1082.480 55.430 1082.740 55.750 ;
        RECT 2063.200 55.430 2063.460 55.750 ;
        RECT 2063.260 3.050 2063.400 55.430 ;
        RECT 2063.200 2.730 2063.460 3.050 ;
        RECT 2066.420 2.730 2066.680 3.050 ;
        RECT 2066.480 2.400 2066.620 2.730 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1086.130 1589.740 1086.450 1589.800 ;
        RECT 1089.350 1589.740 1089.670 1589.800 ;
        RECT 1086.130 1589.600 1089.670 1589.740 ;
        RECT 1086.130 1589.540 1086.450 1589.600 ;
        RECT 1089.350 1589.540 1089.670 1589.600 ;
        RECT 1089.350 56.000 1089.670 56.060 ;
        RECT 2084.330 56.000 2084.650 56.060 ;
        RECT 1089.350 55.860 2084.650 56.000 ;
        RECT 1089.350 55.800 1089.670 55.860 ;
        RECT 2084.330 55.800 2084.650 55.860 ;
      LAYER via ;
        RECT 1086.160 1589.540 1086.420 1589.800 ;
        RECT 1089.380 1589.540 1089.640 1589.800 ;
        RECT 1089.380 55.800 1089.640 56.060 ;
        RECT 2084.360 55.800 2084.620 56.060 ;
      LAYER met2 ;
        RECT 1086.160 1600.000 1086.440 1604.000 ;
        RECT 1086.220 1589.830 1086.360 1600.000 ;
        RECT 1086.160 1589.510 1086.420 1589.830 ;
        RECT 1089.380 1589.510 1089.640 1589.830 ;
        RECT 1089.440 56.090 1089.580 1589.510 ;
        RECT 1089.380 55.770 1089.640 56.090 ;
        RECT 2084.360 55.770 2084.620 56.090 ;
        RECT 2084.420 2.400 2084.560 55.770 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1093.030 1588.040 1093.350 1588.100 ;
        RECT 1096.250 1588.040 1096.570 1588.100 ;
        RECT 1093.030 1587.900 1096.570 1588.040 ;
        RECT 1093.030 1587.840 1093.350 1587.900 ;
        RECT 1096.250 1587.840 1096.570 1587.900 ;
        RECT 1096.250 56.340 1096.570 56.400 ;
        RECT 2097.670 56.340 2097.990 56.400 ;
        RECT 1096.250 56.200 2097.990 56.340 ;
        RECT 1096.250 56.140 1096.570 56.200 ;
        RECT 2097.670 56.140 2097.990 56.200 ;
        RECT 2097.670 2.960 2097.990 3.020 ;
        RECT 2101.810 2.960 2102.130 3.020 ;
        RECT 2097.670 2.820 2102.130 2.960 ;
        RECT 2097.670 2.760 2097.990 2.820 ;
        RECT 2101.810 2.760 2102.130 2.820 ;
      LAYER via ;
        RECT 1093.060 1587.840 1093.320 1588.100 ;
        RECT 1096.280 1587.840 1096.540 1588.100 ;
        RECT 1096.280 56.140 1096.540 56.400 ;
        RECT 2097.700 56.140 2097.960 56.400 ;
        RECT 2097.700 2.760 2097.960 3.020 ;
        RECT 2101.840 2.760 2102.100 3.020 ;
      LAYER met2 ;
        RECT 1093.060 1600.000 1093.340 1604.000 ;
        RECT 1093.120 1588.130 1093.260 1600.000 ;
        RECT 1093.060 1587.810 1093.320 1588.130 ;
        RECT 1096.280 1587.810 1096.540 1588.130 ;
        RECT 1096.340 56.430 1096.480 1587.810 ;
        RECT 1096.280 56.110 1096.540 56.430 ;
        RECT 2097.700 56.110 2097.960 56.430 ;
        RECT 2097.760 3.050 2097.900 56.110 ;
        RECT 2097.700 2.730 2097.960 3.050 ;
        RECT 2101.840 2.730 2102.100 3.050 ;
        RECT 2101.900 2.400 2102.040 2.730 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1099.930 1589.740 1100.250 1589.800 ;
        RECT 1103.150 1589.740 1103.470 1589.800 ;
        RECT 1099.930 1589.600 1103.470 1589.740 ;
        RECT 1099.930 1589.540 1100.250 1589.600 ;
        RECT 1103.150 1589.540 1103.470 1589.600 ;
        RECT 1103.150 56.680 1103.470 56.740 ;
        RECT 2118.370 56.680 2118.690 56.740 ;
        RECT 1103.150 56.540 2118.690 56.680 ;
        RECT 1103.150 56.480 1103.470 56.540 ;
        RECT 2118.370 56.480 2118.690 56.540 ;
        RECT 2118.370 2.960 2118.690 3.020 ;
        RECT 2119.750 2.960 2120.070 3.020 ;
        RECT 2118.370 2.820 2120.070 2.960 ;
        RECT 2118.370 2.760 2118.690 2.820 ;
        RECT 2119.750 2.760 2120.070 2.820 ;
      LAYER via ;
        RECT 1099.960 1589.540 1100.220 1589.800 ;
        RECT 1103.180 1589.540 1103.440 1589.800 ;
        RECT 1103.180 56.480 1103.440 56.740 ;
        RECT 2118.400 56.480 2118.660 56.740 ;
        RECT 2118.400 2.760 2118.660 3.020 ;
        RECT 2119.780 2.760 2120.040 3.020 ;
      LAYER met2 ;
        RECT 1099.960 1600.000 1100.240 1604.000 ;
        RECT 1100.020 1589.830 1100.160 1600.000 ;
        RECT 1099.960 1589.510 1100.220 1589.830 ;
        RECT 1103.180 1589.510 1103.440 1589.830 ;
        RECT 1103.240 56.770 1103.380 1589.510 ;
        RECT 1103.180 56.450 1103.440 56.770 ;
        RECT 2118.400 56.450 2118.660 56.770 ;
        RECT 2118.460 3.050 2118.600 56.450 ;
        RECT 2118.400 2.730 2118.660 3.050 ;
        RECT 2119.780 2.730 2120.040 3.050 ;
        RECT 2119.840 2.400 2119.980 2.730 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1106.370 1588.040 1106.690 1588.100 ;
        RECT 1109.590 1588.040 1109.910 1588.100 ;
        RECT 1106.370 1587.900 1109.910 1588.040 ;
        RECT 1106.370 1587.840 1106.690 1587.900 ;
        RECT 1109.590 1587.840 1109.910 1587.900 ;
        RECT 1109.590 57.020 1109.910 57.080 ;
        RECT 2132.170 57.020 2132.490 57.080 ;
        RECT 1109.590 56.880 2132.490 57.020 ;
        RECT 1109.590 56.820 1109.910 56.880 ;
        RECT 2132.170 56.820 2132.490 56.880 ;
        RECT 2132.170 2.960 2132.490 3.020 ;
        RECT 2137.690 2.960 2138.010 3.020 ;
        RECT 2132.170 2.820 2138.010 2.960 ;
        RECT 2132.170 2.760 2132.490 2.820 ;
        RECT 2137.690 2.760 2138.010 2.820 ;
      LAYER via ;
        RECT 1106.400 1587.840 1106.660 1588.100 ;
        RECT 1109.620 1587.840 1109.880 1588.100 ;
        RECT 1109.620 56.820 1109.880 57.080 ;
        RECT 2132.200 56.820 2132.460 57.080 ;
        RECT 2132.200 2.760 2132.460 3.020 ;
        RECT 2137.720 2.760 2137.980 3.020 ;
      LAYER met2 ;
        RECT 1106.400 1600.000 1106.680 1604.000 ;
        RECT 1106.460 1588.130 1106.600 1600.000 ;
        RECT 1106.400 1587.810 1106.660 1588.130 ;
        RECT 1109.620 1587.810 1109.880 1588.130 ;
        RECT 1109.680 57.110 1109.820 1587.810 ;
        RECT 1109.620 56.790 1109.880 57.110 ;
        RECT 2132.200 56.790 2132.460 57.110 ;
        RECT 2132.260 3.050 2132.400 56.790 ;
        RECT 2132.200 2.730 2132.460 3.050 ;
        RECT 2137.720 2.730 2137.980 3.050 ;
        RECT 2137.780 2.400 2137.920 2.730 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1113.270 1589.740 1113.590 1589.800 ;
        RECT 1116.950 1589.740 1117.270 1589.800 ;
        RECT 1113.270 1589.600 1117.270 1589.740 ;
        RECT 1113.270 1589.540 1113.590 1589.600 ;
        RECT 1116.950 1589.540 1117.270 1589.600 ;
        RECT 1116.950 57.360 1117.270 57.420 ;
        RECT 2152.870 57.360 2153.190 57.420 ;
        RECT 1116.950 57.220 2153.190 57.360 ;
        RECT 1116.950 57.160 1117.270 57.220 ;
        RECT 2152.870 57.160 2153.190 57.220 ;
        RECT 2152.870 2.960 2153.190 3.020 ;
        RECT 2155.630 2.960 2155.950 3.020 ;
        RECT 2152.870 2.820 2155.950 2.960 ;
        RECT 2152.870 2.760 2153.190 2.820 ;
        RECT 2155.630 2.760 2155.950 2.820 ;
      LAYER via ;
        RECT 1113.300 1589.540 1113.560 1589.800 ;
        RECT 1116.980 1589.540 1117.240 1589.800 ;
        RECT 1116.980 57.160 1117.240 57.420 ;
        RECT 2152.900 57.160 2153.160 57.420 ;
        RECT 2152.900 2.760 2153.160 3.020 ;
        RECT 2155.660 2.760 2155.920 3.020 ;
      LAYER met2 ;
        RECT 1113.300 1600.000 1113.580 1604.000 ;
        RECT 1113.360 1589.830 1113.500 1600.000 ;
        RECT 1113.300 1589.510 1113.560 1589.830 ;
        RECT 1116.980 1589.510 1117.240 1589.830 ;
        RECT 1117.040 57.450 1117.180 1589.510 ;
        RECT 1116.980 57.130 1117.240 57.450 ;
        RECT 2152.900 57.130 2153.160 57.450 ;
        RECT 2152.960 3.050 2153.100 57.130 ;
        RECT 2152.900 2.730 2153.160 3.050 ;
        RECT 2155.660 2.730 2155.920 3.050 ;
        RECT 2155.720 2.400 2155.860 2.730 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1120.170 1587.700 1120.490 1587.760 ;
        RECT 1123.390 1587.700 1123.710 1587.760 ;
        RECT 1120.170 1587.560 1123.710 1587.700 ;
        RECT 1120.170 1587.500 1120.490 1587.560 ;
        RECT 1123.390 1587.500 1123.710 1587.560 ;
        RECT 1123.390 57.700 1123.710 57.760 ;
        RECT 2166.670 57.700 2166.990 57.760 ;
        RECT 1123.390 57.560 2166.990 57.700 ;
        RECT 1123.390 57.500 1123.710 57.560 ;
        RECT 2166.670 57.500 2166.990 57.560 ;
        RECT 2166.670 17.580 2166.990 17.640 ;
        RECT 2173.110 17.580 2173.430 17.640 ;
        RECT 2166.670 17.440 2173.430 17.580 ;
        RECT 2166.670 17.380 2166.990 17.440 ;
        RECT 2173.110 17.380 2173.430 17.440 ;
      LAYER via ;
        RECT 1120.200 1587.500 1120.460 1587.760 ;
        RECT 1123.420 1587.500 1123.680 1587.760 ;
        RECT 1123.420 57.500 1123.680 57.760 ;
        RECT 2166.700 57.500 2166.960 57.760 ;
        RECT 2166.700 17.380 2166.960 17.640 ;
        RECT 2173.140 17.380 2173.400 17.640 ;
      LAYER met2 ;
        RECT 1120.200 1600.000 1120.480 1604.000 ;
        RECT 1120.260 1587.790 1120.400 1600.000 ;
        RECT 1120.200 1587.470 1120.460 1587.790 ;
        RECT 1123.420 1587.470 1123.680 1587.790 ;
        RECT 1123.480 57.790 1123.620 1587.470 ;
        RECT 1123.420 57.470 1123.680 57.790 ;
        RECT 2166.700 57.470 2166.960 57.790 ;
        RECT 2166.760 17.670 2166.900 57.470 ;
        RECT 2166.700 17.350 2166.960 17.670 ;
        RECT 2173.140 17.350 2173.400 17.670 ;
        RECT 2173.200 2.400 2173.340 17.350 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1126.610 1589.740 1126.930 1589.800 ;
        RECT 1130.750 1589.740 1131.070 1589.800 ;
        RECT 1126.610 1589.600 1131.070 1589.740 ;
        RECT 1126.610 1589.540 1126.930 1589.600 ;
        RECT 1130.750 1589.540 1131.070 1589.600 ;
        RECT 1130.750 58.040 1131.070 58.100 ;
        RECT 2187.370 58.040 2187.690 58.100 ;
        RECT 1130.750 57.900 2187.690 58.040 ;
        RECT 1130.750 57.840 1131.070 57.900 ;
        RECT 2187.370 57.840 2187.690 57.900 ;
      LAYER via ;
        RECT 1126.640 1589.540 1126.900 1589.800 ;
        RECT 1130.780 1589.540 1131.040 1589.800 ;
        RECT 1130.780 57.840 1131.040 58.100 ;
        RECT 2187.400 57.840 2187.660 58.100 ;
      LAYER met2 ;
        RECT 1126.640 1600.000 1126.920 1604.000 ;
        RECT 1126.700 1589.830 1126.840 1600.000 ;
        RECT 1126.640 1589.510 1126.900 1589.830 ;
        RECT 1130.780 1589.510 1131.040 1589.830 ;
        RECT 1130.840 58.130 1130.980 1589.510 ;
        RECT 1130.780 57.810 1131.040 58.130 ;
        RECT 2187.400 57.810 2187.660 58.130 ;
        RECT 2187.460 3.130 2187.600 57.810 ;
        RECT 2187.460 2.990 2190.820 3.130 ;
        RECT 2190.680 2.960 2190.820 2.990 ;
        RECT 2190.680 2.820 2191.280 2.960 ;
        RECT 2191.140 2.400 2191.280 2.820 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1133.510 1589.740 1133.830 1589.800 ;
        RECT 1137.650 1589.740 1137.970 1589.800 ;
        RECT 1133.510 1589.600 1137.970 1589.740 ;
        RECT 1133.510 1589.540 1133.830 1589.600 ;
        RECT 1137.650 1589.540 1137.970 1589.600 ;
        RECT 1137.650 58.380 1137.970 58.440 ;
        RECT 2208.070 58.380 2208.390 58.440 ;
        RECT 1137.650 58.240 2208.390 58.380 ;
        RECT 1137.650 58.180 1137.970 58.240 ;
        RECT 2208.070 58.180 2208.390 58.240 ;
        RECT 2208.070 2.960 2208.390 3.020 ;
        RECT 2208.990 2.960 2209.310 3.020 ;
        RECT 2208.070 2.820 2209.310 2.960 ;
        RECT 2208.070 2.760 2208.390 2.820 ;
        RECT 2208.990 2.760 2209.310 2.820 ;
      LAYER via ;
        RECT 1133.540 1589.540 1133.800 1589.800 ;
        RECT 1137.680 1589.540 1137.940 1589.800 ;
        RECT 1137.680 58.180 1137.940 58.440 ;
        RECT 2208.100 58.180 2208.360 58.440 ;
        RECT 2208.100 2.760 2208.360 3.020 ;
        RECT 2209.020 2.760 2209.280 3.020 ;
      LAYER met2 ;
        RECT 1133.540 1600.000 1133.820 1604.000 ;
        RECT 1133.600 1589.830 1133.740 1600.000 ;
        RECT 1133.540 1589.510 1133.800 1589.830 ;
        RECT 1137.680 1589.510 1137.940 1589.830 ;
        RECT 1137.740 58.470 1137.880 1589.510 ;
        RECT 1137.680 58.150 1137.940 58.470 ;
        RECT 2208.100 58.150 2208.360 58.470 ;
        RECT 2208.160 3.050 2208.300 58.150 ;
        RECT 2208.100 2.730 2208.360 3.050 ;
        RECT 2209.020 2.730 2209.280 3.050 ;
        RECT 2209.080 2.400 2209.220 2.730 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1139.950 1589.740 1140.270 1589.800 ;
        RECT 1144.550 1589.740 1144.870 1589.800 ;
        RECT 1139.950 1589.600 1144.870 1589.740 ;
        RECT 1139.950 1589.540 1140.270 1589.600 ;
        RECT 1144.550 1589.540 1144.870 1589.600 ;
        RECT 1144.550 62.120 1144.870 62.180 ;
        RECT 2221.870 62.120 2222.190 62.180 ;
        RECT 1144.550 61.980 2222.190 62.120 ;
        RECT 1144.550 61.920 1144.870 61.980 ;
        RECT 2221.870 61.920 2222.190 61.980 ;
        RECT 2221.870 2.960 2222.190 3.020 ;
        RECT 2226.930 2.960 2227.250 3.020 ;
        RECT 2221.870 2.820 2227.250 2.960 ;
        RECT 2221.870 2.760 2222.190 2.820 ;
        RECT 2226.930 2.760 2227.250 2.820 ;
      LAYER via ;
        RECT 1139.980 1589.540 1140.240 1589.800 ;
        RECT 1144.580 1589.540 1144.840 1589.800 ;
        RECT 1144.580 61.920 1144.840 62.180 ;
        RECT 2221.900 61.920 2222.160 62.180 ;
        RECT 2221.900 2.760 2222.160 3.020 ;
        RECT 2226.960 2.760 2227.220 3.020 ;
      LAYER met2 ;
        RECT 1139.980 1600.000 1140.260 1604.000 ;
        RECT 1140.040 1589.830 1140.180 1600.000 ;
        RECT 1139.980 1589.510 1140.240 1589.830 ;
        RECT 1144.580 1589.510 1144.840 1589.830 ;
        RECT 1144.640 62.210 1144.780 1589.510 ;
        RECT 1144.580 61.890 1144.840 62.210 ;
        RECT 2221.900 61.890 2222.160 62.210 ;
        RECT 2221.960 3.050 2222.100 61.890 ;
        RECT 2221.900 2.730 2222.160 3.050 ;
        RECT 2226.960 2.730 2227.220 3.050 ;
        RECT 2227.020 2.400 2227.160 2.730 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 610.105 18.785 610.275 20.995 ;
        RECT 616.545 18.275 616.715 18.955 ;
        RECT 616.545 18.105 617.635 18.275 ;
        RECT 639.545 16.745 639.715 18.275 ;
      LAYER mcon ;
        RECT 610.105 20.825 610.275 20.995 ;
        RECT 616.545 18.785 616.715 18.955 ;
        RECT 617.465 18.105 617.635 18.275 ;
        RECT 639.545 18.105 639.715 18.275 ;
      LAYER met1 ;
        RECT 594.850 1587.360 595.170 1587.420 ;
        RECT 599.450 1587.360 599.770 1587.420 ;
        RECT 594.850 1587.220 599.770 1587.360 ;
        RECT 594.850 1587.160 595.170 1587.220 ;
        RECT 599.450 1587.160 599.770 1587.220 ;
        RECT 599.450 20.980 599.770 21.040 ;
        RECT 610.045 20.980 610.335 21.025 ;
        RECT 599.450 20.840 610.335 20.980 ;
        RECT 599.450 20.780 599.770 20.840 ;
        RECT 610.045 20.795 610.335 20.840 ;
        RECT 610.045 18.940 610.335 18.985 ;
        RECT 616.485 18.940 616.775 18.985 ;
        RECT 610.045 18.800 616.775 18.940 ;
        RECT 610.045 18.755 610.335 18.800 ;
        RECT 616.485 18.755 616.775 18.800 ;
        RECT 617.405 18.260 617.695 18.305 ;
        RECT 639.485 18.260 639.775 18.305 ;
        RECT 617.405 18.120 639.775 18.260 ;
        RECT 617.405 18.075 617.695 18.120 ;
        RECT 639.485 18.075 639.775 18.120 ;
        RECT 639.485 16.900 639.775 16.945 ;
        RECT 639.485 16.760 740.900 16.900 ;
        RECT 639.485 16.715 639.775 16.760 ;
        RECT 740.760 16.560 740.900 16.760 ;
        RECT 781.610 16.560 781.930 16.620 ;
        RECT 740.760 16.420 781.930 16.560 ;
        RECT 781.610 16.360 781.930 16.420 ;
      LAYER via ;
        RECT 594.880 1587.160 595.140 1587.420 ;
        RECT 599.480 1587.160 599.740 1587.420 ;
        RECT 599.480 20.780 599.740 21.040 ;
        RECT 781.640 16.360 781.900 16.620 ;
      LAYER met2 ;
        RECT 594.880 1600.000 595.160 1604.000 ;
        RECT 594.940 1587.450 595.080 1600.000 ;
        RECT 594.880 1587.130 595.140 1587.450 ;
        RECT 599.480 1587.130 599.740 1587.450 ;
        RECT 599.540 21.070 599.680 1587.130 ;
        RECT 599.480 20.750 599.740 21.070 ;
        RECT 781.640 16.330 781.900 16.650 ;
        RECT 781.700 2.400 781.840 16.330 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1146.850 1588.040 1147.170 1588.100 ;
        RECT 1150.990 1588.040 1151.310 1588.100 ;
        RECT 1146.850 1587.900 1151.310 1588.040 ;
        RECT 1146.850 1587.840 1147.170 1587.900 ;
        RECT 1150.990 1587.840 1151.310 1587.900 ;
        RECT 1150.990 61.780 1151.310 61.840 ;
        RECT 2242.570 61.780 2242.890 61.840 ;
        RECT 1150.990 61.640 2242.890 61.780 ;
        RECT 1150.990 61.580 1151.310 61.640 ;
        RECT 2242.570 61.580 2242.890 61.640 ;
        RECT 2242.570 2.960 2242.890 3.020 ;
        RECT 2244.870 2.960 2245.190 3.020 ;
        RECT 2242.570 2.820 2245.190 2.960 ;
        RECT 2242.570 2.760 2242.890 2.820 ;
        RECT 2244.870 2.760 2245.190 2.820 ;
      LAYER via ;
        RECT 1146.880 1587.840 1147.140 1588.100 ;
        RECT 1151.020 1587.840 1151.280 1588.100 ;
        RECT 1151.020 61.580 1151.280 61.840 ;
        RECT 2242.600 61.580 2242.860 61.840 ;
        RECT 2242.600 2.760 2242.860 3.020 ;
        RECT 2244.900 2.760 2245.160 3.020 ;
      LAYER met2 ;
        RECT 1146.880 1600.000 1147.160 1604.000 ;
        RECT 1146.940 1588.130 1147.080 1600.000 ;
        RECT 1146.880 1587.810 1147.140 1588.130 ;
        RECT 1151.020 1587.810 1151.280 1588.130 ;
        RECT 1151.080 61.870 1151.220 1587.810 ;
        RECT 1151.020 61.550 1151.280 61.870 ;
        RECT 2242.600 61.550 2242.860 61.870 ;
        RECT 2242.660 3.050 2242.800 61.550 ;
        RECT 2242.600 2.730 2242.860 3.050 ;
        RECT 2244.900 2.730 2245.160 3.050 ;
        RECT 2244.960 2.400 2245.100 2.730 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1153.750 1588.040 1154.070 1588.100 ;
        RECT 1158.350 1588.040 1158.670 1588.100 ;
        RECT 1153.750 1587.900 1158.670 1588.040 ;
        RECT 1153.750 1587.840 1154.070 1587.900 ;
        RECT 1158.350 1587.840 1158.670 1587.900 ;
        RECT 1158.350 61.440 1158.670 61.500 ;
        RECT 2256.370 61.440 2256.690 61.500 ;
        RECT 1158.350 61.300 2256.690 61.440 ;
        RECT 1158.350 61.240 1158.670 61.300 ;
        RECT 2256.370 61.240 2256.690 61.300 ;
        RECT 2256.370 17.580 2256.690 17.640 ;
        RECT 2262.350 17.580 2262.670 17.640 ;
        RECT 2256.370 17.440 2262.670 17.580 ;
        RECT 2256.370 17.380 2256.690 17.440 ;
        RECT 2262.350 17.380 2262.670 17.440 ;
      LAYER via ;
        RECT 1153.780 1587.840 1154.040 1588.100 ;
        RECT 1158.380 1587.840 1158.640 1588.100 ;
        RECT 1158.380 61.240 1158.640 61.500 ;
        RECT 2256.400 61.240 2256.660 61.500 ;
        RECT 2256.400 17.380 2256.660 17.640 ;
        RECT 2262.380 17.380 2262.640 17.640 ;
      LAYER met2 ;
        RECT 1153.780 1600.000 1154.060 1604.000 ;
        RECT 1153.840 1588.130 1153.980 1600.000 ;
        RECT 1153.780 1587.810 1154.040 1588.130 ;
        RECT 1158.380 1587.810 1158.640 1588.130 ;
        RECT 1158.440 61.530 1158.580 1587.810 ;
        RECT 1158.380 61.210 1158.640 61.530 ;
        RECT 2256.400 61.210 2256.660 61.530 ;
        RECT 2256.460 17.670 2256.600 61.210 ;
        RECT 2256.400 17.350 2256.660 17.670 ;
        RECT 2262.380 17.350 2262.640 17.670 ;
        RECT 2262.440 2.400 2262.580 17.350 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1160.190 1588.040 1160.510 1588.100 ;
        RECT 1164.790 1588.040 1165.110 1588.100 ;
        RECT 1160.190 1587.900 1165.110 1588.040 ;
        RECT 1160.190 1587.840 1160.510 1587.900 ;
        RECT 1164.790 1587.840 1165.110 1587.900 ;
        RECT 1164.790 61.100 1165.110 61.160 ;
        RECT 2277.070 61.100 2277.390 61.160 ;
        RECT 1164.790 60.960 2277.390 61.100 ;
        RECT 1164.790 60.900 1165.110 60.960 ;
        RECT 2277.070 60.900 2277.390 60.960 ;
        RECT 2277.070 2.960 2277.390 3.020 ;
        RECT 2280.290 2.960 2280.610 3.020 ;
        RECT 2277.070 2.820 2280.610 2.960 ;
        RECT 2277.070 2.760 2277.390 2.820 ;
        RECT 2280.290 2.760 2280.610 2.820 ;
      LAYER via ;
        RECT 1160.220 1587.840 1160.480 1588.100 ;
        RECT 1164.820 1587.840 1165.080 1588.100 ;
        RECT 1164.820 60.900 1165.080 61.160 ;
        RECT 2277.100 60.900 2277.360 61.160 ;
        RECT 2277.100 2.760 2277.360 3.020 ;
        RECT 2280.320 2.760 2280.580 3.020 ;
      LAYER met2 ;
        RECT 1160.220 1600.000 1160.500 1604.000 ;
        RECT 1160.280 1588.130 1160.420 1600.000 ;
        RECT 1160.220 1587.810 1160.480 1588.130 ;
        RECT 1164.820 1587.810 1165.080 1588.130 ;
        RECT 1164.880 61.190 1165.020 1587.810 ;
        RECT 1164.820 60.870 1165.080 61.190 ;
        RECT 2277.100 60.870 2277.360 61.190 ;
        RECT 2277.160 3.050 2277.300 60.870 ;
        RECT 2277.100 2.730 2277.360 3.050 ;
        RECT 2280.320 2.730 2280.580 3.050 ;
        RECT 2280.380 2.400 2280.520 2.730 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1167.090 1588.040 1167.410 1588.100 ;
        RECT 1172.150 1588.040 1172.470 1588.100 ;
        RECT 1167.090 1587.900 1172.470 1588.040 ;
        RECT 1167.090 1587.840 1167.410 1587.900 ;
        RECT 1172.150 1587.840 1172.470 1587.900 ;
        RECT 1172.150 60.760 1172.470 60.820 ;
        RECT 2298.230 60.760 2298.550 60.820 ;
        RECT 1172.150 60.620 2298.550 60.760 ;
        RECT 1172.150 60.560 1172.470 60.620 ;
        RECT 2298.230 60.560 2298.550 60.620 ;
      LAYER via ;
        RECT 1167.120 1587.840 1167.380 1588.100 ;
        RECT 1172.180 1587.840 1172.440 1588.100 ;
        RECT 1172.180 60.560 1172.440 60.820 ;
        RECT 2298.260 60.560 2298.520 60.820 ;
      LAYER met2 ;
        RECT 1167.120 1600.000 1167.400 1604.000 ;
        RECT 1167.180 1588.130 1167.320 1600.000 ;
        RECT 1167.120 1587.810 1167.380 1588.130 ;
        RECT 1172.180 1587.810 1172.440 1588.130 ;
        RECT 1172.240 60.850 1172.380 1587.810 ;
        RECT 1172.180 60.530 1172.440 60.850 ;
        RECT 2298.260 60.530 2298.520 60.850 ;
        RECT 2298.320 2.400 2298.460 60.530 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1173.990 1588.040 1174.310 1588.100 ;
        RECT 1178.590 1588.040 1178.910 1588.100 ;
        RECT 1173.990 1587.900 1178.910 1588.040 ;
        RECT 1173.990 1587.840 1174.310 1587.900 ;
        RECT 1178.590 1587.840 1178.910 1587.900 ;
        RECT 1178.590 60.420 1178.910 60.480 ;
        RECT 2311.570 60.420 2311.890 60.480 ;
        RECT 1178.590 60.280 2311.890 60.420 ;
        RECT 1178.590 60.220 1178.910 60.280 ;
        RECT 2311.570 60.220 2311.890 60.280 ;
        RECT 2311.570 2.960 2311.890 3.020 ;
        RECT 2316.170 2.960 2316.490 3.020 ;
        RECT 2311.570 2.820 2316.490 2.960 ;
        RECT 2311.570 2.760 2311.890 2.820 ;
        RECT 2316.170 2.760 2316.490 2.820 ;
      LAYER via ;
        RECT 1174.020 1587.840 1174.280 1588.100 ;
        RECT 1178.620 1587.840 1178.880 1588.100 ;
        RECT 1178.620 60.220 1178.880 60.480 ;
        RECT 2311.600 60.220 2311.860 60.480 ;
        RECT 2311.600 2.760 2311.860 3.020 ;
        RECT 2316.200 2.760 2316.460 3.020 ;
      LAYER met2 ;
        RECT 1174.020 1600.000 1174.300 1604.000 ;
        RECT 1174.080 1588.130 1174.220 1600.000 ;
        RECT 1174.020 1587.810 1174.280 1588.130 ;
        RECT 1178.620 1587.810 1178.880 1588.130 ;
        RECT 1178.680 60.510 1178.820 1587.810 ;
        RECT 1178.620 60.190 1178.880 60.510 ;
        RECT 2311.600 60.190 2311.860 60.510 ;
        RECT 2311.660 3.050 2311.800 60.190 ;
        RECT 2311.600 2.730 2311.860 3.050 ;
        RECT 2316.200 2.730 2316.460 3.050 ;
        RECT 2316.260 2.400 2316.400 2.730 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1180.430 1588.040 1180.750 1588.100 ;
        RECT 1185.950 1588.040 1186.270 1588.100 ;
        RECT 1180.430 1587.900 1186.270 1588.040 ;
        RECT 1180.430 1587.840 1180.750 1587.900 ;
        RECT 1185.950 1587.840 1186.270 1587.900 ;
        RECT 1185.950 60.080 1186.270 60.140 ;
        RECT 2332.270 60.080 2332.590 60.140 ;
        RECT 1185.950 59.940 2332.590 60.080 ;
        RECT 1185.950 59.880 1186.270 59.940 ;
        RECT 2332.270 59.880 2332.590 59.940 ;
        RECT 2332.270 2.960 2332.590 3.020 ;
        RECT 2334.110 2.960 2334.430 3.020 ;
        RECT 2332.270 2.820 2334.430 2.960 ;
        RECT 2332.270 2.760 2332.590 2.820 ;
        RECT 2334.110 2.760 2334.430 2.820 ;
      LAYER via ;
        RECT 1180.460 1587.840 1180.720 1588.100 ;
        RECT 1185.980 1587.840 1186.240 1588.100 ;
        RECT 1185.980 59.880 1186.240 60.140 ;
        RECT 2332.300 59.880 2332.560 60.140 ;
        RECT 2332.300 2.760 2332.560 3.020 ;
        RECT 2334.140 2.760 2334.400 3.020 ;
      LAYER met2 ;
        RECT 1180.460 1600.000 1180.740 1604.000 ;
        RECT 1180.520 1588.130 1180.660 1600.000 ;
        RECT 1180.460 1587.810 1180.720 1588.130 ;
        RECT 1185.980 1587.810 1186.240 1588.130 ;
        RECT 1186.040 60.170 1186.180 1587.810 ;
        RECT 1185.980 59.850 1186.240 60.170 ;
        RECT 2332.300 59.850 2332.560 60.170 ;
        RECT 2332.360 3.050 2332.500 59.850 ;
        RECT 2332.300 2.730 2332.560 3.050 ;
        RECT 2334.140 2.730 2334.400 3.050 ;
        RECT 2334.200 2.400 2334.340 2.730 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1187.330 1588.040 1187.650 1588.100 ;
        RECT 1192.390 1588.040 1192.710 1588.100 ;
        RECT 1187.330 1587.900 1192.710 1588.040 ;
        RECT 1187.330 1587.840 1187.650 1587.900 ;
        RECT 1192.390 1587.840 1192.710 1587.900 ;
        RECT 1192.390 59.740 1192.710 59.800 ;
        RECT 2346.070 59.740 2346.390 59.800 ;
        RECT 1192.390 59.600 2346.390 59.740 ;
        RECT 1192.390 59.540 1192.710 59.600 ;
        RECT 2346.070 59.540 2346.390 59.600 ;
        RECT 2346.070 2.960 2346.390 3.020 ;
        RECT 2351.590 2.960 2351.910 3.020 ;
        RECT 2346.070 2.820 2351.910 2.960 ;
        RECT 2346.070 2.760 2346.390 2.820 ;
        RECT 2351.590 2.760 2351.910 2.820 ;
      LAYER via ;
        RECT 1187.360 1587.840 1187.620 1588.100 ;
        RECT 1192.420 1587.840 1192.680 1588.100 ;
        RECT 1192.420 59.540 1192.680 59.800 ;
        RECT 2346.100 59.540 2346.360 59.800 ;
        RECT 2346.100 2.760 2346.360 3.020 ;
        RECT 2351.620 2.760 2351.880 3.020 ;
      LAYER met2 ;
        RECT 1187.360 1600.000 1187.640 1604.000 ;
        RECT 1187.420 1588.130 1187.560 1600.000 ;
        RECT 1187.360 1587.810 1187.620 1588.130 ;
        RECT 1192.420 1587.810 1192.680 1588.130 ;
        RECT 1192.480 59.830 1192.620 1587.810 ;
        RECT 1192.420 59.510 1192.680 59.830 ;
        RECT 2346.100 59.510 2346.360 59.830 ;
        RECT 2346.160 3.050 2346.300 59.510 ;
        RECT 2346.100 2.730 2346.360 3.050 ;
        RECT 2351.620 2.730 2351.880 3.050 ;
        RECT 2351.680 2.400 2351.820 2.730 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1194.230 1588.040 1194.550 1588.100 ;
        RECT 1199.750 1588.040 1200.070 1588.100 ;
        RECT 1194.230 1587.900 1200.070 1588.040 ;
        RECT 1194.230 1587.840 1194.550 1587.900 ;
        RECT 1199.750 1587.840 1200.070 1587.900 ;
        RECT 1199.750 59.400 1200.070 59.460 ;
        RECT 2366.770 59.400 2367.090 59.460 ;
        RECT 1199.750 59.260 2367.090 59.400 ;
        RECT 1199.750 59.200 1200.070 59.260 ;
        RECT 2366.770 59.200 2367.090 59.260 ;
      LAYER via ;
        RECT 1194.260 1587.840 1194.520 1588.100 ;
        RECT 1199.780 1587.840 1200.040 1588.100 ;
        RECT 1199.780 59.200 1200.040 59.460 ;
        RECT 2366.800 59.200 2367.060 59.460 ;
      LAYER met2 ;
        RECT 1194.260 1600.000 1194.540 1604.000 ;
        RECT 1194.320 1588.130 1194.460 1600.000 ;
        RECT 1194.260 1587.810 1194.520 1588.130 ;
        RECT 1199.780 1587.810 1200.040 1588.130 ;
        RECT 1199.840 59.490 1199.980 1587.810 ;
        RECT 1199.780 59.170 1200.040 59.490 ;
        RECT 2366.800 59.170 2367.060 59.490 ;
        RECT 2366.860 3.130 2367.000 59.170 ;
        RECT 2366.860 2.990 2369.300 3.130 ;
        RECT 2369.160 2.960 2369.300 2.990 ;
        RECT 2369.160 2.820 2369.760 2.960 ;
        RECT 2369.620 2.400 2369.760 2.820 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1200.670 1588.040 1200.990 1588.100 ;
        RECT 1206.190 1588.040 1206.510 1588.100 ;
        RECT 1200.670 1587.900 1206.510 1588.040 ;
        RECT 1200.670 1587.840 1200.990 1587.900 ;
        RECT 1206.190 1587.840 1206.510 1587.900 ;
        RECT 1206.190 59.060 1206.510 59.120 ;
        RECT 2387.470 59.060 2387.790 59.120 ;
        RECT 1206.190 58.920 2387.790 59.060 ;
        RECT 1206.190 58.860 1206.510 58.920 ;
        RECT 2387.470 58.860 2387.790 58.920 ;
      LAYER via ;
        RECT 1200.700 1587.840 1200.960 1588.100 ;
        RECT 1206.220 1587.840 1206.480 1588.100 ;
        RECT 1206.220 58.860 1206.480 59.120 ;
        RECT 2387.500 58.860 2387.760 59.120 ;
      LAYER met2 ;
        RECT 1200.700 1600.000 1200.980 1604.000 ;
        RECT 1200.760 1588.130 1200.900 1600.000 ;
        RECT 1200.700 1587.810 1200.960 1588.130 ;
        RECT 1206.220 1587.810 1206.480 1588.130 ;
        RECT 1206.280 59.150 1206.420 1587.810 ;
        RECT 1206.220 58.830 1206.480 59.150 ;
        RECT 2387.500 58.830 2387.760 59.150 ;
        RECT 2387.560 2.400 2387.700 58.830 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1207.570 1587.700 1207.890 1587.760 ;
        RECT 1213.550 1587.700 1213.870 1587.760 ;
        RECT 1207.570 1587.560 1213.870 1587.700 ;
        RECT 1207.570 1587.500 1207.890 1587.560 ;
        RECT 1213.550 1587.500 1213.870 1587.560 ;
        RECT 1213.550 58.720 1213.870 58.780 ;
        RECT 2401.270 58.720 2401.590 58.780 ;
        RECT 1213.550 58.580 2401.590 58.720 ;
        RECT 1213.550 58.520 1213.870 58.580 ;
        RECT 2401.270 58.520 2401.590 58.580 ;
      LAYER via ;
        RECT 1207.600 1587.500 1207.860 1587.760 ;
        RECT 1213.580 1587.500 1213.840 1587.760 ;
        RECT 1213.580 58.520 1213.840 58.780 ;
        RECT 2401.300 58.520 2401.560 58.780 ;
      LAYER met2 ;
        RECT 1207.600 1600.000 1207.880 1604.000 ;
        RECT 1207.660 1587.790 1207.800 1600.000 ;
        RECT 1207.600 1587.470 1207.860 1587.790 ;
        RECT 1213.580 1587.470 1213.840 1587.790 ;
        RECT 1213.640 58.810 1213.780 1587.470 ;
        RECT 1213.580 58.490 1213.840 58.810 ;
        RECT 2401.300 58.490 2401.560 58.810 ;
        RECT 2401.360 17.410 2401.500 58.490 ;
        RECT 2401.360 17.270 2405.640 17.410 ;
        RECT 2405.500 2.400 2405.640 17.270 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 601.290 1587.360 601.610 1587.420 ;
        RECT 606.350 1587.360 606.670 1587.420 ;
        RECT 601.290 1587.220 606.670 1587.360 ;
        RECT 601.290 1587.160 601.610 1587.220 ;
        RECT 606.350 1587.160 606.670 1587.220 ;
        RECT 606.350 19.960 606.670 20.020 ;
        RECT 799.550 19.960 799.870 20.020 ;
        RECT 606.350 19.820 799.870 19.960 ;
        RECT 606.350 19.760 606.670 19.820 ;
        RECT 799.550 19.760 799.870 19.820 ;
      LAYER via ;
        RECT 601.320 1587.160 601.580 1587.420 ;
        RECT 606.380 1587.160 606.640 1587.420 ;
        RECT 606.380 19.760 606.640 20.020 ;
        RECT 799.580 19.760 799.840 20.020 ;
      LAYER met2 ;
        RECT 601.320 1600.000 601.600 1604.000 ;
        RECT 601.380 1587.450 601.520 1600.000 ;
        RECT 601.320 1587.130 601.580 1587.450 ;
        RECT 606.380 1587.130 606.640 1587.450 ;
        RECT 606.440 20.050 606.580 1587.130 ;
        RECT 606.380 19.730 606.640 20.050 ;
        RECT 799.580 19.730 799.840 20.050 ;
        RECT 799.640 2.400 799.780 19.730 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 542.870 1592.120 543.190 1592.180 ;
        RECT 643.150 1592.120 643.470 1592.180 ;
        RECT 542.870 1591.980 643.470 1592.120 ;
        RECT 542.870 1591.920 543.190 1591.980 ;
        RECT 643.150 1591.920 643.470 1591.980 ;
        RECT 643.150 2.960 643.470 3.020 ;
        RECT 644.990 2.960 645.310 3.020 ;
        RECT 643.150 2.820 645.310 2.960 ;
        RECT 643.150 2.760 643.470 2.820 ;
        RECT 644.990 2.760 645.310 2.820 ;
      LAYER via ;
        RECT 542.900 1591.920 543.160 1592.180 ;
        RECT 643.180 1591.920 643.440 1592.180 ;
        RECT 643.180 2.760 643.440 3.020 ;
        RECT 645.020 2.760 645.280 3.020 ;
      LAYER met2 ;
        RECT 542.900 1600.000 543.180 1604.000 ;
        RECT 542.960 1592.210 543.100 1600.000 ;
        RECT 542.900 1591.890 543.160 1592.210 ;
        RECT 643.180 1591.890 643.440 1592.210 ;
        RECT 643.240 3.050 643.380 1591.890 ;
        RECT 643.180 2.730 643.440 3.050 ;
        RECT 645.020 2.730 645.280 3.050 ;
        RECT 645.080 2.400 645.220 2.730 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1216.310 1588.040 1216.630 1588.100 ;
        RECT 1220.910 1588.040 1221.230 1588.100 ;
        RECT 1216.310 1587.900 1221.230 1588.040 ;
        RECT 1216.310 1587.840 1216.630 1587.900 ;
        RECT 1220.910 1587.840 1221.230 1587.900 ;
      LAYER via ;
        RECT 1216.340 1587.840 1216.600 1588.100 ;
        RECT 1220.940 1587.840 1221.200 1588.100 ;
      LAYER met2 ;
        RECT 1216.340 1600.000 1216.620 1604.000 ;
        RECT 1216.400 1588.130 1216.540 1600.000 ;
        RECT 1216.340 1587.810 1216.600 1588.130 ;
        RECT 1220.940 1587.810 1221.200 1588.130 ;
        RECT 1221.000 61.045 1221.140 1587.810 ;
        RECT 1220.930 60.675 1221.210 61.045 ;
        RECT 2429.350 60.675 2429.630 61.045 ;
        RECT 2429.420 17.410 2429.560 60.675 ;
        RECT 2428.960 17.270 2429.560 17.410 ;
        RECT 2428.960 2.400 2429.100 17.270 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
      LAYER via2 ;
        RECT 1220.930 60.720 1221.210 61.000 ;
        RECT 2429.350 60.720 2429.630 61.000 ;
      LAYER met3 ;
        RECT 1220.905 61.010 1221.235 61.025 ;
        RECT 2429.325 61.010 2429.655 61.025 ;
        RECT 1220.905 60.710 2429.655 61.010 ;
        RECT 1220.905 60.695 1221.235 60.710 ;
        RECT 2429.325 60.695 2429.655 60.710 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1223.210 1587.700 1223.530 1587.760 ;
        RECT 1227.810 1587.700 1228.130 1587.760 ;
        RECT 1223.210 1587.560 1228.130 1587.700 ;
        RECT 1223.210 1587.500 1223.530 1587.560 ;
        RECT 1227.810 1587.500 1228.130 1587.560 ;
      LAYER via ;
        RECT 1223.240 1587.500 1223.500 1587.760 ;
        RECT 1227.840 1587.500 1228.100 1587.760 ;
      LAYER met2 ;
        RECT 1223.240 1600.000 1223.520 1604.000 ;
        RECT 1223.300 1587.790 1223.440 1600.000 ;
        RECT 1223.240 1587.470 1223.500 1587.790 ;
        RECT 1227.840 1587.470 1228.100 1587.790 ;
        RECT 1227.900 60.365 1228.040 1587.470 ;
        RECT 1227.830 59.995 1228.110 60.365 ;
        RECT 2442.690 59.995 2442.970 60.365 ;
        RECT 2442.760 17.410 2442.900 59.995 ;
        RECT 2442.760 17.270 2447.040 17.410 ;
        RECT 2446.900 2.400 2447.040 17.270 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
      LAYER via2 ;
        RECT 1227.830 60.040 1228.110 60.320 ;
        RECT 2442.690 60.040 2442.970 60.320 ;
      LAYER met3 ;
        RECT 1227.805 60.330 1228.135 60.345 ;
        RECT 2442.665 60.330 2442.995 60.345 ;
        RECT 1227.805 60.030 2442.995 60.330 ;
        RECT 1227.805 60.015 1228.135 60.030 ;
        RECT 2442.665 60.015 2442.995 60.030 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1230.110 1588.040 1230.430 1588.100 ;
        RECT 1234.710 1588.040 1235.030 1588.100 ;
        RECT 1230.110 1587.900 1235.030 1588.040 ;
        RECT 1230.110 1587.840 1230.430 1587.900 ;
        RECT 1234.710 1587.840 1235.030 1587.900 ;
      LAYER via ;
        RECT 1230.140 1587.840 1230.400 1588.100 ;
        RECT 1234.740 1587.840 1235.000 1588.100 ;
      LAYER met2 ;
        RECT 1230.140 1600.000 1230.420 1604.000 ;
        RECT 1230.200 1588.130 1230.340 1600.000 ;
        RECT 1230.140 1587.810 1230.400 1588.130 ;
        RECT 1234.740 1587.810 1235.000 1588.130 ;
        RECT 1234.800 59.685 1234.940 1587.810 ;
        RECT 1234.730 59.315 1235.010 59.685 ;
        RECT 2463.390 59.315 2463.670 59.685 ;
        RECT 2463.460 3.130 2463.600 59.315 ;
        RECT 2463.460 2.990 2464.520 3.130 ;
        RECT 2464.380 2.960 2464.520 2.990 ;
        RECT 2464.380 2.820 2464.980 2.960 ;
        RECT 2464.840 2.400 2464.980 2.820 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
      LAYER via2 ;
        RECT 1234.730 59.360 1235.010 59.640 ;
        RECT 2463.390 59.360 2463.670 59.640 ;
      LAYER met3 ;
        RECT 1234.705 59.650 1235.035 59.665 ;
        RECT 2463.365 59.650 2463.695 59.665 ;
        RECT 1234.705 59.350 2463.695 59.650 ;
        RECT 1234.705 59.335 1235.035 59.350 ;
        RECT 2463.365 59.335 2463.695 59.350 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1236.550 1588.040 1236.870 1588.100 ;
        RECT 1241.150 1588.040 1241.470 1588.100 ;
        RECT 1236.550 1587.900 1241.470 1588.040 ;
        RECT 1236.550 1587.840 1236.870 1587.900 ;
        RECT 1241.150 1587.840 1241.470 1587.900 ;
        RECT 2477.170 2.960 2477.490 3.020 ;
        RECT 2482.690 2.960 2483.010 3.020 ;
        RECT 2477.170 2.820 2483.010 2.960 ;
        RECT 2477.170 2.760 2477.490 2.820 ;
        RECT 2482.690 2.760 2483.010 2.820 ;
      LAYER via ;
        RECT 1236.580 1587.840 1236.840 1588.100 ;
        RECT 1241.180 1587.840 1241.440 1588.100 ;
        RECT 2477.200 2.760 2477.460 3.020 ;
        RECT 2482.720 2.760 2482.980 3.020 ;
      LAYER met2 ;
        RECT 1236.580 1600.000 1236.860 1604.000 ;
        RECT 1236.640 1588.130 1236.780 1600.000 ;
        RECT 1236.580 1587.810 1236.840 1588.130 ;
        RECT 1241.180 1587.810 1241.440 1588.130 ;
        RECT 1241.240 59.005 1241.380 1587.810 ;
        RECT 1241.170 58.635 1241.450 59.005 ;
        RECT 2477.190 58.635 2477.470 59.005 ;
        RECT 2477.260 3.050 2477.400 58.635 ;
        RECT 2477.200 2.730 2477.460 3.050 ;
        RECT 2482.720 2.730 2482.980 3.050 ;
        RECT 2482.780 2.400 2482.920 2.730 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
      LAYER via2 ;
        RECT 1241.170 58.680 1241.450 58.960 ;
        RECT 2477.190 58.680 2477.470 58.960 ;
      LAYER met3 ;
        RECT 1241.145 58.970 1241.475 58.985 ;
        RECT 2477.165 58.970 2477.495 58.985 ;
        RECT 1241.145 58.670 2477.495 58.970 ;
        RECT 1241.145 58.655 1241.475 58.670 ;
        RECT 2477.165 58.655 2477.495 58.670 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1243.450 1590.760 1243.770 1590.820 ;
        RECT 1248.050 1590.760 1248.370 1590.820 ;
        RECT 1243.450 1590.620 1248.370 1590.760 ;
        RECT 1243.450 1590.560 1243.770 1590.620 ;
        RECT 1248.050 1590.560 1248.370 1590.620 ;
        RECT 2497.870 2.960 2498.190 3.020 ;
        RECT 2500.630 2.960 2500.950 3.020 ;
        RECT 2497.870 2.820 2500.950 2.960 ;
        RECT 2497.870 2.760 2498.190 2.820 ;
        RECT 2500.630 2.760 2500.950 2.820 ;
      LAYER via ;
        RECT 1243.480 1590.560 1243.740 1590.820 ;
        RECT 1248.080 1590.560 1248.340 1590.820 ;
        RECT 2497.900 2.760 2498.160 3.020 ;
        RECT 2500.660 2.760 2500.920 3.020 ;
      LAYER met2 ;
        RECT 1243.480 1600.000 1243.760 1604.000 ;
        RECT 1243.540 1590.850 1243.680 1600.000 ;
        RECT 1243.480 1590.530 1243.740 1590.850 ;
        RECT 1248.080 1590.530 1248.340 1590.850 ;
        RECT 1248.140 58.325 1248.280 1590.530 ;
        RECT 1248.070 57.955 1248.350 58.325 ;
        RECT 2497.890 57.955 2498.170 58.325 ;
        RECT 2497.960 3.050 2498.100 57.955 ;
        RECT 2497.900 2.730 2498.160 3.050 ;
        RECT 2500.660 2.730 2500.920 3.050 ;
        RECT 2500.720 2.400 2500.860 2.730 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
      LAYER via2 ;
        RECT 1248.070 58.000 1248.350 58.280 ;
        RECT 2497.890 58.000 2498.170 58.280 ;
      LAYER met3 ;
        RECT 1248.045 58.290 1248.375 58.305 ;
        RECT 2497.865 58.290 2498.195 58.305 ;
        RECT 1248.045 57.990 2498.195 58.290 ;
        RECT 1248.045 57.975 1248.375 57.990 ;
        RECT 2497.865 57.975 2498.195 57.990 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1250.350 1590.760 1250.670 1590.820 ;
        RECT 1254.950 1590.760 1255.270 1590.820 ;
        RECT 1250.350 1590.620 1255.270 1590.760 ;
        RECT 1250.350 1590.560 1250.670 1590.620 ;
        RECT 1254.950 1590.560 1255.270 1590.620 ;
        RECT 2511.670 17.580 2511.990 17.640 ;
        RECT 2518.110 17.580 2518.430 17.640 ;
        RECT 2511.670 17.440 2518.430 17.580 ;
        RECT 2511.670 17.380 2511.990 17.440 ;
        RECT 2518.110 17.380 2518.430 17.440 ;
      LAYER via ;
        RECT 1250.380 1590.560 1250.640 1590.820 ;
        RECT 1254.980 1590.560 1255.240 1590.820 ;
        RECT 2511.700 17.380 2511.960 17.640 ;
        RECT 2518.140 17.380 2518.400 17.640 ;
      LAYER met2 ;
        RECT 1250.380 1600.000 1250.660 1604.000 ;
        RECT 1250.440 1590.850 1250.580 1600.000 ;
        RECT 1250.380 1590.530 1250.640 1590.850 ;
        RECT 1254.980 1590.530 1255.240 1590.850 ;
        RECT 1255.040 75.325 1255.180 1590.530 ;
        RECT 1254.970 74.955 1255.250 75.325 ;
        RECT 2511.690 74.955 2511.970 75.325 ;
        RECT 2511.760 17.670 2511.900 74.955 ;
        RECT 2511.700 17.350 2511.960 17.670 ;
        RECT 2518.140 17.350 2518.400 17.670 ;
        RECT 2518.200 2.400 2518.340 17.350 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
      LAYER via2 ;
        RECT 1254.970 75.000 1255.250 75.280 ;
        RECT 2511.690 75.000 2511.970 75.280 ;
      LAYER met3 ;
        RECT 1254.945 75.290 1255.275 75.305 ;
        RECT 2511.665 75.290 2511.995 75.305 ;
        RECT 1254.945 74.990 2511.995 75.290 ;
        RECT 1254.945 74.975 1255.275 74.990 ;
        RECT 2511.665 74.975 2511.995 74.990 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1256.790 1590.760 1257.110 1590.820 ;
        RECT 1261.850 1590.760 1262.170 1590.820 ;
        RECT 1256.790 1590.620 1262.170 1590.760 ;
        RECT 1256.790 1590.560 1257.110 1590.620 ;
        RECT 1261.850 1590.560 1262.170 1590.620 ;
        RECT 2532.370 2.960 2532.690 3.020 ;
        RECT 2536.050 2.960 2536.370 3.020 ;
        RECT 2532.370 2.820 2536.370 2.960 ;
        RECT 2532.370 2.760 2532.690 2.820 ;
        RECT 2536.050 2.760 2536.370 2.820 ;
      LAYER via ;
        RECT 1256.820 1590.560 1257.080 1590.820 ;
        RECT 1261.880 1590.560 1262.140 1590.820 ;
        RECT 2532.400 2.760 2532.660 3.020 ;
        RECT 2536.080 2.760 2536.340 3.020 ;
      LAYER met2 ;
        RECT 1256.820 1600.000 1257.100 1604.000 ;
        RECT 1256.880 1590.850 1257.020 1600.000 ;
        RECT 1256.820 1590.530 1257.080 1590.850 ;
        RECT 1261.880 1590.530 1262.140 1590.850 ;
        RECT 1261.940 74.645 1262.080 1590.530 ;
        RECT 1261.870 74.275 1262.150 74.645 ;
        RECT 2532.390 74.275 2532.670 74.645 ;
        RECT 2532.460 3.050 2532.600 74.275 ;
        RECT 2532.400 2.730 2532.660 3.050 ;
        RECT 2536.080 2.730 2536.340 3.050 ;
        RECT 2536.140 2.400 2536.280 2.730 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
      LAYER via2 ;
        RECT 1261.870 74.320 1262.150 74.600 ;
        RECT 2532.390 74.320 2532.670 74.600 ;
      LAYER met3 ;
        RECT 1261.845 74.610 1262.175 74.625 ;
        RECT 2532.365 74.610 2532.695 74.625 ;
        RECT 1261.845 74.310 2532.695 74.610 ;
        RECT 1261.845 74.295 1262.175 74.310 ;
        RECT 2532.365 74.295 2532.695 74.310 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1263.690 1590.760 1264.010 1590.820 ;
        RECT 1268.290 1590.760 1268.610 1590.820 ;
        RECT 1263.690 1590.620 1268.610 1590.760 ;
        RECT 1263.690 1590.560 1264.010 1590.620 ;
        RECT 1268.290 1590.560 1268.610 1590.620 ;
        RECT 2553.070 2.960 2553.390 3.020 ;
        RECT 2553.990 2.960 2554.310 3.020 ;
        RECT 2553.070 2.820 2554.310 2.960 ;
        RECT 2553.070 2.760 2553.390 2.820 ;
        RECT 2553.990 2.760 2554.310 2.820 ;
      LAYER via ;
        RECT 1263.720 1590.560 1263.980 1590.820 ;
        RECT 1268.320 1590.560 1268.580 1590.820 ;
        RECT 2553.100 2.760 2553.360 3.020 ;
        RECT 2554.020 2.760 2554.280 3.020 ;
      LAYER met2 ;
        RECT 1263.720 1600.000 1264.000 1604.000 ;
        RECT 1263.780 1590.850 1263.920 1600.000 ;
        RECT 1263.720 1590.530 1263.980 1590.850 ;
        RECT 1268.320 1590.530 1268.580 1590.850 ;
        RECT 1268.380 73.965 1268.520 1590.530 ;
        RECT 1268.310 73.595 1268.590 73.965 ;
        RECT 2553.090 73.595 2553.370 73.965 ;
        RECT 2553.160 3.050 2553.300 73.595 ;
        RECT 2553.100 2.730 2553.360 3.050 ;
        RECT 2554.020 2.730 2554.280 3.050 ;
        RECT 2554.080 2.400 2554.220 2.730 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
      LAYER via2 ;
        RECT 1268.310 73.640 1268.590 73.920 ;
        RECT 2553.090 73.640 2553.370 73.920 ;
      LAYER met3 ;
        RECT 1268.285 73.930 1268.615 73.945 ;
        RECT 2553.065 73.930 2553.395 73.945 ;
        RECT 1268.285 73.630 2553.395 73.930 ;
        RECT 1268.285 73.615 1268.615 73.630 ;
        RECT 2553.065 73.615 2553.395 73.630 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1270.130 1590.760 1270.450 1590.820 ;
        RECT 1275.190 1590.760 1275.510 1590.820 ;
        RECT 1270.130 1590.620 1275.510 1590.760 ;
        RECT 1270.130 1590.560 1270.450 1590.620 ;
        RECT 1275.190 1590.560 1275.510 1590.620 ;
        RECT 2566.870 2.960 2567.190 3.020 ;
        RECT 2571.930 2.960 2572.250 3.020 ;
        RECT 2566.870 2.820 2572.250 2.960 ;
        RECT 2566.870 2.760 2567.190 2.820 ;
        RECT 2571.930 2.760 2572.250 2.820 ;
      LAYER via ;
        RECT 1270.160 1590.560 1270.420 1590.820 ;
        RECT 1275.220 1590.560 1275.480 1590.820 ;
        RECT 2566.900 2.760 2567.160 3.020 ;
        RECT 2571.960 2.760 2572.220 3.020 ;
      LAYER met2 ;
        RECT 1270.160 1600.000 1270.440 1604.000 ;
        RECT 1270.220 1590.850 1270.360 1600.000 ;
        RECT 1270.160 1590.530 1270.420 1590.850 ;
        RECT 1275.220 1590.530 1275.480 1590.850 ;
        RECT 1275.280 73.285 1275.420 1590.530 ;
        RECT 1275.210 72.915 1275.490 73.285 ;
        RECT 2566.890 72.915 2567.170 73.285 ;
        RECT 2566.960 3.050 2567.100 72.915 ;
        RECT 2566.900 2.730 2567.160 3.050 ;
        RECT 2571.960 2.730 2572.220 3.050 ;
        RECT 2572.020 2.400 2572.160 2.730 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
      LAYER via2 ;
        RECT 1275.210 72.960 1275.490 73.240 ;
        RECT 2566.890 72.960 2567.170 73.240 ;
      LAYER met3 ;
        RECT 1275.185 73.250 1275.515 73.265 ;
        RECT 2566.865 73.250 2567.195 73.265 ;
        RECT 1275.185 72.950 2567.195 73.250 ;
        RECT 1275.185 72.935 1275.515 72.950 ;
        RECT 2566.865 72.935 2567.195 72.950 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1277.030 1590.760 1277.350 1590.820 ;
        RECT 1282.090 1590.760 1282.410 1590.820 ;
        RECT 1277.030 1590.620 1282.410 1590.760 ;
        RECT 1277.030 1590.560 1277.350 1590.620 ;
        RECT 1282.090 1590.560 1282.410 1590.620 ;
        RECT 1282.090 67.900 1282.410 67.960 ;
        RECT 2587.570 67.900 2587.890 67.960 ;
        RECT 1282.090 67.760 2587.890 67.900 ;
        RECT 1282.090 67.700 1282.410 67.760 ;
        RECT 2587.570 67.700 2587.890 67.760 ;
      LAYER via ;
        RECT 1277.060 1590.560 1277.320 1590.820 ;
        RECT 1282.120 1590.560 1282.380 1590.820 ;
        RECT 1282.120 67.700 1282.380 67.960 ;
        RECT 2587.600 67.700 2587.860 67.960 ;
      LAYER met2 ;
        RECT 1277.060 1600.000 1277.340 1604.000 ;
        RECT 1277.120 1590.850 1277.260 1600.000 ;
        RECT 1277.060 1590.530 1277.320 1590.850 ;
        RECT 1282.120 1590.530 1282.380 1590.850 ;
        RECT 1282.180 67.990 1282.320 1590.530 ;
        RECT 1282.120 67.670 1282.380 67.990 ;
        RECT 2587.600 67.670 2587.860 67.990 ;
        RECT 2587.660 3.130 2587.800 67.670 ;
        RECT 2587.660 2.990 2589.640 3.130 ;
        RECT 2589.500 2.400 2589.640 2.990 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 762.365 1588.565 762.535 1590.775 ;
      LAYER mcon ;
        RECT 762.365 1590.605 762.535 1590.775 ;
      LAYER met1 ;
        RECT 610.490 1590.760 610.810 1590.820 ;
        RECT 762.305 1590.760 762.595 1590.805 ;
        RECT 610.490 1590.620 762.595 1590.760 ;
        RECT 610.490 1590.560 610.810 1590.620 ;
        RECT 762.305 1590.575 762.595 1590.620 ;
        RECT 762.305 1588.720 762.595 1588.765 ;
        RECT 797.250 1588.720 797.570 1588.780 ;
        RECT 762.305 1588.580 797.570 1588.720 ;
        RECT 762.305 1588.535 762.595 1588.580 ;
        RECT 797.250 1588.520 797.570 1588.580 ;
        RECT 797.250 19.280 797.570 19.340 ;
        RECT 823.470 19.280 823.790 19.340 ;
        RECT 797.250 19.140 823.790 19.280 ;
        RECT 797.250 19.080 797.570 19.140 ;
        RECT 823.470 19.080 823.790 19.140 ;
      LAYER via ;
        RECT 610.520 1590.560 610.780 1590.820 ;
        RECT 797.280 1588.520 797.540 1588.780 ;
        RECT 797.280 19.080 797.540 19.340 ;
        RECT 823.500 19.080 823.760 19.340 ;
      LAYER met2 ;
        RECT 610.520 1600.000 610.800 1604.000 ;
        RECT 610.580 1590.850 610.720 1600.000 ;
        RECT 610.520 1590.530 610.780 1590.850 ;
        RECT 797.280 1588.490 797.540 1588.810 ;
        RECT 797.340 19.370 797.480 1588.490 ;
        RECT 797.280 19.050 797.540 19.370 ;
        RECT 823.500 19.050 823.760 19.370 ;
        RECT 823.560 2.400 823.700 19.050 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1283.930 1590.760 1284.250 1590.820 ;
        RECT 1288.990 1590.760 1289.310 1590.820 ;
        RECT 1283.930 1590.620 1289.310 1590.760 ;
        RECT 1283.930 1590.560 1284.250 1590.620 ;
        RECT 1288.990 1590.560 1289.310 1590.620 ;
        RECT 1288.990 67.560 1289.310 67.620 ;
        RECT 2601.370 67.560 2601.690 67.620 ;
        RECT 1288.990 67.420 2601.690 67.560 ;
        RECT 1288.990 67.360 1289.310 67.420 ;
        RECT 2601.370 67.360 2601.690 67.420 ;
        RECT 2601.370 17.580 2601.690 17.640 ;
        RECT 2607.350 17.580 2607.670 17.640 ;
        RECT 2601.370 17.440 2607.670 17.580 ;
        RECT 2601.370 17.380 2601.690 17.440 ;
        RECT 2607.350 17.380 2607.670 17.440 ;
      LAYER via ;
        RECT 1283.960 1590.560 1284.220 1590.820 ;
        RECT 1289.020 1590.560 1289.280 1590.820 ;
        RECT 1289.020 67.360 1289.280 67.620 ;
        RECT 2601.400 67.360 2601.660 67.620 ;
        RECT 2601.400 17.380 2601.660 17.640 ;
        RECT 2607.380 17.380 2607.640 17.640 ;
      LAYER met2 ;
        RECT 1283.960 1600.000 1284.240 1604.000 ;
        RECT 1284.020 1590.850 1284.160 1600.000 ;
        RECT 1283.960 1590.530 1284.220 1590.850 ;
        RECT 1289.020 1590.530 1289.280 1590.850 ;
        RECT 1289.080 67.650 1289.220 1590.530 ;
        RECT 1289.020 67.330 1289.280 67.650 ;
        RECT 2601.400 67.330 2601.660 67.650 ;
        RECT 2601.460 17.670 2601.600 67.330 ;
        RECT 2601.400 17.350 2601.660 17.670 ;
        RECT 2607.380 17.350 2607.640 17.670 ;
        RECT 2607.440 2.400 2607.580 17.350 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1290.370 1590.760 1290.690 1590.820 ;
        RECT 1295.890 1590.760 1296.210 1590.820 ;
        RECT 1290.370 1590.620 1296.210 1590.760 ;
        RECT 1290.370 1590.560 1290.690 1590.620 ;
        RECT 1295.890 1590.560 1296.210 1590.620 ;
        RECT 1295.890 67.220 1296.210 67.280 ;
        RECT 2622.070 67.220 2622.390 67.280 ;
        RECT 1295.890 67.080 2622.390 67.220 ;
        RECT 1295.890 67.020 1296.210 67.080 ;
        RECT 2622.070 67.020 2622.390 67.080 ;
        RECT 2622.070 2.960 2622.390 3.020 ;
        RECT 2625.290 2.960 2625.610 3.020 ;
        RECT 2622.070 2.820 2625.610 2.960 ;
        RECT 2622.070 2.760 2622.390 2.820 ;
        RECT 2625.290 2.760 2625.610 2.820 ;
      LAYER via ;
        RECT 1290.400 1590.560 1290.660 1590.820 ;
        RECT 1295.920 1590.560 1296.180 1590.820 ;
        RECT 1295.920 67.020 1296.180 67.280 ;
        RECT 2622.100 67.020 2622.360 67.280 ;
        RECT 2622.100 2.760 2622.360 3.020 ;
        RECT 2625.320 2.760 2625.580 3.020 ;
      LAYER met2 ;
        RECT 1290.400 1600.000 1290.680 1604.000 ;
        RECT 1290.460 1590.850 1290.600 1600.000 ;
        RECT 1290.400 1590.530 1290.660 1590.850 ;
        RECT 1295.920 1590.530 1296.180 1590.850 ;
        RECT 1295.980 67.310 1296.120 1590.530 ;
        RECT 1295.920 66.990 1296.180 67.310 ;
        RECT 2622.100 66.990 2622.360 67.310 ;
        RECT 2622.160 3.050 2622.300 66.990 ;
        RECT 2622.100 2.730 2622.360 3.050 ;
        RECT 2625.320 2.730 2625.580 3.050 ;
        RECT 2625.380 2.400 2625.520 2.730 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1297.270 1587.700 1297.590 1587.760 ;
        RECT 1302.790 1587.700 1303.110 1587.760 ;
        RECT 1297.270 1587.560 1303.110 1587.700 ;
        RECT 1297.270 1587.500 1297.590 1587.560 ;
        RECT 1302.790 1587.500 1303.110 1587.560 ;
        RECT 1302.790 66.880 1303.110 66.940 ;
        RECT 2642.770 66.880 2643.090 66.940 ;
        RECT 1302.790 66.740 2643.090 66.880 ;
        RECT 1302.790 66.680 1303.110 66.740 ;
        RECT 2642.770 66.680 2643.090 66.740 ;
      LAYER via ;
        RECT 1297.300 1587.500 1297.560 1587.760 ;
        RECT 1302.820 1587.500 1303.080 1587.760 ;
        RECT 1302.820 66.680 1303.080 66.940 ;
        RECT 2642.800 66.680 2643.060 66.940 ;
      LAYER met2 ;
        RECT 1297.300 1600.000 1297.580 1604.000 ;
        RECT 1297.360 1587.790 1297.500 1600.000 ;
        RECT 1297.300 1587.470 1297.560 1587.790 ;
        RECT 1302.820 1587.470 1303.080 1587.790 ;
        RECT 1302.880 66.970 1303.020 1587.470 ;
        RECT 1302.820 66.650 1303.080 66.970 ;
        RECT 2642.800 66.650 2643.060 66.970 ;
        RECT 2642.860 17.410 2643.000 66.650 ;
        RECT 2642.860 17.270 2643.460 17.410 ;
        RECT 2643.320 2.400 2643.460 17.270 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1304.170 1589.400 1304.490 1589.460 ;
        RECT 1309.690 1589.400 1310.010 1589.460 ;
        RECT 1304.170 1589.260 1310.010 1589.400 ;
        RECT 1304.170 1589.200 1304.490 1589.260 ;
        RECT 1309.690 1589.200 1310.010 1589.260 ;
        RECT 1309.690 66.540 1310.010 66.600 ;
        RECT 2656.570 66.540 2656.890 66.600 ;
        RECT 1309.690 66.400 2656.890 66.540 ;
        RECT 1309.690 66.340 1310.010 66.400 ;
        RECT 2656.570 66.340 2656.890 66.400 ;
      LAYER via ;
        RECT 1304.200 1589.200 1304.460 1589.460 ;
        RECT 1309.720 1589.200 1309.980 1589.460 ;
        RECT 1309.720 66.340 1309.980 66.600 ;
        RECT 2656.600 66.340 2656.860 66.600 ;
      LAYER met2 ;
        RECT 1304.200 1600.000 1304.480 1604.000 ;
        RECT 1304.260 1589.490 1304.400 1600.000 ;
        RECT 1304.200 1589.170 1304.460 1589.490 ;
        RECT 1309.720 1589.170 1309.980 1589.490 ;
        RECT 1309.780 66.630 1309.920 1589.170 ;
        RECT 1309.720 66.310 1309.980 66.630 ;
        RECT 2656.600 66.310 2656.860 66.630 ;
        RECT 2656.660 17.410 2656.800 66.310 ;
        RECT 2656.660 17.270 2661.400 17.410 ;
        RECT 2661.260 2.400 2661.400 17.270 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1309.230 1590.760 1309.550 1590.820 ;
        RECT 1310.610 1590.760 1310.930 1590.820 ;
        RECT 1309.230 1590.620 1310.930 1590.760 ;
        RECT 1309.230 1590.560 1309.550 1590.620 ;
        RECT 1310.610 1590.560 1310.930 1590.620 ;
        RECT 1309.230 66.200 1309.550 66.260 ;
        RECT 2677.270 66.200 2677.590 66.260 ;
        RECT 1309.230 66.060 2677.590 66.200 ;
        RECT 1309.230 66.000 1309.550 66.060 ;
        RECT 2677.270 66.000 2677.590 66.060 ;
      LAYER via ;
        RECT 1309.260 1590.560 1309.520 1590.820 ;
        RECT 1310.640 1590.560 1310.900 1590.820 ;
        RECT 1309.260 66.000 1309.520 66.260 ;
        RECT 2677.300 66.000 2677.560 66.260 ;
      LAYER met2 ;
        RECT 1310.640 1600.000 1310.920 1604.000 ;
        RECT 1310.700 1590.850 1310.840 1600.000 ;
        RECT 1309.260 1590.530 1309.520 1590.850 ;
        RECT 1310.640 1590.530 1310.900 1590.850 ;
        RECT 1309.320 66.290 1309.460 1590.530 ;
        RECT 1309.260 65.970 1309.520 66.290 ;
        RECT 2677.300 65.970 2677.560 66.290 ;
        RECT 2677.360 17.410 2677.500 65.970 ;
        RECT 2677.360 17.270 2678.880 17.410 ;
        RECT 2678.740 2.400 2678.880 17.270 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1316.590 1590.760 1316.910 1590.820 ;
        RECT 1317.510 1590.760 1317.830 1590.820 ;
        RECT 1316.590 1590.620 1317.830 1590.760 ;
        RECT 1316.590 1590.560 1316.910 1590.620 ;
        RECT 1317.510 1590.560 1317.830 1590.620 ;
        RECT 1316.590 65.860 1316.910 65.920 ;
        RECT 2691.070 65.860 2691.390 65.920 ;
        RECT 1316.590 65.720 2691.390 65.860 ;
        RECT 1316.590 65.660 1316.910 65.720 ;
        RECT 2691.070 65.660 2691.390 65.720 ;
        RECT 2691.070 2.960 2691.390 3.020 ;
        RECT 2696.590 2.960 2696.910 3.020 ;
        RECT 2691.070 2.820 2696.910 2.960 ;
        RECT 2691.070 2.760 2691.390 2.820 ;
        RECT 2696.590 2.760 2696.910 2.820 ;
      LAYER via ;
        RECT 1316.620 1590.560 1316.880 1590.820 ;
        RECT 1317.540 1590.560 1317.800 1590.820 ;
        RECT 1316.620 65.660 1316.880 65.920 ;
        RECT 2691.100 65.660 2691.360 65.920 ;
        RECT 2691.100 2.760 2691.360 3.020 ;
        RECT 2696.620 2.760 2696.880 3.020 ;
      LAYER met2 ;
        RECT 1317.540 1600.000 1317.820 1604.000 ;
        RECT 1317.600 1590.850 1317.740 1600.000 ;
        RECT 1316.620 1590.530 1316.880 1590.850 ;
        RECT 1317.540 1590.530 1317.800 1590.850 ;
        RECT 1316.680 65.950 1316.820 1590.530 ;
        RECT 1316.620 65.630 1316.880 65.950 ;
        RECT 2691.100 65.630 2691.360 65.950 ;
        RECT 2691.160 3.050 2691.300 65.630 ;
        RECT 2691.100 2.730 2691.360 3.050 ;
        RECT 2696.620 2.730 2696.880 3.050 ;
        RECT 2696.680 2.400 2696.820 2.730 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1323.490 1590.760 1323.810 1590.820 ;
        RECT 1324.410 1590.760 1324.730 1590.820 ;
        RECT 1323.490 1590.620 1324.730 1590.760 ;
        RECT 1323.490 1590.560 1323.810 1590.620 ;
        RECT 1324.410 1590.560 1324.730 1590.620 ;
        RECT 1323.490 65.520 1323.810 65.580 ;
        RECT 2711.770 65.520 2712.090 65.580 ;
        RECT 1323.490 65.380 2712.090 65.520 ;
        RECT 1323.490 65.320 1323.810 65.380 ;
        RECT 2711.770 65.320 2712.090 65.380 ;
        RECT 2711.770 2.960 2712.090 3.020 ;
        RECT 2714.530 2.960 2714.850 3.020 ;
        RECT 2711.770 2.820 2714.850 2.960 ;
        RECT 2711.770 2.760 2712.090 2.820 ;
        RECT 2714.530 2.760 2714.850 2.820 ;
      LAYER via ;
        RECT 1323.520 1590.560 1323.780 1590.820 ;
        RECT 1324.440 1590.560 1324.700 1590.820 ;
        RECT 1323.520 65.320 1323.780 65.580 ;
        RECT 2711.800 65.320 2712.060 65.580 ;
        RECT 2711.800 2.760 2712.060 3.020 ;
        RECT 2714.560 2.760 2714.820 3.020 ;
      LAYER met2 ;
        RECT 1324.440 1600.000 1324.720 1604.000 ;
        RECT 1324.500 1590.850 1324.640 1600.000 ;
        RECT 1323.520 1590.530 1323.780 1590.850 ;
        RECT 1324.440 1590.530 1324.700 1590.850 ;
        RECT 1323.580 65.610 1323.720 1590.530 ;
        RECT 1323.520 65.290 1323.780 65.610 ;
        RECT 2711.800 65.290 2712.060 65.610 ;
        RECT 2711.860 3.050 2712.000 65.290 ;
        RECT 2711.800 2.730 2712.060 3.050 ;
        RECT 2714.560 2.730 2714.820 3.050 ;
        RECT 2714.620 2.400 2714.760 2.730 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1330.880 1600.000 1331.160 1604.000 ;
        RECT 1330.940 67.845 1331.080 1600.000 ;
        RECT 1330.870 67.475 1331.150 67.845 ;
        RECT 2732.490 67.475 2732.770 67.845 ;
        RECT 2732.560 2.400 2732.700 67.475 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
      LAYER via2 ;
        RECT 1330.870 67.520 1331.150 67.800 ;
        RECT 2732.490 67.520 2732.770 67.800 ;
      LAYER met3 ;
        RECT 1330.845 67.810 1331.175 67.825 ;
        RECT 2732.465 67.810 2732.795 67.825 ;
        RECT 1330.845 67.510 2732.795 67.810 ;
        RECT 1330.845 67.495 1331.175 67.510 ;
        RECT 2732.465 67.495 2732.795 67.510 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2746.270 2.960 2746.590 3.020 ;
        RECT 2750.410 2.960 2750.730 3.020 ;
        RECT 2746.270 2.820 2750.730 2.960 ;
        RECT 2746.270 2.760 2746.590 2.820 ;
        RECT 2750.410 2.760 2750.730 2.820 ;
      LAYER via ;
        RECT 2746.300 2.760 2746.560 3.020 ;
        RECT 2750.440 2.760 2750.700 3.020 ;
      LAYER met2 ;
        RECT 1337.780 1600.450 1338.060 1604.000 ;
        RECT 1337.380 1600.310 1338.060 1600.450 ;
        RECT 1337.380 67.165 1337.520 1600.310 ;
        RECT 1337.780 1600.000 1338.060 1600.310 ;
        RECT 1337.310 66.795 1337.590 67.165 ;
        RECT 2746.290 66.795 2746.570 67.165 ;
        RECT 2746.360 3.050 2746.500 66.795 ;
        RECT 2746.300 2.730 2746.560 3.050 ;
        RECT 2750.440 2.730 2750.700 3.050 ;
        RECT 2750.500 2.400 2750.640 2.730 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
      LAYER via2 ;
        RECT 1337.310 66.840 1337.590 67.120 ;
        RECT 2746.290 66.840 2746.570 67.120 ;
      LAYER met3 ;
        RECT 1337.285 67.130 1337.615 67.145 ;
        RECT 2746.265 67.130 2746.595 67.145 ;
        RECT 1337.285 66.830 2746.595 67.130 ;
        RECT 1337.285 66.815 1337.615 66.830 ;
        RECT 2746.265 66.815 2746.595 66.830 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1344.680 1600.450 1344.960 1604.000 ;
        RECT 1344.280 1600.310 1344.960 1600.450 ;
        RECT 1344.280 66.485 1344.420 1600.310 ;
        RECT 1344.680 1600.000 1344.960 1600.310 ;
        RECT 1344.210 66.115 1344.490 66.485 ;
        RECT 2766.990 66.115 2767.270 66.485 ;
        RECT 2767.060 3.130 2767.200 66.115 ;
        RECT 2767.060 2.990 2768.120 3.130 ;
        RECT 2767.980 2.400 2768.120 2.990 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
      LAYER via2 ;
        RECT 1344.210 66.160 1344.490 66.440 ;
        RECT 2766.990 66.160 2767.270 66.440 ;
      LAYER met3 ;
        RECT 1344.185 66.450 1344.515 66.465 ;
        RECT 2766.965 66.450 2767.295 66.465 ;
        RECT 1344.185 66.150 2767.295 66.450 ;
        RECT 1344.185 66.135 1344.515 66.150 ;
        RECT 2766.965 66.135 2767.295 66.150 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 633.565 14.025 633.735 18.615 ;
        RECT 687.845 14.025 688.015 19.635 ;
      LAYER mcon ;
        RECT 687.845 19.465 688.015 19.635 ;
        RECT 633.565 18.445 633.735 18.615 ;
      LAYER met1 ;
        RECT 617.390 1588.040 617.710 1588.100 ;
        RECT 620.610 1588.040 620.930 1588.100 ;
        RECT 617.390 1587.900 620.930 1588.040 ;
        RECT 617.390 1587.840 617.710 1587.900 ;
        RECT 620.610 1587.840 620.930 1587.900 ;
        RECT 687.785 19.620 688.075 19.665 ;
        RECT 840.950 19.620 841.270 19.680 ;
        RECT 687.785 19.480 841.270 19.620 ;
        RECT 687.785 19.435 688.075 19.480 ;
        RECT 840.950 19.420 841.270 19.480 ;
        RECT 620.610 18.600 620.930 18.660 ;
        RECT 633.505 18.600 633.795 18.645 ;
        RECT 620.610 18.460 633.795 18.600 ;
        RECT 620.610 18.400 620.930 18.460 ;
        RECT 633.505 18.415 633.795 18.460 ;
        RECT 633.505 14.180 633.795 14.225 ;
        RECT 647.750 14.180 648.070 14.240 ;
        RECT 633.505 14.040 648.070 14.180 ;
        RECT 633.505 13.995 633.795 14.040 ;
        RECT 647.750 13.980 648.070 14.040 ;
        RECT 669.830 14.180 670.150 14.240 ;
        RECT 687.785 14.180 688.075 14.225 ;
        RECT 669.830 14.040 688.075 14.180 ;
        RECT 669.830 13.980 670.150 14.040 ;
        RECT 687.785 13.995 688.075 14.040 ;
      LAYER via ;
        RECT 617.420 1587.840 617.680 1588.100 ;
        RECT 620.640 1587.840 620.900 1588.100 ;
        RECT 840.980 19.420 841.240 19.680 ;
        RECT 620.640 18.400 620.900 18.660 ;
        RECT 647.780 13.980 648.040 14.240 ;
        RECT 669.860 13.980 670.120 14.240 ;
      LAYER met2 ;
        RECT 617.420 1600.000 617.700 1604.000 ;
        RECT 617.480 1588.130 617.620 1600.000 ;
        RECT 617.420 1587.810 617.680 1588.130 ;
        RECT 620.640 1587.810 620.900 1588.130 ;
        RECT 620.700 18.690 620.840 1587.810 ;
        RECT 840.980 19.390 841.240 19.710 ;
        RECT 620.640 18.370 620.900 18.690 ;
        RECT 647.780 14.125 648.040 14.270 ;
        RECT 669.860 14.125 670.120 14.270 ;
        RECT 647.770 13.755 648.050 14.125 ;
        RECT 669.850 13.755 670.130 14.125 ;
        RECT 841.040 2.400 841.180 19.390 ;
        RECT 840.830 -4.800 841.390 2.400 ;
      LAYER via2 ;
        RECT 647.770 13.800 648.050 14.080 ;
        RECT 669.850 13.800 670.130 14.080 ;
      LAYER met3 ;
        RECT 647.745 14.090 648.075 14.105 ;
        RECT 669.825 14.090 670.155 14.105 ;
        RECT 647.745 13.790 670.155 14.090 ;
        RECT 647.745 13.775 648.075 13.790 ;
        RECT 669.825 13.775 670.155 13.790 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2780.770 2.960 2781.090 3.020 ;
        RECT 2785.830 2.960 2786.150 3.020 ;
        RECT 2780.770 2.820 2786.150 2.960 ;
        RECT 2780.770 2.760 2781.090 2.820 ;
        RECT 2785.830 2.760 2786.150 2.820 ;
      LAYER via ;
        RECT 2780.800 2.760 2781.060 3.020 ;
        RECT 2785.860 2.760 2786.120 3.020 ;
      LAYER met2 ;
        RECT 1351.120 1600.000 1351.400 1604.000 ;
        RECT 1351.180 65.805 1351.320 1600.000 ;
        RECT 1351.110 65.435 1351.390 65.805 ;
        RECT 2780.790 65.435 2781.070 65.805 ;
        RECT 2780.860 3.050 2781.000 65.435 ;
        RECT 2780.800 2.730 2781.060 3.050 ;
        RECT 2785.860 2.730 2786.120 3.050 ;
        RECT 2785.920 2.400 2786.060 2.730 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
      LAYER via2 ;
        RECT 1351.110 65.480 1351.390 65.760 ;
        RECT 2780.790 65.480 2781.070 65.760 ;
      LAYER met3 ;
        RECT 1351.085 65.770 1351.415 65.785 ;
        RECT 2780.765 65.770 2781.095 65.785 ;
        RECT 1351.085 65.470 2781.095 65.770 ;
        RECT 1351.085 65.455 1351.415 65.470 ;
        RECT 2780.765 65.455 2781.095 65.470 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.020 1600.000 1358.300 1604.000 ;
        RECT 1358.080 65.125 1358.220 1600.000 ;
        RECT 1358.010 64.755 1358.290 65.125 ;
        RECT 2801.490 64.755 2801.770 65.125 ;
        RECT 2801.560 17.410 2801.700 64.755 ;
        RECT 2801.560 17.270 2804.000 17.410 ;
        RECT 2803.860 2.400 2804.000 17.270 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
      LAYER via2 ;
        RECT 1358.010 64.800 1358.290 65.080 ;
        RECT 2801.490 64.800 2801.770 65.080 ;
      LAYER met3 ;
        RECT 1357.985 65.090 1358.315 65.105 ;
        RECT 2801.465 65.090 2801.795 65.105 ;
        RECT 1357.985 64.790 2801.795 65.090 ;
        RECT 1357.985 64.775 1358.315 64.790 ;
        RECT 2801.465 64.775 2801.795 64.790 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1386.585 1590.265 1386.755 1592.475 ;
      LAYER mcon ;
        RECT 1386.585 1592.305 1386.755 1592.475 ;
      LAYER met1 ;
        RECT 1364.430 1592.460 1364.750 1592.520 ;
        RECT 1386.525 1592.460 1386.815 1592.505 ;
        RECT 1364.430 1592.320 1386.815 1592.460 ;
        RECT 1364.430 1592.260 1364.750 1592.320 ;
        RECT 1386.525 1592.275 1386.815 1592.320 ;
        RECT 1386.525 1590.420 1386.815 1590.465 ;
        RECT 2647.370 1590.420 2647.690 1590.480 ;
        RECT 1386.525 1590.280 2647.690 1590.420 ;
        RECT 1386.525 1590.235 1386.815 1590.280 ;
        RECT 2647.370 1590.220 2647.690 1590.280 ;
        RECT 2647.370 17.580 2647.690 17.640 ;
        RECT 2821.710 17.580 2822.030 17.640 ;
        RECT 2647.370 17.440 2822.030 17.580 ;
        RECT 2647.370 17.380 2647.690 17.440 ;
        RECT 2821.710 17.380 2822.030 17.440 ;
      LAYER via ;
        RECT 1364.460 1592.260 1364.720 1592.520 ;
        RECT 2647.400 1590.220 2647.660 1590.480 ;
        RECT 2647.400 17.380 2647.660 17.640 ;
        RECT 2821.740 17.380 2822.000 17.640 ;
      LAYER met2 ;
        RECT 1364.460 1600.000 1364.740 1604.000 ;
        RECT 1364.520 1592.550 1364.660 1600.000 ;
        RECT 1364.460 1592.230 1364.720 1592.550 ;
        RECT 2647.400 1590.190 2647.660 1590.510 ;
        RECT 2647.460 17.670 2647.600 1590.190 ;
        RECT 2647.400 17.350 2647.660 17.670 ;
        RECT 2821.740 17.350 2822.000 17.670 ;
        RECT 2821.800 2.400 2821.940 17.350 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1371.790 80.140 1372.110 80.200 ;
        RECT 2835.970 80.140 2836.290 80.200 ;
        RECT 1371.790 80.000 2836.290 80.140 ;
        RECT 1371.790 79.940 1372.110 80.000 ;
        RECT 2835.970 79.940 2836.290 80.000 ;
      LAYER via ;
        RECT 1371.820 79.940 1372.080 80.200 ;
        RECT 2836.000 79.940 2836.260 80.200 ;
      LAYER met2 ;
        RECT 1371.360 1600.450 1371.640 1604.000 ;
        RECT 1371.360 1600.310 1372.020 1600.450 ;
        RECT 1371.360 1600.000 1371.640 1600.310 ;
        RECT 1371.880 80.230 1372.020 1600.310 ;
        RECT 1371.820 79.910 1372.080 80.230 ;
        RECT 2836.000 79.910 2836.260 80.230 ;
        RECT 2836.060 17.410 2836.200 79.910 ;
        RECT 2836.060 17.270 2839.420 17.410 ;
        RECT 2839.280 2.400 2839.420 17.270 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1378.230 1590.760 1378.550 1590.820 ;
        RECT 2646.910 1590.760 2647.230 1590.820 ;
        RECT 1378.230 1590.620 2647.230 1590.760 ;
        RECT 1378.230 1590.560 1378.550 1590.620 ;
        RECT 2646.910 1590.560 2647.230 1590.620 ;
        RECT 2646.910 17.240 2647.230 17.300 ;
        RECT 2857.130 17.240 2857.450 17.300 ;
        RECT 2646.910 17.100 2857.450 17.240 ;
        RECT 2646.910 17.040 2647.230 17.100 ;
        RECT 2857.130 17.040 2857.450 17.100 ;
      LAYER via ;
        RECT 1378.260 1590.560 1378.520 1590.820 ;
        RECT 2646.940 1590.560 2647.200 1590.820 ;
        RECT 2646.940 17.040 2647.200 17.300 ;
        RECT 2857.160 17.040 2857.420 17.300 ;
      LAYER met2 ;
        RECT 1378.260 1600.000 1378.540 1604.000 ;
        RECT 1378.320 1590.850 1378.460 1600.000 ;
        RECT 1378.260 1590.530 1378.520 1590.850 ;
        RECT 2646.940 1590.530 2647.200 1590.850 ;
        RECT 2647.000 17.330 2647.140 1590.530 ;
        RECT 2646.940 17.010 2647.200 17.330 ;
        RECT 2857.160 17.010 2857.420 17.330 ;
        RECT 2857.220 2.400 2857.360 17.010 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1385.590 79.800 1385.910 79.860 ;
        RECT 2870.470 79.800 2870.790 79.860 ;
        RECT 1385.590 79.660 2870.790 79.800 ;
        RECT 1385.590 79.600 1385.910 79.660 ;
        RECT 2870.470 79.600 2870.790 79.660 ;
      LAYER via ;
        RECT 1385.620 79.600 1385.880 79.860 ;
        RECT 2870.500 79.600 2870.760 79.860 ;
      LAYER met2 ;
        RECT 1384.700 1600.450 1384.980 1604.000 ;
        RECT 1384.700 1600.310 1385.820 1600.450 ;
        RECT 1384.700 1600.000 1384.980 1600.310 ;
        RECT 1385.680 79.890 1385.820 1600.310 ;
        RECT 1385.620 79.570 1385.880 79.890 ;
        RECT 2870.500 79.570 2870.760 79.890 ;
        RECT 2870.560 17.410 2870.700 79.570 ;
        RECT 2870.560 17.270 2875.300 17.410 ;
        RECT 2875.160 2.400 2875.300 17.270 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1392.490 79.460 1392.810 79.520 ;
        RECT 2891.170 79.460 2891.490 79.520 ;
        RECT 1392.490 79.320 2891.490 79.460 ;
        RECT 1392.490 79.260 1392.810 79.320 ;
        RECT 2891.170 79.260 2891.490 79.320 ;
      LAYER via ;
        RECT 1392.520 79.260 1392.780 79.520 ;
        RECT 2891.200 79.260 2891.460 79.520 ;
      LAYER met2 ;
        RECT 1391.600 1600.450 1391.880 1604.000 ;
        RECT 1391.600 1600.310 1392.720 1600.450 ;
        RECT 1391.600 1600.000 1391.880 1600.310 ;
        RECT 1392.580 79.550 1392.720 1600.310 ;
        RECT 1392.520 79.230 1392.780 79.550 ;
        RECT 2891.200 79.230 2891.460 79.550 ;
        RECT 2891.260 3.130 2891.400 79.230 ;
        RECT 2891.260 2.990 2893.240 3.130 ;
        RECT 2893.100 2.400 2893.240 2.990 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1398.500 1600.000 1398.780 1604.000 ;
        RECT 1398.560 1591.725 1398.700 1600.000 ;
        RECT 1398.490 1591.355 1398.770 1591.725 ;
        RECT 1609.170 16.475 1609.450 16.845 ;
        RECT 2910.970 16.475 2911.250 16.845 ;
        RECT 1609.240 15.485 1609.380 16.475 ;
        RECT 1609.170 15.115 1609.450 15.485 ;
        RECT 2911.040 2.400 2911.180 16.475 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 1398.490 1591.400 1398.770 1591.680 ;
        RECT 1609.170 16.520 1609.450 16.800 ;
        RECT 2910.970 16.520 2911.250 16.800 ;
        RECT 1609.170 15.160 1609.450 15.440 ;
      LAYER met3 ;
        RECT 1398.465 1591.690 1398.795 1591.705 ;
        RECT 1603.830 1591.690 1604.210 1591.700 ;
        RECT 1398.465 1591.390 1604.210 1591.690 ;
        RECT 1398.465 1591.375 1398.795 1591.390 ;
        RECT 1603.830 1591.380 1604.210 1591.390 ;
        RECT 1609.145 16.810 1609.475 16.825 ;
        RECT 2910.945 16.810 2911.275 16.825 ;
        RECT 1609.145 16.510 2911.275 16.810 ;
        RECT 1609.145 16.495 1609.475 16.510 ;
        RECT 2910.945 16.495 2911.275 16.510 ;
        RECT 1603.830 15.450 1604.210 15.460 ;
        RECT 1609.145 15.450 1609.475 15.465 ;
        RECT 1603.830 15.150 1609.475 15.450 ;
        RECT 1603.830 15.140 1604.210 15.150 ;
        RECT 1609.145 15.135 1609.475 15.150 ;
      LAYER via3 ;
        RECT 1603.860 1591.380 1604.180 1591.700 ;
        RECT 1603.860 15.140 1604.180 15.460 ;
      LAYER met4 ;
        RECT 1603.855 1591.375 1604.185 1591.705 ;
        RECT 1603.870 15.465 1604.170 1591.375 ;
        RECT 1603.855 15.135 1604.185 15.465 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 803.765 1545.725 803.935 1592.475 ;
        RECT 803.765 386.325 803.935 434.435 ;
        RECT 810.205 14.875 810.375 15.555 ;
        RECT 810.205 14.705 811.295 14.875 ;
      LAYER mcon ;
        RECT 803.765 1592.305 803.935 1592.475 ;
        RECT 803.765 434.265 803.935 434.435 ;
        RECT 810.205 15.385 810.375 15.555 ;
        RECT 811.125 14.705 811.295 14.875 ;
      LAYER met1 ;
        RECT 623.830 1592.460 624.150 1592.520 ;
        RECT 803.705 1592.460 803.995 1592.505 ;
        RECT 623.830 1592.320 803.995 1592.460 ;
        RECT 623.830 1592.260 624.150 1592.320 ;
        RECT 803.705 1592.275 803.995 1592.320 ;
        RECT 803.690 1545.880 804.010 1545.940 ;
        RECT 803.495 1545.740 804.010 1545.880 ;
        RECT 803.690 1545.680 804.010 1545.740 ;
        RECT 802.770 966.180 803.090 966.240 ;
        RECT 803.690 966.180 804.010 966.240 ;
        RECT 802.770 966.040 804.010 966.180 ;
        RECT 802.770 965.980 803.090 966.040 ;
        RECT 803.690 965.980 804.010 966.040 ;
        RECT 803.690 434.420 804.010 434.480 ;
        RECT 803.495 434.280 804.010 434.420 ;
        RECT 803.690 434.220 804.010 434.280 ;
        RECT 803.690 386.480 804.010 386.540 ;
        RECT 803.495 386.340 804.010 386.480 ;
        RECT 803.690 386.280 804.010 386.340 ;
        RECT 803.230 96.800 803.550 96.860 ;
        RECT 803.690 96.800 804.010 96.860 ;
        RECT 803.230 96.660 804.010 96.800 ;
        RECT 803.230 96.600 803.550 96.660 ;
        RECT 803.690 96.600 804.010 96.660 ;
        RECT 803.690 15.540 804.010 15.600 ;
        RECT 810.145 15.540 810.435 15.585 ;
        RECT 803.690 15.400 810.435 15.540 ;
        RECT 803.690 15.340 804.010 15.400 ;
        RECT 810.145 15.355 810.435 15.400 ;
        RECT 811.065 14.860 811.355 14.905 ;
        RECT 858.890 14.860 859.210 14.920 ;
        RECT 811.065 14.720 859.210 14.860 ;
        RECT 811.065 14.675 811.355 14.720 ;
        RECT 858.890 14.660 859.210 14.720 ;
      LAYER via ;
        RECT 623.860 1592.260 624.120 1592.520 ;
        RECT 803.720 1545.680 803.980 1545.940 ;
        RECT 802.800 965.980 803.060 966.240 ;
        RECT 803.720 965.980 803.980 966.240 ;
        RECT 803.720 434.220 803.980 434.480 ;
        RECT 803.720 386.280 803.980 386.540 ;
        RECT 803.260 96.600 803.520 96.860 ;
        RECT 803.720 96.600 803.980 96.860 ;
        RECT 803.720 15.340 803.980 15.600 ;
        RECT 858.920 14.660 859.180 14.920 ;
      LAYER met2 ;
        RECT 623.860 1600.000 624.140 1604.000 ;
        RECT 623.920 1592.550 624.060 1600.000 ;
        RECT 623.860 1592.230 624.120 1592.550 ;
        RECT 803.720 1545.650 803.980 1545.970 ;
        RECT 803.780 1014.405 803.920 1545.650 ;
        RECT 802.790 1014.035 803.070 1014.405 ;
        RECT 803.710 1014.035 803.990 1014.405 ;
        RECT 802.860 966.270 803.000 1014.035 ;
        RECT 802.800 965.950 803.060 966.270 ;
        RECT 803.720 965.950 803.980 966.270 ;
        RECT 803.780 434.510 803.920 965.950 ;
        RECT 803.720 434.190 803.980 434.510 ;
        RECT 803.720 386.250 803.980 386.570 ;
        RECT 803.780 144.570 803.920 386.250 ;
        RECT 803.320 144.430 803.920 144.570 ;
        RECT 803.320 96.890 803.460 144.430 ;
        RECT 803.260 96.570 803.520 96.890 ;
        RECT 803.720 96.570 803.980 96.890 ;
        RECT 803.780 15.630 803.920 96.570 ;
        RECT 803.720 15.310 803.980 15.630 ;
        RECT 858.920 14.630 859.180 14.950 ;
        RECT 858.980 2.400 859.120 14.630 ;
        RECT 858.770 -4.800 859.330 2.400 ;
      LAYER via2 ;
        RECT 802.790 1014.080 803.070 1014.360 ;
        RECT 803.710 1014.080 803.990 1014.360 ;
      LAYER met3 ;
        RECT 802.765 1014.370 803.095 1014.385 ;
        RECT 803.685 1014.370 804.015 1014.385 ;
        RECT 802.765 1014.070 804.015 1014.370 ;
        RECT 802.765 1014.055 803.095 1014.070 ;
        RECT 803.685 1014.055 804.015 1014.070 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 630.730 1591.780 631.050 1591.840 ;
        RECT 824.390 1591.780 824.710 1591.840 ;
        RECT 630.730 1591.640 824.710 1591.780 ;
        RECT 630.730 1591.580 631.050 1591.640 ;
        RECT 824.390 1591.580 824.710 1591.640 ;
        RECT 824.390 15.540 824.710 15.600 ;
        RECT 876.830 15.540 877.150 15.600 ;
        RECT 824.390 15.400 877.150 15.540 ;
        RECT 824.390 15.340 824.710 15.400 ;
        RECT 876.830 15.340 877.150 15.400 ;
      LAYER via ;
        RECT 630.760 1591.580 631.020 1591.840 ;
        RECT 824.420 1591.580 824.680 1591.840 ;
        RECT 824.420 15.340 824.680 15.600 ;
        RECT 876.860 15.340 877.120 15.600 ;
      LAYER met2 ;
        RECT 630.760 1600.000 631.040 1604.000 ;
        RECT 630.820 1591.870 630.960 1600.000 ;
        RECT 630.760 1591.550 631.020 1591.870 ;
        RECT 824.420 1591.550 824.680 1591.870 ;
        RECT 824.480 15.630 824.620 1591.550 ;
        RECT 824.420 15.310 824.680 15.630 ;
        RECT 876.860 15.310 877.120 15.630 ;
        RECT 876.920 2.400 877.060 15.310 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 637.170 1591.440 637.490 1591.500 ;
        RECT 831.750 1591.440 832.070 1591.500 ;
        RECT 637.170 1591.300 832.070 1591.440 ;
        RECT 637.170 1591.240 637.490 1591.300 ;
        RECT 831.750 1591.240 832.070 1591.300 ;
        RECT 831.750 16.900 832.070 16.960 ;
        RECT 894.770 16.900 895.090 16.960 ;
        RECT 831.750 16.760 895.090 16.900 ;
        RECT 831.750 16.700 832.070 16.760 ;
        RECT 894.770 16.700 895.090 16.760 ;
      LAYER via ;
        RECT 637.200 1591.240 637.460 1591.500 ;
        RECT 831.780 1591.240 832.040 1591.500 ;
        RECT 831.780 16.700 832.040 16.960 ;
        RECT 894.800 16.700 895.060 16.960 ;
      LAYER met2 ;
        RECT 637.200 1600.000 637.480 1604.000 ;
        RECT 637.260 1591.530 637.400 1600.000 ;
        RECT 637.200 1591.210 637.460 1591.530 ;
        RECT 831.780 1591.210 832.040 1591.530 ;
        RECT 831.840 16.990 831.980 1591.210 ;
        RECT 831.780 16.670 832.040 16.990 ;
        RECT 894.800 16.670 895.060 16.990 ;
        RECT 894.860 2.400 895.000 16.670 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 669.445 14.025 669.615 18.615 ;
        RECT 741.205 16.745 741.375 18.615 ;
        RECT 810.665 16.745 810.835 18.615 ;
      LAYER mcon ;
        RECT 669.445 18.445 669.615 18.615 ;
        RECT 741.205 18.445 741.375 18.615 ;
        RECT 810.665 18.445 810.835 18.615 ;
      LAYER met1 ;
        RECT 644.070 1587.360 644.390 1587.420 ;
        RECT 648.210 1587.360 648.530 1587.420 ;
        RECT 644.070 1587.220 648.530 1587.360 ;
        RECT 644.070 1587.160 644.390 1587.220 ;
        RECT 648.210 1587.160 648.530 1587.220 ;
        RECT 912.710 19.960 913.030 20.020 ;
        RECT 883.820 19.820 913.030 19.960 ;
        RECT 883.820 19.620 883.960 19.820 ;
        RECT 912.710 19.760 913.030 19.820 ;
        RECT 883.360 19.480 883.960 19.620 ;
        RECT 883.360 18.940 883.500 19.480 ;
        RECT 858.980 18.800 883.500 18.940 ;
        RECT 669.385 18.600 669.675 18.645 ;
        RECT 741.145 18.600 741.435 18.645 ;
        RECT 669.385 18.460 741.435 18.600 ;
        RECT 669.385 18.415 669.675 18.460 ;
        RECT 741.145 18.415 741.435 18.460 ;
        RECT 810.605 18.600 810.895 18.645 ;
        RECT 858.980 18.600 859.120 18.800 ;
        RECT 810.605 18.460 859.120 18.600 ;
        RECT 810.605 18.415 810.895 18.460 ;
        RECT 741.145 16.900 741.435 16.945 ;
        RECT 810.605 16.900 810.895 16.945 ;
        RECT 741.145 16.760 810.895 16.900 ;
        RECT 741.145 16.715 741.435 16.760 ;
        RECT 810.605 16.715 810.895 16.760 ;
        RECT 648.210 14.180 648.530 14.240 ;
        RECT 669.385 14.180 669.675 14.225 ;
        RECT 648.210 14.040 669.675 14.180 ;
        RECT 648.210 13.980 648.530 14.040 ;
        RECT 669.385 13.995 669.675 14.040 ;
      LAYER via ;
        RECT 644.100 1587.160 644.360 1587.420 ;
        RECT 648.240 1587.160 648.500 1587.420 ;
        RECT 912.740 19.760 913.000 20.020 ;
        RECT 648.240 13.980 648.500 14.240 ;
      LAYER met2 ;
        RECT 644.100 1600.000 644.380 1604.000 ;
        RECT 644.160 1587.450 644.300 1600.000 ;
        RECT 644.100 1587.130 644.360 1587.450 ;
        RECT 648.240 1587.130 648.500 1587.450 ;
        RECT 648.300 14.270 648.440 1587.130 ;
        RECT 912.740 19.730 913.000 20.050 ;
        RECT 648.240 13.950 648.500 14.270 ;
        RECT 912.800 2.400 912.940 19.730 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 879.665 19.805 883.055 19.975 ;
        RECT 849.305 18.955 849.475 19.635 ;
        RECT 849.305 18.785 850.395 18.955 ;
        RECT 858.505 18.615 858.675 18.955 ;
        RECT 858.505 18.445 859.595 18.615 ;
        RECT 879.665 18.445 879.835 19.805 ;
        RECT 883.345 19.295 883.515 19.975 ;
        RECT 883.345 19.125 884.435 19.295 ;
        RECT 884.265 15.045 884.435 19.125 ;
        RECT 906.805 15.045 906.975 16.235 ;
      LAYER mcon ;
        RECT 882.885 19.805 883.055 19.975 ;
        RECT 883.345 19.805 883.515 19.975 ;
        RECT 849.305 19.465 849.475 19.635 ;
        RECT 850.225 18.785 850.395 18.955 ;
        RECT 858.505 18.785 858.675 18.955 ;
        RECT 859.425 18.445 859.595 18.615 ;
        RECT 906.805 16.065 906.975 16.235 ;
      LAYER met1 ;
        RECT 650.970 1592.120 651.290 1592.180 ;
        RECT 838.190 1592.120 838.510 1592.180 ;
        RECT 650.970 1591.980 838.510 1592.120 ;
        RECT 650.970 1591.920 651.290 1591.980 ;
        RECT 838.190 1591.920 838.510 1591.980 ;
        RECT 838.190 19.960 838.510 20.020 ;
        RECT 882.825 19.960 883.115 20.005 ;
        RECT 883.285 19.960 883.575 20.005 ;
        RECT 838.190 19.820 841.640 19.960 ;
        RECT 838.190 19.760 838.510 19.820 ;
        RECT 841.500 19.620 841.640 19.820 ;
        RECT 882.825 19.820 883.575 19.960 ;
        RECT 882.825 19.775 883.115 19.820 ;
        RECT 883.285 19.775 883.575 19.820 ;
        RECT 849.245 19.620 849.535 19.665 ;
        RECT 841.500 19.480 849.535 19.620 ;
        RECT 849.245 19.435 849.535 19.480 ;
        RECT 850.165 18.940 850.455 18.985 ;
        RECT 858.445 18.940 858.735 18.985 ;
        RECT 850.165 18.800 858.735 18.940 ;
        RECT 850.165 18.755 850.455 18.800 ;
        RECT 858.445 18.755 858.735 18.800 ;
        RECT 859.365 18.600 859.655 18.645 ;
        RECT 879.605 18.600 879.895 18.645 ;
        RECT 859.365 18.460 879.895 18.600 ;
        RECT 859.365 18.415 859.655 18.460 ;
        RECT 879.605 18.415 879.895 18.460 ;
        RECT 906.745 16.220 907.035 16.265 ;
        RECT 930.190 16.220 930.510 16.280 ;
        RECT 906.745 16.080 930.510 16.220 ;
        RECT 906.745 16.035 907.035 16.080 ;
        RECT 930.190 16.020 930.510 16.080 ;
        RECT 884.205 15.200 884.495 15.245 ;
        RECT 906.745 15.200 907.035 15.245 ;
        RECT 884.205 15.060 907.035 15.200 ;
        RECT 884.205 15.015 884.495 15.060 ;
        RECT 906.745 15.015 907.035 15.060 ;
      LAYER via ;
        RECT 651.000 1591.920 651.260 1592.180 ;
        RECT 838.220 1591.920 838.480 1592.180 ;
        RECT 838.220 19.760 838.480 20.020 ;
        RECT 930.220 16.020 930.480 16.280 ;
      LAYER met2 ;
        RECT 651.000 1600.000 651.280 1604.000 ;
        RECT 651.060 1592.210 651.200 1600.000 ;
        RECT 651.000 1591.890 651.260 1592.210 ;
        RECT 838.220 1591.890 838.480 1592.210 ;
        RECT 838.280 20.050 838.420 1591.890 ;
        RECT 838.220 19.730 838.480 20.050 ;
        RECT 930.220 15.990 930.480 16.310 ;
        RECT 930.280 2.400 930.420 15.990 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 657.410 1587.360 657.730 1587.420 ;
        RECT 662.010 1587.360 662.330 1587.420 ;
        RECT 657.410 1587.220 662.330 1587.360 ;
        RECT 657.410 1587.160 657.730 1587.220 ;
        RECT 662.010 1587.160 662.330 1587.220 ;
        RECT 662.010 18.260 662.330 18.320 ;
        RECT 948.130 18.260 948.450 18.320 ;
        RECT 662.010 18.120 663.620 18.260 ;
        RECT 662.010 18.060 662.330 18.120 ;
        RECT 663.480 17.920 663.620 18.120 ;
        RECT 686.940 18.120 948.450 18.260 ;
        RECT 686.940 17.920 687.080 18.120 ;
        RECT 948.130 18.060 948.450 18.120 ;
        RECT 663.480 17.780 687.080 17.920 ;
      LAYER via ;
        RECT 657.440 1587.160 657.700 1587.420 ;
        RECT 662.040 1587.160 662.300 1587.420 ;
        RECT 662.040 18.060 662.300 18.320 ;
        RECT 948.160 18.060 948.420 18.320 ;
      LAYER met2 ;
        RECT 657.440 1600.000 657.720 1604.000 ;
        RECT 657.500 1587.450 657.640 1600.000 ;
        RECT 657.440 1587.130 657.700 1587.450 ;
        RECT 662.040 1587.130 662.300 1587.450 ;
        RECT 662.100 18.350 662.240 1587.130 ;
        RECT 662.040 18.030 662.300 18.350 ;
        RECT 948.160 18.030 948.420 18.350 ;
        RECT 948.220 2.400 948.360 18.030 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 936.245 18.275 936.415 20.315 ;
        RECT 931.645 18.105 936.415 18.275 ;
        RECT 709.465 17.085 709.635 17.935 ;
        RECT 931.645 17.765 931.815 18.105 ;
      LAYER mcon ;
        RECT 936.245 20.145 936.415 20.315 ;
        RECT 709.465 17.765 709.635 17.935 ;
      LAYER met1 ;
        RECT 664.310 1587.360 664.630 1587.420 ;
        RECT 668.910 1587.360 669.230 1587.420 ;
        RECT 664.310 1587.220 669.230 1587.360 ;
        RECT 664.310 1587.160 664.630 1587.220 ;
        RECT 668.910 1587.160 669.230 1587.220 ;
        RECT 936.185 20.300 936.475 20.345 ;
        RECT 966.070 20.300 966.390 20.360 ;
        RECT 936.185 20.160 966.390 20.300 ;
        RECT 936.185 20.115 936.475 20.160 ;
        RECT 966.070 20.100 966.390 20.160 ;
        RECT 709.405 17.920 709.695 17.965 ;
        RECT 931.585 17.920 931.875 17.965 ;
        RECT 709.405 17.780 931.875 17.920 ;
        RECT 709.405 17.735 709.695 17.780 ;
        RECT 931.585 17.735 931.875 17.780 ;
        RECT 668.450 17.240 668.770 17.300 ;
        RECT 709.405 17.240 709.695 17.285 ;
        RECT 668.450 17.100 709.695 17.240 ;
        RECT 668.450 17.040 668.770 17.100 ;
        RECT 709.405 17.055 709.695 17.100 ;
      LAYER via ;
        RECT 664.340 1587.160 664.600 1587.420 ;
        RECT 668.940 1587.160 669.200 1587.420 ;
        RECT 966.100 20.100 966.360 20.360 ;
        RECT 668.480 17.040 668.740 17.300 ;
      LAYER met2 ;
        RECT 664.340 1600.000 664.620 1604.000 ;
        RECT 664.400 1587.450 664.540 1600.000 ;
        RECT 664.340 1587.130 664.600 1587.450 ;
        RECT 668.940 1587.130 669.200 1587.450 ;
        RECT 669.000 31.010 669.140 1587.130 ;
        RECT 668.540 30.870 669.140 31.010 ;
        RECT 668.540 17.330 668.680 30.870 ;
        RECT 966.100 20.070 966.360 20.390 ;
        RECT 668.480 17.010 668.740 17.330 ;
        RECT 966.160 2.400 966.300 20.070 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 946.825 17.765 946.995 19.635 ;
      LAYER mcon ;
        RECT 946.825 19.465 946.995 19.635 ;
      LAYER met1 ;
        RECT 671.210 1592.800 671.530 1592.860 ;
        RECT 845.090 1592.800 845.410 1592.860 ;
        RECT 671.210 1592.660 845.410 1592.800 ;
        RECT 671.210 1592.600 671.530 1592.660 ;
        RECT 845.090 1592.600 845.410 1592.660 ;
        RECT 845.090 19.960 845.410 20.020 ;
        RECT 882.350 19.960 882.670 20.020 ;
        RECT 845.090 19.820 882.670 19.960 ;
        RECT 845.090 19.760 845.410 19.820 ;
        RECT 882.350 19.760 882.670 19.820 ;
        RECT 884.190 19.620 884.510 19.680 ;
        RECT 946.765 19.620 947.055 19.665 ;
        RECT 884.190 19.480 947.055 19.620 ;
        RECT 884.190 19.420 884.510 19.480 ;
        RECT 946.765 19.435 947.055 19.480 ;
        RECT 946.765 17.920 947.055 17.965 ;
        RECT 984.010 17.920 984.330 17.980 ;
        RECT 946.765 17.780 984.330 17.920 ;
        RECT 946.765 17.735 947.055 17.780 ;
        RECT 984.010 17.720 984.330 17.780 ;
      LAYER via ;
        RECT 671.240 1592.600 671.500 1592.860 ;
        RECT 845.120 1592.600 845.380 1592.860 ;
        RECT 845.120 19.760 845.380 20.020 ;
        RECT 882.380 19.760 882.640 20.020 ;
        RECT 884.220 19.420 884.480 19.680 ;
        RECT 984.040 17.720 984.300 17.980 ;
      LAYER met2 ;
        RECT 671.240 1600.000 671.520 1604.000 ;
        RECT 671.300 1592.890 671.440 1600.000 ;
        RECT 671.240 1592.570 671.500 1592.890 ;
        RECT 845.120 1592.570 845.380 1592.890 ;
        RECT 845.180 20.050 845.320 1592.570 ;
        RECT 882.370 20.555 882.650 20.925 ;
        RECT 884.210 20.555 884.490 20.925 ;
        RECT 882.440 20.050 882.580 20.555 ;
        RECT 845.120 19.730 845.380 20.050 ;
        RECT 882.380 19.730 882.640 20.050 ;
        RECT 884.280 19.710 884.420 20.555 ;
        RECT 884.220 19.390 884.480 19.710 ;
        RECT 984.040 17.690 984.300 18.010 ;
        RECT 984.100 2.400 984.240 17.690 ;
        RECT 983.890 -4.800 984.450 2.400 ;
      LAYER via2 ;
        RECT 882.370 20.600 882.650 20.880 ;
        RECT 884.210 20.600 884.490 20.880 ;
      LAYER met3 ;
        RECT 882.345 20.890 882.675 20.905 ;
        RECT 884.185 20.890 884.515 20.905 ;
        RECT 882.345 20.590 884.515 20.890 ;
        RECT 882.345 20.575 882.675 20.590 ;
        RECT 884.185 20.575 884.515 20.590 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.150 17.920 551.470 17.980 ;
        RECT 662.930 17.920 663.250 17.980 ;
        RECT 551.150 17.780 663.250 17.920 ;
        RECT 551.150 17.720 551.470 17.780 ;
        RECT 662.930 17.720 663.250 17.780 ;
      LAYER via ;
        RECT 551.180 17.720 551.440 17.980 ;
        RECT 662.960 17.720 663.220 17.980 ;
      LAYER met2 ;
        RECT 549.800 1600.450 550.080 1604.000 ;
        RECT 549.800 1600.310 551.380 1600.450 ;
        RECT 549.800 1600.000 550.080 1600.310 ;
        RECT 551.240 18.010 551.380 1600.310 ;
        RECT 551.180 17.690 551.440 18.010 ;
        RECT 662.960 17.690 663.220 18.010 ;
        RECT 663.020 2.400 663.160 17.690 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 689.225 1586.865 689.395 1587.715 ;
        RECT 690.605 1587.545 690.775 1589.415 ;
        RECT 760.985 1589.245 761.155 1590.095 ;
        RECT 954.645 18.615 954.815 19.295 ;
        RECT 954.645 18.445 955.735 18.615 ;
      LAYER mcon ;
        RECT 760.985 1589.925 761.155 1590.095 ;
        RECT 690.605 1589.245 690.775 1589.415 ;
        RECT 689.225 1587.545 689.395 1587.715 ;
        RECT 954.645 19.125 954.815 19.295 ;
        RECT 955.565 18.445 955.735 18.615 ;
      LAYER met1 ;
        RECT 760.925 1590.080 761.215 1590.125 ;
        RECT 831.290 1590.080 831.610 1590.140 ;
        RECT 760.925 1589.940 831.610 1590.080 ;
        RECT 760.925 1589.895 761.215 1589.940 ;
        RECT 831.290 1589.880 831.610 1589.940 ;
        RECT 690.545 1589.400 690.835 1589.445 ;
        RECT 760.925 1589.400 761.215 1589.445 ;
        RECT 690.545 1589.260 761.215 1589.400 ;
        RECT 690.545 1589.215 690.835 1589.260 ;
        RECT 760.925 1589.215 761.215 1589.260 ;
        RECT 689.165 1587.700 689.455 1587.745 ;
        RECT 690.545 1587.700 690.835 1587.745 ;
        RECT 689.165 1587.560 690.835 1587.700 ;
        RECT 689.165 1587.515 689.455 1587.560 ;
        RECT 690.545 1587.515 690.835 1587.560 ;
        RECT 679.490 1587.020 679.810 1587.080 ;
        RECT 689.165 1587.020 689.455 1587.065 ;
        RECT 679.490 1586.880 689.455 1587.020 ;
        RECT 679.490 1586.820 679.810 1586.880 ;
        RECT 689.165 1586.835 689.455 1586.880 ;
        RECT 831.290 19.280 831.610 19.340 ;
        RECT 882.810 19.280 883.130 19.340 ;
        RECT 831.290 19.140 883.130 19.280 ;
        RECT 831.290 19.080 831.610 19.140 ;
        RECT 882.810 19.080 883.130 19.140 ;
        RECT 883.730 19.280 884.050 19.340 ;
        RECT 954.585 19.280 954.875 19.325 ;
        RECT 883.730 19.140 954.875 19.280 ;
        RECT 883.730 19.080 884.050 19.140 ;
        RECT 954.585 19.095 954.875 19.140 ;
        RECT 955.505 18.600 955.795 18.645 ;
        RECT 1001.950 18.600 1002.270 18.660 ;
        RECT 955.505 18.460 1002.270 18.600 ;
        RECT 955.505 18.415 955.795 18.460 ;
        RECT 1001.950 18.400 1002.270 18.460 ;
      LAYER via ;
        RECT 831.320 1589.880 831.580 1590.140 ;
        RECT 679.520 1586.820 679.780 1587.080 ;
        RECT 831.320 19.080 831.580 19.340 ;
        RECT 882.840 19.080 883.100 19.340 ;
        RECT 883.760 19.080 884.020 19.340 ;
        RECT 1001.980 18.400 1002.240 18.660 ;
      LAYER met2 ;
        RECT 677.680 1600.450 677.960 1604.000 ;
        RECT 677.680 1600.310 679.720 1600.450 ;
        RECT 677.680 1600.000 677.960 1600.310 ;
        RECT 679.580 1587.110 679.720 1600.310 ;
        RECT 831.320 1589.850 831.580 1590.170 ;
        RECT 679.520 1586.790 679.780 1587.110 ;
        RECT 831.380 19.370 831.520 1589.850 ;
        RECT 882.830 21.235 883.110 21.605 ;
        RECT 883.750 21.235 884.030 21.605 ;
        RECT 882.900 19.370 883.040 21.235 ;
        RECT 883.820 19.370 883.960 21.235 ;
        RECT 831.320 19.050 831.580 19.370 ;
        RECT 882.840 19.050 883.100 19.370 ;
        RECT 883.760 19.050 884.020 19.370 ;
        RECT 1001.980 18.370 1002.240 18.690 ;
        RECT 1002.040 2.400 1002.180 18.370 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
      LAYER via2 ;
        RECT 882.830 21.280 883.110 21.560 ;
        RECT 883.750 21.280 884.030 21.560 ;
      LAYER met3 ;
        RECT 882.805 21.570 883.135 21.585 ;
        RECT 883.725 21.570 884.055 21.585 ;
        RECT 882.805 21.270 884.055 21.570 ;
        RECT 882.805 21.255 883.135 21.270 ;
        RECT 883.725 21.255 884.055 21.270 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 683.170 1535.340 683.490 1535.400 ;
        RECT 689.610 1535.340 689.930 1535.400 ;
        RECT 683.170 1535.200 689.930 1535.340 ;
        RECT 683.170 1535.140 683.490 1535.200 ;
        RECT 689.610 1535.140 689.930 1535.200 ;
        RECT 689.610 17.580 689.930 17.640 ;
        RECT 1019.430 17.580 1019.750 17.640 ;
        RECT 689.610 17.440 1019.750 17.580 ;
        RECT 689.610 17.380 689.930 17.440 ;
        RECT 1019.430 17.380 1019.750 17.440 ;
      LAYER via ;
        RECT 683.200 1535.140 683.460 1535.400 ;
        RECT 689.640 1535.140 689.900 1535.400 ;
        RECT 689.640 17.380 689.900 17.640 ;
        RECT 1019.460 17.380 1019.720 17.640 ;
      LAYER met2 ;
        RECT 684.580 1600.450 684.860 1604.000 ;
        RECT 683.260 1600.310 684.860 1600.450 ;
        RECT 683.260 1535.430 683.400 1600.310 ;
        RECT 684.580 1600.000 684.860 1600.310 ;
        RECT 683.200 1535.110 683.460 1535.430 ;
        RECT 689.640 1535.110 689.900 1535.430 ;
        RECT 689.700 17.670 689.840 1535.110 ;
        RECT 689.640 17.350 689.900 17.670 ;
        RECT 1019.460 17.350 1019.720 17.670 ;
        RECT 1019.520 2.400 1019.660 17.350 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 709.925 14.365 710.095 17.255 ;
      LAYER mcon ;
        RECT 709.925 17.085 710.095 17.255 ;
      LAYER met1 ;
        RECT 691.450 1587.700 691.770 1587.760 ;
        RECT 696.510 1587.700 696.830 1587.760 ;
        RECT 691.450 1587.560 696.830 1587.700 ;
        RECT 691.450 1587.500 691.770 1587.560 ;
        RECT 696.510 1587.500 696.830 1587.560 ;
        RECT 709.865 17.240 710.155 17.285 ;
        RECT 1037.370 17.240 1037.690 17.300 ;
        RECT 709.865 17.100 1037.690 17.240 ;
        RECT 709.865 17.055 710.155 17.100 ;
        RECT 1037.370 17.040 1037.690 17.100 ;
        RECT 696.510 14.520 696.830 14.580 ;
        RECT 709.865 14.520 710.155 14.565 ;
        RECT 696.510 14.380 710.155 14.520 ;
        RECT 696.510 14.320 696.830 14.380 ;
        RECT 709.865 14.335 710.155 14.380 ;
      LAYER via ;
        RECT 691.480 1587.500 691.740 1587.760 ;
        RECT 696.540 1587.500 696.800 1587.760 ;
        RECT 1037.400 17.040 1037.660 17.300 ;
        RECT 696.540 14.320 696.800 14.580 ;
      LAYER met2 ;
        RECT 691.480 1600.000 691.760 1604.000 ;
        RECT 691.540 1587.790 691.680 1600.000 ;
        RECT 691.480 1587.470 691.740 1587.790 ;
        RECT 696.540 1587.470 696.800 1587.790 ;
        RECT 696.600 14.610 696.740 1587.470 ;
        RECT 1037.400 17.010 1037.660 17.330 ;
        RECT 696.540 14.290 696.800 14.610 ;
        RECT 1037.460 2.400 1037.600 17.010 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 696.970 1535.340 697.290 1535.400 ;
        RECT 703.410 1535.340 703.730 1535.400 ;
        RECT 696.970 1535.200 703.730 1535.340 ;
        RECT 696.970 1535.140 697.290 1535.200 ;
        RECT 703.410 1535.140 703.730 1535.200 ;
      LAYER via ;
        RECT 697.000 1535.140 697.260 1535.400 ;
        RECT 703.440 1535.140 703.700 1535.400 ;
      LAYER met2 ;
        RECT 697.920 1600.450 698.200 1604.000 ;
        RECT 697.060 1600.310 698.200 1600.450 ;
        RECT 697.060 1535.430 697.200 1600.310 ;
        RECT 697.920 1600.000 698.200 1600.310 ;
        RECT 697.000 1535.110 697.260 1535.430 ;
        RECT 703.440 1535.110 703.700 1535.430 ;
        RECT 703.500 20.245 703.640 1535.110 ;
        RECT 703.430 19.875 703.710 20.245 ;
        RECT 1055.330 19.875 1055.610 20.245 ;
        RECT 1055.400 2.400 1055.540 19.875 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
      LAYER via2 ;
        RECT 703.430 19.920 703.710 20.200 ;
        RECT 1055.330 19.920 1055.610 20.200 ;
      LAYER met3 ;
        RECT 703.405 20.210 703.735 20.225 ;
        RECT 1055.305 20.210 1055.635 20.225 ;
        RECT 703.405 19.910 1055.635 20.210 ;
        RECT 703.405 19.895 703.735 19.910 ;
        RECT 1055.305 19.895 1055.635 19.910 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 704.330 1535.340 704.650 1535.400 ;
        RECT 710.310 1535.340 710.630 1535.400 ;
        RECT 704.330 1535.200 710.630 1535.340 ;
        RECT 704.330 1535.140 704.650 1535.200 ;
        RECT 710.310 1535.140 710.630 1535.200 ;
      LAYER via ;
        RECT 704.360 1535.140 704.620 1535.400 ;
        RECT 710.340 1535.140 710.600 1535.400 ;
      LAYER met2 ;
        RECT 704.820 1600.450 705.100 1604.000 ;
        RECT 704.420 1600.310 705.100 1600.450 ;
        RECT 704.420 1535.430 704.560 1600.310 ;
        RECT 704.820 1600.000 705.100 1600.310 ;
        RECT 704.360 1535.110 704.620 1535.430 ;
        RECT 710.340 1535.110 710.600 1535.430 ;
        RECT 710.400 19.565 710.540 1535.110 ;
        RECT 710.330 19.195 710.610 19.565 ;
        RECT 1073.270 19.195 1073.550 19.565 ;
        RECT 1073.340 2.400 1073.480 19.195 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
      LAYER via2 ;
        RECT 710.330 19.240 710.610 19.520 ;
        RECT 1073.270 19.240 1073.550 19.520 ;
      LAYER met3 ;
        RECT 710.305 19.530 710.635 19.545 ;
        RECT 1073.245 19.530 1073.575 19.545 ;
        RECT 710.305 19.230 1073.575 19.530 ;
        RECT 710.305 19.215 710.635 19.230 ;
        RECT 1073.245 19.215 1073.575 19.230 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 711.230 1587.700 711.550 1587.760 ;
        RECT 717.210 1587.700 717.530 1587.760 ;
        RECT 711.230 1587.560 717.530 1587.700 ;
        RECT 711.230 1587.500 711.550 1587.560 ;
        RECT 717.210 1587.500 717.530 1587.560 ;
      LAYER via ;
        RECT 711.260 1587.500 711.520 1587.760 ;
        RECT 717.240 1587.500 717.500 1587.760 ;
      LAYER met2 ;
        RECT 711.260 1600.000 711.540 1604.000 ;
        RECT 711.320 1587.790 711.460 1600.000 ;
        RECT 711.260 1587.470 711.520 1587.790 ;
        RECT 717.240 1587.470 717.500 1587.790 ;
        RECT 717.300 18.885 717.440 1587.470 ;
        RECT 717.230 18.515 717.510 18.885 ;
        RECT 1090.750 18.515 1091.030 18.885 ;
        RECT 1090.820 2.400 1090.960 18.515 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
      LAYER via2 ;
        RECT 717.230 18.560 717.510 18.840 ;
        RECT 1090.750 18.560 1091.030 18.840 ;
      LAYER met3 ;
        RECT 717.205 18.850 717.535 18.865 ;
        RECT 1090.725 18.850 1091.055 18.865 ;
        RECT 717.205 18.550 1091.055 18.850 ;
        RECT 717.205 18.535 717.535 18.550 ;
        RECT 1090.725 18.535 1091.055 18.550 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 718.130 1535.340 718.450 1535.400 ;
        RECT 724.110 1535.340 724.430 1535.400 ;
        RECT 718.130 1535.200 724.430 1535.340 ;
        RECT 718.130 1535.140 718.450 1535.200 ;
        RECT 724.110 1535.140 724.430 1535.200 ;
      LAYER via ;
        RECT 718.160 1535.140 718.420 1535.400 ;
        RECT 724.140 1535.140 724.400 1535.400 ;
      LAYER met2 ;
        RECT 718.160 1600.000 718.440 1604.000 ;
        RECT 718.220 1535.430 718.360 1600.000 ;
        RECT 718.160 1535.110 718.420 1535.430 ;
        RECT 724.140 1535.110 724.400 1535.430 ;
        RECT 724.200 16.845 724.340 1535.110 ;
        RECT 724.130 16.475 724.410 16.845 ;
        RECT 1108.690 16.475 1108.970 16.845 ;
        RECT 1108.760 2.400 1108.900 16.475 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
      LAYER via2 ;
        RECT 724.130 16.520 724.410 16.800 ;
        RECT 1108.690 16.520 1108.970 16.800 ;
      LAYER met3 ;
        RECT 724.105 16.810 724.435 16.825 ;
        RECT 1108.665 16.810 1108.995 16.825 ;
        RECT 724.105 16.510 1108.995 16.810 ;
        RECT 724.105 16.495 724.435 16.510 ;
        RECT 1108.665 16.495 1108.995 16.510 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 761.905 1589.585 762.075 1593.155 ;
        RECT 810.665 1588.225 810.835 1589.755 ;
      LAYER mcon ;
        RECT 761.905 1592.985 762.075 1593.155 ;
        RECT 810.665 1589.585 810.835 1589.755 ;
      LAYER met1 ;
        RECT 725.030 1593.140 725.350 1593.200 ;
        RECT 761.845 1593.140 762.135 1593.185 ;
        RECT 725.030 1593.000 762.135 1593.140 ;
        RECT 725.030 1592.940 725.350 1593.000 ;
        RECT 761.845 1592.955 762.135 1593.000 ;
        RECT 761.845 1589.740 762.135 1589.785 ;
        RECT 810.605 1589.740 810.895 1589.785 ;
        RECT 761.845 1589.600 810.895 1589.740 ;
        RECT 761.845 1589.555 762.135 1589.600 ;
        RECT 810.605 1589.555 810.895 1589.600 ;
        RECT 810.605 1588.380 810.895 1588.425 ;
        RECT 858.890 1588.380 859.210 1588.440 ;
        RECT 810.605 1588.240 859.210 1588.380 ;
        RECT 810.605 1588.195 810.895 1588.240 ;
        RECT 858.890 1588.180 859.210 1588.240 ;
        RECT 883.730 14.860 884.050 14.920 ;
        RECT 1126.610 14.860 1126.930 14.920 ;
        RECT 883.730 14.720 1126.930 14.860 ;
        RECT 883.730 14.660 884.050 14.720 ;
        RECT 1126.610 14.660 1126.930 14.720 ;
      LAYER via ;
        RECT 725.060 1592.940 725.320 1593.200 ;
        RECT 858.920 1588.180 859.180 1588.440 ;
        RECT 883.760 14.660 884.020 14.920 ;
        RECT 1126.640 14.660 1126.900 14.920 ;
      LAYER met2 ;
        RECT 725.060 1600.000 725.340 1604.000 ;
        RECT 725.120 1593.230 725.260 1600.000 ;
        RECT 725.060 1592.910 725.320 1593.230 ;
        RECT 858.920 1588.150 859.180 1588.470 ;
        RECT 858.980 15.485 859.120 1588.150 ;
        RECT 858.910 15.115 859.190 15.485 ;
        RECT 883.750 15.115 884.030 15.485 ;
        RECT 883.820 14.950 883.960 15.115 ;
        RECT 883.760 14.630 884.020 14.950 ;
        RECT 1126.640 14.630 1126.900 14.950 ;
        RECT 1126.700 2.400 1126.840 14.630 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
      LAYER via2 ;
        RECT 858.910 15.160 859.190 15.440 ;
        RECT 883.750 15.160 884.030 15.440 ;
      LAYER met3 ;
        RECT 858.885 15.450 859.215 15.465 ;
        RECT 883.725 15.450 884.055 15.465 ;
        RECT 858.885 15.150 884.055 15.450 ;
        RECT 858.885 15.135 859.215 15.150 ;
        RECT 883.725 15.135 884.055 15.150 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 731.470 1587.360 731.790 1587.420 ;
        RECT 737.450 1587.360 737.770 1587.420 ;
        RECT 731.470 1587.220 737.770 1587.360 ;
        RECT 731.470 1587.160 731.790 1587.220 ;
        RECT 737.450 1587.160 737.770 1587.220 ;
        RECT 737.450 39.000 737.770 39.060 ;
        RECT 1144.550 39.000 1144.870 39.060 ;
        RECT 737.450 38.860 1144.870 39.000 ;
        RECT 737.450 38.800 737.770 38.860 ;
        RECT 1144.550 38.800 1144.870 38.860 ;
      LAYER via ;
        RECT 731.500 1587.160 731.760 1587.420 ;
        RECT 737.480 1587.160 737.740 1587.420 ;
        RECT 737.480 38.800 737.740 39.060 ;
        RECT 1144.580 38.800 1144.840 39.060 ;
      LAYER met2 ;
        RECT 731.500 1600.000 731.780 1604.000 ;
        RECT 731.560 1587.450 731.700 1600.000 ;
        RECT 731.500 1587.130 731.760 1587.450 ;
        RECT 737.480 1587.130 737.740 1587.450 ;
        RECT 737.540 39.090 737.680 1587.130 ;
        RECT 737.480 38.770 737.740 39.090 ;
        RECT 1144.580 38.770 1144.840 39.090 ;
        RECT 1144.640 2.400 1144.780 38.770 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 738.370 1589.740 738.690 1589.800 ;
        RECT 744.350 1589.740 744.670 1589.800 ;
        RECT 738.370 1589.600 744.670 1589.740 ;
        RECT 738.370 1589.540 738.690 1589.600 ;
        RECT 744.350 1589.540 744.670 1589.600 ;
        RECT 744.350 38.320 744.670 38.380 ;
        RECT 1162.490 38.320 1162.810 38.380 ;
        RECT 744.350 38.180 1162.810 38.320 ;
        RECT 744.350 38.120 744.670 38.180 ;
        RECT 1162.490 38.120 1162.810 38.180 ;
      LAYER via ;
        RECT 738.400 1589.540 738.660 1589.800 ;
        RECT 744.380 1589.540 744.640 1589.800 ;
        RECT 744.380 38.120 744.640 38.380 ;
        RECT 1162.520 38.120 1162.780 38.380 ;
      LAYER met2 ;
        RECT 738.400 1600.000 738.680 1604.000 ;
        RECT 738.460 1589.830 738.600 1600.000 ;
        RECT 738.400 1589.510 738.660 1589.830 ;
        RECT 744.380 1589.510 744.640 1589.830 ;
        RECT 744.440 38.410 744.580 1589.510 ;
        RECT 744.380 38.090 744.640 38.410 ;
        RECT 1162.520 38.090 1162.780 38.410 ;
        RECT 1162.580 2.400 1162.720 38.090 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 558.510 17.580 558.830 17.640 ;
        RECT 680.410 17.580 680.730 17.640 ;
        RECT 558.510 17.440 680.730 17.580 ;
        RECT 558.510 17.380 558.830 17.440 ;
        RECT 680.410 17.380 680.730 17.440 ;
      LAYER via ;
        RECT 558.540 17.380 558.800 17.640 ;
        RECT 680.440 17.380 680.700 17.640 ;
      LAYER met2 ;
        RECT 556.700 1600.450 556.980 1604.000 ;
        RECT 556.700 1600.310 558.740 1600.450 ;
        RECT 556.700 1600.000 556.980 1600.310 ;
        RECT 558.600 17.670 558.740 1600.310 ;
        RECT 558.540 17.350 558.800 17.670 ;
        RECT 680.440 17.350 680.700 17.670 ;
        RECT 680.500 2.400 680.640 17.350 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 756.845 1587.545 757.015 1589.075 ;
        RECT 776.625 1587.545 776.795 1589.075 ;
      LAYER mcon ;
        RECT 756.845 1588.905 757.015 1589.075 ;
        RECT 776.625 1588.905 776.795 1589.075 ;
      LAYER met1 ;
        RECT 745.270 1589.060 745.590 1589.120 ;
        RECT 756.785 1589.060 757.075 1589.105 ;
        RECT 745.270 1588.920 757.075 1589.060 ;
        RECT 745.270 1588.860 745.590 1588.920 ;
        RECT 756.785 1588.875 757.075 1588.920 ;
        RECT 776.565 1589.060 776.855 1589.105 ;
        RECT 865.790 1589.060 866.110 1589.120 ;
        RECT 776.565 1588.920 866.110 1589.060 ;
        RECT 776.565 1588.875 776.855 1588.920 ;
        RECT 865.790 1588.860 866.110 1588.920 ;
        RECT 756.785 1587.700 757.075 1587.745 ;
        RECT 776.565 1587.700 776.855 1587.745 ;
        RECT 756.785 1587.560 776.855 1587.700 ;
        RECT 756.785 1587.515 757.075 1587.560 ;
        RECT 776.565 1587.515 776.855 1587.560 ;
        RECT 1179.970 15.540 1180.290 15.600 ;
        RECT 883.820 15.400 1180.290 15.540 ;
        RECT 883.820 15.200 883.960 15.400 ;
        RECT 1179.970 15.340 1180.290 15.400 ;
        RECT 883.360 15.060 883.960 15.200 ;
        RECT 865.790 14.860 866.110 14.920 ;
        RECT 883.360 14.860 883.500 15.060 ;
        RECT 865.790 14.720 883.500 14.860 ;
        RECT 865.790 14.660 866.110 14.720 ;
      LAYER via ;
        RECT 745.300 1588.860 745.560 1589.120 ;
        RECT 865.820 1588.860 866.080 1589.120 ;
        RECT 1180.000 15.340 1180.260 15.600 ;
        RECT 865.820 14.660 866.080 14.920 ;
      LAYER met2 ;
        RECT 745.300 1600.000 745.580 1604.000 ;
        RECT 745.360 1589.150 745.500 1600.000 ;
        RECT 745.300 1588.830 745.560 1589.150 ;
        RECT 865.820 1588.830 866.080 1589.150 ;
        RECT 865.880 14.950 866.020 1588.830 ;
        RECT 1180.000 15.310 1180.260 15.630 ;
        RECT 865.820 14.630 866.080 14.950 ;
        RECT 1180.060 2.400 1180.200 15.310 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 907.725 15.045 907.895 30.515 ;
      LAYER mcon ;
        RECT 907.725 30.345 907.895 30.515 ;
      LAYER met1 ;
        RECT 751.710 1593.820 752.030 1593.880 ;
        RECT 879.130 1593.820 879.450 1593.880 ;
        RECT 751.710 1593.680 879.450 1593.820 ;
        RECT 751.710 1593.620 752.030 1593.680 ;
        RECT 879.130 1593.620 879.450 1593.680 ;
        RECT 879.590 30.500 879.910 30.560 ;
        RECT 907.665 30.500 907.955 30.545 ;
        RECT 879.590 30.360 907.955 30.500 ;
        RECT 879.590 30.300 879.910 30.360 ;
        RECT 907.665 30.315 907.955 30.360 ;
        RECT 907.665 15.200 907.955 15.245 ;
        RECT 1197.910 15.200 1198.230 15.260 ;
        RECT 907.665 15.060 1198.230 15.200 ;
        RECT 907.665 15.015 907.955 15.060 ;
        RECT 1197.910 15.000 1198.230 15.060 ;
      LAYER via ;
        RECT 751.740 1593.620 752.000 1593.880 ;
        RECT 879.160 1593.620 879.420 1593.880 ;
        RECT 879.620 30.300 879.880 30.560 ;
        RECT 1197.940 15.000 1198.200 15.260 ;
      LAYER met2 ;
        RECT 751.740 1600.000 752.020 1604.000 ;
        RECT 751.800 1593.910 751.940 1600.000 ;
        RECT 751.740 1593.590 752.000 1593.910 ;
        RECT 879.160 1593.590 879.420 1593.910 ;
        RECT 879.220 1590.930 879.360 1593.590 ;
        RECT 879.220 1590.790 879.820 1590.930 ;
        RECT 879.680 30.590 879.820 1590.790 ;
        RECT 879.620 30.270 879.880 30.590 ;
        RECT 1197.940 14.970 1198.200 15.290 ;
        RECT 1198.000 2.400 1198.140 14.970 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 758.150 44.440 758.470 44.500 ;
        RECT 1215.850 44.440 1216.170 44.500 ;
        RECT 758.150 44.300 1216.170 44.440 ;
        RECT 758.150 44.240 758.470 44.300 ;
        RECT 1215.850 44.240 1216.170 44.300 ;
      LAYER via ;
        RECT 758.180 44.240 758.440 44.500 ;
        RECT 1215.880 44.240 1216.140 44.500 ;
      LAYER met2 ;
        RECT 758.640 1600.450 758.920 1604.000 ;
        RECT 758.240 1600.310 758.920 1600.450 ;
        RECT 758.240 44.530 758.380 1600.310 ;
        RECT 758.640 1600.000 758.920 1600.310 ;
        RECT 758.180 44.210 758.440 44.530 ;
        RECT 1215.880 44.210 1216.140 44.530 ;
        RECT 1215.940 2.400 1216.080 44.210 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 907.265 15.725 907.435 18.955 ;
      LAYER mcon ;
        RECT 907.265 18.785 907.435 18.955 ;
      LAYER met1 ;
        RECT 765.510 1589.400 765.830 1589.460 ;
        RECT 880.050 1589.400 880.370 1589.460 ;
        RECT 765.510 1589.260 880.370 1589.400 ;
        RECT 765.510 1589.200 765.830 1589.260 ;
        RECT 880.050 1589.200 880.370 1589.260 ;
        RECT 907.205 18.940 907.495 18.985 ;
        RECT 883.820 18.800 907.495 18.940 ;
        RECT 880.050 18.600 880.370 18.660 ;
        RECT 883.820 18.600 883.960 18.800 ;
        RECT 907.205 18.755 907.495 18.800 ;
        RECT 880.050 18.460 883.960 18.600 ;
        RECT 880.050 18.400 880.370 18.460 ;
        RECT 907.205 15.880 907.495 15.925 ;
        RECT 1233.790 15.880 1234.110 15.940 ;
        RECT 907.205 15.740 1234.110 15.880 ;
        RECT 907.205 15.695 907.495 15.740 ;
        RECT 1233.790 15.680 1234.110 15.740 ;
      LAYER via ;
        RECT 765.540 1589.200 765.800 1589.460 ;
        RECT 880.080 1589.200 880.340 1589.460 ;
        RECT 880.080 18.400 880.340 18.660 ;
        RECT 1233.820 15.680 1234.080 15.940 ;
      LAYER met2 ;
        RECT 765.540 1600.000 765.820 1604.000 ;
        RECT 765.600 1589.490 765.740 1600.000 ;
        RECT 765.540 1589.170 765.800 1589.490 ;
        RECT 880.080 1589.170 880.340 1589.490 ;
        RECT 880.140 18.690 880.280 1589.170 ;
        RECT 880.080 18.370 880.340 18.690 ;
        RECT 1233.820 15.650 1234.080 15.970 ;
        RECT 1233.880 2.400 1234.020 15.650 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 771.950 47.840 772.270 47.900 ;
        RECT 1251.730 47.840 1252.050 47.900 ;
        RECT 771.950 47.700 1252.050 47.840 ;
        RECT 771.950 47.640 772.270 47.700 ;
        RECT 1251.730 47.640 1252.050 47.700 ;
      LAYER via ;
        RECT 771.980 47.640 772.240 47.900 ;
        RECT 1251.760 47.640 1252.020 47.900 ;
      LAYER met2 ;
        RECT 771.980 1600.000 772.260 1604.000 ;
        RECT 772.040 47.930 772.180 1600.000 ;
        RECT 771.980 47.610 772.240 47.930 ;
        RECT 1251.760 47.610 1252.020 47.930 ;
        RECT 1251.820 2.400 1251.960 47.610 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 927.505 16.235 927.675 18.955 ;
        RECT 927.505 16.065 930.895 16.235 ;
      LAYER mcon ;
        RECT 927.505 18.785 927.675 18.955 ;
        RECT 930.725 16.065 930.895 16.235 ;
      LAYER met1 ;
        RECT 778.850 1593.140 779.170 1593.200 ;
        RECT 892.930 1593.140 893.250 1593.200 ;
        RECT 778.850 1593.000 893.250 1593.140 ;
        RECT 778.850 1592.940 779.170 1593.000 ;
        RECT 892.930 1592.940 893.250 1593.000 ;
        RECT 907.650 18.940 907.970 19.000 ;
        RECT 927.445 18.940 927.735 18.985 ;
        RECT 907.650 18.800 927.735 18.940 ;
        RECT 907.650 18.740 907.970 18.800 ;
        RECT 927.445 18.755 927.735 18.800 ;
        RECT 930.665 16.220 930.955 16.265 ;
        RECT 1269.210 16.220 1269.530 16.280 ;
        RECT 930.665 16.080 1269.530 16.220 ;
        RECT 930.665 16.035 930.955 16.080 ;
        RECT 1269.210 16.020 1269.530 16.080 ;
      LAYER via ;
        RECT 778.880 1592.940 779.140 1593.200 ;
        RECT 892.960 1592.940 893.220 1593.200 ;
        RECT 907.680 18.740 907.940 19.000 ;
        RECT 1269.240 16.020 1269.500 16.280 ;
      LAYER met2 ;
        RECT 778.880 1600.000 779.160 1604.000 ;
        RECT 778.940 1593.230 779.080 1600.000 ;
        RECT 778.880 1592.910 779.140 1593.230 ;
        RECT 892.960 1592.910 893.220 1593.230 ;
        RECT 893.020 1590.250 893.160 1592.910 ;
        RECT 893.020 1590.110 893.620 1590.250 ;
        RECT 893.480 20.925 893.620 1590.110 ;
        RECT 893.410 20.555 893.690 20.925 ;
        RECT 907.670 20.555 907.950 20.925 ;
        RECT 907.740 19.030 907.880 20.555 ;
        RECT 907.680 18.710 907.940 19.030 ;
        RECT 1269.240 15.990 1269.500 16.310 ;
        RECT 1269.300 2.400 1269.440 15.990 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
      LAYER via2 ;
        RECT 893.410 20.600 893.690 20.880 ;
        RECT 907.670 20.600 907.950 20.880 ;
      LAYER met3 ;
        RECT 893.385 20.890 893.715 20.905 ;
        RECT 907.645 20.890 907.975 20.905 ;
        RECT 893.385 20.590 907.975 20.890 ;
        RECT 893.385 20.575 893.715 20.590 ;
        RECT 907.645 20.575 907.975 20.590 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 785.750 46.820 786.070 46.880 ;
        RECT 1287.150 46.820 1287.470 46.880 ;
        RECT 785.750 46.680 1287.470 46.820 ;
        RECT 785.750 46.620 786.070 46.680 ;
        RECT 1287.150 46.620 1287.470 46.680 ;
      LAYER via ;
        RECT 785.780 46.620 786.040 46.880 ;
        RECT 1287.180 46.620 1287.440 46.880 ;
      LAYER met2 ;
        RECT 785.320 1600.450 785.600 1604.000 ;
        RECT 785.320 1600.310 785.980 1600.450 ;
        RECT 785.320 1600.000 785.600 1600.310 ;
        RECT 785.840 46.910 785.980 1600.310 ;
        RECT 785.780 46.590 786.040 46.910 ;
        RECT 1287.180 46.590 1287.440 46.910 ;
        RECT 1287.240 2.400 1287.380 46.590 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 792.190 46.480 792.510 46.540 ;
        RECT 1305.090 46.480 1305.410 46.540 ;
        RECT 792.190 46.340 1305.410 46.480 ;
        RECT 792.190 46.280 792.510 46.340 ;
        RECT 1305.090 46.280 1305.410 46.340 ;
      LAYER via ;
        RECT 792.220 46.280 792.480 46.540 ;
        RECT 1305.120 46.280 1305.380 46.540 ;
      LAYER met2 ;
        RECT 792.220 1600.000 792.500 1604.000 ;
        RECT 792.280 46.570 792.420 1600.000 ;
        RECT 792.220 46.250 792.480 46.570 ;
        RECT 1305.120 46.250 1305.380 46.570 ;
        RECT 1305.180 2.400 1305.320 46.250 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 799.090 46.140 799.410 46.200 ;
        RECT 1323.030 46.140 1323.350 46.200 ;
        RECT 799.090 46.000 1323.350 46.140 ;
        RECT 799.090 45.940 799.410 46.000 ;
        RECT 1323.030 45.940 1323.350 46.000 ;
      LAYER via ;
        RECT 799.120 45.940 799.380 46.200 ;
        RECT 1323.060 45.940 1323.320 46.200 ;
      LAYER met2 ;
        RECT 799.120 1600.000 799.400 1604.000 ;
        RECT 799.180 46.230 799.320 1600.000 ;
        RECT 799.120 45.910 799.380 46.230 ;
        RECT 1323.060 45.910 1323.320 46.230 ;
        RECT 1323.120 2.400 1323.260 45.910 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 805.990 45.800 806.310 45.860 ;
        RECT 1340.510 45.800 1340.830 45.860 ;
        RECT 805.990 45.660 1340.830 45.800 ;
        RECT 805.990 45.600 806.310 45.660 ;
        RECT 1340.510 45.600 1340.830 45.660 ;
      LAYER via ;
        RECT 806.020 45.600 806.280 45.860 ;
        RECT 1340.540 45.600 1340.800 45.860 ;
      LAYER met2 ;
        RECT 805.560 1600.450 805.840 1604.000 ;
        RECT 805.560 1600.310 806.220 1600.450 ;
        RECT 805.560 1600.000 805.840 1600.310 ;
        RECT 806.080 45.890 806.220 1600.310 ;
        RECT 806.020 45.570 806.280 45.890 ;
        RECT 1340.540 45.570 1340.800 45.890 ;
        RECT 1340.600 2.400 1340.740 45.570 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 14.860 565.730 14.920 ;
        RECT 698.350 14.860 698.670 14.920 ;
        RECT 565.410 14.720 698.670 14.860 ;
        RECT 565.410 14.660 565.730 14.720 ;
        RECT 698.350 14.660 698.670 14.720 ;
      LAYER via ;
        RECT 565.440 14.660 565.700 14.920 ;
        RECT 698.380 14.660 698.640 14.920 ;
      LAYER met2 ;
        RECT 563.140 1600.450 563.420 1604.000 ;
        RECT 563.140 1600.310 565.180 1600.450 ;
        RECT 563.140 1600.000 563.420 1600.310 ;
        RECT 565.040 1588.210 565.180 1600.310 ;
        RECT 565.040 1588.070 565.640 1588.210 ;
        RECT 565.500 14.950 565.640 1588.070 ;
        RECT 565.440 14.630 565.700 14.950 ;
        RECT 698.380 14.630 698.640 14.950 ;
        RECT 698.440 2.400 698.580 14.630 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 913.245 16.745 913.415 19.975 ;
        RECT 931.185 16.745 931.355 19.975 ;
      LAYER mcon ;
        RECT 913.245 19.805 913.415 19.975 ;
        RECT 931.185 19.805 931.355 19.975 ;
      LAYER met1 ;
        RECT 812.430 1588.720 812.750 1588.780 ;
        RECT 900.290 1588.720 900.610 1588.780 ;
        RECT 812.430 1588.580 900.610 1588.720 ;
        RECT 812.430 1588.520 812.750 1588.580 ;
        RECT 900.290 1588.520 900.610 1588.580 ;
        RECT 913.185 19.960 913.475 20.005 ;
        RECT 931.125 19.960 931.415 20.005 ;
        RECT 913.185 19.820 931.415 19.960 ;
        RECT 913.185 19.775 913.475 19.820 ;
        RECT 931.125 19.775 931.415 19.820 ;
        RECT 900.290 16.900 900.610 16.960 ;
        RECT 913.185 16.900 913.475 16.945 ;
        RECT 900.290 16.760 913.475 16.900 ;
        RECT 900.290 16.700 900.610 16.760 ;
        RECT 913.185 16.715 913.475 16.760 ;
        RECT 931.125 16.900 931.415 16.945 ;
        RECT 1358.450 16.900 1358.770 16.960 ;
        RECT 931.125 16.760 1358.770 16.900 ;
        RECT 931.125 16.715 931.415 16.760 ;
        RECT 1358.450 16.700 1358.770 16.760 ;
      LAYER via ;
        RECT 812.460 1588.520 812.720 1588.780 ;
        RECT 900.320 1588.520 900.580 1588.780 ;
        RECT 900.320 16.700 900.580 16.960 ;
        RECT 1358.480 16.700 1358.740 16.960 ;
      LAYER met2 ;
        RECT 812.460 1600.000 812.740 1604.000 ;
        RECT 812.520 1588.810 812.660 1600.000 ;
        RECT 812.460 1588.490 812.720 1588.810 ;
        RECT 900.320 1588.490 900.580 1588.810 ;
        RECT 900.380 16.990 900.520 1588.490 ;
        RECT 900.320 16.670 900.580 16.990 ;
        RECT 1358.480 16.670 1358.740 16.990 ;
        RECT 1358.540 2.400 1358.680 16.670 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 819.330 1593.480 819.650 1593.540 ;
        RECT 1231.490 1593.480 1231.810 1593.540 ;
        RECT 819.330 1593.340 1231.810 1593.480 ;
        RECT 819.330 1593.280 819.650 1593.340 ;
        RECT 1231.490 1593.280 1231.810 1593.340 ;
        RECT 1231.490 14.520 1231.810 14.580 ;
        RECT 1376.390 14.520 1376.710 14.580 ;
        RECT 1231.490 14.380 1376.710 14.520 ;
        RECT 1231.490 14.320 1231.810 14.380 ;
        RECT 1376.390 14.320 1376.710 14.380 ;
      LAYER via ;
        RECT 819.360 1593.280 819.620 1593.540 ;
        RECT 1231.520 1593.280 1231.780 1593.540 ;
        RECT 1231.520 14.320 1231.780 14.580 ;
        RECT 1376.420 14.320 1376.680 14.580 ;
      LAYER met2 ;
        RECT 819.360 1600.000 819.640 1604.000 ;
        RECT 819.420 1593.570 819.560 1600.000 ;
        RECT 819.360 1593.250 819.620 1593.570 ;
        RECT 1231.520 1593.250 1231.780 1593.570 ;
        RECT 1231.580 14.610 1231.720 1593.250 ;
        RECT 1231.520 14.290 1231.780 14.610 ;
        RECT 1376.420 14.290 1376.680 14.610 ;
        RECT 1376.480 2.400 1376.620 14.290 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 848.845 1590.605 849.015 1591.795 ;
        RECT 1243.065 1588.565 1243.235 1590.775 ;
      LAYER mcon ;
        RECT 848.845 1591.625 849.015 1591.795 ;
        RECT 1243.065 1590.605 1243.235 1590.775 ;
      LAYER met1 ;
        RECT 825.770 1591.780 826.090 1591.840 ;
        RECT 848.785 1591.780 849.075 1591.825 ;
        RECT 825.770 1591.640 849.075 1591.780 ;
        RECT 825.770 1591.580 826.090 1591.640 ;
        RECT 848.785 1591.595 849.075 1591.640 ;
        RECT 848.785 1590.760 849.075 1590.805 ;
        RECT 1243.005 1590.760 1243.295 1590.805 ;
        RECT 848.785 1590.620 1243.295 1590.760 ;
        RECT 848.785 1590.575 849.075 1590.620 ;
        RECT 1243.005 1590.575 1243.295 1590.620 ;
        RECT 1243.005 1588.720 1243.295 1588.765 ;
        RECT 1266.450 1588.720 1266.770 1588.780 ;
        RECT 1243.005 1588.580 1266.770 1588.720 ;
        RECT 1243.005 1588.535 1243.295 1588.580 ;
        RECT 1266.450 1588.520 1266.770 1588.580 ;
        RECT 1266.450 14.860 1266.770 14.920 ;
        RECT 1394.330 14.860 1394.650 14.920 ;
        RECT 1266.450 14.720 1394.650 14.860 ;
        RECT 1266.450 14.660 1266.770 14.720 ;
        RECT 1394.330 14.660 1394.650 14.720 ;
      LAYER via ;
        RECT 825.800 1591.580 826.060 1591.840 ;
        RECT 1266.480 1588.520 1266.740 1588.780 ;
        RECT 1266.480 14.660 1266.740 14.920 ;
        RECT 1394.360 14.660 1394.620 14.920 ;
      LAYER met2 ;
        RECT 825.800 1600.000 826.080 1604.000 ;
        RECT 825.860 1591.870 826.000 1600.000 ;
        RECT 825.800 1591.550 826.060 1591.870 ;
        RECT 1266.480 1588.490 1266.740 1588.810 ;
        RECT 1266.540 14.950 1266.680 1588.490 ;
        RECT 1266.480 14.630 1266.740 14.950 ;
        RECT 1394.360 14.630 1394.620 14.950 ;
        RECT 1394.420 2.400 1394.560 14.630 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 914.090 1588.380 914.410 1588.440 ;
        RECT 859.440 1588.240 914.410 1588.380 ;
        RECT 832.670 1587.700 832.990 1587.760 ;
        RECT 859.440 1587.700 859.580 1588.240 ;
        RECT 914.090 1588.180 914.410 1588.240 ;
        RECT 832.670 1587.560 859.580 1587.700 ;
        RECT 832.670 1587.500 832.990 1587.560 ;
        RECT 914.090 16.900 914.410 16.960 ;
        RECT 930.650 16.900 930.970 16.960 ;
        RECT 914.090 16.760 930.970 16.900 ;
        RECT 914.090 16.700 914.410 16.760 ;
        RECT 930.650 16.700 930.970 16.760 ;
        RECT 932.030 16.560 932.350 16.620 ;
        RECT 1412.270 16.560 1412.590 16.620 ;
        RECT 932.030 16.420 1412.590 16.560 ;
        RECT 932.030 16.360 932.350 16.420 ;
        RECT 1412.270 16.360 1412.590 16.420 ;
      LAYER via ;
        RECT 832.700 1587.500 832.960 1587.760 ;
        RECT 914.120 1588.180 914.380 1588.440 ;
        RECT 914.120 16.700 914.380 16.960 ;
        RECT 930.680 16.700 930.940 16.960 ;
        RECT 932.060 16.360 932.320 16.620 ;
        RECT 1412.300 16.360 1412.560 16.620 ;
      LAYER met2 ;
        RECT 832.700 1600.000 832.980 1604.000 ;
        RECT 832.760 1587.790 832.900 1600.000 ;
        RECT 914.120 1588.150 914.380 1588.470 ;
        RECT 832.700 1587.470 832.960 1587.790 ;
        RECT 914.180 16.990 914.320 1588.150 ;
        RECT 914.120 16.670 914.380 16.990 ;
        RECT 930.680 16.670 930.940 16.990 ;
        RECT 930.740 16.165 930.880 16.670 ;
        RECT 932.060 16.330 932.320 16.650 ;
        RECT 1412.300 16.330 1412.560 16.650 ;
        RECT 932.120 16.165 932.260 16.330 ;
        RECT 930.670 15.795 930.950 16.165 ;
        RECT 932.050 15.795 932.330 16.165 ;
        RECT 1412.360 2.400 1412.500 16.330 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
      LAYER via2 ;
        RECT 930.670 15.840 930.950 16.120 ;
        RECT 932.050 15.840 932.330 16.120 ;
      LAYER met3 ;
        RECT 930.645 16.130 930.975 16.145 ;
        RECT 932.025 16.130 932.355 16.145 ;
        RECT 930.645 15.830 932.355 16.130 ;
        RECT 930.645 15.815 930.975 15.830 ;
        RECT 932.025 15.815 932.355 15.830 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1341.965 1589.245 1342.135 1590.435 ;
      LAYER mcon ;
        RECT 1341.965 1590.265 1342.135 1590.435 ;
      LAYER met1 ;
        RECT 843.340 1590.620 848.540 1590.760 ;
        RECT 839.570 1590.080 839.890 1590.140 ;
        RECT 843.340 1590.080 843.480 1590.620 ;
        RECT 848.400 1590.420 848.540 1590.620 ;
        RECT 1341.905 1590.420 1342.195 1590.465 ;
        RECT 848.400 1590.280 1342.195 1590.420 ;
        RECT 1341.905 1590.235 1342.195 1590.280 ;
        RECT 839.570 1589.940 843.480 1590.080 ;
        RECT 839.570 1589.880 839.890 1589.940 ;
        RECT 1341.905 1589.400 1342.195 1589.445 ;
        RECT 1355.690 1589.400 1356.010 1589.460 ;
        RECT 1341.905 1589.260 1356.010 1589.400 ;
        RECT 1341.905 1589.215 1342.195 1589.260 ;
        RECT 1355.690 1589.200 1356.010 1589.260 ;
        RECT 1429.750 14.520 1430.070 14.580 ;
        RECT 1387.520 14.380 1430.070 14.520 ;
        RECT 1355.690 14.180 1356.010 14.240 ;
        RECT 1387.520 14.180 1387.660 14.380 ;
        RECT 1429.750 14.320 1430.070 14.380 ;
        RECT 1355.690 14.040 1387.660 14.180 ;
        RECT 1355.690 13.980 1356.010 14.040 ;
      LAYER via ;
        RECT 839.600 1589.880 839.860 1590.140 ;
        RECT 1355.720 1589.200 1355.980 1589.460 ;
        RECT 1355.720 13.980 1355.980 14.240 ;
        RECT 1429.780 14.320 1430.040 14.580 ;
      LAYER met2 ;
        RECT 839.600 1600.000 839.880 1604.000 ;
        RECT 839.660 1590.170 839.800 1600.000 ;
        RECT 839.600 1589.850 839.860 1590.170 ;
        RECT 1355.720 1589.170 1355.980 1589.490 ;
        RECT 1355.780 14.270 1355.920 1589.170 ;
        RECT 1429.780 14.290 1430.040 14.610 ;
        RECT 1355.720 13.950 1355.980 14.270 ;
        RECT 1429.840 2.400 1429.980 14.290 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 954.185 19.805 954.815 19.975 ;
        RECT 965.685 19.805 967.235 19.975 ;
        RECT 954.185 18.445 954.355 19.805 ;
      LAYER mcon ;
        RECT 954.645 19.805 954.815 19.975 ;
        RECT 967.065 19.805 967.235 19.975 ;
      LAYER met1 ;
        RECT 846.010 1590.080 846.330 1590.140 ;
        RECT 846.010 1589.940 904.660 1590.080 ;
        RECT 846.010 1589.880 846.330 1589.940 ;
        RECT 904.520 1589.740 904.660 1589.940 ;
        RECT 920.990 1589.740 921.310 1589.800 ;
        RECT 904.520 1589.600 921.310 1589.740 ;
        RECT 920.990 1589.540 921.310 1589.600 ;
        RECT 954.585 19.960 954.875 20.005 ;
        RECT 965.625 19.960 965.915 20.005 ;
        RECT 954.585 19.820 965.915 19.960 ;
        RECT 954.585 19.775 954.875 19.820 ;
        RECT 965.625 19.775 965.915 19.820 ;
        RECT 967.005 19.960 967.295 20.005 ;
        RECT 1447.690 19.960 1448.010 20.020 ;
        RECT 967.005 19.820 1448.010 19.960 ;
        RECT 967.005 19.775 967.295 19.820 ;
        RECT 1447.690 19.760 1448.010 19.820 ;
        RECT 920.990 18.600 921.310 18.660 ;
        RECT 954.125 18.600 954.415 18.645 ;
        RECT 920.990 18.460 954.415 18.600 ;
        RECT 920.990 18.400 921.310 18.460 ;
        RECT 954.125 18.415 954.415 18.460 ;
      LAYER via ;
        RECT 846.040 1589.880 846.300 1590.140 ;
        RECT 921.020 1589.540 921.280 1589.800 ;
        RECT 1447.720 19.760 1447.980 20.020 ;
        RECT 921.020 18.400 921.280 18.660 ;
      LAYER met2 ;
        RECT 846.040 1600.000 846.320 1604.000 ;
        RECT 846.100 1590.170 846.240 1600.000 ;
        RECT 846.040 1589.850 846.300 1590.170 ;
        RECT 921.020 1589.510 921.280 1589.830 ;
        RECT 921.080 18.690 921.220 1589.510 ;
        RECT 1447.720 19.730 1447.980 20.050 ;
        RECT 921.020 18.370 921.280 18.690 ;
        RECT 1447.780 2.400 1447.920 19.730 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1357.605 1589.245 1357.775 1592.475 ;
        RECT 1389.805 15.215 1389.975 16.915 ;
        RECT 1390.725 15.215 1390.895 15.555 ;
        RECT 1412.805 15.385 1412.975 16.575 ;
        RECT 1389.805 15.045 1390.895 15.215 ;
      LAYER mcon ;
        RECT 1357.605 1592.305 1357.775 1592.475 ;
        RECT 1389.805 16.745 1389.975 16.915 ;
        RECT 1412.805 16.405 1412.975 16.575 ;
        RECT 1390.725 15.385 1390.895 15.555 ;
      LAYER met1 ;
        RECT 852.910 1592.460 853.230 1592.520 ;
        RECT 1357.545 1592.460 1357.835 1592.505 ;
        RECT 852.910 1592.320 1357.835 1592.460 ;
        RECT 852.910 1592.260 853.230 1592.320 ;
        RECT 1357.545 1592.275 1357.835 1592.320 ;
        RECT 1357.545 1589.400 1357.835 1589.445 ;
        RECT 1376.390 1589.400 1376.710 1589.460 ;
        RECT 1357.545 1589.260 1376.710 1589.400 ;
        RECT 1357.545 1589.215 1357.835 1589.260 ;
        RECT 1376.390 1589.200 1376.710 1589.260 ;
        RECT 1376.390 16.900 1376.710 16.960 ;
        RECT 1389.745 16.900 1390.035 16.945 ;
        RECT 1376.390 16.760 1390.035 16.900 ;
        RECT 1376.390 16.700 1376.710 16.760 ;
        RECT 1389.745 16.715 1390.035 16.760 ;
        RECT 1412.745 16.560 1413.035 16.605 ;
        RECT 1465.630 16.560 1465.950 16.620 ;
        RECT 1412.745 16.420 1465.950 16.560 ;
        RECT 1412.745 16.375 1413.035 16.420 ;
        RECT 1465.630 16.360 1465.950 16.420 ;
        RECT 1390.665 15.540 1390.955 15.585 ;
        RECT 1412.745 15.540 1413.035 15.585 ;
        RECT 1390.665 15.400 1413.035 15.540 ;
        RECT 1390.665 15.355 1390.955 15.400 ;
        RECT 1412.745 15.355 1413.035 15.400 ;
      LAYER via ;
        RECT 852.940 1592.260 853.200 1592.520 ;
        RECT 1376.420 1589.200 1376.680 1589.460 ;
        RECT 1376.420 16.700 1376.680 16.960 ;
        RECT 1465.660 16.360 1465.920 16.620 ;
      LAYER met2 ;
        RECT 852.940 1600.000 853.220 1604.000 ;
        RECT 853.000 1592.550 853.140 1600.000 ;
        RECT 852.940 1592.230 853.200 1592.550 ;
        RECT 1376.420 1589.170 1376.680 1589.490 ;
        RECT 1376.480 16.990 1376.620 1589.170 ;
        RECT 1376.420 16.670 1376.680 16.990 ;
        RECT 1465.660 16.330 1465.920 16.650 ;
        RECT 1465.720 2.400 1465.860 16.330 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 859.810 1592.120 860.130 1592.180 ;
        RECT 1397.090 1592.120 1397.410 1592.180 ;
        RECT 859.810 1591.980 1397.410 1592.120 ;
        RECT 859.810 1591.920 860.130 1591.980 ;
        RECT 1397.090 1591.920 1397.410 1591.980 ;
        RECT 1397.090 14.180 1397.410 14.240 ;
        RECT 1483.570 14.180 1483.890 14.240 ;
        RECT 1397.090 14.040 1483.890 14.180 ;
        RECT 1397.090 13.980 1397.410 14.040 ;
        RECT 1483.570 13.980 1483.890 14.040 ;
      LAYER via ;
        RECT 859.840 1591.920 860.100 1592.180 ;
        RECT 1397.120 1591.920 1397.380 1592.180 ;
        RECT 1397.120 13.980 1397.380 14.240 ;
        RECT 1483.600 13.980 1483.860 14.240 ;
      LAYER met2 ;
        RECT 859.840 1600.000 860.120 1604.000 ;
        RECT 859.900 1592.210 860.040 1600.000 ;
        RECT 859.840 1591.890 860.100 1592.210 ;
        RECT 1397.120 1591.890 1397.380 1592.210 ;
        RECT 1397.180 14.270 1397.320 1591.890 ;
        RECT 1397.120 13.950 1397.380 14.270 ;
        RECT 1483.600 13.950 1483.860 14.270 ;
        RECT 1483.660 2.400 1483.800 13.950 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 935.325 18.785 935.495 20.655 ;
      LAYER mcon ;
        RECT 935.325 20.485 935.495 20.655 ;
      LAYER met1 ;
        RECT 903.600 1589.600 904.200 1589.740 ;
        RECT 903.600 1589.400 903.740 1589.600 ;
        RECT 903.140 1589.260 903.740 1589.400 ;
        RECT 904.060 1589.400 904.200 1589.600 ;
        RECT 927.890 1589.400 928.210 1589.460 ;
        RECT 904.060 1589.260 928.210 1589.400 ;
        RECT 866.250 1589.060 866.570 1589.120 ;
        RECT 903.140 1589.060 903.280 1589.260 ;
        RECT 927.890 1589.200 928.210 1589.260 ;
        RECT 866.250 1588.920 903.280 1589.060 ;
        RECT 866.250 1588.860 866.570 1588.920 ;
        RECT 935.265 20.640 935.555 20.685 ;
        RECT 1501.510 20.640 1501.830 20.700 ;
        RECT 935.265 20.500 1501.830 20.640 ;
        RECT 935.265 20.455 935.555 20.500 ;
        RECT 1501.510 20.440 1501.830 20.500 ;
        RECT 927.890 18.940 928.210 19.000 ;
        RECT 935.265 18.940 935.555 18.985 ;
        RECT 927.890 18.800 935.555 18.940 ;
        RECT 927.890 18.740 928.210 18.800 ;
        RECT 935.265 18.755 935.555 18.800 ;
      LAYER via ;
        RECT 866.280 1588.860 866.540 1589.120 ;
        RECT 927.920 1589.200 928.180 1589.460 ;
        RECT 1501.540 20.440 1501.800 20.700 ;
        RECT 927.920 18.740 928.180 19.000 ;
      LAYER met2 ;
        RECT 866.280 1600.000 866.560 1604.000 ;
        RECT 866.340 1589.150 866.480 1600.000 ;
        RECT 927.920 1589.170 928.180 1589.490 ;
        RECT 866.280 1588.830 866.540 1589.150 ;
        RECT 927.980 19.030 928.120 1589.170 ;
        RECT 1501.540 20.410 1501.800 20.730 ;
        RECT 927.920 18.710 928.180 19.030 ;
        RECT 1501.600 2.400 1501.740 20.410 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 873.150 1591.780 873.470 1591.840 ;
        RECT 1431.590 1591.780 1431.910 1591.840 ;
        RECT 873.150 1591.640 1431.910 1591.780 ;
        RECT 873.150 1591.580 873.470 1591.640 ;
        RECT 1431.590 1591.580 1431.910 1591.640 ;
        RECT 1431.590 14.520 1431.910 14.580 ;
        RECT 1518.990 14.520 1519.310 14.580 ;
        RECT 1431.590 14.380 1519.310 14.520 ;
        RECT 1431.590 14.320 1431.910 14.380 ;
        RECT 1518.990 14.320 1519.310 14.380 ;
      LAYER via ;
        RECT 873.180 1591.580 873.440 1591.840 ;
        RECT 1431.620 1591.580 1431.880 1591.840 ;
        RECT 1431.620 14.320 1431.880 14.580 ;
        RECT 1519.020 14.320 1519.280 14.580 ;
      LAYER met2 ;
        RECT 873.180 1600.000 873.460 1604.000 ;
        RECT 873.240 1591.870 873.380 1600.000 ;
        RECT 873.180 1591.550 873.440 1591.870 ;
        RECT 1431.620 1591.550 1431.880 1591.870 ;
        RECT 1431.680 14.610 1431.820 1591.550 ;
        RECT 1431.620 14.290 1431.880 14.610 ;
        RECT 1519.020 14.290 1519.280 14.610 ;
        RECT 1519.080 2.400 1519.220 14.290 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 571.390 15.880 571.710 15.940 ;
        RECT 716.290 15.880 716.610 15.940 ;
        RECT 571.390 15.740 716.610 15.880 ;
        RECT 571.390 15.680 571.710 15.740 ;
        RECT 716.290 15.680 716.610 15.740 ;
      LAYER via ;
        RECT 571.420 15.680 571.680 15.940 ;
        RECT 716.320 15.680 716.580 15.940 ;
      LAYER met2 ;
        RECT 570.040 1600.450 570.320 1604.000 ;
        RECT 570.040 1600.310 571.620 1600.450 ;
        RECT 570.040 1600.000 570.320 1600.310 ;
        RECT 571.480 15.970 571.620 1600.310 ;
        RECT 571.420 15.650 571.680 15.970 ;
        RECT 716.320 15.650 716.580 15.970 ;
        RECT 716.380 2.400 716.520 15.650 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 879.590 1591.440 879.910 1591.500 ;
        RECT 1521.290 1591.440 1521.610 1591.500 ;
        RECT 879.590 1591.300 1521.610 1591.440 ;
        RECT 879.590 1591.240 879.910 1591.300 ;
        RECT 1521.290 1591.240 1521.610 1591.300 ;
        RECT 1521.290 20.640 1521.610 20.700 ;
        RECT 1536.930 20.640 1537.250 20.700 ;
        RECT 1521.290 20.500 1537.250 20.640 ;
        RECT 1521.290 20.440 1521.610 20.500 ;
        RECT 1536.930 20.440 1537.250 20.500 ;
      LAYER via ;
        RECT 879.620 1591.240 879.880 1591.500 ;
        RECT 1521.320 1591.240 1521.580 1591.500 ;
        RECT 1521.320 20.440 1521.580 20.700 ;
        RECT 1536.960 20.440 1537.220 20.700 ;
      LAYER met2 ;
        RECT 879.620 1600.000 879.900 1604.000 ;
        RECT 879.680 1591.530 879.820 1600.000 ;
        RECT 879.620 1591.210 879.880 1591.530 ;
        RECT 1521.320 1591.210 1521.580 1591.530 ;
        RECT 1521.380 20.730 1521.520 1591.210 ;
        RECT 1521.320 20.410 1521.580 20.730 ;
        RECT 1536.960 20.410 1537.220 20.730 ;
        RECT 1537.020 2.400 1537.160 20.410 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 886.490 1592.800 886.810 1592.860 ;
        RECT 945.370 1592.800 945.690 1592.860 ;
        RECT 886.490 1592.660 945.690 1592.800 ;
        RECT 886.490 1592.600 886.810 1592.660 ;
        RECT 945.370 1592.600 945.690 1592.660 ;
        RECT 945.370 1588.380 945.690 1588.440 ;
        RECT 949.050 1588.380 949.370 1588.440 ;
        RECT 945.370 1588.240 949.370 1588.380 ;
        RECT 945.370 1588.180 945.690 1588.240 ;
        RECT 949.050 1588.180 949.370 1588.240 ;
        RECT 1554.870 20.300 1555.190 20.360 ;
        RECT 966.620 20.160 1555.190 20.300 ;
        RECT 949.050 19.620 949.370 19.680 ;
        RECT 966.620 19.620 966.760 20.160 ;
        RECT 1554.870 20.100 1555.190 20.160 ;
        RECT 949.050 19.480 966.760 19.620 ;
        RECT 949.050 19.420 949.370 19.480 ;
      LAYER via ;
        RECT 886.520 1592.600 886.780 1592.860 ;
        RECT 945.400 1592.600 945.660 1592.860 ;
        RECT 945.400 1588.180 945.660 1588.440 ;
        RECT 949.080 1588.180 949.340 1588.440 ;
        RECT 949.080 19.420 949.340 19.680 ;
        RECT 1554.900 20.100 1555.160 20.360 ;
      LAYER met2 ;
        RECT 886.520 1600.000 886.800 1604.000 ;
        RECT 886.580 1592.890 886.720 1600.000 ;
        RECT 886.520 1592.570 886.780 1592.890 ;
        RECT 945.400 1592.570 945.660 1592.890 ;
        RECT 945.460 1588.470 945.600 1592.570 ;
        RECT 945.400 1588.150 945.660 1588.470 ;
        RECT 949.080 1588.150 949.340 1588.470 ;
        RECT 949.140 19.710 949.280 1588.150 ;
        RECT 1554.900 20.070 1555.160 20.390 ;
        RECT 949.080 19.390 949.340 19.710 ;
        RECT 1554.960 2.400 1555.100 20.070 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 893.420 1600.000 893.700 1604.000 ;
        RECT 893.480 1591.045 893.620 1600.000 ;
        RECT 893.410 1590.675 893.690 1591.045 ;
        RECT 1572.830 16.475 1573.110 16.845 ;
        RECT 1572.900 2.400 1573.040 16.475 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
      LAYER via2 ;
        RECT 893.410 1590.720 893.690 1591.000 ;
        RECT 1572.830 16.520 1573.110 16.800 ;
      LAYER met3 ;
        RECT 893.385 1591.010 893.715 1591.025 ;
        RECT 1555.990 1591.010 1556.370 1591.020 ;
        RECT 893.385 1590.710 1556.370 1591.010 ;
        RECT 893.385 1590.695 893.715 1590.710 ;
        RECT 1555.990 1590.700 1556.370 1590.710 ;
        RECT 1555.990 16.810 1556.370 16.820 ;
        RECT 1572.805 16.810 1573.135 16.825 ;
        RECT 1555.990 16.510 1573.135 16.810 ;
        RECT 1555.990 16.500 1556.370 16.510 ;
        RECT 1572.805 16.495 1573.135 16.510 ;
      LAYER via3 ;
        RECT 1556.020 1590.700 1556.340 1591.020 ;
        RECT 1556.020 16.500 1556.340 16.820 ;
      LAYER met4 ;
        RECT 1556.015 1590.695 1556.345 1591.025 ;
        RECT 1556.030 16.825 1556.330 1590.695 ;
        RECT 1556.015 16.495 1556.345 16.825 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 899.830 1587.360 900.150 1587.420 ;
        RECT 902.590 1587.360 902.910 1587.420 ;
        RECT 899.830 1587.220 902.910 1587.360 ;
        RECT 899.830 1587.160 900.150 1587.220 ;
        RECT 902.590 1587.160 902.910 1587.220 ;
        RECT 902.590 77.760 902.910 77.820 ;
        RECT 1587.070 77.760 1587.390 77.820 ;
        RECT 902.590 77.620 1587.390 77.760 ;
        RECT 902.590 77.560 902.910 77.620 ;
        RECT 1587.070 77.560 1587.390 77.620 ;
        RECT 1587.070 2.960 1587.390 3.020 ;
        RECT 1590.290 2.960 1590.610 3.020 ;
        RECT 1587.070 2.820 1590.610 2.960 ;
        RECT 1587.070 2.760 1587.390 2.820 ;
        RECT 1590.290 2.760 1590.610 2.820 ;
      LAYER via ;
        RECT 899.860 1587.160 900.120 1587.420 ;
        RECT 902.620 1587.160 902.880 1587.420 ;
        RECT 902.620 77.560 902.880 77.820 ;
        RECT 1587.100 77.560 1587.360 77.820 ;
        RECT 1587.100 2.760 1587.360 3.020 ;
        RECT 1590.320 2.760 1590.580 3.020 ;
      LAYER met2 ;
        RECT 899.860 1600.000 900.140 1604.000 ;
        RECT 899.920 1587.450 900.060 1600.000 ;
        RECT 899.860 1587.130 900.120 1587.450 ;
        RECT 902.620 1587.130 902.880 1587.450 ;
        RECT 902.680 77.850 902.820 1587.130 ;
        RECT 902.620 77.530 902.880 77.850 ;
        RECT 1587.100 77.530 1587.360 77.850 ;
        RECT 1587.160 3.050 1587.300 77.530 ;
        RECT 1587.100 2.730 1587.360 3.050 ;
        RECT 1590.320 2.730 1590.580 3.050 ;
        RECT 1590.380 2.400 1590.520 2.730 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 906.760 1600.000 907.040 1604.000 ;
        RECT 906.820 1590.365 906.960 1600.000 ;
        RECT 906.750 1589.995 907.030 1590.365 ;
        RECT 1608.250 16.475 1608.530 16.845 ;
        RECT 1608.320 2.400 1608.460 16.475 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
      LAYER via2 ;
        RECT 906.750 1590.040 907.030 1590.320 ;
        RECT 1608.250 16.520 1608.530 16.800 ;
      LAYER met3 ;
        RECT 906.725 1590.330 907.055 1590.345 ;
        RECT 1607.510 1590.330 1607.890 1590.340 ;
        RECT 906.725 1590.030 1607.890 1590.330 ;
        RECT 906.725 1590.015 907.055 1590.030 ;
        RECT 1607.510 1590.020 1607.890 1590.030 ;
        RECT 1607.510 16.810 1607.890 16.820 ;
        RECT 1608.225 16.810 1608.555 16.825 ;
        RECT 1607.510 16.510 1608.555 16.810 ;
        RECT 1607.510 16.500 1607.890 16.510 ;
        RECT 1608.225 16.495 1608.555 16.510 ;
      LAYER via3 ;
        RECT 1607.540 1590.020 1607.860 1590.340 ;
        RECT 1607.540 16.500 1607.860 16.820 ;
      LAYER met4 ;
        RECT 1607.535 1590.015 1607.865 1590.345 ;
        RECT 1607.550 16.825 1607.850 1590.015 ;
        RECT 1607.535 16.495 1607.865 16.825 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 949.585 1587.885 949.755 1589.075 ;
      LAYER mcon ;
        RECT 949.585 1588.905 949.755 1589.075 ;
      LAYER met1 ;
        RECT 949.525 1589.060 949.815 1589.105 ;
        RECT 1252.190 1589.060 1252.510 1589.120 ;
        RECT 949.525 1588.920 1252.510 1589.060 ;
        RECT 949.525 1588.875 949.815 1588.920 ;
        RECT 1252.190 1588.860 1252.510 1588.920 ;
        RECT 913.630 1588.040 913.950 1588.100 ;
        RECT 949.525 1588.040 949.815 1588.085 ;
        RECT 913.630 1587.900 949.815 1588.040 ;
        RECT 913.630 1587.840 913.950 1587.900 ;
        RECT 949.525 1587.855 949.815 1587.900 ;
        RECT 1252.190 15.200 1252.510 15.260 ;
        RECT 1626.170 15.200 1626.490 15.260 ;
        RECT 1252.190 15.060 1626.490 15.200 ;
        RECT 1252.190 15.000 1252.510 15.060 ;
        RECT 1626.170 15.000 1626.490 15.060 ;
      LAYER via ;
        RECT 1252.220 1588.860 1252.480 1589.120 ;
        RECT 913.660 1587.840 913.920 1588.100 ;
        RECT 1252.220 15.000 1252.480 15.260 ;
        RECT 1626.200 15.000 1626.460 15.260 ;
      LAYER met2 ;
        RECT 913.660 1600.000 913.940 1604.000 ;
        RECT 913.720 1588.130 913.860 1600.000 ;
        RECT 1252.220 1588.830 1252.480 1589.150 ;
        RECT 913.660 1587.810 913.920 1588.130 ;
        RECT 1252.280 15.290 1252.420 1588.830 ;
        RECT 1252.220 14.970 1252.480 15.290 ;
        RECT 1626.200 14.970 1626.460 15.290 ;
        RECT 1626.260 2.400 1626.400 14.970 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 921.450 1589.740 921.770 1589.800 ;
        RECT 921.450 1589.600 935.480 1589.740 ;
        RECT 921.450 1589.540 921.770 1589.600 ;
        RECT 935.340 1589.400 935.480 1589.600 ;
        RECT 1265.530 1589.400 1265.850 1589.460 ;
        RECT 935.340 1589.260 1265.850 1589.400 ;
        RECT 1265.530 1589.200 1265.850 1589.260 ;
        RECT 1265.990 15.880 1266.310 15.940 ;
        RECT 1644.110 15.880 1644.430 15.940 ;
        RECT 1265.990 15.740 1644.430 15.880 ;
        RECT 1265.990 15.680 1266.310 15.740 ;
        RECT 1644.110 15.680 1644.430 15.740 ;
      LAYER via ;
        RECT 921.480 1589.540 921.740 1589.800 ;
        RECT 1265.560 1589.200 1265.820 1589.460 ;
        RECT 1266.020 15.680 1266.280 15.940 ;
        RECT 1644.140 15.680 1644.400 15.940 ;
      LAYER met2 ;
        RECT 920.100 1600.450 920.380 1604.000 ;
        RECT 920.100 1600.310 921.680 1600.450 ;
        RECT 920.100 1600.000 920.380 1600.310 ;
        RECT 921.540 1589.830 921.680 1600.310 ;
        RECT 921.480 1589.510 921.740 1589.830 ;
        RECT 1265.560 1589.170 1265.820 1589.490 ;
        RECT 1265.620 1588.890 1265.760 1589.170 ;
        RECT 1265.620 1588.750 1266.220 1588.890 ;
        RECT 1266.080 15.970 1266.220 1588.750 ;
        RECT 1266.020 15.650 1266.280 15.970 ;
        RECT 1644.140 15.650 1644.400 15.970 ;
        RECT 1644.200 2.400 1644.340 15.650 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 926.970 1589.060 927.290 1589.120 ;
        RECT 948.590 1589.060 948.910 1589.120 ;
        RECT 926.970 1588.920 948.910 1589.060 ;
        RECT 926.970 1588.860 927.290 1588.920 ;
        RECT 948.590 1588.860 948.910 1588.920 ;
        RECT 1662.050 19.620 1662.370 19.680 ;
        RECT 967.080 19.480 1662.370 19.620 ;
        RECT 967.080 19.280 967.220 19.480 ;
        RECT 1662.050 19.420 1662.370 19.480 ;
        RECT 955.120 19.140 967.220 19.280 ;
        RECT 952.270 18.940 952.590 19.000 ;
        RECT 955.120 18.940 955.260 19.140 ;
        RECT 952.270 18.800 955.260 18.940 ;
        RECT 952.270 18.740 952.590 18.800 ;
        RECT 948.590 18.260 948.910 18.320 ;
        RECT 951.350 18.260 951.670 18.320 ;
        RECT 948.590 18.120 951.670 18.260 ;
        RECT 948.590 18.060 948.910 18.120 ;
        RECT 951.350 18.060 951.670 18.120 ;
      LAYER via ;
        RECT 927.000 1588.860 927.260 1589.120 ;
        RECT 948.620 1588.860 948.880 1589.120 ;
        RECT 1662.080 19.420 1662.340 19.680 ;
        RECT 952.300 18.740 952.560 19.000 ;
        RECT 948.620 18.060 948.880 18.320 ;
        RECT 951.380 18.060 951.640 18.320 ;
      LAYER met2 ;
        RECT 927.000 1600.000 927.280 1604.000 ;
        RECT 927.060 1589.150 927.200 1600.000 ;
        RECT 927.000 1588.830 927.260 1589.150 ;
        RECT 948.620 1588.830 948.880 1589.150 ;
        RECT 948.680 18.350 948.820 1588.830 ;
        RECT 1662.080 19.390 1662.340 19.710 ;
        RECT 952.300 18.770 952.560 19.030 ;
        RECT 951.440 18.710 952.560 18.770 ;
        RECT 951.440 18.630 952.500 18.710 ;
        RECT 951.440 18.350 951.580 18.630 ;
        RECT 948.620 18.030 948.880 18.350 ;
        RECT 951.380 18.030 951.640 18.350 ;
        RECT 1662.140 2.400 1662.280 19.390 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 933.870 1593.140 934.190 1593.200 ;
        RECT 969.290 1593.140 969.610 1593.200 ;
        RECT 933.870 1593.000 969.610 1593.140 ;
        RECT 933.870 1592.940 934.190 1593.000 ;
        RECT 969.290 1592.940 969.610 1593.000 ;
        RECT 969.290 19.280 969.610 19.340 ;
        RECT 1679.530 19.280 1679.850 19.340 ;
        RECT 969.290 19.140 1679.850 19.280 ;
        RECT 969.290 19.080 969.610 19.140 ;
        RECT 1679.530 19.080 1679.850 19.140 ;
      LAYER via ;
        RECT 933.900 1592.940 934.160 1593.200 ;
        RECT 969.320 1592.940 969.580 1593.200 ;
        RECT 969.320 19.080 969.580 19.340 ;
        RECT 1679.560 19.080 1679.820 19.340 ;
      LAYER met2 ;
        RECT 933.900 1600.000 934.180 1604.000 ;
        RECT 933.960 1593.230 934.100 1600.000 ;
        RECT 933.900 1592.910 934.160 1593.230 ;
        RECT 969.320 1592.910 969.580 1593.230 ;
        RECT 969.380 19.370 969.520 1592.910 ;
        RECT 969.320 19.050 969.580 19.370 ;
        RECT 1679.560 19.050 1679.820 19.370 ;
        RECT 1679.620 2.400 1679.760 19.050 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1242.605 1587.885 1242.775 1588.735 ;
      LAYER mcon ;
        RECT 1242.605 1588.565 1242.775 1588.735 ;
      LAYER met1 ;
        RECT 940.310 1588.720 940.630 1588.780 ;
        RECT 1242.545 1588.720 1242.835 1588.765 ;
        RECT 940.310 1588.580 1242.835 1588.720 ;
        RECT 940.310 1588.520 940.630 1588.580 ;
        RECT 1242.545 1588.535 1242.835 1588.580 ;
        RECT 1242.545 1588.040 1242.835 1588.085 ;
        RECT 1279.790 1588.040 1280.110 1588.100 ;
        RECT 1242.545 1587.900 1280.110 1588.040 ;
        RECT 1242.545 1587.855 1242.835 1587.900 ;
        RECT 1279.790 1587.840 1280.110 1587.900 ;
        RECT 1279.790 16.220 1280.110 16.280 ;
        RECT 1697.470 16.220 1697.790 16.280 ;
        RECT 1279.790 16.080 1697.790 16.220 ;
        RECT 1279.790 16.020 1280.110 16.080 ;
        RECT 1697.470 16.020 1697.790 16.080 ;
      LAYER via ;
        RECT 940.340 1588.520 940.600 1588.780 ;
        RECT 1279.820 1587.840 1280.080 1588.100 ;
        RECT 1279.820 16.020 1280.080 16.280 ;
        RECT 1697.500 16.020 1697.760 16.280 ;
      LAYER met2 ;
        RECT 940.340 1600.000 940.620 1604.000 ;
        RECT 940.400 1588.810 940.540 1600.000 ;
        RECT 940.340 1588.490 940.600 1588.810 ;
        RECT 1279.820 1587.810 1280.080 1588.130 ;
        RECT 1279.880 16.310 1280.020 1587.810 ;
        RECT 1279.820 15.990 1280.080 16.310 ;
        RECT 1697.500 15.990 1697.760 16.310 ;
        RECT 1697.560 2.400 1697.700 15.990 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 576.940 1600.450 577.220 1604.000 ;
        RECT 576.940 1600.310 578.980 1600.450 ;
        RECT 576.940 1600.000 577.220 1600.310 ;
        RECT 578.840 14.805 578.980 1600.310 ;
        RECT 578.770 14.435 579.050 14.805 ;
        RECT 734.250 14.435 734.530 14.805 ;
        RECT 734.320 2.400 734.460 14.435 ;
        RECT 734.110 -4.800 734.670 2.400 ;
      LAYER via2 ;
        RECT 578.770 14.480 579.050 14.760 ;
        RECT 734.250 14.480 734.530 14.760 ;
      LAYER met3 ;
        RECT 578.745 14.770 579.075 14.785 ;
        RECT 734.225 14.770 734.555 14.785 ;
        RECT 578.745 14.470 734.555 14.770 ;
        RECT 578.745 14.455 579.075 14.470 ;
        RECT 734.225 14.455 734.555 14.470 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 950.890 62.460 951.210 62.520 ;
        RECT 1711.270 62.460 1711.590 62.520 ;
        RECT 950.890 62.320 1711.590 62.460 ;
        RECT 950.890 62.260 951.210 62.320 ;
        RECT 1711.270 62.260 1711.590 62.320 ;
        RECT 1711.270 2.960 1711.590 3.020 ;
        RECT 1715.410 2.960 1715.730 3.020 ;
        RECT 1711.270 2.820 1715.730 2.960 ;
        RECT 1711.270 2.760 1711.590 2.820 ;
        RECT 1715.410 2.760 1715.730 2.820 ;
      LAYER via ;
        RECT 950.920 62.260 951.180 62.520 ;
        RECT 1711.300 62.260 1711.560 62.520 ;
        RECT 1711.300 2.760 1711.560 3.020 ;
        RECT 1715.440 2.760 1715.700 3.020 ;
      LAYER met2 ;
        RECT 947.240 1600.450 947.520 1604.000 ;
        RECT 947.240 1600.310 949.280 1600.450 ;
        RECT 947.240 1600.000 947.520 1600.310 ;
        RECT 949.140 1589.570 949.280 1600.310 ;
        RECT 949.140 1589.430 951.120 1589.570 ;
        RECT 950.980 62.550 951.120 1589.430 ;
        RECT 950.920 62.230 951.180 62.550 ;
        RECT 1711.300 62.230 1711.560 62.550 ;
        RECT 1711.360 3.050 1711.500 62.230 ;
        RECT 1711.300 2.730 1711.560 3.050 ;
        RECT 1715.440 2.730 1715.700 3.050 ;
        RECT 1715.500 2.400 1715.640 2.730 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 953.650 1588.380 953.970 1588.440 ;
        RECT 958.710 1588.380 959.030 1588.440 ;
        RECT 953.650 1588.240 959.030 1588.380 ;
        RECT 953.650 1588.180 953.970 1588.240 ;
        RECT 958.710 1588.180 959.030 1588.240 ;
        RECT 958.710 18.940 959.030 19.000 ;
        RECT 1733.350 18.940 1733.670 19.000 ;
        RECT 958.710 18.800 1733.670 18.940 ;
        RECT 958.710 18.740 959.030 18.800 ;
        RECT 1733.350 18.740 1733.670 18.800 ;
      LAYER via ;
        RECT 953.680 1588.180 953.940 1588.440 ;
        RECT 958.740 1588.180 959.000 1588.440 ;
        RECT 958.740 18.740 959.000 19.000 ;
        RECT 1733.380 18.740 1733.640 19.000 ;
      LAYER met2 ;
        RECT 953.680 1600.000 953.960 1604.000 ;
        RECT 953.740 1588.470 953.880 1600.000 ;
        RECT 953.680 1588.150 953.940 1588.470 ;
        RECT 958.740 1588.150 959.000 1588.470 ;
        RECT 958.800 19.030 958.940 1588.150 ;
        RECT 958.740 18.710 959.000 19.030 ;
        RECT 1733.380 18.710 1733.640 19.030 ;
        RECT 1733.440 2.400 1733.580 18.710 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 960.550 1590.080 960.870 1590.140 ;
        RECT 964.690 1590.080 965.010 1590.140 ;
        RECT 960.550 1589.940 965.010 1590.080 ;
        RECT 960.550 1589.880 960.870 1589.940 ;
        RECT 964.690 1589.880 965.010 1589.940 ;
        RECT 964.690 62.800 965.010 62.860 ;
        RECT 1745.770 62.800 1746.090 62.860 ;
        RECT 964.690 62.660 1746.090 62.800 ;
        RECT 964.690 62.600 965.010 62.660 ;
        RECT 1745.770 62.600 1746.090 62.660 ;
      LAYER via ;
        RECT 960.580 1589.880 960.840 1590.140 ;
        RECT 964.720 1589.880 964.980 1590.140 ;
        RECT 964.720 62.600 964.980 62.860 ;
        RECT 1745.800 62.600 1746.060 62.860 ;
      LAYER met2 ;
        RECT 960.580 1600.000 960.860 1604.000 ;
        RECT 960.640 1590.170 960.780 1600.000 ;
        RECT 960.580 1589.850 960.840 1590.170 ;
        RECT 964.720 1589.850 964.980 1590.170 ;
        RECT 964.780 62.890 964.920 1589.850 ;
        RECT 964.720 62.570 964.980 62.890 ;
        RECT 1745.800 62.570 1746.060 62.890 ;
        RECT 1745.860 16.730 1746.000 62.570 ;
        RECT 1745.860 16.590 1751.520 16.730 ;
        RECT 1751.380 2.400 1751.520 16.590 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 967.450 1592.800 967.770 1592.860 ;
        RECT 1445.390 1592.800 1445.710 1592.860 ;
        RECT 967.450 1592.660 1445.710 1592.800 ;
        RECT 967.450 1592.600 967.770 1592.660 ;
        RECT 1445.390 1592.600 1445.710 1592.660 ;
        RECT 1445.390 14.860 1445.710 14.920 ;
        RECT 1768.770 14.860 1769.090 14.920 ;
        RECT 1445.390 14.720 1769.090 14.860 ;
        RECT 1445.390 14.660 1445.710 14.720 ;
        RECT 1768.770 14.660 1769.090 14.720 ;
      LAYER via ;
        RECT 967.480 1592.600 967.740 1592.860 ;
        RECT 1445.420 1592.600 1445.680 1592.860 ;
        RECT 1445.420 14.660 1445.680 14.920 ;
        RECT 1768.800 14.660 1769.060 14.920 ;
      LAYER met2 ;
        RECT 967.480 1600.000 967.760 1604.000 ;
        RECT 967.540 1592.890 967.680 1600.000 ;
        RECT 967.480 1592.570 967.740 1592.890 ;
        RECT 1445.420 1592.570 1445.680 1592.890 ;
        RECT 1445.480 14.950 1445.620 1592.570 ;
        RECT 1445.420 14.630 1445.680 14.950 ;
        RECT 1768.800 14.630 1769.060 14.950 ;
        RECT 1768.860 2.400 1769.000 14.630 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 973.890 1590.080 974.210 1590.140 ;
        RECT 978.490 1590.080 978.810 1590.140 ;
        RECT 973.890 1589.940 978.810 1590.080 ;
        RECT 973.890 1589.880 974.210 1589.940 ;
        RECT 978.490 1589.880 978.810 1589.940 ;
        RECT 978.490 63.140 978.810 63.200 ;
        RECT 1780.270 63.140 1780.590 63.200 ;
        RECT 978.490 63.000 1780.590 63.140 ;
        RECT 978.490 62.940 978.810 63.000 ;
        RECT 1780.270 62.940 1780.590 63.000 ;
        RECT 1780.270 18.600 1780.590 18.660 ;
        RECT 1786.710 18.600 1787.030 18.660 ;
        RECT 1780.270 18.460 1787.030 18.600 ;
        RECT 1780.270 18.400 1780.590 18.460 ;
        RECT 1786.710 18.400 1787.030 18.460 ;
      LAYER via ;
        RECT 973.920 1589.880 974.180 1590.140 ;
        RECT 978.520 1589.880 978.780 1590.140 ;
        RECT 978.520 62.940 978.780 63.200 ;
        RECT 1780.300 62.940 1780.560 63.200 ;
        RECT 1780.300 18.400 1780.560 18.660 ;
        RECT 1786.740 18.400 1787.000 18.660 ;
      LAYER met2 ;
        RECT 973.920 1600.000 974.200 1604.000 ;
        RECT 973.980 1590.170 974.120 1600.000 ;
        RECT 973.920 1589.850 974.180 1590.170 ;
        RECT 978.520 1589.850 978.780 1590.170 ;
        RECT 978.580 63.230 978.720 1589.850 ;
        RECT 978.520 62.910 978.780 63.230 ;
        RECT 1780.300 62.910 1780.560 63.230 ;
        RECT 1780.360 18.690 1780.500 62.910 ;
        RECT 1780.300 18.370 1780.560 18.690 ;
        RECT 1786.740 18.370 1787.000 18.690 ;
        RECT 1786.800 2.400 1786.940 18.370 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 980.790 1589.740 981.110 1589.800 ;
        RECT 986.310 1589.740 986.630 1589.800 ;
        RECT 980.790 1589.600 986.630 1589.740 ;
        RECT 980.790 1589.540 981.110 1589.600 ;
        RECT 986.310 1589.540 986.630 1589.600 ;
        RECT 1804.650 18.940 1804.970 19.000 ;
        RECT 1779.900 18.800 1804.970 18.940 ;
        RECT 1779.900 18.600 1780.040 18.800 ;
        RECT 1804.650 18.740 1804.970 18.800 ;
        RECT 1005.720 18.460 1780.040 18.600 ;
        RECT 986.310 18.260 986.630 18.320 ;
        RECT 1005.720 18.260 1005.860 18.460 ;
        RECT 986.310 18.120 1005.860 18.260 ;
        RECT 986.310 18.060 986.630 18.120 ;
      LAYER via ;
        RECT 980.820 1589.540 981.080 1589.800 ;
        RECT 986.340 1589.540 986.600 1589.800 ;
        RECT 1804.680 18.740 1804.940 19.000 ;
        RECT 986.340 18.060 986.600 18.320 ;
      LAYER met2 ;
        RECT 980.820 1600.000 981.100 1604.000 ;
        RECT 980.880 1589.830 981.020 1600.000 ;
        RECT 980.820 1589.510 981.080 1589.830 ;
        RECT 986.340 1589.510 986.600 1589.830 ;
        RECT 986.400 18.350 986.540 1589.510 ;
        RECT 1804.680 18.710 1804.940 19.030 ;
        RECT 986.340 18.030 986.600 18.350 ;
        RECT 1804.740 2.400 1804.880 18.710 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 987.690 1590.080 988.010 1590.140 ;
        RECT 992.290 1590.080 992.610 1590.140 ;
        RECT 987.690 1589.940 992.610 1590.080 ;
        RECT 987.690 1589.880 988.010 1589.940 ;
        RECT 992.290 1589.880 992.610 1589.940 ;
        RECT 992.290 63.480 992.610 63.540 ;
        RECT 1821.670 63.480 1821.990 63.540 ;
        RECT 992.290 63.340 1821.990 63.480 ;
        RECT 992.290 63.280 992.610 63.340 ;
        RECT 1821.670 63.280 1821.990 63.340 ;
        RECT 1821.670 2.960 1821.990 3.020 ;
        RECT 1822.590 2.960 1822.910 3.020 ;
        RECT 1821.670 2.820 1822.910 2.960 ;
        RECT 1821.670 2.760 1821.990 2.820 ;
        RECT 1822.590 2.760 1822.910 2.820 ;
      LAYER via ;
        RECT 987.720 1589.880 987.980 1590.140 ;
        RECT 992.320 1589.880 992.580 1590.140 ;
        RECT 992.320 63.280 992.580 63.540 ;
        RECT 1821.700 63.280 1821.960 63.540 ;
        RECT 1821.700 2.760 1821.960 3.020 ;
        RECT 1822.620 2.760 1822.880 3.020 ;
      LAYER met2 ;
        RECT 987.720 1600.000 988.000 1604.000 ;
        RECT 987.780 1590.170 987.920 1600.000 ;
        RECT 987.720 1589.850 987.980 1590.170 ;
        RECT 992.320 1589.850 992.580 1590.170 ;
        RECT 992.380 63.570 992.520 1589.850 ;
        RECT 992.320 63.250 992.580 63.570 ;
        RECT 1821.700 63.250 1821.960 63.570 ;
        RECT 1821.760 3.050 1821.900 63.250 ;
        RECT 1821.700 2.730 1821.960 3.050 ;
        RECT 1822.620 2.730 1822.880 3.050 ;
        RECT 1822.680 2.400 1822.820 2.730 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 994.130 1593.140 994.450 1593.200 ;
        RECT 1459.190 1593.140 1459.510 1593.200 ;
        RECT 994.130 1593.000 1459.510 1593.140 ;
        RECT 994.130 1592.940 994.450 1593.000 ;
        RECT 1459.190 1592.940 1459.510 1593.000 ;
        RECT 1459.190 15.540 1459.510 15.600 ;
        RECT 1840.070 15.540 1840.390 15.600 ;
        RECT 1459.190 15.400 1840.390 15.540 ;
        RECT 1459.190 15.340 1459.510 15.400 ;
        RECT 1840.070 15.340 1840.390 15.400 ;
      LAYER via ;
        RECT 994.160 1592.940 994.420 1593.200 ;
        RECT 1459.220 1592.940 1459.480 1593.200 ;
        RECT 1459.220 15.340 1459.480 15.600 ;
        RECT 1840.100 15.340 1840.360 15.600 ;
      LAYER met2 ;
        RECT 994.160 1600.000 994.440 1604.000 ;
        RECT 994.220 1593.230 994.360 1600.000 ;
        RECT 994.160 1592.910 994.420 1593.230 ;
        RECT 1459.220 1592.910 1459.480 1593.230 ;
        RECT 1459.280 15.630 1459.420 1592.910 ;
        RECT 1459.220 15.310 1459.480 15.630 ;
        RECT 1840.100 15.310 1840.360 15.630 ;
        RECT 1840.160 2.400 1840.300 15.310 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1001.030 1590.080 1001.350 1590.140 ;
        RECT 1006.090 1590.080 1006.410 1590.140 ;
        RECT 1001.030 1589.940 1006.410 1590.080 ;
        RECT 1001.030 1589.880 1001.350 1589.940 ;
        RECT 1006.090 1589.880 1006.410 1589.940 ;
        RECT 1006.090 63.820 1006.410 63.880 ;
        RECT 1856.170 63.820 1856.490 63.880 ;
        RECT 1006.090 63.680 1856.490 63.820 ;
        RECT 1006.090 63.620 1006.410 63.680 ;
        RECT 1856.170 63.620 1856.490 63.680 ;
      LAYER via ;
        RECT 1001.060 1589.880 1001.320 1590.140 ;
        RECT 1006.120 1589.880 1006.380 1590.140 ;
        RECT 1006.120 63.620 1006.380 63.880 ;
        RECT 1856.200 63.620 1856.460 63.880 ;
      LAYER met2 ;
        RECT 1001.060 1600.000 1001.340 1604.000 ;
        RECT 1001.120 1590.170 1001.260 1600.000 ;
        RECT 1001.060 1589.850 1001.320 1590.170 ;
        RECT 1006.120 1589.850 1006.380 1590.170 ;
        RECT 1006.180 63.910 1006.320 1589.850 ;
        RECT 1006.120 63.590 1006.380 63.910 ;
        RECT 1856.200 63.590 1856.460 63.910 ;
        RECT 1856.260 3.130 1856.400 63.590 ;
        RECT 1856.260 2.990 1858.240 3.130 ;
        RECT 1858.100 2.400 1858.240 2.990 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.930 1590.080 1008.250 1590.140 ;
        RECT 1012.990 1590.080 1013.310 1590.140 ;
        RECT 1007.930 1589.940 1013.310 1590.080 ;
        RECT 1007.930 1589.880 1008.250 1589.940 ;
        RECT 1012.990 1589.880 1013.310 1589.940 ;
        RECT 1012.990 64.160 1013.310 64.220 ;
        RECT 1869.970 64.160 1870.290 64.220 ;
        RECT 1012.990 64.020 1870.290 64.160 ;
        RECT 1012.990 63.960 1013.310 64.020 ;
        RECT 1869.970 63.960 1870.290 64.020 ;
        RECT 1869.970 18.600 1870.290 18.660 ;
        RECT 1875.950 18.600 1876.270 18.660 ;
        RECT 1869.970 18.460 1876.270 18.600 ;
        RECT 1869.970 18.400 1870.290 18.460 ;
        RECT 1875.950 18.400 1876.270 18.460 ;
      LAYER via ;
        RECT 1007.960 1589.880 1008.220 1590.140 ;
        RECT 1013.020 1589.880 1013.280 1590.140 ;
        RECT 1013.020 63.960 1013.280 64.220 ;
        RECT 1870.000 63.960 1870.260 64.220 ;
        RECT 1870.000 18.400 1870.260 18.660 ;
        RECT 1875.980 18.400 1876.240 18.660 ;
      LAYER met2 ;
        RECT 1007.960 1600.000 1008.240 1604.000 ;
        RECT 1008.020 1590.170 1008.160 1600.000 ;
        RECT 1007.960 1589.850 1008.220 1590.170 ;
        RECT 1013.020 1589.850 1013.280 1590.170 ;
        RECT 1013.080 64.250 1013.220 1589.850 ;
        RECT 1013.020 63.930 1013.280 64.250 ;
        RECT 1870.000 63.930 1870.260 64.250 ;
        RECT 1870.060 18.690 1870.200 63.930 ;
        RECT 1870.000 18.370 1870.260 18.690 ;
        RECT 1875.980 18.370 1876.240 18.690 ;
        RECT 1876.040 2.400 1876.180 18.370 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 741.205 20.485 741.835 20.655 ;
        RECT 741.665 18.445 741.835 20.485 ;
      LAYER met1 ;
        RECT 586.110 20.640 586.430 20.700 ;
        RECT 741.145 20.640 741.435 20.685 ;
        RECT 586.110 20.500 741.435 20.640 ;
        RECT 586.110 20.440 586.430 20.500 ;
        RECT 741.145 20.455 741.435 20.500 ;
        RECT 741.605 18.600 741.895 18.645 ;
        RECT 752.170 18.600 752.490 18.660 ;
        RECT 741.605 18.460 752.490 18.600 ;
        RECT 741.605 18.415 741.895 18.460 ;
        RECT 752.170 18.400 752.490 18.460 ;
      LAYER via ;
        RECT 586.140 20.440 586.400 20.700 ;
        RECT 752.200 18.400 752.460 18.660 ;
      LAYER met2 ;
        RECT 583.380 1600.450 583.660 1604.000 ;
        RECT 583.380 1600.310 585.420 1600.450 ;
        RECT 583.380 1600.000 583.660 1600.310 ;
        RECT 585.280 1580.050 585.420 1600.310 ;
        RECT 585.280 1579.910 586.340 1580.050 ;
        RECT 586.200 20.730 586.340 1579.910 ;
        RECT 586.140 20.410 586.400 20.730 ;
        RECT 752.200 18.370 752.460 18.690 ;
        RECT 752.260 2.400 752.400 18.370 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1014.370 1590.080 1014.690 1590.140 ;
        RECT 1019.890 1590.080 1020.210 1590.140 ;
        RECT 1014.370 1589.940 1020.210 1590.080 ;
        RECT 1014.370 1589.880 1014.690 1589.940 ;
        RECT 1019.890 1589.880 1020.210 1589.940 ;
        RECT 1019.890 64.500 1020.210 64.560 ;
        RECT 1890.670 64.500 1890.990 64.560 ;
        RECT 1019.890 64.360 1890.990 64.500 ;
        RECT 1019.890 64.300 1020.210 64.360 ;
        RECT 1890.670 64.300 1890.990 64.360 ;
        RECT 1890.670 2.960 1890.990 3.020 ;
        RECT 1893.890 2.960 1894.210 3.020 ;
        RECT 1890.670 2.820 1894.210 2.960 ;
        RECT 1890.670 2.760 1890.990 2.820 ;
        RECT 1893.890 2.760 1894.210 2.820 ;
      LAYER via ;
        RECT 1014.400 1589.880 1014.660 1590.140 ;
        RECT 1019.920 1589.880 1020.180 1590.140 ;
        RECT 1019.920 64.300 1020.180 64.560 ;
        RECT 1890.700 64.300 1890.960 64.560 ;
        RECT 1890.700 2.760 1890.960 3.020 ;
        RECT 1893.920 2.760 1894.180 3.020 ;
      LAYER met2 ;
        RECT 1014.400 1600.000 1014.680 1604.000 ;
        RECT 1014.460 1590.170 1014.600 1600.000 ;
        RECT 1014.400 1589.850 1014.660 1590.170 ;
        RECT 1019.920 1589.850 1020.180 1590.170 ;
        RECT 1019.980 64.590 1020.120 1589.850 ;
        RECT 1019.920 64.270 1020.180 64.590 ;
        RECT 1890.700 64.270 1890.960 64.590 ;
        RECT 1890.760 3.050 1890.900 64.270 ;
        RECT 1890.700 2.730 1890.960 3.050 ;
        RECT 1893.920 2.730 1894.180 3.050 ;
        RECT 1893.980 2.400 1894.120 2.730 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1390.265 15.385 1390.435 16.915 ;
      LAYER mcon ;
        RECT 1390.265 16.745 1390.435 16.915 ;
      LAYER met1 ;
        RECT 1356.150 1588.380 1356.470 1588.440 ;
        RECT 1048.500 1588.240 1356.470 1588.380 ;
        RECT 1021.270 1587.700 1021.590 1587.760 ;
        RECT 1048.500 1587.700 1048.640 1588.240 ;
        RECT 1356.150 1588.180 1356.470 1588.240 ;
        RECT 1021.270 1587.560 1048.640 1587.700 ;
        RECT 1021.270 1587.500 1021.590 1587.560 ;
        RECT 1390.205 16.900 1390.495 16.945 ;
        RECT 1911.830 16.900 1912.150 16.960 ;
        RECT 1390.205 16.760 1912.150 16.900 ;
        RECT 1390.205 16.715 1390.495 16.760 ;
        RECT 1911.830 16.700 1912.150 16.760 ;
        RECT 1356.150 15.540 1356.470 15.600 ;
        RECT 1390.205 15.540 1390.495 15.585 ;
        RECT 1356.150 15.400 1390.495 15.540 ;
        RECT 1356.150 15.340 1356.470 15.400 ;
        RECT 1390.205 15.355 1390.495 15.400 ;
      LAYER via ;
        RECT 1021.300 1587.500 1021.560 1587.760 ;
        RECT 1356.180 1588.180 1356.440 1588.440 ;
        RECT 1911.860 16.700 1912.120 16.960 ;
        RECT 1356.180 15.340 1356.440 15.600 ;
      LAYER met2 ;
        RECT 1021.300 1600.000 1021.580 1604.000 ;
        RECT 1021.360 1587.790 1021.500 1600.000 ;
        RECT 1356.180 1588.150 1356.440 1588.470 ;
        RECT 1021.300 1587.470 1021.560 1587.790 ;
        RECT 1356.240 15.630 1356.380 1588.150 ;
        RECT 1911.860 16.670 1912.120 16.990 ;
        RECT 1356.180 15.310 1356.440 15.630 ;
        RECT 1911.920 2.400 1912.060 16.670 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1026.790 1590.080 1027.110 1590.140 ;
        RECT 1027.710 1590.080 1028.030 1590.140 ;
        RECT 1026.790 1589.940 1028.030 1590.080 ;
        RECT 1026.790 1589.880 1027.110 1589.940 ;
        RECT 1027.710 1589.880 1028.030 1589.940 ;
        RECT 1026.790 64.840 1027.110 64.900 ;
        RECT 1925.170 64.840 1925.490 64.900 ;
        RECT 1026.790 64.700 1925.490 64.840 ;
        RECT 1026.790 64.640 1027.110 64.700 ;
        RECT 1925.170 64.640 1925.490 64.700 ;
      LAYER via ;
        RECT 1026.820 1589.880 1027.080 1590.140 ;
        RECT 1027.740 1589.880 1028.000 1590.140 ;
        RECT 1026.820 64.640 1027.080 64.900 ;
        RECT 1925.200 64.640 1925.460 64.900 ;
      LAYER met2 ;
        RECT 1027.740 1600.000 1028.020 1604.000 ;
        RECT 1027.800 1590.170 1027.940 1600.000 ;
        RECT 1026.820 1589.850 1027.080 1590.170 ;
        RECT 1027.740 1589.850 1028.000 1590.170 ;
        RECT 1026.880 64.930 1027.020 1589.850 ;
        RECT 1026.820 64.610 1027.080 64.930 ;
        RECT 1925.200 64.610 1925.460 64.930 ;
        RECT 1925.260 16.730 1925.400 64.610 ;
        RECT 1925.260 16.590 1929.540 16.730 ;
        RECT 1929.400 2.400 1929.540 16.590 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1034.610 18.260 1034.930 18.320 ;
        RECT 1947.250 18.260 1947.570 18.320 ;
        RECT 1034.610 18.120 1947.570 18.260 ;
        RECT 1034.610 18.060 1034.930 18.120 ;
        RECT 1947.250 18.060 1947.570 18.120 ;
      LAYER via ;
        RECT 1034.640 18.060 1034.900 18.320 ;
        RECT 1947.280 18.060 1947.540 18.320 ;
      LAYER met2 ;
        RECT 1034.640 1600.000 1034.920 1604.000 ;
        RECT 1034.700 18.350 1034.840 1600.000 ;
        RECT 1034.640 18.030 1034.900 18.350 ;
        RECT 1947.280 18.030 1947.540 18.350 ;
        RECT 1947.340 2.400 1947.480 18.030 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.050 65.180 1041.370 65.240 ;
        RECT 1959.670 65.180 1959.990 65.240 ;
        RECT 1041.050 65.040 1959.990 65.180 ;
        RECT 1041.050 64.980 1041.370 65.040 ;
        RECT 1959.670 64.980 1959.990 65.040 ;
      LAYER via ;
        RECT 1041.080 64.980 1041.340 65.240 ;
        RECT 1959.700 64.980 1959.960 65.240 ;
      LAYER met2 ;
        RECT 1041.540 1600.450 1041.820 1604.000 ;
        RECT 1041.140 1600.310 1041.820 1600.450 ;
        RECT 1041.140 65.270 1041.280 1600.310 ;
        RECT 1041.540 1600.000 1041.820 1600.310 ;
        RECT 1041.080 64.950 1041.340 65.270 ;
        RECT 1959.700 64.950 1959.960 65.270 ;
        RECT 1959.760 16.730 1959.900 64.950 ;
        RECT 1959.760 16.590 1965.420 16.730 ;
        RECT 1965.280 2.400 1965.420 16.590 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1048.410 17.920 1048.730 17.980 ;
        RECT 1983.130 17.920 1983.450 17.980 ;
        RECT 1048.410 17.780 1983.450 17.920 ;
        RECT 1048.410 17.720 1048.730 17.780 ;
        RECT 1983.130 17.720 1983.450 17.780 ;
      LAYER via ;
        RECT 1048.440 17.720 1048.700 17.980 ;
        RECT 1983.160 17.720 1983.420 17.980 ;
      LAYER met2 ;
        RECT 1047.980 1600.450 1048.260 1604.000 ;
        RECT 1047.980 1600.310 1048.640 1600.450 ;
        RECT 1047.980 1600.000 1048.260 1600.310 ;
        RECT 1048.500 18.010 1048.640 1600.310 ;
        RECT 1048.440 17.690 1048.700 18.010 ;
        RECT 1983.160 17.690 1983.420 18.010 ;
        RECT 1983.220 2.400 1983.360 17.690 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1088.060 1594.020 1096.940 1594.160 ;
        RECT 1054.850 1593.820 1055.170 1593.880 ;
        RECT 1088.060 1593.820 1088.200 1594.020 ;
        RECT 1054.850 1593.680 1088.200 1593.820 ;
        RECT 1096.800 1593.820 1096.940 1594.020 ;
        RECT 1466.090 1593.820 1466.410 1593.880 ;
        RECT 1096.800 1593.680 1466.410 1593.820 ;
        RECT 1054.850 1593.620 1055.170 1593.680 ;
        RECT 1466.090 1593.620 1466.410 1593.680 ;
        RECT 1466.090 16.560 1466.410 16.620 ;
        RECT 2001.070 16.560 2001.390 16.620 ;
        RECT 1466.090 16.420 2001.390 16.560 ;
        RECT 1466.090 16.360 1466.410 16.420 ;
        RECT 2001.070 16.360 2001.390 16.420 ;
      LAYER via ;
        RECT 1054.880 1593.620 1055.140 1593.880 ;
        RECT 1466.120 1593.620 1466.380 1593.880 ;
        RECT 1466.120 16.360 1466.380 16.620 ;
        RECT 2001.100 16.360 2001.360 16.620 ;
      LAYER met2 ;
        RECT 1054.880 1600.000 1055.160 1604.000 ;
        RECT 1054.940 1593.910 1055.080 1600.000 ;
        RECT 1054.880 1593.590 1055.140 1593.910 ;
        RECT 1466.120 1593.590 1466.380 1593.910 ;
        RECT 1466.180 16.650 1466.320 1593.590 ;
        RECT 1466.120 16.330 1466.380 16.650 ;
        RECT 2001.100 16.330 2001.360 16.650 ;
        RECT 2001.160 2.400 2001.300 16.330 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1061.750 68.920 1062.070 68.980 ;
        RECT 2014.870 68.920 2015.190 68.980 ;
        RECT 1061.750 68.780 2015.190 68.920 ;
        RECT 1061.750 68.720 1062.070 68.780 ;
        RECT 2014.870 68.720 2015.190 68.780 ;
      LAYER via ;
        RECT 1061.780 68.720 1062.040 68.980 ;
        RECT 2014.900 68.720 2015.160 68.980 ;
      LAYER met2 ;
        RECT 1061.780 1600.000 1062.060 1604.000 ;
        RECT 1061.840 69.010 1061.980 1600.000 ;
        RECT 1061.780 68.690 1062.040 69.010 ;
        RECT 2014.900 68.690 2015.160 69.010 ;
        RECT 2014.960 17.410 2015.100 68.690 ;
        RECT 2014.960 17.270 2018.780 17.410 ;
        RECT 2018.640 2.400 2018.780 17.270 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1068.190 78.100 1068.510 78.160 ;
        RECT 2035.570 78.100 2035.890 78.160 ;
        RECT 1068.190 77.960 2035.890 78.100 ;
        RECT 1068.190 77.900 1068.510 77.960 ;
        RECT 2035.570 77.900 2035.890 77.960 ;
      LAYER via ;
        RECT 1068.220 77.900 1068.480 78.160 ;
        RECT 2035.600 77.900 2035.860 78.160 ;
      LAYER met2 ;
        RECT 1068.220 1600.000 1068.500 1604.000 ;
        RECT 1068.280 78.190 1068.420 1600.000 ;
        RECT 1068.220 77.870 1068.480 78.190 ;
        RECT 2035.600 77.870 2035.860 78.190 ;
        RECT 2035.660 17.410 2035.800 77.870 ;
        RECT 2035.660 17.270 2036.720 17.410 ;
        RECT 2036.580 2.400 2036.720 17.270 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.010 17.580 1076.330 17.640 ;
        RECT 2054.430 17.580 2054.750 17.640 ;
        RECT 1076.010 17.440 2054.750 17.580 ;
        RECT 1076.010 17.380 1076.330 17.440 ;
        RECT 2054.430 17.380 2054.750 17.440 ;
      LAYER via ;
        RECT 1076.040 17.380 1076.300 17.640 ;
        RECT 2054.460 17.380 2054.720 17.640 ;
      LAYER met2 ;
        RECT 1075.120 1600.450 1075.400 1604.000 ;
        RECT 1075.120 1600.310 1076.240 1600.450 ;
        RECT 1075.120 1600.000 1075.400 1600.310 ;
        RECT 1076.100 17.670 1076.240 1600.310 ;
        RECT 1076.040 17.350 1076.300 17.670 ;
        RECT 2054.460 17.350 2054.720 17.670 ;
        RECT 2054.520 2.400 2054.660 17.350 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 590.280 1600.450 590.560 1604.000 ;
        RECT 590.280 1600.310 592.320 1600.450 ;
        RECT 590.280 1600.000 590.560 1600.310 ;
        RECT 592.180 1580.050 592.320 1600.310 ;
        RECT 592.180 1579.910 593.240 1580.050 ;
        RECT 593.100 15.485 593.240 1579.910 ;
        RECT 593.030 15.115 593.310 15.485 ;
        RECT 769.670 15.115 769.950 15.485 ;
        RECT 769.740 2.400 769.880 15.115 ;
        RECT 769.530 -4.800 770.090 2.400 ;
      LAYER via2 ;
        RECT 593.030 15.160 593.310 15.440 ;
        RECT 769.670 15.160 769.950 15.440 ;
      LAYER met3 ;
        RECT 593.005 15.450 593.335 15.465 ;
        RECT 769.645 15.450 769.975 15.465 ;
        RECT 593.005 15.150 769.975 15.450 ;
        RECT 593.005 15.135 593.335 15.150 ;
        RECT 769.645 15.135 769.975 15.150 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1081.990 68.580 1082.310 68.640 ;
        RECT 2070.070 68.580 2070.390 68.640 ;
        RECT 1081.990 68.440 2070.390 68.580 ;
        RECT 1081.990 68.380 1082.310 68.440 ;
        RECT 2070.070 68.380 2070.390 68.440 ;
      LAYER via ;
        RECT 1082.020 68.380 1082.280 68.640 ;
        RECT 2070.100 68.380 2070.360 68.640 ;
      LAYER met2 ;
        RECT 1082.020 1600.000 1082.300 1604.000 ;
        RECT 1082.080 68.670 1082.220 1600.000 ;
        RECT 1082.020 68.350 1082.280 68.670 ;
        RECT 2070.100 68.350 2070.360 68.670 ;
        RECT 2070.160 3.130 2070.300 68.350 ;
        RECT 2070.160 2.990 2072.600 3.130 ;
        RECT 2072.460 2.400 2072.600 2.990 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1096.325 1589.925 1096.495 1593.835 ;
      LAYER mcon ;
        RECT 1096.325 1593.665 1096.495 1593.835 ;
      LAYER met1 ;
        RECT 1088.430 1593.820 1088.750 1593.880 ;
        RECT 1096.265 1593.820 1096.555 1593.865 ;
        RECT 1088.430 1593.680 1096.555 1593.820 ;
        RECT 1088.430 1593.620 1088.750 1593.680 ;
        RECT 1096.265 1593.635 1096.555 1593.680 ;
        RECT 1096.265 1590.080 1096.555 1590.125 ;
        RECT 1479.890 1590.080 1480.210 1590.140 ;
        RECT 1096.265 1589.940 1480.210 1590.080 ;
        RECT 1096.265 1589.895 1096.555 1589.940 ;
        RECT 1479.890 1589.880 1480.210 1589.940 ;
        RECT 1479.890 19.960 1480.210 20.020 ;
        RECT 2089.850 19.960 2090.170 20.020 ;
        RECT 1479.890 19.820 2090.170 19.960 ;
        RECT 1479.890 19.760 1480.210 19.820 ;
        RECT 2089.850 19.760 2090.170 19.820 ;
      LAYER via ;
        RECT 1088.460 1593.620 1088.720 1593.880 ;
        RECT 1479.920 1589.880 1480.180 1590.140 ;
        RECT 1479.920 19.760 1480.180 20.020 ;
        RECT 2089.880 19.760 2090.140 20.020 ;
      LAYER met2 ;
        RECT 1088.460 1600.000 1088.740 1604.000 ;
        RECT 1088.520 1593.910 1088.660 1600.000 ;
        RECT 1088.460 1593.590 1088.720 1593.910 ;
        RECT 1479.920 1589.850 1480.180 1590.170 ;
        RECT 1479.980 20.050 1480.120 1589.850 ;
        RECT 1479.920 19.730 1480.180 20.050 ;
        RECT 2089.880 19.730 2090.140 20.050 ;
        RECT 2089.940 2.400 2090.080 19.730 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1095.790 78.440 1096.110 78.500 ;
        RECT 2104.570 78.440 2104.890 78.500 ;
        RECT 1095.790 78.300 2104.890 78.440 ;
        RECT 1095.790 78.240 1096.110 78.300 ;
        RECT 2104.570 78.240 2104.890 78.300 ;
        RECT 2104.570 2.960 2104.890 3.020 ;
        RECT 2107.790 2.960 2108.110 3.020 ;
        RECT 2104.570 2.820 2108.110 2.960 ;
        RECT 2104.570 2.760 2104.890 2.820 ;
        RECT 2107.790 2.760 2108.110 2.820 ;
      LAYER via ;
        RECT 1095.820 78.240 1096.080 78.500 ;
        RECT 2104.600 78.240 2104.860 78.500 ;
        RECT 2104.600 2.760 2104.860 3.020 ;
        RECT 2107.820 2.760 2108.080 3.020 ;
      LAYER met2 ;
        RECT 1095.360 1600.450 1095.640 1604.000 ;
        RECT 1095.360 1600.310 1096.020 1600.450 ;
        RECT 1095.360 1600.000 1095.640 1600.310 ;
        RECT 1095.880 78.530 1096.020 1600.310 ;
        RECT 1095.820 78.210 1096.080 78.530 ;
        RECT 2104.600 78.210 2104.860 78.530 ;
        RECT 2104.660 3.050 2104.800 78.210 ;
        RECT 2104.600 2.730 2104.860 3.050 ;
        RECT 2107.820 2.730 2108.080 3.050 ;
        RECT 2107.880 2.400 2108.020 2.730 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1102.690 68.240 1103.010 68.300 ;
        RECT 2125.270 68.240 2125.590 68.300 ;
        RECT 1102.690 68.100 2125.590 68.240 ;
        RECT 1102.690 68.040 1103.010 68.100 ;
        RECT 2125.270 68.040 2125.590 68.100 ;
      LAYER via ;
        RECT 1102.720 68.040 1102.980 68.300 ;
        RECT 2125.300 68.040 2125.560 68.300 ;
      LAYER met2 ;
        RECT 1102.260 1600.450 1102.540 1604.000 ;
        RECT 1102.260 1600.310 1102.920 1600.450 ;
        RECT 1102.260 1600.000 1102.540 1600.310 ;
        RECT 1102.780 68.330 1102.920 1600.310 ;
        RECT 1102.720 68.010 1102.980 68.330 ;
        RECT 2125.300 68.010 2125.560 68.330 ;
        RECT 2125.360 3.130 2125.500 68.010 ;
        RECT 2125.360 2.990 2125.960 3.130 ;
        RECT 2125.820 2.400 2125.960 2.990 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.510 17.240 1110.830 17.300 ;
        RECT 2143.670 17.240 2143.990 17.300 ;
        RECT 1110.510 17.100 2143.990 17.240 ;
        RECT 1110.510 17.040 1110.830 17.100 ;
        RECT 2143.670 17.040 2143.990 17.100 ;
      LAYER via ;
        RECT 1110.540 17.040 1110.800 17.300 ;
        RECT 2143.700 17.040 2143.960 17.300 ;
      LAYER met2 ;
        RECT 1108.700 1600.450 1108.980 1604.000 ;
        RECT 1108.700 1600.310 1110.740 1600.450 ;
        RECT 1108.700 1600.000 1108.980 1600.310 ;
        RECT 1110.600 17.330 1110.740 1600.310 ;
        RECT 1110.540 17.010 1110.800 17.330 ;
        RECT 2143.700 17.010 2143.960 17.330 ;
        RECT 2143.760 2.400 2143.900 17.010 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1116.490 75.380 1116.810 75.440 ;
        RECT 2159.770 75.380 2160.090 75.440 ;
        RECT 1116.490 75.240 2160.090 75.380 ;
        RECT 1116.490 75.180 1116.810 75.240 ;
        RECT 2159.770 75.180 2160.090 75.240 ;
      LAYER via ;
        RECT 1116.520 75.180 1116.780 75.440 ;
        RECT 2159.800 75.180 2160.060 75.440 ;
      LAYER met2 ;
        RECT 1115.600 1600.450 1115.880 1604.000 ;
        RECT 1115.600 1600.310 1116.720 1600.450 ;
        RECT 1115.600 1600.000 1115.880 1600.310 ;
        RECT 1116.580 75.470 1116.720 1600.310 ;
        RECT 1116.520 75.150 1116.780 75.470 ;
        RECT 2159.800 75.150 2160.060 75.470 ;
        RECT 2159.860 3.130 2160.000 75.150 ;
        RECT 2159.860 2.990 2161.380 3.130 ;
        RECT 2161.240 2.960 2161.380 2.990 ;
        RECT 2161.240 2.820 2161.840 2.960 ;
        RECT 2161.700 2.400 2161.840 2.820 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1145.085 1587.885 1145.255 1589.755 ;
      LAYER mcon ;
        RECT 1145.085 1589.585 1145.255 1589.755 ;
      LAYER met1 ;
        RECT 1145.025 1589.740 1145.315 1589.785 ;
        RECT 1480.350 1589.740 1480.670 1589.800 ;
        RECT 1145.025 1589.600 1480.670 1589.740 ;
        RECT 1145.025 1589.555 1145.315 1589.600 ;
        RECT 1480.350 1589.540 1480.670 1589.600 ;
        RECT 1122.010 1588.040 1122.330 1588.100 ;
        RECT 1145.025 1588.040 1145.315 1588.085 ;
        RECT 1122.010 1587.900 1145.315 1588.040 ;
        RECT 1122.010 1587.840 1122.330 1587.900 ;
        RECT 1145.025 1587.855 1145.315 1587.900 ;
      LAYER via ;
        RECT 1480.380 1589.540 1480.640 1589.800 ;
        RECT 1122.040 1587.840 1122.300 1588.100 ;
      LAYER met2 ;
        RECT 1122.040 1600.000 1122.320 1604.000 ;
        RECT 1122.100 1588.130 1122.240 1600.000 ;
        RECT 1480.380 1589.510 1480.640 1589.830 ;
        RECT 1122.040 1587.810 1122.300 1588.130 ;
        RECT 1480.440 16.165 1480.580 1589.510 ;
        RECT 1480.370 15.795 1480.650 16.165 ;
        RECT 2179.110 15.795 2179.390 16.165 ;
        RECT 2179.180 2.400 2179.320 15.795 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
      LAYER via2 ;
        RECT 1480.370 15.840 1480.650 16.120 ;
        RECT 2179.110 15.840 2179.390 16.120 ;
      LAYER met3 ;
        RECT 1480.345 16.130 1480.675 16.145 ;
        RECT 2179.085 16.130 2179.415 16.145 ;
        RECT 1480.345 15.830 2179.415 16.130 ;
        RECT 1480.345 15.815 1480.675 15.830 ;
        RECT 2179.085 15.815 2179.415 15.830 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1130.290 75.040 1130.610 75.100 ;
        RECT 2194.270 75.040 2194.590 75.100 ;
        RECT 1130.290 74.900 2194.590 75.040 ;
        RECT 1130.290 74.840 1130.610 74.900 ;
        RECT 2194.270 74.840 2194.590 74.900 ;
        RECT 2194.270 2.960 2194.590 3.020 ;
        RECT 2197.030 2.960 2197.350 3.020 ;
        RECT 2194.270 2.820 2197.350 2.960 ;
        RECT 2194.270 2.760 2194.590 2.820 ;
        RECT 2197.030 2.760 2197.350 2.820 ;
      LAYER via ;
        RECT 1130.320 74.840 1130.580 75.100 ;
        RECT 2194.300 74.840 2194.560 75.100 ;
        RECT 2194.300 2.760 2194.560 3.020 ;
        RECT 2197.060 2.760 2197.320 3.020 ;
      LAYER met2 ;
        RECT 1128.940 1600.450 1129.220 1604.000 ;
        RECT 1128.940 1600.310 1130.520 1600.450 ;
        RECT 1128.940 1600.000 1129.220 1600.310 ;
        RECT 1130.380 75.130 1130.520 1600.310 ;
        RECT 1130.320 74.810 1130.580 75.130 ;
        RECT 2194.300 74.810 2194.560 75.130 ;
        RECT 2194.360 3.050 2194.500 74.810 ;
        RECT 2194.300 2.730 2194.560 3.050 ;
        RECT 2197.060 2.730 2197.320 3.050 ;
        RECT 2197.120 2.400 2197.260 2.730 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1137.190 78.780 1137.510 78.840 ;
        RECT 2214.970 78.780 2215.290 78.840 ;
        RECT 1137.190 78.640 2215.290 78.780 ;
        RECT 1137.190 78.580 1137.510 78.640 ;
        RECT 2214.970 78.580 2215.290 78.640 ;
      LAYER via ;
        RECT 1137.220 78.580 1137.480 78.840 ;
        RECT 2215.000 78.580 2215.260 78.840 ;
      LAYER met2 ;
        RECT 1135.840 1600.450 1136.120 1604.000 ;
        RECT 1135.840 1600.310 1137.420 1600.450 ;
        RECT 1135.840 1600.000 1136.120 1600.310 ;
        RECT 1137.280 78.870 1137.420 1600.310 ;
        RECT 1137.220 78.550 1137.480 78.870 ;
        RECT 2215.000 78.550 2215.260 78.870 ;
        RECT 2215.060 2.400 2215.200 78.550 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1144.090 74.700 1144.410 74.760 ;
        RECT 2228.770 74.700 2229.090 74.760 ;
        RECT 1144.090 74.560 2229.090 74.700 ;
        RECT 1144.090 74.500 1144.410 74.560 ;
        RECT 2228.770 74.500 2229.090 74.560 ;
        RECT 2228.770 2.960 2229.090 3.020 ;
        RECT 2232.910 2.960 2233.230 3.020 ;
        RECT 2228.770 2.820 2233.230 2.960 ;
        RECT 2228.770 2.760 2229.090 2.820 ;
        RECT 2232.910 2.760 2233.230 2.820 ;
      LAYER via ;
        RECT 1144.120 74.500 1144.380 74.760 ;
        RECT 2228.800 74.500 2229.060 74.760 ;
        RECT 2228.800 2.760 2229.060 3.020 ;
        RECT 2232.940 2.760 2233.200 3.020 ;
      LAYER met2 ;
        RECT 1142.280 1600.450 1142.560 1604.000 ;
        RECT 1142.280 1600.310 1144.320 1600.450 ;
        RECT 1142.280 1600.000 1142.560 1600.310 ;
        RECT 1144.180 74.790 1144.320 1600.310 ;
        RECT 1144.120 74.470 1144.380 74.790 ;
        RECT 2228.800 74.470 2229.060 74.790 ;
        RECT 2228.860 3.050 2229.000 74.470 ;
        RECT 2228.800 2.730 2229.060 3.050 ;
        RECT 2232.940 2.730 2233.200 3.050 ;
        RECT 2233.000 2.400 2233.140 2.730 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 634.945 1587.205 635.115 1588.395 ;
        RECT 665.305 18.615 665.475 18.955 ;
        RECT 666.225 18.615 666.395 19.635 ;
        RECT 665.305 18.445 666.395 18.615 ;
        RECT 687.385 17.765 687.555 19.635 ;
        RECT 709.005 15.385 709.175 17.935 ;
        RECT 738.445 15.385 738.615 16.235 ;
        RECT 762.365 15.895 762.535 16.235 ;
        RECT 762.365 15.725 764.375 15.895 ;
      LAYER mcon ;
        RECT 634.945 1588.225 635.115 1588.395 ;
        RECT 666.225 19.465 666.395 19.635 ;
        RECT 665.305 18.785 665.475 18.955 ;
        RECT 687.385 19.465 687.555 19.635 ;
        RECT 709.005 17.765 709.175 17.935 ;
        RECT 738.445 16.065 738.615 16.235 ;
        RECT 762.365 16.065 762.535 16.235 ;
        RECT 764.205 15.725 764.375 15.895 ;
      LAYER met1 ;
        RECT 597.150 1588.380 597.470 1588.440 ;
        RECT 634.885 1588.380 635.175 1588.425 ;
        RECT 597.150 1588.240 635.175 1588.380 ;
        RECT 597.150 1588.180 597.470 1588.240 ;
        RECT 634.885 1588.195 635.175 1588.240 ;
        RECT 651.890 1587.700 652.210 1587.760 ;
        RECT 643.700 1587.560 652.210 1587.700 ;
        RECT 634.885 1587.360 635.175 1587.405 ;
        RECT 643.700 1587.360 643.840 1587.560 ;
        RECT 651.890 1587.500 652.210 1587.560 ;
        RECT 634.885 1587.220 643.840 1587.360 ;
        RECT 634.885 1587.175 635.175 1587.220 ;
        RECT 666.165 19.620 666.455 19.665 ;
        RECT 687.325 19.620 687.615 19.665 ;
        RECT 666.165 19.480 687.615 19.620 ;
        RECT 666.165 19.435 666.455 19.480 ;
        RECT 687.325 19.435 687.615 19.480 ;
        RECT 665.245 18.940 665.535 18.985 ;
        RECT 657.500 18.800 665.535 18.940 ;
        RECT 651.890 18.260 652.210 18.320 ;
        RECT 657.500 18.260 657.640 18.800 ;
        RECT 665.245 18.755 665.535 18.800 ;
        RECT 651.890 18.120 657.640 18.260 ;
        RECT 651.890 18.060 652.210 18.120 ;
        RECT 687.325 17.920 687.615 17.965 ;
        RECT 708.945 17.920 709.235 17.965 ;
        RECT 687.325 17.780 709.235 17.920 ;
        RECT 687.325 17.735 687.615 17.780 ;
        RECT 708.945 17.735 709.235 17.780 ;
        RECT 738.385 16.220 738.675 16.265 ;
        RECT 762.305 16.220 762.595 16.265 ;
        RECT 738.385 16.080 762.595 16.220 ;
        RECT 738.385 16.035 738.675 16.080 ;
        RECT 762.305 16.035 762.595 16.080 ;
        RECT 764.145 15.880 764.435 15.925 ;
        RECT 787.590 15.880 787.910 15.940 ;
        RECT 764.145 15.740 787.910 15.880 ;
        RECT 764.145 15.695 764.435 15.740 ;
        RECT 787.590 15.680 787.910 15.740 ;
        RECT 708.945 15.540 709.235 15.585 ;
        RECT 738.385 15.540 738.675 15.585 ;
        RECT 708.945 15.400 738.675 15.540 ;
        RECT 708.945 15.355 709.235 15.400 ;
        RECT 738.385 15.355 738.675 15.400 ;
      LAYER via ;
        RECT 597.180 1588.180 597.440 1588.440 ;
        RECT 651.920 1587.500 652.180 1587.760 ;
        RECT 651.920 18.060 652.180 18.320 ;
        RECT 787.620 15.680 787.880 15.940 ;
      LAYER met2 ;
        RECT 597.180 1600.000 597.460 1604.000 ;
        RECT 597.240 1588.470 597.380 1600.000 ;
        RECT 597.180 1588.150 597.440 1588.470 ;
        RECT 651.920 1587.470 652.180 1587.790 ;
        RECT 651.980 18.350 652.120 1587.470 ;
        RECT 651.920 18.030 652.180 18.350 ;
        RECT 787.620 15.650 787.880 15.970 ;
        RECT 787.680 2.400 787.820 15.650 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1149.150 1587.700 1149.470 1587.760 ;
        RECT 1151.910 1587.700 1152.230 1587.760 ;
        RECT 1149.150 1587.560 1152.230 1587.700 ;
        RECT 1149.150 1587.500 1149.470 1587.560 ;
        RECT 1151.910 1587.500 1152.230 1587.560 ;
      LAYER via ;
        RECT 1149.180 1587.500 1149.440 1587.760 ;
        RECT 1151.940 1587.500 1152.200 1587.760 ;
      LAYER met2 ;
        RECT 1149.180 1600.000 1149.460 1604.000 ;
        RECT 1149.240 1587.790 1149.380 1600.000 ;
        RECT 1149.180 1587.470 1149.440 1587.790 ;
        RECT 1151.940 1587.470 1152.200 1587.790 ;
        RECT 1152.000 20.245 1152.140 1587.470 ;
        RECT 1151.930 19.875 1152.210 20.245 ;
        RECT 2250.870 19.875 2251.150 20.245 ;
        RECT 2250.940 2.400 2251.080 19.875 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
      LAYER via2 ;
        RECT 1151.930 19.920 1152.210 20.200 ;
        RECT 2250.870 19.920 2251.150 20.200 ;
      LAYER met3 ;
        RECT 1151.905 20.210 1152.235 20.225 ;
        RECT 2250.845 20.210 2251.175 20.225 ;
        RECT 1151.905 19.910 2251.175 20.210 ;
        RECT 1151.905 19.895 1152.235 19.910 ;
        RECT 2250.845 19.895 2251.175 19.910 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1157.890 74.360 1158.210 74.420 ;
        RECT 2263.270 74.360 2263.590 74.420 ;
        RECT 1157.890 74.220 2263.590 74.360 ;
        RECT 1157.890 74.160 1158.210 74.220 ;
        RECT 2263.270 74.160 2263.590 74.220 ;
        RECT 2263.270 2.960 2263.590 3.020 ;
        RECT 2268.330 2.960 2268.650 3.020 ;
        RECT 2263.270 2.820 2268.650 2.960 ;
        RECT 2263.270 2.760 2263.590 2.820 ;
        RECT 2268.330 2.760 2268.650 2.820 ;
      LAYER via ;
        RECT 1157.920 74.160 1158.180 74.420 ;
        RECT 2263.300 74.160 2263.560 74.420 ;
        RECT 2263.300 2.760 2263.560 3.020 ;
        RECT 2268.360 2.760 2268.620 3.020 ;
      LAYER met2 ;
        RECT 1156.080 1600.450 1156.360 1604.000 ;
        RECT 1156.080 1600.310 1158.120 1600.450 ;
        RECT 1156.080 1600.000 1156.360 1600.310 ;
        RECT 1157.980 74.450 1158.120 1600.310 ;
        RECT 1157.920 74.130 1158.180 74.450 ;
        RECT 2263.300 74.130 2263.560 74.450 ;
        RECT 2263.360 3.050 2263.500 74.130 ;
        RECT 2263.300 2.730 2263.560 3.050 ;
        RECT 2268.360 2.730 2268.620 3.050 ;
        RECT 2268.420 2.400 2268.560 2.730 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.490 1587.700 1162.810 1587.760 ;
        RECT 1165.710 1587.700 1166.030 1587.760 ;
        RECT 1162.490 1587.560 1166.030 1587.700 ;
        RECT 1162.490 1587.500 1162.810 1587.560 ;
        RECT 1165.710 1587.500 1166.030 1587.560 ;
      LAYER via ;
        RECT 1162.520 1587.500 1162.780 1587.760 ;
        RECT 1165.740 1587.500 1166.000 1587.760 ;
      LAYER met2 ;
        RECT 1162.520 1600.000 1162.800 1604.000 ;
        RECT 1162.580 1587.790 1162.720 1600.000 ;
        RECT 1162.520 1587.470 1162.780 1587.790 ;
        RECT 1165.740 1587.470 1166.000 1587.790 ;
        RECT 1165.800 19.565 1165.940 1587.470 ;
        RECT 1165.730 19.195 1166.010 19.565 ;
        RECT 2286.290 19.195 2286.570 19.565 ;
        RECT 2286.360 2.400 2286.500 19.195 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
      LAYER via2 ;
        RECT 1165.730 19.240 1166.010 19.520 ;
        RECT 2286.290 19.240 2286.570 19.520 ;
      LAYER met3 ;
        RECT 1165.705 19.530 1166.035 19.545 ;
        RECT 2286.265 19.530 2286.595 19.545 ;
        RECT 1165.705 19.230 2286.595 19.530 ;
        RECT 1165.705 19.215 1166.035 19.230 ;
        RECT 2286.265 19.215 2286.595 19.230 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1171.690 74.020 1172.010 74.080 ;
        RECT 2297.770 74.020 2298.090 74.080 ;
        RECT 1171.690 73.880 2298.090 74.020 ;
        RECT 1171.690 73.820 1172.010 73.880 ;
        RECT 2297.770 73.820 2298.090 73.880 ;
        RECT 2297.770 17.580 2298.090 17.640 ;
        RECT 2304.210 17.580 2304.530 17.640 ;
        RECT 2297.770 17.440 2304.530 17.580 ;
        RECT 2297.770 17.380 2298.090 17.440 ;
        RECT 2304.210 17.380 2304.530 17.440 ;
      LAYER via ;
        RECT 1171.720 73.820 1171.980 74.080 ;
        RECT 2297.800 73.820 2298.060 74.080 ;
        RECT 2297.800 17.380 2298.060 17.640 ;
        RECT 2304.240 17.380 2304.500 17.640 ;
      LAYER met2 ;
        RECT 1169.420 1601.130 1169.700 1604.000 ;
        RECT 1169.420 1600.990 1171.460 1601.130 ;
        RECT 1169.420 1600.000 1169.700 1600.990 ;
        RECT 1171.320 1590.250 1171.460 1600.990 ;
        RECT 1171.320 1590.110 1171.920 1590.250 ;
        RECT 1171.780 74.110 1171.920 1590.110 ;
        RECT 1171.720 73.790 1171.980 74.110 ;
        RECT 2297.800 73.790 2298.060 74.110 ;
        RECT 2297.860 17.670 2298.000 73.790 ;
        RECT 2297.800 17.350 2298.060 17.670 ;
        RECT 2304.240 17.350 2304.500 17.670 ;
        RECT 2304.300 2.400 2304.440 17.350 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1176.290 1587.700 1176.610 1587.760 ;
        RECT 1179.510 1587.700 1179.830 1587.760 ;
        RECT 1176.290 1587.560 1179.830 1587.700 ;
        RECT 1176.290 1587.500 1176.610 1587.560 ;
        RECT 1179.510 1587.500 1179.830 1587.560 ;
      LAYER via ;
        RECT 1176.320 1587.500 1176.580 1587.760 ;
        RECT 1179.540 1587.500 1179.800 1587.760 ;
      LAYER met2 ;
        RECT 1176.320 1600.000 1176.600 1604.000 ;
        RECT 1176.380 1587.790 1176.520 1600.000 ;
        RECT 1176.320 1587.470 1176.580 1587.790 ;
        RECT 1179.540 1587.470 1179.800 1587.790 ;
        RECT 1179.600 18.885 1179.740 1587.470 ;
        RECT 1179.530 18.515 1179.810 18.885 ;
        RECT 2322.170 18.515 2322.450 18.885 ;
        RECT 2322.240 2.400 2322.380 18.515 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
      LAYER via2 ;
        RECT 1179.530 18.560 1179.810 18.840 ;
        RECT 2322.170 18.560 2322.450 18.840 ;
      LAYER met3 ;
        RECT 1179.505 18.850 1179.835 18.865 ;
        RECT 2322.145 18.850 2322.475 18.865 ;
        RECT 1179.505 18.550 2322.475 18.850 ;
        RECT 1179.505 18.535 1179.835 18.550 ;
        RECT 2322.145 18.535 2322.475 18.550 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1182.730 1587.700 1183.050 1587.760 ;
        RECT 1185.490 1587.700 1185.810 1587.760 ;
        RECT 1182.730 1587.560 1185.810 1587.700 ;
        RECT 1182.730 1587.500 1183.050 1587.560 ;
        RECT 1185.490 1587.500 1185.810 1587.560 ;
        RECT 1185.490 73.680 1185.810 73.740 ;
        RECT 2339.170 73.680 2339.490 73.740 ;
        RECT 1185.490 73.540 2339.490 73.680 ;
        RECT 1185.490 73.480 1185.810 73.540 ;
        RECT 2339.170 73.480 2339.490 73.540 ;
      LAYER via ;
        RECT 1182.760 1587.500 1183.020 1587.760 ;
        RECT 1185.520 1587.500 1185.780 1587.760 ;
        RECT 1185.520 73.480 1185.780 73.740 ;
        RECT 2339.200 73.480 2339.460 73.740 ;
      LAYER met2 ;
        RECT 1182.760 1600.000 1183.040 1604.000 ;
        RECT 1182.820 1587.790 1182.960 1600.000 ;
        RECT 1182.760 1587.470 1183.020 1587.790 ;
        RECT 1185.520 1587.470 1185.780 1587.790 ;
        RECT 1185.580 73.770 1185.720 1587.470 ;
        RECT 1185.520 73.450 1185.780 73.770 ;
        RECT 2339.200 73.450 2339.460 73.770 ;
        RECT 2339.260 3.130 2339.400 73.450 ;
        RECT 2339.260 2.990 2339.860 3.130 ;
        RECT 2339.720 2.400 2339.860 2.990 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1189.630 1587.700 1189.950 1587.760 ;
        RECT 1193.310 1587.700 1193.630 1587.760 ;
        RECT 1189.630 1587.560 1193.630 1587.700 ;
        RECT 1189.630 1587.500 1189.950 1587.560 ;
        RECT 1193.310 1587.500 1193.630 1587.560 ;
      LAYER via ;
        RECT 1189.660 1587.500 1189.920 1587.760 ;
        RECT 1193.340 1587.500 1193.600 1587.760 ;
      LAYER met2 ;
        RECT 1189.660 1600.000 1189.940 1604.000 ;
        RECT 1189.720 1587.790 1189.860 1600.000 ;
        RECT 1189.660 1587.470 1189.920 1587.790 ;
        RECT 1193.340 1587.470 1193.600 1587.790 ;
        RECT 1193.400 18.205 1193.540 1587.470 ;
        RECT 1193.330 17.835 1193.610 18.205 ;
        RECT 2357.590 17.835 2357.870 18.205 ;
        RECT 2357.660 2.400 2357.800 17.835 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
      LAYER via2 ;
        RECT 1193.330 17.880 1193.610 18.160 ;
        RECT 2357.590 17.880 2357.870 18.160 ;
      LAYER met3 ;
        RECT 1193.305 18.170 1193.635 18.185 ;
        RECT 2357.565 18.170 2357.895 18.185 ;
        RECT 1193.305 17.870 2357.895 18.170 ;
        RECT 1193.305 17.855 1193.635 17.870 ;
        RECT 2357.565 17.855 2357.895 17.870 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1196.070 1587.700 1196.390 1587.760 ;
        RECT 1199.290 1587.700 1199.610 1587.760 ;
        RECT 1196.070 1587.560 1199.610 1587.700 ;
        RECT 1196.070 1587.500 1196.390 1587.560 ;
        RECT 1199.290 1587.500 1199.610 1587.560 ;
        RECT 1199.290 73.340 1199.610 73.400 ;
        RECT 2373.670 73.340 2373.990 73.400 ;
        RECT 1199.290 73.200 2373.990 73.340 ;
        RECT 1199.290 73.140 1199.610 73.200 ;
        RECT 2373.670 73.140 2373.990 73.200 ;
      LAYER via ;
        RECT 1196.100 1587.500 1196.360 1587.760 ;
        RECT 1199.320 1587.500 1199.580 1587.760 ;
        RECT 1199.320 73.140 1199.580 73.400 ;
        RECT 2373.700 73.140 2373.960 73.400 ;
      LAYER met2 ;
        RECT 1196.100 1600.000 1196.380 1604.000 ;
        RECT 1196.160 1587.790 1196.300 1600.000 ;
        RECT 1196.100 1587.470 1196.360 1587.790 ;
        RECT 1199.320 1587.470 1199.580 1587.790 ;
        RECT 1199.380 73.430 1199.520 1587.470 ;
        RECT 1199.320 73.110 1199.580 73.430 ;
        RECT 2373.700 73.110 2373.960 73.430 ;
        RECT 2373.760 3.130 2373.900 73.110 ;
        RECT 2373.760 2.990 2375.280 3.130 ;
        RECT 2375.140 2.960 2375.280 2.990 ;
        RECT 2375.140 2.820 2375.740 2.960 ;
        RECT 2375.600 2.400 2375.740 2.820 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1202.970 1587.700 1203.290 1587.760 ;
        RECT 1207.110 1587.700 1207.430 1587.760 ;
        RECT 1202.970 1587.560 1207.430 1587.700 ;
        RECT 1202.970 1587.500 1203.290 1587.560 ;
        RECT 1207.110 1587.500 1207.430 1587.560 ;
      LAYER via ;
        RECT 1203.000 1587.500 1203.260 1587.760 ;
        RECT 1207.140 1587.500 1207.400 1587.760 ;
      LAYER met2 ;
        RECT 1203.000 1600.000 1203.280 1604.000 ;
        RECT 1203.060 1587.790 1203.200 1600.000 ;
        RECT 1203.000 1587.470 1203.260 1587.790 ;
        RECT 1207.140 1587.470 1207.400 1587.790 ;
        RECT 1207.200 17.525 1207.340 1587.470 ;
        RECT 1207.130 17.155 1207.410 17.525 ;
        RECT 2393.470 17.155 2393.750 17.525 ;
        RECT 2393.540 2.400 2393.680 17.155 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
      LAYER via2 ;
        RECT 1207.130 17.200 1207.410 17.480 ;
        RECT 2393.470 17.200 2393.750 17.480 ;
      LAYER met3 ;
        RECT 1207.105 17.490 1207.435 17.505 ;
        RECT 2393.445 17.490 2393.775 17.505 ;
        RECT 1207.105 17.190 2393.775 17.490 ;
        RECT 1207.105 17.175 1207.435 17.190 ;
        RECT 2393.445 17.175 2393.775 17.190 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1209.870 1588.040 1210.190 1588.100 ;
        RECT 1213.090 1588.040 1213.410 1588.100 ;
        RECT 1209.870 1587.900 1213.410 1588.040 ;
        RECT 1209.870 1587.840 1210.190 1587.900 ;
        RECT 1213.090 1587.840 1213.410 1587.900 ;
        RECT 1213.090 73.000 1213.410 73.060 ;
        RECT 2408.170 73.000 2408.490 73.060 ;
        RECT 1213.090 72.860 2408.490 73.000 ;
        RECT 1213.090 72.800 1213.410 72.860 ;
        RECT 2408.170 72.800 2408.490 72.860 ;
      LAYER via ;
        RECT 1209.900 1587.840 1210.160 1588.100 ;
        RECT 1213.120 1587.840 1213.380 1588.100 ;
        RECT 1213.120 72.800 1213.380 73.060 ;
        RECT 2408.200 72.800 2408.460 73.060 ;
      LAYER met2 ;
        RECT 1209.900 1600.000 1210.180 1604.000 ;
        RECT 1209.960 1588.130 1210.100 1600.000 ;
        RECT 1209.900 1587.810 1210.160 1588.130 ;
        RECT 1213.120 1587.810 1213.380 1588.130 ;
        RECT 1213.180 73.090 1213.320 1587.810 ;
        RECT 1213.120 72.770 1213.380 73.090 ;
        RECT 2408.200 72.770 2408.460 73.090 ;
        RECT 2408.260 17.410 2408.400 72.770 ;
        RECT 2408.260 17.270 2411.620 17.410 ;
        RECT 2411.480 2.400 2411.620 17.270 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 763.285 1588.225 763.455 1590.435 ;
      LAYER mcon ;
        RECT 763.285 1590.265 763.455 1590.435 ;
      LAYER met1 ;
        RECT 603.590 1590.420 603.910 1590.480 ;
        RECT 763.225 1590.420 763.515 1590.465 ;
        RECT 603.590 1590.280 763.515 1590.420 ;
        RECT 603.590 1590.220 603.910 1590.280 ;
        RECT 763.225 1590.235 763.515 1590.280 ;
        RECT 801.850 1588.720 802.170 1588.780 ;
        RECT 797.800 1588.580 802.170 1588.720 ;
        RECT 763.225 1588.380 763.515 1588.425 ;
        RECT 797.800 1588.380 797.940 1588.580 ;
        RECT 801.850 1588.520 802.170 1588.580 ;
        RECT 763.225 1588.240 797.940 1588.380 ;
        RECT 763.225 1588.195 763.515 1588.240 ;
        RECT 801.850 62.120 802.170 62.180 ;
        RECT 805.530 62.120 805.850 62.180 ;
        RECT 801.850 61.980 805.850 62.120 ;
        RECT 801.850 61.920 802.170 61.980 ;
        RECT 805.530 61.920 805.850 61.980 ;
      LAYER via ;
        RECT 603.620 1590.220 603.880 1590.480 ;
        RECT 801.880 1588.520 802.140 1588.780 ;
        RECT 801.880 61.920 802.140 62.180 ;
        RECT 805.560 61.920 805.820 62.180 ;
      LAYER met2 ;
        RECT 603.620 1600.000 603.900 1604.000 ;
        RECT 603.680 1590.510 603.820 1600.000 ;
        RECT 603.620 1590.190 603.880 1590.510 ;
        RECT 801.880 1588.490 802.140 1588.810 ;
        RECT 801.940 62.210 802.080 1588.490 ;
        RECT 801.880 61.890 802.140 62.210 ;
        RECT 805.560 61.890 805.820 62.210 ;
        RECT 805.620 2.400 805.760 61.890 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1159.345 2791.145 1160.435 2791.315 ;
        RECT 1604.165 2791.145 1604.335 2792.675 ;
        RECT 303.745 1590.945 304.835 1591.115 ;
        RECT 303.745 1590.435 303.915 1590.945 ;
        RECT 303.285 1590.265 303.915 1590.435 ;
      LAYER mcon ;
        RECT 1604.165 2792.505 1604.335 2792.675 ;
        RECT 1160.265 2791.145 1160.435 2791.315 ;
        RECT 304.665 1590.945 304.835 1591.115 ;
      LAYER met1 ;
        RECT 1604.105 2792.660 1604.395 2792.705 ;
        RECT 1917.810 2792.660 1918.130 2792.720 ;
        RECT 2215.430 2792.660 2215.750 2792.720 ;
        RECT 1604.105 2792.520 2215.750 2792.660 ;
        RECT 1604.105 2792.475 1604.395 2792.520 ;
        RECT 1917.810 2792.460 1918.130 2792.520 ;
        RECT 2215.430 2792.460 2215.750 2792.520 ;
        RECT 972.050 2791.300 972.370 2791.360 ;
        RECT 1159.285 2791.300 1159.575 2791.345 ;
        RECT 972.050 2791.160 1159.575 2791.300 ;
        RECT 972.050 2791.100 972.370 2791.160 ;
        RECT 1159.285 2791.115 1159.575 2791.160 ;
        RECT 1160.205 2791.300 1160.495 2791.345 ;
        RECT 1568.670 2791.300 1568.990 2791.360 ;
        RECT 1604.105 2791.300 1604.395 2791.345 ;
        RECT 1160.205 2791.160 1604.395 2791.300 ;
        RECT 1160.205 2791.115 1160.495 2791.160 ;
        RECT 1568.670 2791.100 1568.990 2791.160 ;
        RECT 1604.105 2791.115 1604.395 2791.160 ;
        RECT 1917.810 2066.420 1918.130 2066.480 ;
        RECT 2024.990 2066.420 2025.310 2066.480 ;
        RECT 1917.810 2066.280 2025.310 2066.420 ;
        RECT 1917.810 2066.220 1918.130 2066.280 ;
        RECT 2024.990 2066.220 2025.310 2066.280 ;
        RECT 2024.990 2063.360 2025.310 2063.420 ;
        RECT 2566.870 2063.360 2567.190 2063.420 ;
        RECT 2024.990 2063.220 2567.190 2063.360 ;
        RECT 2024.990 2063.160 2025.310 2063.220 ;
        RECT 2566.870 2063.160 2567.190 2063.220 ;
        RECT 1566.370 1593.820 1566.690 1593.880 ;
        RECT 2024.990 1593.820 2025.310 1593.880 ;
        RECT 2215.430 1593.820 2215.750 1593.880 ;
        RECT 1566.370 1593.680 2215.750 1593.820 ;
        RECT 1566.370 1593.620 1566.690 1593.680 ;
        RECT 2024.990 1593.620 2025.310 1593.680 ;
        RECT 2215.430 1593.620 2215.750 1593.680 ;
        RECT 304.605 1591.100 304.895 1591.145 ;
        RECT 1566.370 1591.100 1566.690 1591.160 ;
        RECT 304.605 1590.960 1566.690 1591.100 ;
        RECT 304.605 1590.915 304.895 1590.960 ;
        RECT 1566.370 1590.900 1566.690 1590.960 ;
        RECT 301.830 1590.420 302.150 1590.480 ;
        RECT 303.225 1590.420 303.515 1590.465 ;
        RECT 301.830 1590.280 303.515 1590.420 ;
        RECT 301.830 1590.220 302.150 1590.280 ;
        RECT 303.225 1590.235 303.515 1590.280 ;
        RECT 2.830 17.240 3.150 17.300 ;
        RECT 299.530 17.240 299.850 17.300 ;
        RECT 2.830 17.100 299.850 17.240 ;
        RECT 2.830 17.040 3.150 17.100 ;
        RECT 299.530 17.040 299.850 17.100 ;
      LAYER via ;
        RECT 1917.840 2792.460 1918.100 2792.720 ;
        RECT 2215.460 2792.460 2215.720 2792.720 ;
        RECT 972.080 2791.100 972.340 2791.360 ;
        RECT 1568.700 2791.100 1568.960 2791.360 ;
        RECT 1917.840 2066.220 1918.100 2066.480 ;
        RECT 2025.020 2066.220 2025.280 2066.480 ;
        RECT 2025.020 2063.160 2025.280 2063.420 ;
        RECT 2566.900 2063.160 2567.160 2063.420 ;
        RECT 1566.400 1593.620 1566.660 1593.880 ;
        RECT 2025.020 1593.620 2025.280 1593.880 ;
        RECT 2215.460 1593.620 2215.720 1593.880 ;
        RECT 1566.400 1590.900 1566.660 1591.160 ;
        RECT 301.860 1590.220 302.120 1590.480 ;
        RECT 2.860 17.040 3.120 17.300 ;
        RECT 299.560 17.040 299.820 17.300 ;
      LAYER met2 ;
        RECT 972.070 2794.275 972.350 2794.645 ;
        RECT 1568.690 2794.275 1568.970 2794.645 ;
        RECT 2215.450 2794.275 2215.730 2794.645 ;
        RECT 972.140 2791.390 972.280 2794.275 ;
        RECT 1568.760 2791.390 1568.900 2794.275 ;
        RECT 2215.520 2792.750 2215.660 2794.275 ;
        RECT 1917.840 2792.430 1918.100 2792.750 ;
        RECT 2215.460 2792.430 2215.720 2792.750 ;
        RECT 972.080 2791.070 972.340 2791.390 ;
        RECT 1568.700 2791.070 1568.960 2791.390 ;
        RECT 972.140 2790.565 972.280 2791.070 ;
        RECT 972.070 2790.195 972.350 2790.565 ;
        RECT 1917.900 2066.510 1918.040 2792.430 ;
        RECT 1917.840 2066.365 1918.100 2066.510 ;
        RECT 1917.830 2065.995 1918.110 2066.365 ;
        RECT 2025.020 2066.190 2025.280 2066.510 ;
        RECT 2025.080 2063.450 2025.220 2066.190 ;
        RECT 2025.020 2063.130 2025.280 2063.450 ;
        RECT 2566.890 2063.275 2567.170 2063.645 ;
        RECT 2566.900 2063.130 2567.160 2063.275 ;
        RECT 300.940 1600.450 301.220 1604.000 ;
        RECT 300.080 1600.310 301.220 1600.450 ;
        RECT 300.080 1589.570 300.220 1600.310 ;
        RECT 300.940 1600.000 301.220 1600.310 ;
        RECT 2025.080 1593.910 2025.220 2063.130 ;
        RECT 1566.400 1593.765 1566.660 1593.910 ;
        RECT 1566.390 1593.395 1566.670 1593.765 ;
        RECT 2025.020 1593.590 2025.280 1593.910 ;
        RECT 2215.460 1593.765 2215.720 1593.910 ;
        RECT 2215.450 1593.395 2215.730 1593.765 ;
        RECT 1566.460 1591.190 1566.600 1593.395 ;
        RECT 1566.400 1590.870 1566.660 1591.190 ;
        RECT 301.860 1590.190 302.120 1590.510 ;
        RECT 301.920 1589.570 302.060 1590.190 ;
        RECT 300.080 1589.430 302.060 1589.570 ;
        RECT 300.080 18.090 300.220 1589.430 ;
        RECT 299.620 17.950 300.220 18.090 ;
        RECT 299.620 17.330 299.760 17.950 ;
        RECT 2.860 17.010 3.120 17.330 ;
        RECT 299.560 17.010 299.820 17.330 ;
        RECT 2.920 2.400 3.060 17.010 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 972.070 2794.320 972.350 2794.600 ;
        RECT 1568.690 2794.320 1568.970 2794.600 ;
        RECT 2215.450 2794.320 2215.730 2794.600 ;
        RECT 972.070 2790.240 972.350 2790.520 ;
        RECT 1917.830 2066.040 1918.110 2066.320 ;
        RECT 2566.890 2063.320 2567.170 2063.600 ;
        RECT 1566.390 1593.440 1566.670 1593.720 ;
        RECT 2215.450 1593.440 2215.730 1593.720 ;
      LAYER met3 ;
        RECT 972.045 2794.620 972.375 2794.625 ;
        RECT 971.790 2794.610 972.375 2794.620 ;
        RECT 971.590 2794.310 972.375 2794.610 ;
        RECT 971.790 2794.300 972.375 2794.310 ;
        RECT 972.045 2794.295 972.375 2794.300 ;
        RECT 1568.665 2794.620 1568.995 2794.625 ;
        RECT 2215.425 2794.620 2215.755 2794.625 ;
        RECT 1568.665 2794.610 1569.250 2794.620 ;
        RECT 2215.425 2794.610 2216.010 2794.620 ;
        RECT 1568.665 2794.310 1569.450 2794.610 ;
        RECT 2215.425 2794.310 2216.210 2794.610 ;
        RECT 1568.665 2794.300 1569.250 2794.310 ;
        RECT 2215.425 2794.300 2216.010 2794.310 ;
        RECT 1568.665 2794.295 1568.995 2794.300 ;
        RECT 2215.425 2794.295 2215.755 2794.300 ;
        RECT 321.350 2790.530 321.730 2790.540 ;
        RECT 972.045 2790.530 972.375 2790.545 ;
        RECT 321.350 2790.230 972.375 2790.530 ;
        RECT 321.350 2790.220 321.730 2790.230 ;
        RECT 972.045 2790.215 972.375 2790.230 ;
        RECT 1917.805 2066.340 1918.135 2066.345 ;
        RECT 1917.550 2066.330 1918.135 2066.340 ;
        RECT 1917.350 2066.030 1918.135 2066.330 ;
        RECT 1917.550 2066.020 1918.135 2066.030 ;
        RECT 1917.805 2066.015 1918.135 2066.020 ;
        RECT 2566.865 2063.620 2567.195 2063.625 ;
        RECT 2566.865 2063.610 2567.450 2063.620 ;
        RECT 2566.640 2063.310 2567.450 2063.610 ;
        RECT 2566.865 2063.300 2567.450 2063.310 ;
        RECT 2566.865 2063.295 2567.195 2063.300 ;
        RECT 1566.365 1593.730 1566.695 1593.745 ;
        RECT 2215.425 1593.740 2215.755 1593.745 ;
        RECT 1567.030 1593.730 1567.410 1593.740 ;
        RECT 1566.365 1593.430 1567.410 1593.730 ;
        RECT 1566.365 1593.415 1566.695 1593.430 ;
        RECT 1567.030 1593.420 1567.410 1593.430 ;
        RECT 2215.425 1593.730 2216.010 1593.740 ;
        RECT 2215.425 1593.430 2216.210 1593.730 ;
        RECT 2215.425 1593.420 2216.010 1593.430 ;
        RECT 2215.425 1593.415 2215.755 1593.420 ;
      LAYER via3 ;
        RECT 971.820 2794.300 972.140 2794.620 ;
        RECT 1568.900 2794.300 1569.220 2794.620 ;
        RECT 2215.660 2794.300 2215.980 2794.620 ;
        RECT 321.380 2790.220 321.700 2790.540 ;
        RECT 1917.580 2066.020 1917.900 2066.340 ;
        RECT 2567.100 2063.300 2567.420 2063.620 ;
        RECT 1567.060 1593.420 1567.380 1593.740 ;
        RECT 2215.660 1593.420 2215.980 1593.740 ;
      LAYER met4 ;
        RECT 319.015 2801.750 319.315 2804.600 ;
        RECT 969.015 2801.750 969.315 2804.600 ;
        RECT 1569.015 2801.750 1569.315 2804.600 ;
        RECT 2219.015 2801.750 2219.315 2804.600 ;
        RECT 319.015 2801.450 321.690 2801.750 ;
        RECT 319.015 2800.000 319.315 2801.450 ;
        RECT 321.390 2790.545 321.690 2801.450 ;
        RECT 969.015 2801.450 972.130 2801.750 ;
        RECT 969.015 2800.000 969.315 2801.450 ;
        RECT 971.830 2794.625 972.130 2801.450 ;
        RECT 1568.910 2800.000 1569.315 2801.750 ;
        RECT 2215.670 2801.450 2219.315 2801.750 ;
        RECT 1568.910 2794.625 1569.210 2800.000 ;
        RECT 2215.670 2794.625 2215.970 2801.450 ;
        RECT 2219.015 2800.000 2219.315 2801.450 ;
        RECT 971.815 2794.295 972.145 2794.625 ;
        RECT 1568.895 2794.295 1569.225 2794.625 ;
        RECT 2215.655 2794.295 2215.985 2794.625 ;
        RECT 321.375 2790.215 321.705 2790.545 ;
        RECT 1917.575 2066.015 1917.905 2066.345 ;
        RECT 1917.590 2058.850 1917.890 2066.015 ;
        RECT 2567.095 2063.295 2567.425 2063.625 ;
        RECT 1917.165 2058.550 1917.890 2058.850 ;
        RECT 1917.165 2051.635 1917.465 2058.550 ;
        RECT 2567.110 2055.450 2567.410 2063.295 ;
        RECT 2567.865 2055.450 2568.165 2056.235 ;
        RECT 2567.110 2055.150 2568.165 2055.450 ;
        RECT 2567.865 2051.635 2568.165 2055.150 ;
        RECT 1568.315 1601.550 1568.615 1604.600 ;
        RECT 2219.015 1601.550 2219.315 1604.600 ;
        RECT 1567.070 1601.250 1568.615 1601.550 ;
        RECT 1567.070 1593.745 1567.370 1601.250 ;
        RECT 1568.315 1600.000 1568.615 1601.250 ;
        RECT 2215.670 1601.250 2219.315 1601.550 ;
        RECT 2215.670 1593.745 2215.970 1601.250 ;
        RECT 2219.015 1600.000 2219.315 1601.250 ;
        RECT 1567.055 1593.415 1567.385 1593.745 ;
        RECT 2215.655 1593.415 2215.985 1593.745 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 296.770 1594.840 297.090 1594.900 ;
        RECT 301.370 1594.840 301.690 1594.900 ;
        RECT 296.770 1594.700 301.690 1594.840 ;
        RECT 296.770 1594.640 297.090 1594.700 ;
        RECT 301.370 1594.640 301.690 1594.700 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 296.770 17.580 297.090 17.640 ;
        RECT 8.350 17.440 297.090 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 296.770 17.380 297.090 17.440 ;
      LAYER via ;
        RECT 296.800 1594.640 297.060 1594.900 ;
        RECT 301.400 1594.640 301.660 1594.900 ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 296.800 17.380 297.060 17.640 ;
      LAYER met2 ;
        RECT 302.780 1600.450 303.060 1604.000 ;
        RECT 301.460 1600.310 303.060 1600.450 ;
        RECT 301.460 1594.930 301.600 1600.310 ;
        RECT 302.780 1600.000 303.060 1600.310 ;
        RECT 296.800 1594.610 297.060 1594.930 ;
        RECT 301.400 1594.610 301.660 1594.930 ;
        RECT 296.860 17.670 297.000 1594.610 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 296.800 17.350 297.060 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.080 1600.450 305.360 1604.000 ;
        RECT 304.220 1600.310 305.360 1600.450 ;
        RECT 304.220 16.845 304.360 1600.310 ;
        RECT 305.080 1600.000 305.360 1600.310 ;
        RECT 14.350 16.475 14.630 16.845 ;
        RECT 304.150 16.475 304.430 16.845 ;
        RECT 14.420 2.400 14.560 16.475 ;
        RECT 14.210 -4.800 14.770 2.400 ;
      LAYER via2 ;
        RECT 14.350 16.520 14.630 16.800 ;
        RECT 304.150 16.520 304.430 16.800 ;
      LAYER met3 ;
        RECT 14.325 16.810 14.655 16.825 ;
        RECT 304.125 16.810 304.455 16.825 ;
        RECT 14.325 16.510 304.455 16.810 ;
        RECT 14.325 16.495 14.655 16.510 ;
        RECT 304.125 16.495 304.455 16.510 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 18.260 38.570 18.320 ;
        RECT 311.030 18.260 311.350 18.320 ;
        RECT 38.250 18.120 311.350 18.260 ;
        RECT 38.250 18.060 38.570 18.120 ;
        RECT 311.030 18.060 311.350 18.120 ;
      LAYER via ;
        RECT 38.280 18.060 38.540 18.320 ;
        RECT 311.060 18.060 311.320 18.320 ;
      LAYER met2 ;
        RECT 314.280 1601.130 314.560 1604.000 ;
        RECT 312.500 1600.990 314.560 1601.130 ;
        RECT 312.500 1580.050 312.640 1600.990 ;
        RECT 314.280 1600.000 314.560 1600.990 ;
        RECT 311.120 1579.910 312.640 1580.050 ;
        RECT 311.120 18.350 311.260 1579.910 ;
        RECT 38.280 18.030 38.540 18.350 ;
        RECT 311.060 18.030 311.320 18.350 ;
        RECT 38.340 2.400 38.480 18.030 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 352.505 15.045 352.675 16.235 ;
      LAYER mcon ;
        RECT 352.505 16.065 352.675 16.235 ;
      LAYER met1 ;
        RECT 352.445 16.220 352.735 16.265 ;
        RECT 269.720 16.080 352.735 16.220 ;
        RECT 240.650 15.880 240.970 15.940 ;
        RECT 269.720 15.880 269.860 16.080 ;
        RECT 352.445 16.035 352.735 16.080 ;
        RECT 240.650 15.740 269.860 15.880 ;
        RECT 240.650 15.680 240.970 15.740 ;
        RECT 352.445 15.200 352.735 15.245 ;
        RECT 386.930 15.200 387.250 15.260 ;
        RECT 352.445 15.060 387.250 15.200 ;
        RECT 352.445 15.015 352.735 15.060 ;
        RECT 386.930 15.000 387.250 15.060 ;
      LAYER via ;
        RECT 240.680 15.680 240.940 15.940 ;
        RECT 386.960 15.000 387.220 15.260 ;
      LAYER met2 ;
        RECT 390.640 1600.450 390.920 1604.000 ;
        RECT 388.860 1600.310 390.920 1600.450 ;
        RECT 388.860 1580.050 389.000 1600.310 ;
        RECT 390.640 1600.000 390.920 1600.310 ;
        RECT 387.020 1579.910 389.000 1580.050 ;
        RECT 240.680 15.650 240.940 15.970 ;
        RECT 240.740 2.400 240.880 15.650 ;
        RECT 387.020 15.290 387.160 1579.910 ;
        RECT 386.960 14.970 387.220 15.290 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 394.365 766.105 394.535 814.215 ;
        RECT 393.905 476.085 394.075 524.195 ;
        RECT 394.365 144.925 394.535 193.035 ;
        RECT 352.045 15.045 352.215 20.655 ;
        RECT 376.885 20.145 377.055 20.995 ;
      LAYER mcon ;
        RECT 394.365 814.045 394.535 814.215 ;
        RECT 393.905 524.025 394.075 524.195 ;
        RECT 394.365 192.865 394.535 193.035 ;
        RECT 376.885 20.825 377.055 20.995 ;
        RECT 352.045 20.485 352.215 20.655 ;
      LAYER met1 ;
        RECT 394.290 1545.880 394.610 1545.940 ;
        RECT 395.210 1545.880 395.530 1545.940 ;
        RECT 394.290 1545.740 395.530 1545.880 ;
        RECT 394.290 1545.680 394.610 1545.740 ;
        RECT 395.210 1545.680 395.530 1545.740 ;
        RECT 394.290 834.740 394.610 835.000 ;
        RECT 394.380 834.320 394.520 834.740 ;
        RECT 394.290 834.060 394.610 834.320 ;
        RECT 394.290 814.200 394.610 814.260 ;
        RECT 394.095 814.060 394.610 814.200 ;
        RECT 394.290 814.000 394.610 814.060 ;
        RECT 394.290 766.260 394.610 766.320 ;
        RECT 394.095 766.120 394.610 766.260 ;
        RECT 394.290 766.060 394.610 766.120 ;
        RECT 393.830 700.100 394.150 700.360 ;
        RECT 393.920 699.960 394.060 700.100 ;
        RECT 394.290 699.960 394.610 700.020 ;
        RECT 393.920 699.820 394.610 699.960 ;
        RECT 394.290 699.760 394.610 699.820 ;
        RECT 393.830 627.680 394.150 627.940 ;
        RECT 393.920 627.200 394.060 627.680 ;
        RECT 394.290 627.200 394.610 627.260 ;
        RECT 393.920 627.060 394.610 627.200 ;
        RECT 394.290 627.000 394.610 627.060 ;
        RECT 393.830 524.180 394.150 524.240 ;
        RECT 393.635 524.040 394.150 524.180 ;
        RECT 393.830 523.980 394.150 524.040 ;
        RECT 393.845 476.240 394.135 476.285 ;
        RECT 394.750 476.240 395.070 476.300 ;
        RECT 393.845 476.100 395.070 476.240 ;
        RECT 393.845 476.055 394.135 476.100 ;
        RECT 394.750 476.040 395.070 476.100 ;
        RECT 393.830 427.960 394.150 428.020 ;
        RECT 394.750 427.960 395.070 428.020 ;
        RECT 393.830 427.820 395.070 427.960 ;
        RECT 393.830 427.760 394.150 427.820 ;
        RECT 394.750 427.760 395.070 427.820 ;
        RECT 393.830 379.680 394.150 379.740 ;
        RECT 394.290 379.680 394.610 379.740 ;
        RECT 393.830 379.540 394.610 379.680 ;
        RECT 393.830 379.480 394.150 379.540 ;
        RECT 394.290 379.480 394.610 379.540 ;
        RECT 394.290 193.020 394.610 193.080 ;
        RECT 394.095 192.880 394.610 193.020 ;
        RECT 394.290 192.820 394.610 192.880 ;
        RECT 394.290 145.080 394.610 145.140 ;
        RECT 394.095 144.940 394.610 145.080 ;
        RECT 394.290 144.880 394.610 144.940 ;
        RECT 376.825 20.980 377.115 21.025 ;
        RECT 352.060 20.840 377.115 20.980 ;
        RECT 352.060 20.685 352.200 20.840 ;
        RECT 376.825 20.795 377.115 20.840 ;
        RECT 351.985 20.455 352.275 20.685 ;
        RECT 376.825 20.300 377.115 20.345 ;
        RECT 393.830 20.300 394.150 20.360 ;
        RECT 376.825 20.160 394.150 20.300 ;
        RECT 376.825 20.115 377.115 20.160 ;
        RECT 393.830 20.100 394.150 20.160 ;
        RECT 258.130 15.200 258.450 15.260 ;
        RECT 351.985 15.200 352.275 15.245 ;
        RECT 258.130 15.060 352.275 15.200 ;
        RECT 258.130 15.000 258.450 15.060 ;
        RECT 351.985 15.015 352.275 15.060 ;
      LAYER via ;
        RECT 394.320 1545.680 394.580 1545.940 ;
        RECT 395.240 1545.680 395.500 1545.940 ;
        RECT 394.320 834.740 394.580 835.000 ;
        RECT 394.320 834.060 394.580 834.320 ;
        RECT 394.320 814.000 394.580 814.260 ;
        RECT 394.320 766.060 394.580 766.320 ;
        RECT 393.860 700.100 394.120 700.360 ;
        RECT 394.320 699.760 394.580 700.020 ;
        RECT 393.860 627.680 394.120 627.940 ;
        RECT 394.320 627.000 394.580 627.260 ;
        RECT 393.860 523.980 394.120 524.240 ;
        RECT 394.780 476.040 395.040 476.300 ;
        RECT 393.860 427.760 394.120 428.020 ;
        RECT 394.780 427.760 395.040 428.020 ;
        RECT 393.860 379.480 394.120 379.740 ;
        RECT 394.320 379.480 394.580 379.740 ;
        RECT 394.320 192.820 394.580 193.080 ;
        RECT 394.320 144.880 394.580 145.140 ;
        RECT 393.860 20.100 394.120 20.360 ;
        RECT 258.160 15.000 258.420 15.260 ;
      LAYER met2 ;
        RECT 397.080 1601.130 397.360 1604.000 ;
        RECT 395.300 1600.990 397.360 1601.130 ;
        RECT 395.300 1545.970 395.440 1600.990 ;
        RECT 397.080 1600.000 397.360 1600.990 ;
        RECT 394.320 1545.650 394.580 1545.970 ;
        RECT 395.240 1545.650 395.500 1545.970 ;
        RECT 394.380 1463.090 394.520 1545.650 ;
        RECT 393.920 1462.950 394.520 1463.090 ;
        RECT 393.920 1462.410 394.060 1462.950 ;
        RECT 393.920 1462.270 394.520 1462.410 ;
        RECT 394.380 1318.250 394.520 1462.270 ;
        RECT 393.920 1318.110 394.520 1318.250 ;
        RECT 393.920 1317.570 394.060 1318.110 ;
        RECT 393.920 1317.430 394.520 1317.570 ;
        RECT 394.380 1221.690 394.520 1317.430 ;
        RECT 393.920 1221.550 394.520 1221.690 ;
        RECT 393.920 1221.010 394.060 1221.550 ;
        RECT 393.920 1220.870 394.520 1221.010 ;
        RECT 394.380 1125.130 394.520 1220.870 ;
        RECT 393.920 1124.990 394.520 1125.130 ;
        RECT 393.920 1124.450 394.060 1124.990 ;
        RECT 393.920 1124.310 394.520 1124.450 ;
        RECT 394.380 1028.570 394.520 1124.310 ;
        RECT 393.920 1028.430 394.520 1028.570 ;
        RECT 393.920 1027.890 394.060 1028.430 ;
        RECT 393.920 1027.750 394.520 1027.890 ;
        RECT 394.380 932.010 394.520 1027.750 ;
        RECT 393.920 931.870 394.520 932.010 ;
        RECT 393.920 931.330 394.060 931.870 ;
        RECT 393.920 931.190 394.520 931.330 ;
        RECT 394.380 835.030 394.520 931.190 ;
        RECT 394.320 834.710 394.580 835.030 ;
        RECT 394.320 834.030 394.580 834.350 ;
        RECT 394.380 814.290 394.520 834.030 ;
        RECT 394.320 813.970 394.580 814.290 ;
        RECT 394.320 766.030 394.580 766.350 ;
        RECT 394.380 724.610 394.520 766.030 ;
        RECT 393.920 724.470 394.520 724.610 ;
        RECT 393.920 700.390 394.060 724.470 ;
        RECT 393.860 700.070 394.120 700.390 ;
        RECT 394.320 699.730 394.580 700.050 ;
        RECT 394.380 628.845 394.520 699.730 ;
        RECT 394.310 628.475 394.590 628.845 ;
        RECT 393.850 627.795 394.130 628.165 ;
        RECT 393.860 627.650 394.120 627.795 ;
        RECT 394.320 626.970 394.580 627.290 ;
        RECT 394.380 532.285 394.520 626.970 ;
        RECT 394.310 531.915 394.590 532.285 ;
        RECT 393.850 531.235 394.130 531.605 ;
        RECT 393.920 524.270 394.060 531.235 ;
        RECT 393.860 523.950 394.120 524.270 ;
        RECT 394.780 476.010 395.040 476.330 ;
        RECT 394.840 428.050 394.980 476.010 ;
        RECT 393.860 427.730 394.120 428.050 ;
        RECT 394.780 427.730 395.040 428.050 ;
        RECT 393.920 379.770 394.060 427.730 ;
        RECT 393.860 379.450 394.120 379.770 ;
        RECT 394.320 379.450 394.580 379.770 ;
        RECT 394.380 193.110 394.520 379.450 ;
        RECT 394.320 192.790 394.580 193.110 ;
        RECT 394.320 144.850 394.580 145.170 ;
        RECT 394.380 62.290 394.520 144.850 ;
        RECT 393.920 62.150 394.520 62.290 ;
        RECT 393.920 20.390 394.060 62.150 ;
        RECT 393.860 20.070 394.120 20.390 ;
        RECT 258.160 14.970 258.420 15.290 ;
        RECT 258.220 2.400 258.360 14.970 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 394.310 628.520 394.590 628.800 ;
        RECT 393.850 627.840 394.130 628.120 ;
        RECT 394.310 531.960 394.590 532.240 ;
        RECT 393.850 531.280 394.130 531.560 ;
      LAYER met3 ;
        RECT 394.285 628.810 394.615 628.825 ;
        RECT 394.070 628.495 394.615 628.810 ;
        RECT 394.070 628.145 394.370 628.495 ;
        RECT 393.825 627.830 394.370 628.145 ;
        RECT 393.825 627.815 394.155 627.830 ;
        RECT 394.285 532.250 394.615 532.265 ;
        RECT 394.070 531.935 394.615 532.250 ;
        RECT 394.070 531.585 394.370 531.935 ;
        RECT 393.825 531.270 394.370 531.585 ;
        RECT 393.825 531.255 394.155 531.270 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 401.265 1483.505 401.435 1507.815 ;
      LAYER mcon ;
        RECT 401.265 1507.645 401.435 1507.815 ;
      LAYER met1 ;
        RECT 401.205 1507.800 401.495 1507.845 ;
        RECT 402.110 1507.800 402.430 1507.860 ;
        RECT 401.205 1507.660 402.430 1507.800 ;
        RECT 401.205 1507.615 401.495 1507.660 ;
        RECT 402.110 1507.600 402.430 1507.660 ;
        RECT 401.190 1483.660 401.510 1483.720 ;
        RECT 400.995 1483.520 401.510 1483.660 ;
        RECT 401.190 1483.460 401.510 1483.520 ;
        RECT 401.190 1441.300 401.510 1441.560 ;
        RECT 401.280 1441.160 401.420 1441.300 ;
        RECT 402.110 1441.160 402.430 1441.220 ;
        RECT 401.280 1441.020 402.430 1441.160 ;
        RECT 402.110 1440.960 402.430 1441.020 ;
        RECT 401.650 1304.140 401.970 1304.200 ;
        RECT 402.110 1304.140 402.430 1304.200 ;
        RECT 401.650 1304.000 402.430 1304.140 ;
        RECT 401.650 1303.940 401.970 1304.000 ;
        RECT 402.110 1303.940 402.430 1304.000 ;
        RECT 401.650 1159.300 401.970 1159.360 ;
        RECT 402.110 1159.300 402.430 1159.360 ;
        RECT 401.650 1159.160 402.430 1159.300 ;
        RECT 401.650 1159.100 401.970 1159.160 ;
        RECT 402.110 1159.100 402.430 1159.160 ;
        RECT 401.650 1062.740 401.970 1062.800 ;
        RECT 402.110 1062.740 402.430 1062.800 ;
        RECT 401.650 1062.600 402.430 1062.740 ;
        RECT 401.650 1062.540 401.970 1062.600 ;
        RECT 402.110 1062.540 402.430 1062.600 ;
        RECT 401.650 1014.120 401.970 1014.180 ;
        RECT 402.110 1014.120 402.430 1014.180 ;
        RECT 401.650 1013.980 402.430 1014.120 ;
        RECT 401.650 1013.920 401.970 1013.980 ;
        RECT 402.110 1013.920 402.430 1013.980 ;
        RECT 401.650 917.560 401.970 917.620 ;
        RECT 402.110 917.560 402.430 917.620 ;
        RECT 401.650 917.420 402.430 917.560 ;
        RECT 401.650 917.360 401.970 917.420 ;
        RECT 402.110 917.360 402.430 917.420 ;
        RECT 401.190 786.660 401.510 786.720 ;
        RECT 402.110 786.660 402.430 786.720 ;
        RECT 401.190 786.520 402.430 786.660 ;
        RECT 401.190 786.460 401.510 786.520 ;
        RECT 402.110 786.460 402.430 786.520 ;
        RECT 401.650 772.720 401.970 772.780 ;
        RECT 402.110 772.720 402.430 772.780 ;
        RECT 401.650 772.580 402.430 772.720 ;
        RECT 401.650 772.520 401.970 772.580 ;
        RECT 402.110 772.520 402.430 772.580 ;
        RECT 401.650 689.900 401.970 690.160 ;
        RECT 401.740 689.760 401.880 689.900 ;
        RECT 402.110 689.760 402.430 689.820 ;
        RECT 401.740 689.620 402.430 689.760 ;
        RECT 402.110 689.560 402.430 689.620 ;
        RECT 401.650 593.340 401.970 593.600 ;
        RECT 401.740 593.200 401.880 593.340 ;
        RECT 402.110 593.200 402.430 593.260 ;
        RECT 401.740 593.060 402.430 593.200 ;
        RECT 402.110 593.000 402.430 593.060 ;
        RECT 401.650 351.940 401.970 352.200 ;
        RECT 401.740 351.520 401.880 351.940 ;
        RECT 401.650 351.260 401.970 351.520 ;
        RECT 401.190 303.520 401.510 303.580 ;
        RECT 402.110 303.520 402.430 303.580 ;
        RECT 401.190 303.380 402.430 303.520 ;
        RECT 401.190 303.320 401.510 303.380 ;
        RECT 402.110 303.320 402.430 303.380 ;
        RECT 401.190 206.960 401.510 207.020 ;
        RECT 402.110 206.960 402.430 207.020 ;
        RECT 401.190 206.820 402.430 206.960 ;
        RECT 401.190 206.760 401.510 206.820 ;
        RECT 402.110 206.760 402.430 206.820 ;
        RECT 401.190 110.400 401.510 110.460 ;
        RECT 402.110 110.400 402.430 110.460 ;
        RECT 401.190 110.260 402.430 110.400 ;
        RECT 401.190 110.200 401.510 110.260 ;
        RECT 402.110 110.200 402.430 110.260 ;
        RECT 276.070 24.040 276.390 24.100 ;
        RECT 402.110 24.040 402.430 24.100 ;
        RECT 276.070 23.900 402.430 24.040 ;
        RECT 276.070 23.840 276.390 23.900 ;
        RECT 402.110 23.840 402.430 23.900 ;
      LAYER via ;
        RECT 402.140 1507.600 402.400 1507.860 ;
        RECT 401.220 1483.460 401.480 1483.720 ;
        RECT 401.220 1441.300 401.480 1441.560 ;
        RECT 402.140 1440.960 402.400 1441.220 ;
        RECT 401.680 1303.940 401.940 1304.200 ;
        RECT 402.140 1303.940 402.400 1304.200 ;
        RECT 401.680 1159.100 401.940 1159.360 ;
        RECT 402.140 1159.100 402.400 1159.360 ;
        RECT 401.680 1062.540 401.940 1062.800 ;
        RECT 402.140 1062.540 402.400 1062.800 ;
        RECT 401.680 1013.920 401.940 1014.180 ;
        RECT 402.140 1013.920 402.400 1014.180 ;
        RECT 401.680 917.360 401.940 917.620 ;
        RECT 402.140 917.360 402.400 917.620 ;
        RECT 401.220 786.460 401.480 786.720 ;
        RECT 402.140 786.460 402.400 786.720 ;
        RECT 401.680 772.520 401.940 772.780 ;
        RECT 402.140 772.520 402.400 772.780 ;
        RECT 401.680 689.900 401.940 690.160 ;
        RECT 402.140 689.560 402.400 689.820 ;
        RECT 401.680 593.340 401.940 593.600 ;
        RECT 402.140 593.000 402.400 593.260 ;
        RECT 401.680 351.940 401.940 352.200 ;
        RECT 401.680 351.260 401.940 351.520 ;
        RECT 401.220 303.320 401.480 303.580 ;
        RECT 402.140 303.320 402.400 303.580 ;
        RECT 401.220 206.760 401.480 207.020 ;
        RECT 402.140 206.760 402.400 207.020 ;
        RECT 401.220 110.200 401.480 110.460 ;
        RECT 402.140 110.200 402.400 110.460 ;
        RECT 276.100 23.840 276.360 24.100 ;
        RECT 402.140 23.840 402.400 24.100 ;
      LAYER met2 ;
        RECT 403.980 1600.450 404.260 1604.000 ;
        RECT 402.200 1600.310 404.260 1600.450 ;
        RECT 402.200 1507.890 402.340 1600.310 ;
        RECT 403.980 1600.000 404.260 1600.310 ;
        RECT 402.140 1507.570 402.400 1507.890 ;
        RECT 401.220 1483.430 401.480 1483.750 ;
        RECT 401.280 1441.590 401.420 1483.430 ;
        RECT 401.220 1441.270 401.480 1441.590 ;
        RECT 402.140 1440.930 402.400 1441.250 ;
        RECT 402.200 1317.570 402.340 1440.930 ;
        RECT 401.740 1317.430 402.340 1317.570 ;
        RECT 401.740 1304.230 401.880 1317.430 ;
        RECT 401.680 1303.910 401.940 1304.230 ;
        RECT 402.140 1303.910 402.400 1304.230 ;
        RECT 402.200 1221.010 402.340 1303.910 ;
        RECT 401.740 1220.870 402.340 1221.010 ;
        RECT 401.740 1159.390 401.880 1220.870 ;
        RECT 401.680 1159.070 401.940 1159.390 ;
        RECT 402.140 1159.070 402.400 1159.390 ;
        RECT 402.200 1124.450 402.340 1159.070 ;
        RECT 401.740 1124.310 402.340 1124.450 ;
        RECT 401.740 1062.830 401.880 1124.310 ;
        RECT 401.680 1062.510 401.940 1062.830 ;
        RECT 402.140 1062.510 402.400 1062.830 ;
        RECT 402.200 1027.890 402.340 1062.510 ;
        RECT 401.740 1027.750 402.340 1027.890 ;
        RECT 401.740 1014.210 401.880 1027.750 ;
        RECT 401.680 1013.890 401.940 1014.210 ;
        RECT 402.140 1013.890 402.400 1014.210 ;
        RECT 402.200 931.330 402.340 1013.890 ;
        RECT 401.740 931.190 402.340 931.330 ;
        RECT 401.740 917.650 401.880 931.190 ;
        RECT 401.680 917.330 401.940 917.650 ;
        RECT 402.140 917.330 402.400 917.650 ;
        RECT 402.200 834.770 402.340 917.330 ;
        RECT 401.740 834.630 402.340 834.770 ;
        RECT 401.740 787.170 401.880 834.630 ;
        RECT 401.280 787.030 401.880 787.170 ;
        RECT 401.280 786.750 401.420 787.030 ;
        RECT 401.220 786.430 401.480 786.750 ;
        RECT 402.140 786.430 402.400 786.750 ;
        RECT 402.200 772.810 402.340 786.430 ;
        RECT 401.680 772.490 401.940 772.810 ;
        RECT 402.140 772.490 402.400 772.810 ;
        RECT 401.740 690.190 401.880 772.490 ;
        RECT 401.680 689.870 401.940 690.190 ;
        RECT 402.140 689.530 402.400 689.850 ;
        RECT 402.200 641.650 402.340 689.530 ;
        RECT 401.740 641.510 402.340 641.650 ;
        RECT 401.740 593.630 401.880 641.510 ;
        RECT 401.680 593.310 401.940 593.630 ;
        RECT 402.140 592.970 402.400 593.290 ;
        RECT 402.200 545.090 402.340 592.970 ;
        RECT 401.740 544.950 402.340 545.090 ;
        RECT 401.740 500.210 401.880 544.950 ;
        RECT 401.740 500.070 402.340 500.210 ;
        RECT 402.200 448.530 402.340 500.070 ;
        RECT 401.740 448.390 402.340 448.530 ;
        RECT 401.740 352.230 401.880 448.390 ;
        RECT 401.680 351.910 401.940 352.230 ;
        RECT 401.680 351.230 401.940 351.550 ;
        RECT 401.740 303.690 401.880 351.230 ;
        RECT 401.280 303.610 401.880 303.690 ;
        RECT 401.220 303.550 401.880 303.610 ;
        RECT 401.220 303.290 401.480 303.550 ;
        RECT 402.140 303.290 402.400 303.610 ;
        RECT 402.200 255.410 402.340 303.290 ;
        RECT 401.740 255.270 402.340 255.410 ;
        RECT 401.740 207.130 401.880 255.270 ;
        RECT 401.280 207.050 401.880 207.130 ;
        RECT 401.220 206.990 401.880 207.050 ;
        RECT 401.220 206.730 401.480 206.990 ;
        RECT 402.140 206.730 402.400 207.050 ;
        RECT 402.200 158.850 402.340 206.730 ;
        RECT 401.740 158.710 402.340 158.850 ;
        RECT 401.740 110.570 401.880 158.710 ;
        RECT 401.280 110.490 401.880 110.570 ;
        RECT 401.220 110.430 401.880 110.490 ;
        RECT 401.220 110.170 401.480 110.430 ;
        RECT 402.140 110.170 402.400 110.490 ;
        RECT 402.200 60.250 402.340 110.170 ;
        RECT 402.200 60.110 402.800 60.250 ;
        RECT 402.660 58.890 402.800 60.110 ;
        RECT 402.200 58.750 402.800 58.890 ;
        RECT 402.200 24.130 402.340 58.750 ;
        RECT 276.100 23.810 276.360 24.130 ;
        RECT 402.140 23.810 402.400 24.130 ;
        RECT 276.160 2.400 276.300 23.810 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 408.625 1393.745 408.795 1418.055 ;
        RECT 408.165 351.305 408.335 386.155 ;
        RECT 375.045 14.025 375.215 15.555 ;
        RECT 397.585 15.385 397.755 18.955 ;
      LAYER mcon ;
        RECT 408.625 1417.885 408.795 1418.055 ;
        RECT 408.165 385.985 408.335 386.155 ;
        RECT 397.585 18.785 397.755 18.955 ;
        RECT 375.045 15.385 375.215 15.555 ;
      LAYER met1 ;
        RECT 408.550 1418.040 408.870 1418.100 ;
        RECT 408.355 1417.900 408.870 1418.040 ;
        RECT 408.550 1417.840 408.870 1417.900 ;
        RECT 408.550 1393.900 408.870 1393.960 ;
        RECT 408.355 1393.760 408.870 1393.900 ;
        RECT 408.550 1393.700 408.870 1393.760 ;
        RECT 409.010 1256.200 409.330 1256.260 ;
        RECT 409.470 1256.200 409.790 1256.260 ;
        RECT 409.010 1256.060 409.790 1256.200 ;
        RECT 409.010 1256.000 409.330 1256.060 ;
        RECT 409.470 1256.000 409.790 1256.060 ;
        RECT 409.010 1159.300 409.330 1159.360 ;
        RECT 409.470 1159.300 409.790 1159.360 ;
        RECT 409.010 1159.160 409.790 1159.300 ;
        RECT 409.010 1159.100 409.330 1159.160 ;
        RECT 409.470 1159.100 409.790 1159.160 ;
        RECT 409.010 1062.740 409.330 1062.800 ;
        RECT 409.470 1062.740 409.790 1062.800 ;
        RECT 409.010 1062.600 409.790 1062.740 ;
        RECT 409.010 1062.540 409.330 1062.600 ;
        RECT 409.470 1062.540 409.790 1062.600 ;
        RECT 409.010 966.180 409.330 966.240 ;
        RECT 409.470 966.180 409.790 966.240 ;
        RECT 409.010 966.040 409.790 966.180 ;
        RECT 409.010 965.980 409.330 966.040 ;
        RECT 409.470 965.980 409.790 966.040 ;
        RECT 409.010 869.620 409.330 869.680 ;
        RECT 409.470 869.620 409.790 869.680 ;
        RECT 409.010 869.480 409.790 869.620 ;
        RECT 409.010 869.420 409.330 869.480 ;
        RECT 409.470 869.420 409.790 869.480 ;
        RECT 408.550 786.660 408.870 786.720 ;
        RECT 409.470 786.660 409.790 786.720 ;
        RECT 408.550 786.520 409.790 786.660 ;
        RECT 408.550 786.460 408.870 786.520 ;
        RECT 409.470 786.460 409.790 786.520 ;
        RECT 409.010 772.720 409.330 772.780 ;
        RECT 409.470 772.720 409.790 772.780 ;
        RECT 409.010 772.580 409.790 772.720 ;
        RECT 409.010 772.520 409.330 772.580 ;
        RECT 409.470 772.520 409.790 772.580 ;
        RECT 409.010 689.900 409.330 690.160 ;
        RECT 409.100 689.760 409.240 689.900 ;
        RECT 409.470 689.760 409.790 689.820 ;
        RECT 409.100 689.620 409.790 689.760 ;
        RECT 409.470 689.560 409.790 689.620 ;
        RECT 409.010 593.340 409.330 593.600 ;
        RECT 409.100 593.200 409.240 593.340 ;
        RECT 409.470 593.200 409.790 593.260 ;
        RECT 409.100 593.060 409.790 593.200 ;
        RECT 409.470 593.000 409.790 593.060 ;
        RECT 408.550 400.760 408.870 400.820 ;
        RECT 408.180 400.620 408.870 400.760 ;
        RECT 408.180 400.140 408.320 400.620 ;
        RECT 408.550 400.560 408.870 400.620 ;
        RECT 408.090 399.880 408.410 400.140 ;
        RECT 408.090 386.140 408.410 386.200 ;
        RECT 407.895 386.000 408.410 386.140 ;
        RECT 408.090 385.940 408.410 386.000 ;
        RECT 408.105 351.460 408.395 351.505 ;
        RECT 408.550 351.460 408.870 351.520 ;
        RECT 408.105 351.320 408.870 351.460 ;
        RECT 408.105 351.275 408.395 351.320 ;
        RECT 408.550 351.260 408.870 351.320 ;
        RECT 408.550 303.520 408.870 303.580 ;
        RECT 409.470 303.520 409.790 303.580 ;
        RECT 408.550 303.380 409.790 303.520 ;
        RECT 408.550 303.320 408.870 303.380 ;
        RECT 409.470 303.320 409.790 303.380 ;
        RECT 408.550 206.960 408.870 207.020 ;
        RECT 409.470 206.960 409.790 207.020 ;
        RECT 408.550 206.820 409.790 206.960 ;
        RECT 408.550 206.760 408.870 206.820 ;
        RECT 409.470 206.760 409.790 206.820 ;
        RECT 409.010 145.080 409.330 145.140 ;
        RECT 409.470 145.080 409.790 145.140 ;
        RECT 409.010 144.940 409.790 145.080 ;
        RECT 409.010 144.880 409.330 144.940 ;
        RECT 409.470 144.880 409.790 144.940 ;
        RECT 408.550 110.400 408.870 110.460 ;
        RECT 409.470 110.400 409.790 110.460 ;
        RECT 408.550 110.260 409.790 110.400 ;
        RECT 408.550 110.200 408.870 110.260 ;
        RECT 409.470 110.200 409.790 110.260 ;
        RECT 397.525 18.940 397.815 18.985 ;
        RECT 409.470 18.940 409.790 19.000 ;
        RECT 397.525 18.800 409.790 18.940 ;
        RECT 397.525 18.755 397.815 18.800 ;
        RECT 409.470 18.740 409.790 18.800 ;
        RECT 374.985 15.540 375.275 15.585 ;
        RECT 397.525 15.540 397.815 15.585 ;
        RECT 374.985 15.400 397.815 15.540 ;
        RECT 374.985 15.355 375.275 15.400 ;
        RECT 397.525 15.355 397.815 15.400 ;
        RECT 294.010 14.180 294.330 14.240 ;
        RECT 374.985 14.180 375.275 14.225 ;
        RECT 294.010 14.040 375.275 14.180 ;
        RECT 294.010 13.980 294.330 14.040 ;
        RECT 374.985 13.995 375.275 14.040 ;
      LAYER via ;
        RECT 408.580 1417.840 408.840 1418.100 ;
        RECT 408.580 1393.700 408.840 1393.960 ;
        RECT 409.040 1256.000 409.300 1256.260 ;
        RECT 409.500 1256.000 409.760 1256.260 ;
        RECT 409.040 1159.100 409.300 1159.360 ;
        RECT 409.500 1159.100 409.760 1159.360 ;
        RECT 409.040 1062.540 409.300 1062.800 ;
        RECT 409.500 1062.540 409.760 1062.800 ;
        RECT 409.040 965.980 409.300 966.240 ;
        RECT 409.500 965.980 409.760 966.240 ;
        RECT 409.040 869.420 409.300 869.680 ;
        RECT 409.500 869.420 409.760 869.680 ;
        RECT 408.580 786.460 408.840 786.720 ;
        RECT 409.500 786.460 409.760 786.720 ;
        RECT 409.040 772.520 409.300 772.780 ;
        RECT 409.500 772.520 409.760 772.780 ;
        RECT 409.040 689.900 409.300 690.160 ;
        RECT 409.500 689.560 409.760 689.820 ;
        RECT 409.040 593.340 409.300 593.600 ;
        RECT 409.500 593.000 409.760 593.260 ;
        RECT 408.580 400.560 408.840 400.820 ;
        RECT 408.120 399.880 408.380 400.140 ;
        RECT 408.120 385.940 408.380 386.200 ;
        RECT 408.580 351.260 408.840 351.520 ;
        RECT 408.580 303.320 408.840 303.580 ;
        RECT 409.500 303.320 409.760 303.580 ;
        RECT 408.580 206.760 408.840 207.020 ;
        RECT 409.500 206.760 409.760 207.020 ;
        RECT 409.040 144.880 409.300 145.140 ;
        RECT 409.500 144.880 409.760 145.140 ;
        RECT 408.580 110.200 408.840 110.460 ;
        RECT 409.500 110.200 409.760 110.460 ;
        RECT 409.500 18.740 409.760 19.000 ;
        RECT 294.040 13.980 294.300 14.240 ;
      LAYER met2 ;
        RECT 410.880 1600.450 411.160 1604.000 ;
        RECT 409.560 1600.310 411.160 1600.450 ;
        RECT 409.560 1497.770 409.700 1600.310 ;
        RECT 410.880 1600.000 411.160 1600.310 ;
        RECT 409.100 1497.630 409.700 1497.770 ;
        RECT 409.100 1467.170 409.240 1497.630 ;
        RECT 408.640 1467.030 409.240 1467.170 ;
        RECT 408.640 1418.130 408.780 1467.030 ;
        RECT 408.580 1417.810 408.840 1418.130 ;
        RECT 408.580 1393.845 408.840 1393.990 ;
        RECT 408.570 1393.475 408.850 1393.845 ;
        RECT 409.490 1351.995 409.770 1352.365 ;
        RECT 409.560 1317.570 409.700 1351.995 ;
        RECT 409.100 1317.430 409.700 1317.570 ;
        RECT 409.100 1256.290 409.240 1317.430 ;
        RECT 409.040 1255.970 409.300 1256.290 ;
        RECT 409.500 1255.970 409.760 1256.290 ;
        RECT 409.560 1221.010 409.700 1255.970 ;
        RECT 409.100 1220.870 409.700 1221.010 ;
        RECT 409.100 1159.390 409.240 1220.870 ;
        RECT 409.040 1159.070 409.300 1159.390 ;
        RECT 409.500 1159.070 409.760 1159.390 ;
        RECT 409.560 1124.450 409.700 1159.070 ;
        RECT 409.100 1124.310 409.700 1124.450 ;
        RECT 409.100 1062.830 409.240 1124.310 ;
        RECT 409.040 1062.510 409.300 1062.830 ;
        RECT 409.500 1062.510 409.760 1062.830 ;
        RECT 409.560 1027.890 409.700 1062.510 ;
        RECT 409.100 1027.750 409.700 1027.890 ;
        RECT 409.100 966.270 409.240 1027.750 ;
        RECT 409.040 965.950 409.300 966.270 ;
        RECT 409.500 965.950 409.760 966.270 ;
        RECT 409.560 931.330 409.700 965.950 ;
        RECT 409.100 931.190 409.700 931.330 ;
        RECT 409.100 869.710 409.240 931.190 ;
        RECT 409.040 869.390 409.300 869.710 ;
        RECT 409.500 869.390 409.760 869.710 ;
        RECT 409.560 834.770 409.700 869.390 ;
        RECT 409.100 834.630 409.700 834.770 ;
        RECT 409.100 787.170 409.240 834.630 ;
        RECT 408.640 787.030 409.240 787.170 ;
        RECT 408.640 786.750 408.780 787.030 ;
        RECT 408.580 786.430 408.840 786.750 ;
        RECT 409.500 786.430 409.760 786.750 ;
        RECT 409.560 772.810 409.700 786.430 ;
        RECT 409.040 772.490 409.300 772.810 ;
        RECT 409.500 772.490 409.760 772.810 ;
        RECT 409.100 690.190 409.240 772.490 ;
        RECT 409.040 689.870 409.300 690.190 ;
        RECT 409.500 689.530 409.760 689.850 ;
        RECT 409.560 641.650 409.700 689.530 ;
        RECT 409.100 641.510 409.700 641.650 ;
        RECT 409.100 593.630 409.240 641.510 ;
        RECT 409.040 593.310 409.300 593.630 ;
        RECT 409.500 592.970 409.760 593.290 ;
        RECT 409.560 545.090 409.700 592.970 ;
        RECT 409.100 544.950 409.700 545.090 ;
        RECT 409.100 500.210 409.240 544.950 ;
        RECT 409.100 500.070 409.700 500.210 ;
        RECT 409.560 448.530 409.700 500.070 ;
        RECT 408.640 448.390 409.700 448.530 ;
        RECT 408.640 400.850 408.780 448.390 ;
        RECT 408.580 400.530 408.840 400.850 ;
        RECT 408.120 399.850 408.380 400.170 ;
        RECT 408.180 386.230 408.320 399.850 ;
        RECT 408.120 385.910 408.380 386.230 ;
        RECT 408.580 351.230 408.840 351.550 ;
        RECT 408.640 303.610 408.780 351.230 ;
        RECT 408.580 303.290 408.840 303.610 ;
        RECT 409.500 303.290 409.760 303.610 ;
        RECT 409.560 255.410 409.700 303.290 ;
        RECT 409.100 255.270 409.700 255.410 ;
        RECT 409.100 207.130 409.240 255.270 ;
        RECT 408.640 207.050 409.240 207.130 ;
        RECT 408.580 206.990 409.240 207.050 ;
        RECT 408.580 206.730 408.840 206.990 ;
        RECT 409.500 206.730 409.760 207.050 ;
        RECT 409.560 145.170 409.700 206.730 ;
        RECT 409.040 144.850 409.300 145.170 ;
        RECT 409.500 144.850 409.760 145.170 ;
        RECT 409.100 110.570 409.240 144.850 ;
        RECT 408.640 110.490 409.240 110.570 ;
        RECT 408.580 110.430 409.240 110.490 ;
        RECT 408.580 110.170 408.840 110.430 ;
        RECT 409.500 110.170 409.760 110.490 ;
        RECT 409.560 60.250 409.700 110.170 ;
        RECT 409.560 60.110 410.160 60.250 ;
        RECT 410.020 58.890 410.160 60.110 ;
        RECT 409.560 58.750 410.160 58.890 ;
        RECT 409.560 19.030 409.700 58.750 ;
        RECT 409.500 18.710 409.760 19.030 ;
        RECT 294.040 13.950 294.300 14.270 ;
        RECT 294.100 2.400 294.240 13.950 ;
        RECT 293.890 -4.800 294.450 2.400 ;
      LAYER via2 ;
        RECT 408.570 1393.520 408.850 1393.800 ;
        RECT 409.490 1352.040 409.770 1352.320 ;
      LAYER met3 ;
        RECT 408.545 1393.820 408.875 1393.825 ;
        RECT 408.545 1393.810 409.130 1393.820 ;
        RECT 408.545 1393.510 409.330 1393.810 ;
        RECT 408.545 1393.500 409.130 1393.510 ;
        RECT 408.545 1393.495 408.875 1393.500 ;
        RECT 408.750 1352.330 409.130 1352.340 ;
        RECT 409.465 1352.330 409.795 1352.345 ;
        RECT 408.750 1352.030 409.795 1352.330 ;
        RECT 408.750 1352.020 409.130 1352.030 ;
        RECT 409.465 1352.015 409.795 1352.030 ;
      LAYER via3 ;
        RECT 408.780 1393.500 409.100 1393.820 ;
        RECT 408.780 1352.020 409.100 1352.340 ;
      LAYER met4 ;
        RECT 408.775 1393.495 409.105 1393.825 ;
        RECT 408.790 1352.345 409.090 1393.495 ;
        RECT 408.775 1352.015 409.105 1352.345 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 376.425 18.785 376.595 19.635 ;
      LAYER mcon ;
        RECT 376.425 19.465 376.595 19.635 ;
      LAYER met1 ;
        RECT 397.050 1589.740 397.370 1589.800 ;
        RECT 417.290 1589.740 417.610 1589.800 ;
        RECT 397.050 1589.600 417.610 1589.740 ;
        RECT 397.050 1589.540 397.370 1589.600 ;
        RECT 417.290 1589.540 417.610 1589.600 ;
        RECT 376.365 19.620 376.655 19.665 ;
        RECT 371.380 19.480 376.655 19.620 ;
        RECT 371.380 19.280 371.520 19.480 ;
        RECT 376.365 19.435 376.655 19.480 ;
        RECT 325.380 19.140 371.520 19.280 ;
        RECT 311.950 18.260 312.270 18.320 ;
        RECT 325.380 18.260 325.520 19.140 ;
        RECT 376.365 18.940 376.655 18.985 ;
        RECT 397.050 18.940 397.370 19.000 ;
        RECT 376.365 18.800 397.370 18.940 ;
        RECT 376.365 18.755 376.655 18.800 ;
        RECT 397.050 18.740 397.370 18.800 ;
        RECT 311.950 18.120 325.520 18.260 ;
        RECT 311.950 18.060 312.270 18.120 ;
      LAYER via ;
        RECT 397.080 1589.540 397.340 1589.800 ;
        RECT 417.320 1589.540 417.580 1589.800 ;
        RECT 311.980 18.060 312.240 18.320 ;
        RECT 397.080 18.740 397.340 19.000 ;
      LAYER met2 ;
        RECT 417.320 1600.000 417.600 1604.000 ;
        RECT 417.380 1589.830 417.520 1600.000 ;
        RECT 397.080 1589.510 397.340 1589.830 ;
        RECT 417.320 1589.510 417.580 1589.830 ;
        RECT 397.140 19.030 397.280 1589.510 ;
        RECT 397.080 18.710 397.340 19.030 ;
        RECT 311.980 18.030 312.240 18.350 ;
        RECT 312.040 2.400 312.180 18.030 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 421.430 1579.880 421.750 1579.940 ;
        RECT 422.350 1579.880 422.670 1579.940 ;
        RECT 421.430 1579.740 422.670 1579.880 ;
        RECT 421.430 1579.680 421.750 1579.740 ;
        RECT 422.350 1579.680 422.670 1579.740 ;
        RECT 329.890 18.260 330.210 18.320 ;
        RECT 421.430 18.260 421.750 18.320 ;
        RECT 329.890 18.120 421.750 18.260 ;
        RECT 329.890 18.060 330.210 18.120 ;
        RECT 421.430 18.060 421.750 18.120 ;
      LAYER via ;
        RECT 421.460 1579.680 421.720 1579.940 ;
        RECT 422.380 1579.680 422.640 1579.940 ;
        RECT 329.920 18.060 330.180 18.320 ;
        RECT 421.460 18.060 421.720 18.320 ;
      LAYER met2 ;
        RECT 424.220 1600.450 424.500 1604.000 ;
        RECT 422.440 1600.310 424.500 1600.450 ;
        RECT 422.440 1579.970 422.580 1600.310 ;
        RECT 424.220 1600.000 424.500 1600.310 ;
        RECT 421.460 1579.650 421.720 1579.970 ;
        RECT 422.380 1579.650 422.640 1579.970 ;
        RECT 421.520 18.350 421.660 1579.650 ;
        RECT 329.920 18.030 330.180 18.350 ;
        RECT 421.460 18.030 421.720 18.350 ;
        RECT 329.980 2.400 330.120 18.030 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 429.785 1490.645 429.955 1538.755 ;
        RECT 429.785 476.085 429.955 524.195 ;
        RECT 429.325 386.325 429.495 434.775 ;
      LAYER mcon ;
        RECT 429.785 1538.585 429.955 1538.755 ;
        RECT 429.785 524.025 429.955 524.195 ;
        RECT 429.325 434.605 429.495 434.775 ;
      LAYER met1 ;
        RECT 430.170 1545.880 430.490 1545.940 ;
        RECT 430.630 1545.880 430.950 1545.940 ;
        RECT 430.170 1545.740 430.950 1545.880 ;
        RECT 430.170 1545.680 430.490 1545.740 ;
        RECT 430.630 1545.680 430.950 1545.740 ;
        RECT 429.725 1538.740 430.015 1538.785 ;
        RECT 430.170 1538.740 430.490 1538.800 ;
        RECT 429.725 1538.600 430.490 1538.740 ;
        RECT 429.725 1538.555 430.015 1538.600 ;
        RECT 430.170 1538.540 430.490 1538.600 ;
        RECT 429.710 1490.800 430.030 1490.860 ;
        RECT 429.515 1490.660 430.030 1490.800 ;
        RECT 429.710 1490.600 430.030 1490.660 ;
        RECT 429.710 1463.060 430.030 1463.320 ;
        RECT 429.800 1462.640 429.940 1463.060 ;
        RECT 429.710 1462.380 430.030 1462.640 ;
        RECT 429.250 1394.240 429.570 1394.300 ;
        RECT 429.710 1394.240 430.030 1394.300 ;
        RECT 429.250 1394.100 430.030 1394.240 ;
        RECT 429.250 1394.040 429.570 1394.100 ;
        RECT 429.710 1394.040 430.030 1394.100 ;
        RECT 429.250 1393.560 429.570 1393.620 ;
        RECT 430.170 1393.560 430.490 1393.620 ;
        RECT 429.250 1393.420 430.490 1393.560 ;
        RECT 429.250 1393.360 429.570 1393.420 ;
        RECT 430.170 1393.360 430.490 1393.420 ;
        RECT 430.170 1386.760 430.490 1386.820 ;
        RECT 430.630 1386.760 430.950 1386.820 ;
        RECT 430.170 1386.620 430.950 1386.760 ;
        RECT 430.170 1386.560 430.490 1386.620 ;
        RECT 430.630 1386.560 430.950 1386.620 ;
        RECT 429.710 1255.860 430.030 1255.920 ;
        RECT 430.630 1255.860 430.950 1255.920 ;
        RECT 429.710 1255.720 430.950 1255.860 ;
        RECT 429.710 1255.660 430.030 1255.720 ;
        RECT 430.630 1255.660 430.950 1255.720 ;
        RECT 429.710 1173.240 430.030 1173.300 ;
        RECT 429.340 1173.100 430.030 1173.240 ;
        RECT 429.340 1172.960 429.480 1173.100 ;
        RECT 429.710 1173.040 430.030 1173.100 ;
        RECT 429.250 1172.700 429.570 1172.960 ;
        RECT 429.710 1014.460 430.030 1014.520 ;
        RECT 430.630 1014.460 430.950 1014.520 ;
        RECT 429.710 1014.320 430.950 1014.460 ;
        RECT 429.710 1014.260 430.030 1014.320 ;
        RECT 430.630 1014.260 430.950 1014.320 ;
        RECT 429.710 980.120 430.030 980.180 ;
        RECT 429.340 979.980 430.030 980.120 ;
        RECT 429.340 979.840 429.480 979.980 ;
        RECT 429.710 979.920 430.030 979.980 ;
        RECT 429.250 979.580 429.570 979.840 ;
        RECT 429.710 917.900 430.030 917.960 ;
        RECT 430.630 917.900 430.950 917.960 ;
        RECT 429.710 917.760 430.950 917.900 ;
        RECT 429.710 917.700 430.030 917.760 ;
        RECT 430.630 917.700 430.950 917.760 ;
        RECT 429.710 883.560 430.030 883.620 ;
        RECT 429.340 883.420 430.030 883.560 ;
        RECT 429.340 883.280 429.480 883.420 ;
        RECT 429.710 883.360 430.030 883.420 ;
        RECT 429.250 883.020 429.570 883.280 ;
        RECT 429.250 786.660 429.570 786.720 ;
        RECT 430.170 786.660 430.490 786.720 ;
        RECT 429.250 786.520 430.490 786.660 ;
        RECT 429.250 786.460 429.570 786.520 ;
        RECT 430.170 786.460 430.490 786.520 ;
        RECT 429.250 724.440 429.570 724.500 ;
        RECT 429.710 724.440 430.030 724.500 ;
        RECT 429.250 724.300 430.030 724.440 ;
        RECT 429.250 724.240 429.570 724.300 ;
        RECT 429.710 724.240 430.030 724.300 ;
        RECT 429.250 627.880 429.570 627.940 ;
        RECT 429.710 627.880 430.030 627.940 ;
        RECT 429.250 627.740 430.030 627.880 ;
        RECT 429.250 627.680 429.570 627.740 ;
        RECT 429.710 627.680 430.030 627.740 ;
        RECT 429.710 531.660 430.030 531.720 ;
        RECT 430.170 531.660 430.490 531.720 ;
        RECT 429.710 531.520 430.490 531.660 ;
        RECT 429.710 531.460 430.030 531.520 ;
        RECT 430.170 531.460 430.490 531.520 ;
        RECT 429.710 524.180 430.030 524.240 ;
        RECT 429.515 524.040 430.030 524.180 ;
        RECT 429.710 523.980 430.030 524.040 ;
        RECT 429.725 476.240 430.015 476.285 ;
        RECT 430.170 476.240 430.490 476.300 ;
        RECT 429.725 476.100 430.490 476.240 ;
        RECT 429.725 476.055 430.015 476.100 ;
        RECT 430.170 476.040 430.490 476.100 ;
        RECT 429.265 434.760 429.555 434.805 ;
        RECT 429.710 434.760 430.030 434.820 ;
        RECT 429.265 434.620 430.030 434.760 ;
        RECT 429.265 434.575 429.555 434.620 ;
        RECT 429.710 434.560 430.030 434.620 ;
        RECT 429.250 386.480 429.570 386.540 ;
        RECT 429.055 386.340 429.570 386.480 ;
        RECT 429.250 386.280 429.570 386.340 ;
        RECT 429.250 144.880 429.570 145.140 ;
        RECT 429.340 144.400 429.480 144.880 ;
        RECT 429.710 144.400 430.030 144.460 ;
        RECT 429.340 144.260 430.030 144.400 ;
        RECT 429.710 144.200 430.030 144.260 ;
        RECT 429.710 131.140 430.030 131.200 ;
        RECT 430.170 131.140 430.490 131.200 ;
        RECT 429.710 131.000 430.490 131.140 ;
        RECT 429.710 130.940 430.030 131.000 ;
        RECT 430.170 130.940 430.490 131.000 ;
        RECT 347.370 16.560 347.690 16.620 ;
        RECT 430.170 16.560 430.490 16.620 ;
        RECT 347.370 16.420 430.490 16.560 ;
        RECT 347.370 16.360 347.690 16.420 ;
        RECT 430.170 16.360 430.490 16.420 ;
      LAYER via ;
        RECT 430.200 1545.680 430.460 1545.940 ;
        RECT 430.660 1545.680 430.920 1545.940 ;
        RECT 430.200 1538.540 430.460 1538.800 ;
        RECT 429.740 1490.600 430.000 1490.860 ;
        RECT 429.740 1463.060 430.000 1463.320 ;
        RECT 429.740 1462.380 430.000 1462.640 ;
        RECT 429.280 1394.040 429.540 1394.300 ;
        RECT 429.740 1394.040 430.000 1394.300 ;
        RECT 429.280 1393.360 429.540 1393.620 ;
        RECT 430.200 1393.360 430.460 1393.620 ;
        RECT 430.200 1386.560 430.460 1386.820 ;
        RECT 430.660 1386.560 430.920 1386.820 ;
        RECT 429.740 1255.660 430.000 1255.920 ;
        RECT 430.660 1255.660 430.920 1255.920 ;
        RECT 429.740 1173.040 430.000 1173.300 ;
        RECT 429.280 1172.700 429.540 1172.960 ;
        RECT 429.740 1014.260 430.000 1014.520 ;
        RECT 430.660 1014.260 430.920 1014.520 ;
        RECT 429.740 979.920 430.000 980.180 ;
        RECT 429.280 979.580 429.540 979.840 ;
        RECT 429.740 917.700 430.000 917.960 ;
        RECT 430.660 917.700 430.920 917.960 ;
        RECT 429.740 883.360 430.000 883.620 ;
        RECT 429.280 883.020 429.540 883.280 ;
        RECT 429.280 786.460 429.540 786.720 ;
        RECT 430.200 786.460 430.460 786.720 ;
        RECT 429.280 724.240 429.540 724.500 ;
        RECT 429.740 724.240 430.000 724.500 ;
        RECT 429.280 627.680 429.540 627.940 ;
        RECT 429.740 627.680 430.000 627.940 ;
        RECT 429.740 531.460 430.000 531.720 ;
        RECT 430.200 531.460 430.460 531.720 ;
        RECT 429.740 523.980 430.000 524.240 ;
        RECT 430.200 476.040 430.460 476.300 ;
        RECT 429.740 434.560 430.000 434.820 ;
        RECT 429.280 386.280 429.540 386.540 ;
        RECT 429.280 144.880 429.540 145.140 ;
        RECT 429.740 144.200 430.000 144.460 ;
        RECT 429.740 130.940 430.000 131.200 ;
        RECT 430.200 130.940 430.460 131.200 ;
        RECT 347.400 16.360 347.660 16.620 ;
        RECT 430.200 16.360 430.460 16.620 ;
      LAYER met2 ;
        RECT 431.120 1600.450 431.400 1604.000 ;
        RECT 430.720 1600.310 431.400 1600.450 ;
        RECT 430.720 1545.970 430.860 1600.310 ;
        RECT 431.120 1600.000 431.400 1600.310 ;
        RECT 430.200 1545.650 430.460 1545.970 ;
        RECT 430.660 1545.650 430.920 1545.970 ;
        RECT 430.260 1538.830 430.400 1545.650 ;
        RECT 430.200 1538.510 430.460 1538.830 ;
        RECT 429.740 1490.570 430.000 1490.890 ;
        RECT 429.800 1463.350 429.940 1490.570 ;
        RECT 429.740 1463.030 430.000 1463.350 ;
        RECT 429.740 1462.350 430.000 1462.670 ;
        RECT 429.800 1394.330 429.940 1462.350 ;
        RECT 429.280 1394.010 429.540 1394.330 ;
        RECT 429.740 1394.010 430.000 1394.330 ;
        RECT 429.340 1393.650 429.480 1394.010 ;
        RECT 429.280 1393.330 429.540 1393.650 ;
        RECT 430.200 1393.330 430.460 1393.650 ;
        RECT 430.260 1386.850 430.400 1393.330 ;
        RECT 430.200 1386.530 430.460 1386.850 ;
        RECT 430.660 1386.530 430.920 1386.850 ;
        RECT 430.720 1255.950 430.860 1386.530 ;
        RECT 429.740 1255.630 430.000 1255.950 ;
        RECT 430.660 1255.630 430.920 1255.950 ;
        RECT 429.800 1173.330 429.940 1255.630 ;
        RECT 429.740 1173.010 430.000 1173.330 ;
        RECT 429.280 1172.670 429.540 1172.990 ;
        RECT 429.340 1062.685 429.480 1172.670 ;
        RECT 429.270 1062.315 429.550 1062.685 ;
        RECT 430.650 1062.315 430.930 1062.685 ;
        RECT 430.720 1014.550 430.860 1062.315 ;
        RECT 429.740 1014.230 430.000 1014.550 ;
        RECT 430.660 1014.230 430.920 1014.550 ;
        RECT 429.800 980.210 429.940 1014.230 ;
        RECT 429.740 979.890 430.000 980.210 ;
        RECT 429.280 979.550 429.540 979.870 ;
        RECT 429.340 966.125 429.480 979.550 ;
        RECT 429.270 965.755 429.550 966.125 ;
        RECT 430.650 965.755 430.930 966.125 ;
        RECT 430.720 917.990 430.860 965.755 ;
        RECT 429.740 917.670 430.000 917.990 ;
        RECT 430.660 917.670 430.920 917.990 ;
        RECT 429.800 883.650 429.940 917.670 ;
        RECT 429.740 883.330 430.000 883.650 ;
        RECT 429.280 882.990 429.540 883.310 ;
        RECT 429.340 786.750 429.480 882.990 ;
        RECT 429.280 786.430 429.540 786.750 ;
        RECT 430.200 786.430 430.460 786.750 ;
        RECT 430.260 738.890 430.400 786.430 ;
        RECT 430.260 738.750 430.860 738.890 ;
        RECT 430.720 724.725 430.860 738.750 ;
        RECT 429.280 724.210 429.540 724.530 ;
        RECT 429.730 724.355 430.010 724.725 ;
        RECT 430.650 724.355 430.930 724.725 ;
        RECT 429.740 724.210 430.000 724.355 ;
        RECT 429.340 676.445 429.480 724.210 ;
        RECT 429.270 676.075 429.550 676.445 ;
        RECT 430.190 676.075 430.470 676.445 ;
        RECT 430.260 642.330 430.400 676.075 ;
        RECT 430.260 642.190 430.860 642.330 ;
        RECT 430.720 628.165 430.860 642.190 ;
        RECT 429.280 627.650 429.540 627.970 ;
        RECT 429.730 627.795 430.010 628.165 ;
        RECT 430.650 627.795 430.930 628.165 ;
        RECT 429.740 627.650 430.000 627.795 ;
        RECT 429.340 579.885 429.480 627.650 ;
        RECT 429.270 579.515 429.550 579.885 ;
        RECT 430.190 579.515 430.470 579.885 ;
        RECT 430.260 531.750 430.400 579.515 ;
        RECT 429.740 531.430 430.000 531.750 ;
        RECT 430.200 531.430 430.460 531.750 ;
        RECT 429.800 524.270 429.940 531.430 ;
        RECT 429.740 523.950 430.000 524.270 ;
        RECT 430.200 476.010 430.460 476.330 ;
        RECT 430.260 448.530 430.400 476.010 ;
        RECT 429.800 448.390 430.400 448.530 ;
        RECT 429.800 434.850 429.940 448.390 ;
        RECT 429.740 434.530 430.000 434.850 ;
        RECT 429.280 386.250 429.540 386.570 ;
        RECT 429.340 145.170 429.480 386.250 ;
        RECT 429.280 144.850 429.540 145.170 ;
        RECT 429.740 144.170 430.000 144.490 ;
        RECT 429.800 131.230 429.940 144.170 ;
        RECT 429.740 130.910 430.000 131.230 ;
        RECT 430.200 130.910 430.460 131.230 ;
        RECT 430.260 16.650 430.400 130.910 ;
        RECT 347.400 16.330 347.660 16.650 ;
        RECT 430.200 16.330 430.460 16.650 ;
        RECT 347.460 2.400 347.600 16.330 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 429.270 1062.360 429.550 1062.640 ;
        RECT 430.650 1062.360 430.930 1062.640 ;
        RECT 429.270 965.800 429.550 966.080 ;
        RECT 430.650 965.800 430.930 966.080 ;
        RECT 429.730 724.400 430.010 724.680 ;
        RECT 430.650 724.400 430.930 724.680 ;
        RECT 429.270 676.120 429.550 676.400 ;
        RECT 430.190 676.120 430.470 676.400 ;
        RECT 429.730 627.840 430.010 628.120 ;
        RECT 430.650 627.840 430.930 628.120 ;
        RECT 429.270 579.560 429.550 579.840 ;
        RECT 430.190 579.560 430.470 579.840 ;
      LAYER met3 ;
        RECT 429.245 1062.650 429.575 1062.665 ;
        RECT 430.625 1062.650 430.955 1062.665 ;
        RECT 429.245 1062.350 430.955 1062.650 ;
        RECT 429.245 1062.335 429.575 1062.350 ;
        RECT 430.625 1062.335 430.955 1062.350 ;
        RECT 429.245 966.090 429.575 966.105 ;
        RECT 430.625 966.090 430.955 966.105 ;
        RECT 429.245 965.790 430.955 966.090 ;
        RECT 429.245 965.775 429.575 965.790 ;
        RECT 430.625 965.775 430.955 965.790 ;
        RECT 429.705 724.690 430.035 724.705 ;
        RECT 430.625 724.690 430.955 724.705 ;
        RECT 429.705 724.390 430.955 724.690 ;
        RECT 429.705 724.375 430.035 724.390 ;
        RECT 430.625 724.375 430.955 724.390 ;
        RECT 429.245 676.410 429.575 676.425 ;
        RECT 430.165 676.410 430.495 676.425 ;
        RECT 429.245 676.110 430.495 676.410 ;
        RECT 429.245 676.095 429.575 676.110 ;
        RECT 430.165 676.095 430.495 676.110 ;
        RECT 429.705 628.130 430.035 628.145 ;
        RECT 430.625 628.130 430.955 628.145 ;
        RECT 429.705 627.830 430.955 628.130 ;
        RECT 429.705 627.815 430.035 627.830 ;
        RECT 430.625 627.815 430.955 627.830 ;
        RECT 429.245 579.850 429.575 579.865 ;
        RECT 430.165 579.850 430.495 579.865 ;
        RECT 429.245 579.550 430.495 579.850 ;
        RECT 429.245 579.535 429.575 579.550 ;
        RECT 430.165 579.535 430.495 579.550 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 396.590 1592.120 396.910 1592.180 ;
        RECT 437.530 1592.120 437.850 1592.180 ;
        RECT 396.590 1591.980 437.850 1592.120 ;
        RECT 396.590 1591.920 396.910 1591.980 ;
        RECT 437.530 1591.920 437.850 1591.980 ;
        RECT 365.310 19.960 365.630 20.020 ;
        RECT 396.590 19.960 396.910 20.020 ;
        RECT 365.310 19.820 396.910 19.960 ;
        RECT 365.310 19.760 365.630 19.820 ;
        RECT 396.590 19.760 396.910 19.820 ;
      LAYER via ;
        RECT 396.620 1591.920 396.880 1592.180 ;
        RECT 437.560 1591.920 437.820 1592.180 ;
        RECT 365.340 19.760 365.600 20.020 ;
        RECT 396.620 19.760 396.880 20.020 ;
      LAYER met2 ;
        RECT 437.560 1600.000 437.840 1604.000 ;
        RECT 437.620 1592.210 437.760 1600.000 ;
        RECT 396.620 1591.890 396.880 1592.210 ;
        RECT 437.560 1591.890 437.820 1592.210 ;
        RECT 396.680 20.050 396.820 1591.890 ;
        RECT 365.340 19.730 365.600 20.050 ;
        RECT 396.620 19.730 396.880 20.050 ;
        RECT 365.400 2.400 365.540 19.730 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 410.850 1587.700 411.170 1587.760 ;
        RECT 444.430 1587.700 444.750 1587.760 ;
        RECT 410.850 1587.560 444.750 1587.700 ;
        RECT 410.850 1587.500 411.170 1587.560 ;
        RECT 444.430 1587.500 444.750 1587.560 ;
        RECT 383.250 17.580 383.570 17.640 ;
        RECT 410.850 17.580 411.170 17.640 ;
        RECT 383.250 17.440 411.170 17.580 ;
        RECT 383.250 17.380 383.570 17.440 ;
        RECT 410.850 17.380 411.170 17.440 ;
      LAYER via ;
        RECT 410.880 1587.500 411.140 1587.760 ;
        RECT 444.460 1587.500 444.720 1587.760 ;
        RECT 383.280 17.380 383.540 17.640 ;
        RECT 410.880 17.380 411.140 17.640 ;
      LAYER met2 ;
        RECT 444.460 1600.000 444.740 1604.000 ;
        RECT 444.520 1587.790 444.660 1600.000 ;
        RECT 410.880 1587.470 411.140 1587.790 ;
        RECT 444.460 1587.470 444.720 1587.790 ;
        RECT 410.940 17.670 411.080 1587.470 ;
        RECT 383.280 17.350 383.540 17.670 ;
        RECT 410.880 17.350 411.140 17.670 ;
        RECT 383.340 2.400 383.480 17.350 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 410.390 1592.460 410.710 1592.520 ;
        RECT 450.870 1592.460 451.190 1592.520 ;
        RECT 410.390 1592.320 451.190 1592.460 ;
        RECT 410.390 1592.260 410.710 1592.320 ;
        RECT 450.870 1592.260 451.190 1592.320 ;
        RECT 401.190 20.640 401.510 20.700 ;
        RECT 410.390 20.640 410.710 20.700 ;
        RECT 401.190 20.500 410.710 20.640 ;
        RECT 401.190 20.440 401.510 20.500 ;
        RECT 410.390 20.440 410.710 20.500 ;
      LAYER via ;
        RECT 410.420 1592.260 410.680 1592.520 ;
        RECT 450.900 1592.260 451.160 1592.520 ;
        RECT 401.220 20.440 401.480 20.700 ;
        RECT 410.420 20.440 410.680 20.700 ;
      LAYER met2 ;
        RECT 450.900 1600.000 451.180 1604.000 ;
        RECT 450.960 1592.550 451.100 1600.000 ;
        RECT 410.420 1592.230 410.680 1592.550 ;
        RECT 450.900 1592.230 451.160 1592.550 ;
        RECT 410.480 20.730 410.620 1592.230 ;
        RECT 401.220 20.410 401.480 20.730 ;
        RECT 410.420 20.410 410.680 20.730 ;
        RECT 401.280 2.400 401.420 20.410 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 301.445 1590.265 301.615 1594.175 ;
        RECT 305.125 1592.645 305.295 1594.175 ;
      LAYER mcon ;
        RECT 301.445 1594.005 301.615 1594.175 ;
        RECT 305.125 1594.005 305.295 1594.175 ;
      LAYER met1 ;
        RECT 301.385 1594.160 301.675 1594.205 ;
        RECT 305.065 1594.160 305.355 1594.205 ;
        RECT 301.385 1594.020 305.355 1594.160 ;
        RECT 301.385 1593.975 301.675 1594.020 ;
        RECT 305.065 1593.975 305.355 1594.020 ;
        RECT 305.065 1592.800 305.355 1592.845 ;
        RECT 322.990 1592.800 323.310 1592.860 ;
        RECT 305.065 1592.660 323.310 1592.800 ;
        RECT 305.065 1592.615 305.355 1592.660 ;
        RECT 322.990 1592.600 323.310 1592.660 ;
        RECT 68.610 1590.420 68.930 1590.480 ;
        RECT 301.385 1590.420 301.675 1590.465 ;
        RECT 68.610 1590.280 301.675 1590.420 ;
        RECT 68.610 1590.220 68.930 1590.280 ;
        RECT 301.385 1590.235 301.675 1590.280 ;
        RECT 62.170 15.880 62.490 15.940 ;
        RECT 68.610 15.880 68.930 15.940 ;
        RECT 62.170 15.740 68.930 15.880 ;
        RECT 62.170 15.680 62.490 15.740 ;
        RECT 68.610 15.680 68.930 15.740 ;
      LAYER via ;
        RECT 323.020 1592.600 323.280 1592.860 ;
        RECT 68.640 1590.220 68.900 1590.480 ;
        RECT 62.200 15.680 62.460 15.940 ;
        RECT 68.640 15.680 68.900 15.940 ;
      LAYER met2 ;
        RECT 323.020 1600.000 323.300 1604.000 ;
        RECT 323.080 1592.890 323.220 1600.000 ;
        RECT 323.020 1592.570 323.280 1592.890 ;
        RECT 68.640 1590.190 68.900 1590.510 ;
        RECT 68.700 15.970 68.840 1590.190 ;
        RECT 62.200 15.650 62.460 15.970 ;
        RECT 68.640 15.650 68.900 15.970 ;
        RECT 62.260 2.400 62.400 15.650 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 424.190 1589.060 424.510 1589.120 ;
        RECT 457.770 1589.060 458.090 1589.120 ;
        RECT 424.190 1588.920 458.090 1589.060 ;
        RECT 424.190 1588.860 424.510 1588.920 ;
        RECT 457.770 1588.860 458.090 1588.920 ;
        RECT 419.130 20.640 419.450 20.700 ;
        RECT 424.190 20.640 424.510 20.700 ;
        RECT 419.130 20.500 424.510 20.640 ;
        RECT 419.130 20.440 419.450 20.500 ;
        RECT 424.190 20.440 424.510 20.500 ;
      LAYER via ;
        RECT 424.220 1588.860 424.480 1589.120 ;
        RECT 457.800 1588.860 458.060 1589.120 ;
        RECT 419.160 20.440 419.420 20.700 ;
        RECT 424.220 20.440 424.480 20.700 ;
      LAYER met2 ;
        RECT 457.800 1600.000 458.080 1604.000 ;
        RECT 457.860 1589.150 458.000 1600.000 ;
        RECT 424.220 1588.830 424.480 1589.150 ;
        RECT 457.800 1588.830 458.060 1589.150 ;
        RECT 424.280 20.730 424.420 1588.830 ;
        RECT 419.160 20.410 419.420 20.730 ;
        RECT 424.220 20.410 424.480 20.730 ;
        RECT 419.220 2.400 419.360 20.410 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 441.210 1590.080 441.530 1590.140 ;
        RECT 464.670 1590.080 464.990 1590.140 ;
        RECT 441.210 1589.940 464.990 1590.080 ;
        RECT 441.210 1589.880 441.530 1589.940 ;
        RECT 464.670 1589.880 464.990 1589.940 ;
        RECT 436.610 17.920 436.930 17.980 ;
        RECT 441.210 17.920 441.530 17.980 ;
        RECT 436.610 17.780 441.530 17.920 ;
        RECT 436.610 17.720 436.930 17.780 ;
        RECT 441.210 17.720 441.530 17.780 ;
      LAYER via ;
        RECT 441.240 1589.880 441.500 1590.140 ;
        RECT 464.700 1589.880 464.960 1590.140 ;
        RECT 436.640 17.720 436.900 17.980 ;
        RECT 441.240 17.720 441.500 17.980 ;
      LAYER met2 ;
        RECT 464.700 1600.000 464.980 1604.000 ;
        RECT 464.760 1590.170 464.900 1600.000 ;
        RECT 441.240 1589.850 441.500 1590.170 ;
        RECT 464.700 1589.850 464.960 1590.170 ;
        RECT 441.300 18.010 441.440 1589.850 ;
        RECT 436.640 17.690 436.900 18.010 ;
        RECT 441.240 17.690 441.500 18.010 ;
        RECT 436.700 2.400 436.840 17.690 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 455.010 1588.040 455.330 1588.100 ;
        RECT 471.110 1588.040 471.430 1588.100 ;
        RECT 455.010 1587.900 471.430 1588.040 ;
        RECT 455.010 1587.840 455.330 1587.900 ;
        RECT 471.110 1587.840 471.430 1587.900 ;
      LAYER via ;
        RECT 455.040 1587.840 455.300 1588.100 ;
        RECT 471.140 1587.840 471.400 1588.100 ;
      LAYER met2 ;
        RECT 471.140 1600.000 471.420 1604.000 ;
        RECT 471.200 1588.130 471.340 1600.000 ;
        RECT 455.040 1587.810 455.300 1588.130 ;
        RECT 471.140 1587.810 471.400 1588.130 ;
        RECT 455.100 3.130 455.240 1587.810 ;
        RECT 454.640 2.990 455.240 3.130 ;
        RECT 454.640 2.400 454.780 2.990 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 19.280 472.810 19.340 ;
        RECT 476.630 19.280 476.950 19.340 ;
        RECT 472.490 19.140 476.950 19.280 ;
        RECT 472.490 19.080 472.810 19.140 ;
        RECT 476.630 19.080 476.950 19.140 ;
      LAYER via ;
        RECT 472.520 19.080 472.780 19.340 ;
        RECT 476.660 19.080 476.920 19.340 ;
      LAYER met2 ;
        RECT 478.040 1600.450 478.320 1604.000 ;
        RECT 476.720 1600.310 478.320 1600.450 ;
        RECT 476.720 19.370 476.860 1600.310 ;
        RECT 478.040 1600.000 478.320 1600.310 ;
        RECT 472.520 19.050 472.780 19.370 ;
        RECT 476.660 19.050 476.920 19.370 ;
        RECT 472.580 2.400 472.720 19.050 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 484.910 1587.360 485.230 1587.420 ;
        RECT 488.590 1587.360 488.910 1587.420 ;
        RECT 484.910 1587.220 488.910 1587.360 ;
        RECT 484.910 1587.160 485.230 1587.220 ;
        RECT 488.590 1587.160 488.910 1587.220 ;
      LAYER via ;
        RECT 484.940 1587.160 485.200 1587.420 ;
        RECT 488.620 1587.160 488.880 1587.420 ;
      LAYER met2 ;
        RECT 484.940 1600.000 485.220 1604.000 ;
        RECT 485.000 1587.450 485.140 1600.000 ;
        RECT 484.940 1587.130 485.200 1587.450 ;
        RECT 488.620 1587.130 488.880 1587.450 ;
        RECT 488.680 16.730 488.820 1587.130 ;
        RECT 488.680 16.590 490.660 16.730 ;
        RECT 490.520 2.400 490.660 16.590 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 491.350 1589.400 491.670 1589.460 ;
        RECT 500.550 1589.400 500.870 1589.460 ;
        RECT 491.350 1589.260 500.870 1589.400 ;
        RECT 491.350 1589.200 491.670 1589.260 ;
        RECT 500.550 1589.200 500.870 1589.260 ;
        RECT 500.550 17.580 500.870 17.640 ;
        RECT 507.910 17.580 508.230 17.640 ;
        RECT 500.550 17.440 508.230 17.580 ;
        RECT 500.550 17.380 500.870 17.440 ;
        RECT 507.910 17.380 508.230 17.440 ;
      LAYER via ;
        RECT 491.380 1589.200 491.640 1589.460 ;
        RECT 500.580 1589.200 500.840 1589.460 ;
        RECT 500.580 17.380 500.840 17.640 ;
        RECT 507.940 17.380 508.200 17.640 ;
      LAYER met2 ;
        RECT 491.380 1600.000 491.660 1604.000 ;
        RECT 491.440 1589.490 491.580 1600.000 ;
        RECT 491.380 1589.170 491.640 1589.490 ;
        RECT 500.580 1589.170 500.840 1589.490 ;
        RECT 500.640 17.670 500.780 1589.170 ;
        RECT 500.580 17.350 500.840 17.670 ;
        RECT 507.940 17.350 508.200 17.670 ;
        RECT 508.000 2.400 508.140 17.350 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 498.250 1593.480 498.570 1593.540 ;
        RECT 525.850 1593.480 526.170 1593.540 ;
        RECT 498.250 1593.340 526.170 1593.480 ;
        RECT 498.250 1593.280 498.570 1593.340 ;
        RECT 525.850 1593.280 526.170 1593.340 ;
      LAYER via ;
        RECT 498.280 1593.280 498.540 1593.540 ;
        RECT 525.880 1593.280 526.140 1593.540 ;
      LAYER met2 ;
        RECT 498.280 1600.000 498.560 1604.000 ;
        RECT 498.340 1593.570 498.480 1600.000 ;
        RECT 498.280 1593.250 498.540 1593.570 ;
        RECT 525.880 1593.250 526.140 1593.570 ;
        RECT 525.940 2.400 526.080 1593.250 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 505.150 1588.720 505.470 1588.780 ;
        RECT 513.890 1588.720 514.210 1588.780 ;
        RECT 505.150 1588.580 514.210 1588.720 ;
        RECT 505.150 1588.520 505.470 1588.580 ;
        RECT 513.890 1588.520 514.210 1588.580 ;
        RECT 513.890 18.260 514.210 18.320 ;
        RECT 543.790 18.260 544.110 18.320 ;
        RECT 513.890 18.120 544.110 18.260 ;
        RECT 513.890 18.060 514.210 18.120 ;
        RECT 543.790 18.060 544.110 18.120 ;
      LAYER via ;
        RECT 505.180 1588.520 505.440 1588.780 ;
        RECT 513.920 1588.520 514.180 1588.780 ;
        RECT 513.920 18.060 514.180 18.320 ;
        RECT 543.820 18.060 544.080 18.320 ;
      LAYER met2 ;
        RECT 505.180 1600.000 505.460 1604.000 ;
        RECT 505.240 1588.810 505.380 1600.000 ;
        RECT 505.180 1588.490 505.440 1588.810 ;
        RECT 513.920 1588.490 514.180 1588.810 ;
        RECT 513.980 18.350 514.120 1588.490 ;
        RECT 513.920 18.030 514.180 18.350 ;
        RECT 543.820 18.030 544.080 18.350 ;
        RECT 543.880 2.400 544.020 18.030 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 511.590 1588.040 511.910 1588.100 ;
        RECT 521.250 1588.040 521.570 1588.100 ;
        RECT 511.590 1587.900 521.570 1588.040 ;
        RECT 511.590 1587.840 511.910 1587.900 ;
        RECT 521.250 1587.840 521.570 1587.900 ;
        RECT 521.250 16.900 521.570 16.960 ;
        RECT 561.730 16.900 562.050 16.960 ;
        RECT 521.250 16.760 562.050 16.900 ;
        RECT 521.250 16.700 521.570 16.760 ;
        RECT 561.730 16.700 562.050 16.760 ;
      LAYER via ;
        RECT 511.620 1587.840 511.880 1588.100 ;
        RECT 521.280 1587.840 521.540 1588.100 ;
        RECT 521.280 16.700 521.540 16.960 ;
        RECT 561.760 16.700 562.020 16.960 ;
      LAYER met2 ;
        RECT 511.620 1600.000 511.900 1604.000 ;
        RECT 511.680 1588.130 511.820 1600.000 ;
        RECT 511.620 1587.810 511.880 1588.130 ;
        RECT 521.280 1587.810 521.540 1588.130 ;
        RECT 521.340 16.990 521.480 1587.810 ;
        RECT 521.280 16.670 521.540 16.990 ;
        RECT 561.760 16.670 562.020 16.990 ;
        RECT 561.820 2.400 561.960 16.670 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 518.490 1587.360 518.810 1587.420 ;
        RECT 523.550 1587.360 523.870 1587.420 ;
        RECT 518.490 1587.220 523.870 1587.360 ;
        RECT 518.490 1587.160 518.810 1587.220 ;
        RECT 523.550 1587.160 523.870 1587.220 ;
        RECT 523.550 18.600 523.870 18.660 ;
        RECT 523.550 18.460 544.480 18.600 ;
        RECT 523.550 18.400 523.870 18.460 ;
        RECT 544.340 18.260 544.480 18.460 ;
        RECT 544.340 18.120 550.460 18.260 ;
        RECT 550.320 17.580 550.460 18.120 ;
        RECT 550.320 17.440 556.440 17.580 ;
        RECT 556.300 17.240 556.440 17.440 ;
        RECT 556.300 17.100 562.880 17.240 ;
        RECT 562.740 16.560 562.880 17.100 ;
        RECT 579.670 16.560 579.990 16.620 ;
        RECT 562.740 16.420 579.990 16.560 ;
        RECT 579.670 16.360 579.990 16.420 ;
      LAYER via ;
        RECT 518.520 1587.160 518.780 1587.420 ;
        RECT 523.580 1587.160 523.840 1587.420 ;
        RECT 523.580 18.400 523.840 18.660 ;
        RECT 579.700 16.360 579.960 16.620 ;
      LAYER met2 ;
        RECT 518.520 1600.000 518.800 1604.000 ;
        RECT 518.580 1587.450 518.720 1600.000 ;
        RECT 518.520 1587.130 518.780 1587.450 ;
        RECT 523.580 1587.130 523.840 1587.450 ;
        RECT 523.640 18.690 523.780 1587.130 ;
        RECT 523.580 18.370 523.840 18.690 ;
        RECT 579.700 16.330 579.960 16.650 ;
        RECT 579.760 2.400 579.900 16.330 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 89.310 1590.760 89.630 1590.820 ;
        RECT 332.190 1590.760 332.510 1590.820 ;
        RECT 89.310 1590.620 332.510 1590.760 ;
        RECT 89.310 1590.560 89.630 1590.620 ;
        RECT 332.190 1590.560 332.510 1590.620 ;
        RECT 86.090 16.900 86.410 16.960 ;
        RECT 89.310 16.900 89.630 16.960 ;
        RECT 86.090 16.760 89.630 16.900 ;
        RECT 86.090 16.700 86.410 16.760 ;
        RECT 89.310 16.700 89.630 16.760 ;
      LAYER via ;
        RECT 89.340 1590.560 89.600 1590.820 ;
        RECT 332.220 1590.560 332.480 1590.820 ;
        RECT 86.120 16.700 86.380 16.960 ;
        RECT 89.340 16.700 89.600 16.960 ;
      LAYER met2 ;
        RECT 332.220 1600.000 332.500 1604.000 ;
        RECT 332.280 1590.850 332.420 1600.000 ;
        RECT 89.340 1590.530 89.600 1590.850 ;
        RECT 332.220 1590.530 332.480 1590.850 ;
        RECT 89.400 16.990 89.540 1590.530 ;
        RECT 86.120 16.670 86.380 16.990 ;
        RECT 89.340 16.670 89.600 16.990 ;
        RECT 86.180 2.400 86.320 16.670 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 562.265 16.745 563.355 16.915 ;
        RECT 562.265 16.405 562.435 16.745 ;
      LAYER mcon ;
        RECT 563.185 16.745 563.355 16.915 ;
      LAYER met1 ;
        RECT 524.930 1590.420 525.250 1590.480 ;
        RECT 528.610 1590.420 528.930 1590.480 ;
        RECT 524.930 1590.280 528.930 1590.420 ;
        RECT 524.930 1590.220 525.250 1590.280 ;
        RECT 528.610 1590.220 528.930 1590.280 ;
        RECT 563.125 16.900 563.415 16.945 ;
        RECT 597.150 16.900 597.470 16.960 ;
        RECT 563.125 16.760 597.470 16.900 ;
        RECT 563.125 16.715 563.415 16.760 ;
        RECT 597.150 16.700 597.470 16.760 ;
        RECT 529.990 16.560 530.310 16.620 ;
        RECT 562.205 16.560 562.495 16.605 ;
        RECT 529.990 16.420 562.495 16.560 ;
        RECT 529.990 16.360 530.310 16.420 ;
        RECT 562.205 16.375 562.495 16.420 ;
      LAYER via ;
        RECT 524.960 1590.220 525.220 1590.480 ;
        RECT 528.640 1590.220 528.900 1590.480 ;
        RECT 597.180 16.700 597.440 16.960 ;
        RECT 530.020 16.360 530.280 16.620 ;
      LAYER met2 ;
        RECT 524.960 1600.000 525.240 1604.000 ;
        RECT 525.020 1590.510 525.160 1600.000 ;
        RECT 524.960 1590.190 525.220 1590.510 ;
        RECT 528.640 1590.190 528.900 1590.510 ;
        RECT 528.700 1582.090 528.840 1590.190 ;
        RECT 528.700 1581.950 530.220 1582.090 ;
        RECT 530.080 16.650 530.220 1581.950 ;
        RECT 597.180 16.670 597.440 16.990 ;
        RECT 530.020 16.330 530.280 16.650 ;
        RECT 597.240 2.400 597.380 16.670 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 604.125 18.445 604.295 19.635 ;
      LAYER mcon ;
        RECT 604.125 19.465 604.295 19.635 ;
      LAYER met1 ;
        RECT 531.830 1588.040 532.150 1588.100 ;
        RECT 537.810 1588.040 538.130 1588.100 ;
        RECT 531.830 1587.900 538.130 1588.040 ;
        RECT 531.830 1587.840 532.150 1587.900 ;
        RECT 537.810 1587.840 538.130 1587.900 ;
        RECT 537.810 19.620 538.130 19.680 ;
        RECT 604.065 19.620 604.355 19.665 ;
        RECT 537.810 19.480 604.355 19.620 ;
        RECT 537.810 19.420 538.130 19.480 ;
        RECT 604.065 19.435 604.355 19.480 ;
        RECT 604.065 18.600 604.355 18.645 ;
        RECT 615.090 18.600 615.410 18.660 ;
        RECT 604.065 18.460 615.410 18.600 ;
        RECT 604.065 18.415 604.355 18.460 ;
        RECT 615.090 18.400 615.410 18.460 ;
      LAYER via ;
        RECT 531.860 1587.840 532.120 1588.100 ;
        RECT 537.840 1587.840 538.100 1588.100 ;
        RECT 537.840 19.420 538.100 19.680 ;
        RECT 615.120 18.400 615.380 18.660 ;
      LAYER met2 ;
        RECT 531.860 1600.000 532.140 1604.000 ;
        RECT 531.920 1588.130 532.060 1600.000 ;
        RECT 531.860 1587.810 532.120 1588.130 ;
        RECT 537.840 1587.810 538.100 1588.130 ;
        RECT 537.900 19.710 538.040 1587.810 ;
        RECT 537.840 19.390 538.100 19.710 ;
        RECT 615.120 18.370 615.380 18.690 ;
        RECT 615.180 2.400 615.320 18.370 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 1591.440 109.870 1591.500 ;
        RECT 303.670 1591.440 303.990 1591.500 ;
        RECT 109.550 1591.300 303.990 1591.440 ;
        RECT 109.550 1591.240 109.870 1591.300 ;
        RECT 303.670 1591.240 303.990 1591.300 ;
        RECT 303.670 1590.420 303.990 1590.480 ;
        RECT 340.930 1590.420 341.250 1590.480 ;
        RECT 303.670 1590.280 341.250 1590.420 ;
        RECT 303.670 1590.220 303.990 1590.280 ;
        RECT 340.930 1590.220 341.250 1590.280 ;
      LAYER via ;
        RECT 109.580 1591.240 109.840 1591.500 ;
        RECT 303.700 1591.240 303.960 1591.500 ;
        RECT 303.700 1590.220 303.960 1590.480 ;
        RECT 340.960 1590.220 341.220 1590.480 ;
      LAYER met2 ;
        RECT 340.960 1600.000 341.240 1604.000 ;
        RECT 109.580 1591.210 109.840 1591.530 ;
        RECT 303.700 1591.210 303.960 1591.530 ;
        RECT 109.640 2.400 109.780 1591.210 ;
        RECT 303.760 1590.510 303.900 1591.210 ;
        RECT 341.020 1590.510 341.160 1600.000 ;
        RECT 303.700 1590.190 303.960 1590.510 ;
        RECT 340.960 1590.190 341.220 1590.510 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 303.745 1592.305 304.375 1592.475 ;
        RECT 304.205 1591.285 304.375 1592.305 ;
      LAYER met1 ;
        RECT 137.610 1592.460 137.930 1592.520 ;
        RECT 303.685 1592.460 303.975 1592.505 ;
        RECT 137.610 1592.320 303.975 1592.460 ;
        RECT 137.610 1592.260 137.930 1592.320 ;
        RECT 303.685 1592.275 303.975 1592.320 ;
        RECT 304.145 1591.440 304.435 1591.485 ;
        RECT 350.130 1591.440 350.450 1591.500 ;
        RECT 304.145 1591.300 350.450 1591.440 ;
        RECT 304.145 1591.255 304.435 1591.300 ;
        RECT 350.130 1591.240 350.450 1591.300 ;
        RECT 133.470 16.900 133.790 16.960 ;
        RECT 137.610 16.900 137.930 16.960 ;
        RECT 133.470 16.760 137.930 16.900 ;
        RECT 133.470 16.700 133.790 16.760 ;
        RECT 137.610 16.700 137.930 16.760 ;
      LAYER via ;
        RECT 137.640 1592.260 137.900 1592.520 ;
        RECT 350.160 1591.240 350.420 1591.500 ;
        RECT 133.500 16.700 133.760 16.960 ;
        RECT 137.640 16.700 137.900 16.960 ;
      LAYER met2 ;
        RECT 350.160 1600.000 350.440 1604.000 ;
        RECT 137.640 1592.230 137.900 1592.550 ;
        RECT 137.700 16.990 137.840 1592.230 ;
        RECT 350.220 1591.530 350.360 1600.000 ;
        RECT 350.160 1591.210 350.420 1591.530 ;
        RECT 133.500 16.670 133.760 16.990 ;
        RECT 137.640 16.670 137.900 16.990 ;
        RECT 133.560 2.400 133.700 16.670 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 150.950 1593.140 151.270 1593.200 ;
        RECT 356.570 1593.140 356.890 1593.200 ;
        RECT 150.950 1593.000 356.890 1593.140 ;
        RECT 150.950 1592.940 151.270 1593.000 ;
        RECT 356.570 1592.940 356.890 1593.000 ;
      LAYER via ;
        RECT 150.980 1592.940 151.240 1593.200 ;
        RECT 356.600 1592.940 356.860 1593.200 ;
      LAYER met2 ;
        RECT 356.600 1600.000 356.880 1604.000 ;
        RECT 356.660 1593.230 356.800 1600.000 ;
        RECT 150.980 1592.910 151.240 1593.230 ;
        RECT 356.600 1592.910 356.860 1593.230 ;
        RECT 151.040 17.410 151.180 1592.910 ;
        RECT 151.040 17.270 151.640 17.410 ;
        RECT 151.500 2.400 151.640 17.270 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 361.245 1449.165 361.415 1463.275 ;
        RECT 361.245 1352.605 361.415 1400.715 ;
        RECT 361.245 1256.045 361.415 1304.155 ;
        RECT 361.245 565.845 361.415 613.955 ;
        RECT 361.245 462.485 361.415 510.595 ;
        RECT 362.165 282.625 362.335 324.275 ;
        RECT 361.705 228.225 361.875 275.995 ;
        RECT 361.705 158.525 361.875 227.715 ;
        RECT 346.065 16.405 346.235 19.975 ;
      LAYER mcon ;
        RECT 361.245 1463.105 361.415 1463.275 ;
        RECT 361.245 1400.545 361.415 1400.715 ;
        RECT 361.245 1303.985 361.415 1304.155 ;
        RECT 361.245 613.785 361.415 613.955 ;
        RECT 361.245 510.425 361.415 510.595 ;
        RECT 362.165 324.105 362.335 324.275 ;
        RECT 361.705 275.825 361.875 275.995 ;
        RECT 361.705 227.545 361.875 227.715 ;
        RECT 346.065 19.805 346.235 19.975 ;
      LAYER met1 ;
        RECT 361.185 1463.260 361.475 1463.305 ;
        RECT 361.630 1463.260 361.950 1463.320 ;
        RECT 361.185 1463.120 361.950 1463.260 ;
        RECT 361.185 1463.075 361.475 1463.120 ;
        RECT 361.630 1463.060 361.950 1463.120 ;
        RECT 361.170 1449.320 361.490 1449.380 ;
        RECT 360.975 1449.180 361.490 1449.320 ;
        RECT 361.170 1449.120 361.490 1449.180 ;
        RECT 361.170 1400.700 361.490 1400.760 ;
        RECT 360.975 1400.560 361.490 1400.700 ;
        RECT 361.170 1400.500 361.490 1400.560 ;
        RECT 361.170 1352.760 361.490 1352.820 ;
        RECT 360.975 1352.620 361.490 1352.760 ;
        RECT 361.170 1352.560 361.490 1352.620 ;
        RECT 361.170 1304.140 361.490 1304.200 ;
        RECT 360.975 1304.000 361.490 1304.140 ;
        RECT 361.170 1303.940 361.490 1304.000 ;
        RECT 361.170 1256.200 361.490 1256.260 ;
        RECT 360.975 1256.060 361.490 1256.200 ;
        RECT 361.170 1256.000 361.490 1256.060 ;
        RECT 360.250 1159.300 360.570 1159.360 ;
        RECT 361.170 1159.300 361.490 1159.360 ;
        RECT 360.250 1159.160 361.490 1159.300 ;
        RECT 360.250 1159.100 360.570 1159.160 ;
        RECT 361.170 1159.100 361.490 1159.160 ;
        RECT 360.250 1062.740 360.570 1062.800 ;
        RECT 361.170 1062.740 361.490 1062.800 ;
        RECT 360.250 1062.600 361.490 1062.740 ;
        RECT 360.250 1062.540 360.570 1062.600 ;
        RECT 361.170 1062.540 361.490 1062.600 ;
        RECT 360.250 966.180 360.570 966.240 ;
        RECT 361.170 966.180 361.490 966.240 ;
        RECT 360.250 966.040 361.490 966.180 ;
        RECT 360.250 965.980 360.570 966.040 ;
        RECT 361.170 965.980 361.490 966.040 ;
        RECT 360.250 869.620 360.570 869.680 ;
        RECT 361.170 869.620 361.490 869.680 ;
        RECT 360.250 869.480 361.490 869.620 ;
        RECT 360.250 869.420 360.570 869.480 ;
        RECT 361.170 869.420 361.490 869.480 ;
        RECT 361.170 613.940 361.490 614.000 ;
        RECT 360.975 613.800 361.490 613.940 ;
        RECT 361.170 613.740 361.490 613.800 ;
        RECT 361.170 566.000 361.490 566.060 ;
        RECT 360.975 565.860 361.490 566.000 ;
        RECT 361.170 565.800 361.490 565.860 ;
        RECT 361.185 510.580 361.475 510.625 ;
        RECT 361.630 510.580 361.950 510.640 ;
        RECT 361.185 510.440 361.950 510.580 ;
        RECT 361.185 510.395 361.475 510.440 ;
        RECT 361.630 510.380 361.950 510.440 ;
        RECT 361.170 462.640 361.490 462.700 ;
        RECT 360.975 462.500 361.490 462.640 ;
        RECT 361.170 462.440 361.490 462.500 ;
        RECT 360.710 331.060 361.030 331.120 ;
        RECT 362.090 331.060 362.410 331.120 ;
        RECT 360.710 330.920 362.410 331.060 ;
        RECT 360.710 330.860 361.030 330.920 ;
        RECT 362.090 330.860 362.410 330.920 ;
        RECT 362.090 324.260 362.410 324.320 ;
        RECT 361.895 324.120 362.410 324.260 ;
        RECT 362.090 324.060 362.410 324.120 ;
        RECT 362.090 282.780 362.410 282.840 ;
        RECT 361.895 282.640 362.410 282.780 ;
        RECT 362.090 282.580 362.410 282.640 ;
        RECT 361.645 275.980 361.935 276.025 ;
        RECT 362.090 275.980 362.410 276.040 ;
        RECT 361.645 275.840 362.410 275.980 ;
        RECT 361.645 275.795 361.935 275.840 ;
        RECT 362.090 275.780 362.410 275.840 ;
        RECT 361.630 228.380 361.950 228.440 ;
        RECT 361.435 228.240 361.950 228.380 ;
        RECT 361.630 228.180 361.950 228.240 ;
        RECT 361.630 227.700 361.950 227.760 ;
        RECT 361.435 227.560 361.950 227.700 ;
        RECT 361.630 227.500 361.950 227.560 ;
        RECT 360.710 158.680 361.030 158.740 ;
        RECT 361.645 158.680 361.935 158.725 ;
        RECT 360.710 158.540 361.935 158.680 ;
        RECT 360.710 158.480 361.030 158.540 ;
        RECT 361.645 158.495 361.935 158.540 ;
        RECT 360.710 137.740 361.030 138.000 ;
        RECT 360.800 137.600 360.940 137.740 ;
        RECT 361.630 137.600 361.950 137.660 ;
        RECT 360.800 137.460 361.950 137.600 ;
        RECT 361.630 137.400 361.950 137.460 ;
        RECT 360.250 48.520 360.570 48.580 ;
        RECT 361.630 48.520 361.950 48.580 ;
        RECT 360.250 48.380 361.950 48.520 ;
        RECT 360.250 48.320 360.570 48.380 ;
        RECT 361.630 48.320 361.950 48.380 ;
        RECT 346.005 19.960 346.295 20.005 ;
        RECT 360.250 19.960 360.570 20.020 ;
        RECT 346.005 19.820 360.570 19.960 ;
        RECT 346.005 19.775 346.295 19.820 ;
        RECT 360.250 19.760 360.570 19.820 ;
        RECT 169.350 16.900 169.670 16.960 ;
        RECT 169.350 16.760 328.280 16.900 ;
        RECT 169.350 16.700 169.670 16.760 ;
        RECT 328.140 16.560 328.280 16.760 ;
        RECT 346.005 16.560 346.295 16.605 ;
        RECT 328.140 16.420 346.295 16.560 ;
        RECT 346.005 16.375 346.295 16.420 ;
      LAYER via ;
        RECT 361.660 1463.060 361.920 1463.320 ;
        RECT 361.200 1449.120 361.460 1449.380 ;
        RECT 361.200 1400.500 361.460 1400.760 ;
        RECT 361.200 1352.560 361.460 1352.820 ;
        RECT 361.200 1303.940 361.460 1304.200 ;
        RECT 361.200 1256.000 361.460 1256.260 ;
        RECT 360.280 1159.100 360.540 1159.360 ;
        RECT 361.200 1159.100 361.460 1159.360 ;
        RECT 360.280 1062.540 360.540 1062.800 ;
        RECT 361.200 1062.540 361.460 1062.800 ;
        RECT 360.280 965.980 360.540 966.240 ;
        RECT 361.200 965.980 361.460 966.240 ;
        RECT 360.280 869.420 360.540 869.680 ;
        RECT 361.200 869.420 361.460 869.680 ;
        RECT 361.200 613.740 361.460 614.000 ;
        RECT 361.200 565.800 361.460 566.060 ;
        RECT 361.660 510.380 361.920 510.640 ;
        RECT 361.200 462.440 361.460 462.700 ;
        RECT 360.740 330.860 361.000 331.120 ;
        RECT 362.120 330.860 362.380 331.120 ;
        RECT 362.120 324.060 362.380 324.320 ;
        RECT 362.120 282.580 362.380 282.840 ;
        RECT 362.120 275.780 362.380 276.040 ;
        RECT 361.660 228.180 361.920 228.440 ;
        RECT 361.660 227.500 361.920 227.760 ;
        RECT 360.740 158.480 361.000 158.740 ;
        RECT 360.740 137.740 361.000 138.000 ;
        RECT 361.660 137.400 361.920 137.660 ;
        RECT 360.280 48.320 360.540 48.580 ;
        RECT 361.660 48.320 361.920 48.580 ;
        RECT 360.280 19.760 360.540 20.020 ;
        RECT 169.380 16.700 169.640 16.960 ;
      LAYER met2 ;
        RECT 363.500 1600.450 363.780 1604.000 ;
        RECT 361.720 1600.310 363.780 1600.450 ;
        RECT 361.720 1463.350 361.860 1600.310 ;
        RECT 363.500 1600.000 363.780 1600.310 ;
        RECT 361.660 1463.030 361.920 1463.350 ;
        RECT 361.200 1449.090 361.460 1449.410 ;
        RECT 361.260 1400.790 361.400 1449.090 ;
        RECT 361.200 1400.470 361.460 1400.790 ;
        RECT 361.200 1352.530 361.460 1352.850 ;
        RECT 361.260 1304.230 361.400 1352.530 ;
        RECT 361.200 1303.910 361.460 1304.230 ;
        RECT 361.200 1255.970 361.460 1256.290 ;
        RECT 361.260 1207.525 361.400 1255.970 ;
        RECT 360.270 1207.155 360.550 1207.525 ;
        RECT 361.190 1207.155 361.470 1207.525 ;
        RECT 360.340 1159.390 360.480 1207.155 ;
        RECT 360.280 1159.070 360.540 1159.390 ;
        RECT 361.200 1159.070 361.460 1159.390 ;
        RECT 361.260 1110.965 361.400 1159.070 ;
        RECT 360.270 1110.595 360.550 1110.965 ;
        RECT 361.190 1110.595 361.470 1110.965 ;
        RECT 360.340 1062.830 360.480 1110.595 ;
        RECT 360.280 1062.510 360.540 1062.830 ;
        RECT 361.200 1062.510 361.460 1062.830 ;
        RECT 361.260 1014.405 361.400 1062.510 ;
        RECT 360.270 1014.035 360.550 1014.405 ;
        RECT 361.190 1014.035 361.470 1014.405 ;
        RECT 360.340 966.270 360.480 1014.035 ;
        RECT 360.280 965.950 360.540 966.270 ;
        RECT 361.200 965.950 361.460 966.270 ;
        RECT 361.260 917.845 361.400 965.950 ;
        RECT 360.270 917.475 360.550 917.845 ;
        RECT 361.190 917.475 361.470 917.845 ;
        RECT 360.340 869.710 360.480 917.475 ;
        RECT 360.280 869.390 360.540 869.710 ;
        RECT 361.200 869.390 361.460 869.710 ;
        RECT 361.260 787.170 361.400 869.390 ;
        RECT 360.800 787.030 361.400 787.170 ;
        RECT 360.800 786.490 360.940 787.030 ;
        RECT 360.800 786.350 361.400 786.490 ;
        RECT 361.260 725.405 361.400 786.350 ;
        RECT 361.190 725.035 361.470 725.405 ;
        RECT 361.190 724.355 361.470 724.725 ;
        RECT 361.260 628.845 361.400 724.355 ;
        RECT 361.190 628.475 361.470 628.845 ;
        RECT 361.190 627.795 361.470 628.165 ;
        RECT 361.260 614.030 361.400 627.795 ;
        RECT 361.200 613.710 361.460 614.030 ;
        RECT 361.200 565.770 361.460 566.090 ;
        RECT 361.260 524.180 361.400 565.770 ;
        RECT 361.260 524.040 361.860 524.180 ;
        RECT 361.720 510.670 361.860 524.040 ;
        RECT 361.660 510.350 361.920 510.670 ;
        RECT 361.200 462.410 361.460 462.730 ;
        RECT 361.260 355.370 361.400 462.410 ;
        RECT 360.800 355.230 361.400 355.370 ;
        RECT 360.800 331.150 360.940 355.230 ;
        RECT 360.740 330.830 361.000 331.150 ;
        RECT 362.120 330.830 362.380 331.150 ;
        RECT 362.180 324.350 362.320 330.830 ;
        RECT 362.120 324.030 362.380 324.350 ;
        RECT 362.120 282.550 362.380 282.870 ;
        RECT 362.180 276.070 362.320 282.550 ;
        RECT 362.120 275.750 362.380 276.070 ;
        RECT 361.660 228.150 361.920 228.470 ;
        RECT 361.720 227.790 361.860 228.150 ;
        RECT 361.660 227.470 361.920 227.790 ;
        RECT 360.740 158.450 361.000 158.770 ;
        RECT 360.800 138.030 360.940 158.450 ;
        RECT 360.740 137.710 361.000 138.030 ;
        RECT 361.660 137.370 361.920 137.690 ;
        RECT 361.720 48.610 361.860 137.370 ;
        RECT 360.280 48.290 360.540 48.610 ;
        RECT 361.660 48.290 361.920 48.610 ;
        RECT 360.340 20.050 360.480 48.290 ;
        RECT 360.280 19.730 360.540 20.050 ;
        RECT 169.380 16.670 169.640 16.990 ;
        RECT 169.440 2.400 169.580 16.670 ;
        RECT 169.230 -4.800 169.790 2.400 ;
      LAYER via2 ;
        RECT 360.270 1207.200 360.550 1207.480 ;
        RECT 361.190 1207.200 361.470 1207.480 ;
        RECT 360.270 1110.640 360.550 1110.920 ;
        RECT 361.190 1110.640 361.470 1110.920 ;
        RECT 360.270 1014.080 360.550 1014.360 ;
        RECT 361.190 1014.080 361.470 1014.360 ;
        RECT 360.270 917.520 360.550 917.800 ;
        RECT 361.190 917.520 361.470 917.800 ;
        RECT 361.190 725.080 361.470 725.360 ;
        RECT 361.190 724.400 361.470 724.680 ;
        RECT 361.190 628.520 361.470 628.800 ;
        RECT 361.190 627.840 361.470 628.120 ;
      LAYER met3 ;
        RECT 360.245 1207.490 360.575 1207.505 ;
        RECT 361.165 1207.490 361.495 1207.505 ;
        RECT 360.245 1207.190 361.495 1207.490 ;
        RECT 360.245 1207.175 360.575 1207.190 ;
        RECT 361.165 1207.175 361.495 1207.190 ;
        RECT 360.245 1110.930 360.575 1110.945 ;
        RECT 361.165 1110.930 361.495 1110.945 ;
        RECT 360.245 1110.630 361.495 1110.930 ;
        RECT 360.245 1110.615 360.575 1110.630 ;
        RECT 361.165 1110.615 361.495 1110.630 ;
        RECT 360.245 1014.370 360.575 1014.385 ;
        RECT 361.165 1014.370 361.495 1014.385 ;
        RECT 360.245 1014.070 361.495 1014.370 ;
        RECT 360.245 1014.055 360.575 1014.070 ;
        RECT 361.165 1014.055 361.495 1014.070 ;
        RECT 360.245 917.810 360.575 917.825 ;
        RECT 361.165 917.810 361.495 917.825 ;
        RECT 360.245 917.510 361.495 917.810 ;
        RECT 360.245 917.495 360.575 917.510 ;
        RECT 361.165 917.495 361.495 917.510 ;
        RECT 361.165 725.370 361.495 725.385 ;
        RECT 361.165 725.070 362.170 725.370 ;
        RECT 361.165 725.055 361.495 725.070 ;
        RECT 361.165 724.690 361.495 724.705 ;
        RECT 361.870 724.690 362.170 725.070 ;
        RECT 361.165 724.390 362.170 724.690 ;
        RECT 361.165 724.375 361.495 724.390 ;
        RECT 361.165 628.810 361.495 628.825 ;
        RECT 361.165 628.510 362.170 628.810 ;
        RECT 361.165 628.495 361.495 628.510 ;
        RECT 361.165 628.130 361.495 628.145 ;
        RECT 361.870 628.130 362.170 628.510 ;
        RECT 361.165 627.830 362.170 628.130 ;
        RECT 361.165 627.815 361.495 627.830 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.810 1589.060 193.130 1589.120 ;
        RECT 370.370 1589.060 370.690 1589.120 ;
        RECT 192.810 1588.920 370.690 1589.060 ;
        RECT 192.810 1588.860 193.130 1588.920 ;
        RECT 370.370 1588.860 370.690 1588.920 ;
        RECT 186.830 20.640 187.150 20.700 ;
        RECT 192.810 20.640 193.130 20.700 ;
        RECT 186.830 20.500 193.130 20.640 ;
        RECT 186.830 20.440 187.150 20.500 ;
        RECT 192.810 20.440 193.130 20.500 ;
      LAYER via ;
        RECT 192.840 1588.860 193.100 1589.120 ;
        RECT 370.400 1588.860 370.660 1589.120 ;
        RECT 186.860 20.440 187.120 20.700 ;
        RECT 192.840 20.440 193.100 20.700 ;
      LAYER met2 ;
        RECT 370.400 1600.000 370.680 1604.000 ;
        RECT 370.460 1589.150 370.600 1600.000 ;
        RECT 192.840 1588.830 193.100 1589.150 ;
        RECT 370.400 1588.830 370.660 1589.150 ;
        RECT 192.900 20.730 193.040 1588.830 ;
        RECT 186.860 20.410 187.120 20.730 ;
        RECT 192.840 20.410 193.100 20.730 ;
        RECT 186.920 2.400 187.060 20.410 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.840 1600.450 377.120 1604.000 ;
        RECT 375.520 1600.310 377.120 1600.450 ;
        RECT 375.520 1580.050 375.660 1600.310 ;
        RECT 376.840 1600.000 377.120 1600.310 ;
        RECT 373.680 1579.910 375.660 1580.050 ;
        RECT 373.680 20.245 373.820 1579.910 ;
        RECT 204.790 19.875 205.070 20.245 ;
        RECT 373.610 19.875 373.890 20.245 ;
        RECT 204.860 2.400 205.000 19.875 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 204.790 19.920 205.070 20.200 ;
        RECT 373.610 19.920 373.890 20.200 ;
      LAYER met3 ;
        RECT 204.765 20.210 205.095 20.225 ;
        RECT 373.585 20.210 373.915 20.225 ;
        RECT 204.765 19.910 373.915 20.210 ;
        RECT 204.765 19.895 205.095 19.910 ;
        RECT 373.585 19.895 373.915 19.910 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 227.310 1588.720 227.630 1588.780 ;
        RECT 383.710 1588.720 384.030 1588.780 ;
        RECT 227.310 1588.580 384.030 1588.720 ;
        RECT 227.310 1588.520 227.630 1588.580 ;
        RECT 383.710 1588.520 384.030 1588.580 ;
        RECT 222.710 16.560 223.030 16.620 ;
        RECT 227.310 16.560 227.630 16.620 ;
        RECT 222.710 16.420 227.630 16.560 ;
        RECT 222.710 16.360 223.030 16.420 ;
        RECT 227.310 16.360 227.630 16.420 ;
      LAYER via ;
        RECT 227.340 1588.520 227.600 1588.780 ;
        RECT 383.740 1588.520 384.000 1588.780 ;
        RECT 222.740 16.360 223.000 16.620 ;
        RECT 227.340 16.360 227.600 16.620 ;
      LAYER met2 ;
        RECT 383.740 1600.000 384.020 1604.000 ;
        RECT 383.800 1588.810 383.940 1600.000 ;
        RECT 227.340 1588.490 227.600 1588.810 ;
        RECT 383.740 1588.490 384.000 1588.810 ;
        RECT 227.400 16.650 227.540 1588.490 ;
        RECT 222.740 16.330 223.000 16.650 ;
        RECT 227.340 16.330 227.600 16.650 ;
        RECT 222.800 2.400 222.940 16.330 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 303.670 1579.880 303.990 1579.940 ;
        RECT 305.510 1579.880 305.830 1579.940 ;
        RECT 303.670 1579.740 305.830 1579.880 ;
        RECT 303.670 1579.680 303.990 1579.740 ;
        RECT 305.510 1579.680 305.830 1579.740 ;
      LAYER via ;
        RECT 303.700 1579.680 303.960 1579.940 ;
        RECT 305.540 1579.680 305.800 1579.940 ;
      LAYER met2 ;
        RECT 307.380 1600.450 307.660 1604.000 ;
        RECT 305.600 1600.310 307.660 1600.450 ;
        RECT 305.600 1579.970 305.740 1600.310 ;
        RECT 307.380 1600.000 307.660 1600.310 ;
        RECT 303.700 1579.650 303.960 1579.970 ;
        RECT 305.540 1579.650 305.800 1579.970 ;
        RECT 303.760 17.525 303.900 1579.650 ;
        RECT 20.330 17.155 20.610 17.525 ;
        RECT 303.690 17.155 303.970 17.525 ;
        RECT 20.400 2.400 20.540 17.155 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 20.330 17.200 20.610 17.480 ;
        RECT 303.690 17.200 303.970 17.480 ;
      LAYER met3 ;
        RECT 20.305 17.490 20.635 17.505 ;
        RECT 303.665 17.490 303.995 17.505 ;
        RECT 20.305 17.190 303.995 17.490 ;
        RECT 20.305 17.175 20.635 17.190 ;
        RECT 303.665 17.175 303.995 17.190 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.230 15.540 44.550 15.600 ;
        RECT 47.910 15.540 48.230 15.600 ;
        RECT 44.230 15.400 48.230 15.540 ;
        RECT 44.230 15.340 44.550 15.400 ;
        RECT 47.910 15.340 48.230 15.400 ;
      LAYER via ;
        RECT 44.260 15.340 44.520 15.600 ;
        RECT 47.940 15.340 48.200 15.600 ;
      LAYER met2 ;
        RECT 316.580 1600.000 316.860 1604.000 ;
        RECT 316.640 1591.045 316.780 1600.000 ;
        RECT 47.930 1590.675 48.210 1591.045 ;
        RECT 316.570 1590.675 316.850 1591.045 ;
        RECT 48.000 15.630 48.140 1590.675 ;
        RECT 44.260 15.310 44.520 15.630 ;
        RECT 47.940 15.310 48.200 15.630 ;
        RECT 44.320 2.400 44.460 15.310 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 47.930 1590.720 48.210 1591.000 ;
        RECT 316.570 1590.720 316.850 1591.000 ;
      LAYER met3 ;
        RECT 47.905 1591.010 48.235 1591.025 ;
        RECT 316.545 1591.010 316.875 1591.025 ;
        RECT 47.905 1590.710 316.875 1591.010 ;
        RECT 47.905 1590.695 48.235 1590.710 ;
        RECT 316.545 1590.695 316.875 1590.710 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 387.925 1497.445 388.095 1545.555 ;
        RECT 387.925 1352.605 388.095 1414.655 ;
        RECT 387.925 1256.045 388.095 1304.155 ;
        RECT 387.925 524.365 388.095 572.475 ;
        RECT 387.465 241.825 387.635 331.075 ;
        RECT 374.585 16.065 375.215 16.235 ;
        RECT 374.585 15.385 374.755 16.065 ;
      LAYER mcon ;
        RECT 387.925 1545.385 388.095 1545.555 ;
        RECT 387.925 1414.485 388.095 1414.655 ;
        RECT 387.925 1303.985 388.095 1304.155 ;
        RECT 387.925 572.305 388.095 572.475 ;
        RECT 387.465 330.905 387.635 331.075 ;
        RECT 375.045 16.065 375.215 16.235 ;
      LAYER met1 ;
        RECT 387.850 1579.540 388.170 1579.600 ;
        RECT 391.070 1579.540 391.390 1579.600 ;
        RECT 387.850 1579.400 391.390 1579.540 ;
        RECT 387.850 1579.340 388.170 1579.400 ;
        RECT 391.070 1579.340 391.390 1579.400 ;
        RECT 387.850 1545.540 388.170 1545.600 ;
        RECT 387.655 1545.400 388.170 1545.540 ;
        RECT 387.850 1545.340 388.170 1545.400 ;
        RECT 387.850 1497.600 388.170 1497.660 ;
        RECT 387.655 1497.460 388.170 1497.600 ;
        RECT 387.850 1497.400 388.170 1497.460 ;
        RECT 387.850 1414.640 388.170 1414.700 ;
        RECT 387.655 1414.500 388.170 1414.640 ;
        RECT 387.850 1414.440 388.170 1414.500 ;
        RECT 387.850 1352.760 388.170 1352.820 ;
        RECT 387.655 1352.620 388.170 1352.760 ;
        RECT 387.850 1352.560 388.170 1352.620 ;
        RECT 387.850 1304.140 388.170 1304.200 ;
        RECT 387.655 1304.000 388.170 1304.140 ;
        RECT 387.850 1303.940 388.170 1304.000 ;
        RECT 387.850 1256.200 388.170 1256.260 ;
        RECT 387.655 1256.060 388.170 1256.200 ;
        RECT 387.850 1256.000 388.170 1256.060 ;
        RECT 388.310 1173.240 388.630 1173.300 ;
        RECT 387.940 1173.100 388.630 1173.240 ;
        RECT 387.940 1172.960 388.080 1173.100 ;
        RECT 388.310 1173.040 388.630 1173.100 ;
        RECT 387.850 1172.700 388.170 1172.960 ;
        RECT 387.850 1062.740 388.170 1062.800 ;
        RECT 388.770 1062.740 389.090 1062.800 ;
        RECT 387.850 1062.600 389.090 1062.740 ;
        RECT 387.850 1062.540 388.170 1062.600 ;
        RECT 388.770 1062.540 389.090 1062.600 ;
        RECT 388.310 980.120 388.630 980.180 ;
        RECT 387.940 979.980 388.630 980.120 ;
        RECT 387.940 979.840 388.080 979.980 ;
        RECT 388.310 979.920 388.630 979.980 ;
        RECT 387.850 979.580 388.170 979.840 ;
        RECT 387.390 883.560 387.710 883.620 ;
        RECT 387.390 883.420 388.080 883.560 ;
        RECT 387.390 883.360 387.710 883.420 ;
        RECT 387.940 883.280 388.080 883.420 ;
        RECT 387.850 883.020 388.170 883.280 ;
        RECT 387.850 676.640 388.170 676.900 ;
        RECT 387.940 676.220 388.080 676.640 ;
        RECT 387.850 675.960 388.170 676.220 ;
        RECT 388.310 669.360 388.630 669.420 ;
        RECT 389.230 669.360 389.550 669.420 ;
        RECT 388.310 669.220 389.550 669.360 ;
        RECT 388.310 669.160 388.630 669.220 ;
        RECT 389.230 669.160 389.550 669.220 ;
        RECT 387.390 620.740 387.710 620.800 ;
        RECT 387.850 620.740 388.170 620.800 ;
        RECT 387.390 620.600 388.170 620.740 ;
        RECT 387.390 620.540 387.710 620.600 ;
        RECT 387.850 620.540 388.170 620.600 ;
        RECT 387.850 572.460 388.170 572.520 ;
        RECT 387.655 572.320 388.170 572.460 ;
        RECT 387.850 572.260 388.170 572.320 ;
        RECT 387.850 524.520 388.170 524.580 ;
        RECT 387.655 524.380 388.170 524.520 ;
        RECT 387.850 524.320 388.170 524.380 ;
        RECT 387.850 338.540 388.170 338.600 ;
        RECT 387.480 338.400 388.170 338.540 ;
        RECT 387.480 338.260 387.620 338.400 ;
        RECT 387.850 338.340 388.170 338.400 ;
        RECT 387.390 338.000 387.710 338.260 ;
        RECT 387.390 331.060 387.710 331.120 ;
        RECT 387.195 330.920 387.710 331.060 ;
        RECT 387.390 330.860 387.710 330.920 ;
        RECT 387.390 241.980 387.710 242.040 ;
        RECT 387.195 241.840 387.710 241.980 ;
        RECT 387.390 241.780 387.710 241.840 ;
        RECT 387.390 234.500 387.710 234.560 ;
        RECT 388.770 234.500 389.090 234.560 ;
        RECT 387.390 234.360 389.090 234.500 ;
        RECT 387.390 234.300 387.710 234.360 ;
        RECT 388.770 234.300 389.090 234.360 ;
        RECT 386.010 144.400 386.330 144.460 ;
        RECT 388.770 144.400 389.090 144.460 ;
        RECT 386.010 144.260 389.090 144.400 ;
        RECT 386.010 144.200 386.330 144.260 ;
        RECT 388.770 144.200 389.090 144.260 ;
        RECT 386.010 96.120 386.330 96.180 ;
        RECT 388.770 96.120 389.090 96.180 ;
        RECT 386.010 95.980 389.090 96.120 ;
        RECT 386.010 95.920 386.330 95.980 ;
        RECT 388.770 95.920 389.090 95.980 ;
        RECT 387.390 48.520 387.710 48.580 ;
        RECT 388.770 48.520 389.090 48.580 ;
        RECT 387.390 48.380 389.090 48.520 ;
        RECT 387.390 48.320 387.710 48.380 ;
        RECT 388.770 48.320 389.090 48.380 ;
        RECT 374.985 16.220 375.275 16.265 ;
        RECT 387.390 16.220 387.710 16.280 ;
        RECT 374.985 16.080 387.710 16.220 ;
        RECT 374.985 16.035 375.275 16.080 ;
        RECT 387.390 16.020 387.710 16.080 ;
        RECT 246.630 15.540 246.950 15.600 ;
        RECT 374.525 15.540 374.815 15.585 ;
        RECT 246.630 15.400 374.815 15.540 ;
        RECT 246.630 15.340 246.950 15.400 ;
        RECT 374.525 15.355 374.815 15.400 ;
      LAYER via ;
        RECT 387.880 1579.340 388.140 1579.600 ;
        RECT 391.100 1579.340 391.360 1579.600 ;
        RECT 387.880 1545.340 388.140 1545.600 ;
        RECT 387.880 1497.400 388.140 1497.660 ;
        RECT 387.880 1414.440 388.140 1414.700 ;
        RECT 387.880 1352.560 388.140 1352.820 ;
        RECT 387.880 1303.940 388.140 1304.200 ;
        RECT 387.880 1256.000 388.140 1256.260 ;
        RECT 388.340 1173.040 388.600 1173.300 ;
        RECT 387.880 1172.700 388.140 1172.960 ;
        RECT 387.880 1062.540 388.140 1062.800 ;
        RECT 388.800 1062.540 389.060 1062.800 ;
        RECT 388.340 979.920 388.600 980.180 ;
        RECT 387.880 979.580 388.140 979.840 ;
        RECT 387.420 883.360 387.680 883.620 ;
        RECT 387.880 883.020 388.140 883.280 ;
        RECT 387.880 676.640 388.140 676.900 ;
        RECT 387.880 675.960 388.140 676.220 ;
        RECT 388.340 669.160 388.600 669.420 ;
        RECT 389.260 669.160 389.520 669.420 ;
        RECT 387.420 620.540 387.680 620.800 ;
        RECT 387.880 620.540 388.140 620.800 ;
        RECT 387.880 572.260 388.140 572.520 ;
        RECT 387.880 524.320 388.140 524.580 ;
        RECT 387.880 338.340 388.140 338.600 ;
        RECT 387.420 338.000 387.680 338.260 ;
        RECT 387.420 330.860 387.680 331.120 ;
        RECT 387.420 241.780 387.680 242.040 ;
        RECT 387.420 234.300 387.680 234.560 ;
        RECT 388.800 234.300 389.060 234.560 ;
        RECT 386.040 144.200 386.300 144.460 ;
        RECT 388.800 144.200 389.060 144.460 ;
        RECT 386.040 95.920 386.300 96.180 ;
        RECT 388.800 95.920 389.060 96.180 ;
        RECT 387.420 48.320 387.680 48.580 ;
        RECT 388.800 48.320 389.060 48.580 ;
        RECT 387.420 16.020 387.680 16.280 ;
        RECT 246.660 15.340 246.920 15.600 ;
      LAYER met2 ;
        RECT 392.940 1600.450 393.220 1604.000 ;
        RECT 391.160 1600.310 393.220 1600.450 ;
        RECT 391.160 1579.630 391.300 1600.310 ;
        RECT 392.940 1600.000 393.220 1600.310 ;
        RECT 387.880 1579.310 388.140 1579.630 ;
        RECT 391.100 1579.310 391.360 1579.630 ;
        RECT 387.940 1545.630 388.080 1579.310 ;
        RECT 387.880 1545.310 388.140 1545.630 ;
        RECT 387.880 1497.370 388.140 1497.690 ;
        RECT 387.940 1414.730 388.080 1497.370 ;
        RECT 387.880 1414.410 388.140 1414.730 ;
        RECT 387.880 1352.530 388.140 1352.850 ;
        RECT 387.940 1304.230 388.080 1352.530 ;
        RECT 387.880 1303.910 388.140 1304.230 ;
        RECT 387.880 1255.970 388.140 1256.290 ;
        RECT 387.940 1207.410 388.080 1255.970 ;
        RECT 387.940 1207.270 388.540 1207.410 ;
        RECT 388.400 1173.330 388.540 1207.270 ;
        RECT 388.340 1173.010 388.600 1173.330 ;
        RECT 387.880 1172.670 388.140 1172.990 ;
        RECT 387.940 1110.965 388.080 1172.670 ;
        RECT 387.870 1110.595 388.150 1110.965 ;
        RECT 388.790 1110.595 389.070 1110.965 ;
        RECT 388.860 1062.830 389.000 1110.595 ;
        RECT 387.880 1062.510 388.140 1062.830 ;
        RECT 388.800 1062.510 389.060 1062.830 ;
        RECT 387.940 1014.290 388.080 1062.510 ;
        RECT 387.940 1014.150 388.540 1014.290 ;
        RECT 388.400 980.210 388.540 1014.150 ;
        RECT 388.340 979.890 388.600 980.210 ;
        RECT 387.880 979.550 388.140 979.870 ;
        RECT 387.940 917.730 388.080 979.550 ;
        RECT 387.480 917.590 388.080 917.730 ;
        RECT 387.480 883.650 387.620 917.590 ;
        RECT 387.420 883.330 387.680 883.650 ;
        RECT 387.880 882.990 388.140 883.310 ;
        RECT 387.940 787.170 388.080 882.990 ;
        RECT 387.480 787.030 388.080 787.170 ;
        RECT 387.480 786.490 387.620 787.030 ;
        RECT 387.480 786.350 388.080 786.490 ;
        RECT 387.940 676.930 388.080 786.350 ;
        RECT 387.880 676.610 388.140 676.930 ;
        RECT 387.880 675.930 388.140 676.250 ;
        RECT 387.940 669.530 388.080 675.930 ;
        RECT 387.940 669.450 388.540 669.530 ;
        RECT 387.940 669.390 388.600 669.450 ;
        RECT 388.340 669.130 388.600 669.390 ;
        RECT 389.260 669.130 389.520 669.450 ;
        RECT 388.400 668.975 388.540 669.130 ;
        RECT 389.320 621.365 389.460 669.130 ;
        RECT 387.410 620.995 387.690 621.365 ;
        RECT 389.250 620.995 389.530 621.365 ;
        RECT 387.480 620.830 387.620 620.995 ;
        RECT 387.420 620.510 387.680 620.830 ;
        RECT 387.880 620.510 388.140 620.830 ;
        RECT 387.940 572.550 388.080 620.510 ;
        RECT 387.880 572.230 388.140 572.550 ;
        RECT 387.880 524.290 388.140 524.610 ;
        RECT 387.940 497.490 388.080 524.290 ;
        RECT 387.940 497.350 388.540 497.490 ;
        RECT 388.400 496.130 388.540 497.350 ;
        RECT 387.940 495.990 388.540 496.130 ;
        RECT 387.940 338.630 388.080 495.990 ;
        RECT 387.880 338.310 388.140 338.630 ;
        RECT 387.420 337.970 387.680 338.290 ;
        RECT 387.480 331.150 387.620 337.970 ;
        RECT 387.420 330.830 387.680 331.150 ;
        RECT 387.420 241.750 387.680 242.070 ;
        RECT 387.480 234.590 387.620 241.750 ;
        RECT 387.420 234.270 387.680 234.590 ;
        RECT 388.800 234.270 389.060 234.590 ;
        RECT 388.860 144.490 389.000 234.270 ;
        RECT 386.040 144.170 386.300 144.490 ;
        RECT 388.800 144.170 389.060 144.490 ;
        RECT 386.100 96.210 386.240 144.170 ;
        RECT 386.040 95.890 386.300 96.210 ;
        RECT 388.800 95.890 389.060 96.210 ;
        RECT 388.860 48.610 389.000 95.890 ;
        RECT 387.420 48.290 387.680 48.610 ;
        RECT 388.800 48.290 389.060 48.610 ;
        RECT 387.480 16.310 387.620 48.290 ;
        RECT 387.420 15.990 387.680 16.310 ;
        RECT 246.660 15.310 246.920 15.630 ;
        RECT 246.720 2.400 246.860 15.310 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 387.870 1110.640 388.150 1110.920 ;
        RECT 388.790 1110.640 389.070 1110.920 ;
        RECT 387.410 621.040 387.690 621.320 ;
        RECT 389.250 621.040 389.530 621.320 ;
      LAYER met3 ;
        RECT 387.845 1110.930 388.175 1110.945 ;
        RECT 388.765 1110.930 389.095 1110.945 ;
        RECT 387.845 1110.630 389.095 1110.930 ;
        RECT 387.845 1110.615 388.175 1110.630 ;
        RECT 388.765 1110.615 389.095 1110.630 ;
        RECT 387.385 621.330 387.715 621.345 ;
        RECT 389.225 621.330 389.555 621.345 ;
        RECT 387.385 621.030 389.555 621.330 ;
        RECT 387.385 621.015 387.715 621.030 ;
        RECT 389.225 621.015 389.555 621.030 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 268.710 1587.700 269.030 1587.760 ;
        RECT 399.350 1587.700 399.670 1587.760 ;
        RECT 268.710 1587.560 399.670 1587.700 ;
        RECT 268.710 1587.500 269.030 1587.560 ;
        RECT 399.350 1587.500 399.670 1587.560 ;
        RECT 264.110 16.560 264.430 16.620 ;
        RECT 268.710 16.560 269.030 16.620 ;
        RECT 264.110 16.420 269.030 16.560 ;
        RECT 264.110 16.360 264.430 16.420 ;
        RECT 268.710 16.360 269.030 16.420 ;
      LAYER via ;
        RECT 268.740 1587.500 269.000 1587.760 ;
        RECT 399.380 1587.500 399.640 1587.760 ;
        RECT 264.140 16.360 264.400 16.620 ;
        RECT 268.740 16.360 269.000 16.620 ;
      LAYER met2 ;
        RECT 399.380 1600.000 399.660 1604.000 ;
        RECT 399.440 1587.790 399.580 1600.000 ;
        RECT 268.740 1587.470 269.000 1587.790 ;
        RECT 399.380 1587.470 399.640 1587.790 ;
        RECT 268.800 16.650 268.940 1587.470 ;
        RECT 264.140 16.330 264.400 16.650 ;
        RECT 268.740 16.330 269.000 16.650 ;
        RECT 264.200 2.400 264.340 16.330 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 400.730 1579.880 401.050 1579.940 ;
        RECT 404.870 1579.880 405.190 1579.940 ;
        RECT 400.730 1579.740 405.190 1579.880 ;
        RECT 400.730 1579.680 401.050 1579.740 ;
        RECT 404.870 1579.680 405.190 1579.740 ;
        RECT 282.050 14.520 282.370 14.580 ;
        RECT 400.730 14.520 401.050 14.580 ;
        RECT 282.050 14.380 401.050 14.520 ;
        RECT 282.050 14.320 282.370 14.380 ;
        RECT 400.730 14.320 401.050 14.380 ;
      LAYER via ;
        RECT 400.760 1579.680 401.020 1579.940 ;
        RECT 404.900 1579.680 405.160 1579.940 ;
        RECT 282.080 14.320 282.340 14.580 ;
        RECT 400.760 14.320 401.020 14.580 ;
      LAYER met2 ;
        RECT 406.280 1600.450 406.560 1604.000 ;
        RECT 404.960 1600.310 406.560 1600.450 ;
        RECT 404.960 1579.970 405.100 1600.310 ;
        RECT 406.280 1600.000 406.560 1600.310 ;
        RECT 400.760 1579.650 401.020 1579.970 ;
        RECT 404.900 1579.650 405.160 1579.970 ;
        RECT 400.820 14.610 400.960 1579.650 ;
        RECT 282.080 14.290 282.340 14.610 ;
        RECT 400.760 14.290 401.020 14.610 ;
        RECT 282.140 2.400 282.280 14.290 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 407.630 1579.880 407.950 1579.940 ;
        RECT 411.310 1579.880 411.630 1579.940 ;
        RECT 407.630 1579.740 411.630 1579.880 ;
        RECT 407.630 1579.680 407.950 1579.740 ;
        RECT 411.310 1579.680 411.630 1579.740 ;
        RECT 299.990 17.580 300.310 17.640 ;
        RECT 299.990 17.440 376.120 17.580 ;
        RECT 299.990 17.380 300.310 17.440 ;
        RECT 375.980 17.240 376.120 17.440 ;
        RECT 407.630 17.240 407.950 17.300 ;
        RECT 375.980 17.100 407.950 17.240 ;
        RECT 407.630 17.040 407.950 17.100 ;
      LAYER via ;
        RECT 407.660 1579.680 407.920 1579.940 ;
        RECT 411.340 1579.680 411.600 1579.940 ;
        RECT 300.020 17.380 300.280 17.640 ;
        RECT 407.660 17.040 407.920 17.300 ;
      LAYER met2 ;
        RECT 412.720 1600.450 413.000 1604.000 ;
        RECT 411.400 1600.310 413.000 1600.450 ;
        RECT 411.400 1579.970 411.540 1600.310 ;
        RECT 412.720 1600.000 413.000 1600.310 ;
        RECT 407.660 1579.650 407.920 1579.970 ;
        RECT 411.340 1579.650 411.600 1579.970 ;
        RECT 300.020 17.350 300.280 17.670 ;
        RECT 300.080 2.400 300.220 17.350 ;
        RECT 407.720 17.330 407.860 1579.650 ;
        RECT 407.660 17.010 407.920 17.330 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 323.525 18.445 325.995 18.615 ;
        RECT 375.505 18.445 375.675 20.315 ;
        RECT 323.525 17.765 323.695 18.445 ;
      LAYER mcon ;
        RECT 375.505 20.145 375.675 20.315 ;
        RECT 325.825 18.445 325.995 18.615 ;
      LAYER met1 ;
        RECT 414.530 1578.520 414.850 1578.580 ;
        RECT 417.750 1578.520 418.070 1578.580 ;
        RECT 414.530 1578.380 418.070 1578.520 ;
        RECT 414.530 1578.320 414.850 1578.380 ;
        RECT 417.750 1578.320 418.070 1578.380 ;
        RECT 376.440 20.500 400.960 20.640 ;
        RECT 375.445 20.300 375.735 20.345 ;
        RECT 376.440 20.300 376.580 20.500 ;
        RECT 375.445 20.160 376.580 20.300 ;
        RECT 400.820 20.300 400.960 20.500 ;
        RECT 414.530 20.300 414.850 20.360 ;
        RECT 400.820 20.160 414.850 20.300 ;
        RECT 375.445 20.115 375.735 20.160 ;
        RECT 414.530 20.100 414.850 20.160 ;
        RECT 325.765 18.600 326.055 18.645 ;
        RECT 375.445 18.600 375.735 18.645 ;
        RECT 325.765 18.460 375.735 18.600 ;
        RECT 325.765 18.415 326.055 18.460 ;
        RECT 375.445 18.415 375.735 18.460 ;
        RECT 317.930 17.920 318.250 17.980 ;
        RECT 323.465 17.920 323.755 17.965 ;
        RECT 317.930 17.780 323.755 17.920 ;
        RECT 317.930 17.720 318.250 17.780 ;
        RECT 323.465 17.735 323.755 17.780 ;
      LAYER via ;
        RECT 414.560 1578.320 414.820 1578.580 ;
        RECT 417.780 1578.320 418.040 1578.580 ;
        RECT 414.560 20.100 414.820 20.360 ;
        RECT 317.960 17.720 318.220 17.980 ;
      LAYER met2 ;
        RECT 419.620 1600.450 419.900 1604.000 ;
        RECT 417.840 1600.310 419.900 1600.450 ;
        RECT 417.840 1578.610 417.980 1600.310 ;
        RECT 419.620 1600.000 419.900 1600.310 ;
        RECT 414.560 1578.290 414.820 1578.610 ;
        RECT 417.780 1578.290 418.040 1578.610 ;
        RECT 414.620 20.390 414.760 1578.290 ;
        RECT 414.560 20.070 414.820 20.390 ;
        RECT 317.960 17.690 318.220 18.010 ;
        RECT 318.020 2.400 318.160 17.690 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 370.905 19.465 371.995 19.635 ;
        RECT 371.825 19.125 371.995 19.465 ;
      LAYER met1 ;
        RECT 389.690 1588.040 390.010 1588.100 ;
        RECT 426.490 1588.040 426.810 1588.100 ;
        RECT 389.690 1587.900 426.810 1588.040 ;
        RECT 389.690 1587.840 390.010 1587.900 ;
        RECT 426.490 1587.840 426.810 1587.900 ;
        RECT 335.870 19.620 336.190 19.680 ;
        RECT 370.845 19.620 371.135 19.665 ;
        RECT 335.870 19.480 371.135 19.620 ;
        RECT 335.870 19.420 336.190 19.480 ;
        RECT 370.845 19.435 371.135 19.480 ;
        RECT 371.765 19.280 372.055 19.325 ;
        RECT 389.690 19.280 390.010 19.340 ;
        RECT 371.765 19.140 390.010 19.280 ;
        RECT 371.765 19.095 372.055 19.140 ;
        RECT 389.690 19.080 390.010 19.140 ;
      LAYER via ;
        RECT 389.720 1587.840 389.980 1588.100 ;
        RECT 426.520 1587.840 426.780 1588.100 ;
        RECT 335.900 19.420 336.160 19.680 ;
        RECT 389.720 19.080 389.980 19.340 ;
      LAYER met2 ;
        RECT 426.520 1600.000 426.800 1604.000 ;
        RECT 426.580 1588.130 426.720 1600.000 ;
        RECT 389.720 1587.810 389.980 1588.130 ;
        RECT 426.520 1587.810 426.780 1588.130 ;
        RECT 335.900 19.390 336.160 19.710 ;
        RECT 335.960 2.400 336.100 19.390 ;
        RECT 389.780 19.370 389.920 1587.810 ;
        RECT 389.720 19.050 389.980 19.370 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 397.125 16.745 397.295 19.975 ;
      LAYER mcon ;
        RECT 397.125 19.805 397.295 19.975 ;
      LAYER met1 ;
        RECT 427.870 1579.880 428.190 1579.940 ;
        RECT 431.550 1579.880 431.870 1579.940 ;
        RECT 427.870 1579.740 431.870 1579.880 ;
        RECT 427.870 1579.680 428.190 1579.740 ;
        RECT 431.550 1579.680 431.870 1579.740 ;
        RECT 397.065 19.960 397.355 20.005 ;
        RECT 427.870 19.960 428.190 20.020 ;
        RECT 397.065 19.820 428.190 19.960 ;
        RECT 397.065 19.775 397.355 19.820 ;
        RECT 427.870 19.760 428.190 19.820 ;
        RECT 353.350 16.900 353.670 16.960 ;
        RECT 397.065 16.900 397.355 16.945 ;
        RECT 353.350 16.760 397.355 16.900 ;
        RECT 353.350 16.700 353.670 16.760 ;
        RECT 397.065 16.715 397.355 16.760 ;
      LAYER via ;
        RECT 427.900 1579.680 428.160 1579.940 ;
        RECT 431.580 1579.680 431.840 1579.940 ;
        RECT 427.900 19.760 428.160 20.020 ;
        RECT 353.380 16.700 353.640 16.960 ;
      LAYER met2 ;
        RECT 432.960 1600.450 433.240 1604.000 ;
        RECT 431.640 1600.310 433.240 1600.450 ;
        RECT 431.640 1579.970 431.780 1600.310 ;
        RECT 432.960 1600.000 433.240 1600.310 ;
        RECT 427.900 1579.650 428.160 1579.970 ;
        RECT 431.580 1579.650 431.840 1579.970 ;
        RECT 427.960 20.050 428.100 1579.650 ;
        RECT 427.900 19.730 428.160 20.050 ;
        RECT 353.380 16.670 353.640 16.990 ;
        RECT 353.440 2.400 353.580 16.670 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 372.285 1497.445 372.455 1545.555 ;
        RECT 372.285 1400.885 372.455 1490.475 ;
        RECT 372.285 766.105 372.455 814.215 ;
        RECT 372.285 669.545 372.455 717.655 ;
        RECT 372.285 476.085 372.455 524.195 ;
        RECT 372.285 282.965 372.455 331.075 ;
        RECT 372.285 186.405 372.455 234.515 ;
        RECT 371.365 48.365 371.535 137.955 ;
      LAYER mcon ;
        RECT 372.285 1545.385 372.455 1545.555 ;
        RECT 372.285 1490.305 372.455 1490.475 ;
        RECT 372.285 814.045 372.455 814.215 ;
        RECT 372.285 717.485 372.455 717.655 ;
        RECT 372.285 524.025 372.455 524.195 ;
        RECT 372.285 330.905 372.455 331.075 ;
        RECT 372.285 234.345 372.455 234.515 ;
        RECT 371.365 137.785 371.535 137.955 ;
      LAYER met1 ;
        RECT 439.830 1590.760 440.150 1590.820 ;
        RECT 420.140 1590.620 440.150 1590.760 ;
        RECT 372.210 1590.420 372.530 1590.480 ;
        RECT 420.140 1590.420 420.280 1590.620 ;
        RECT 439.830 1590.560 440.150 1590.620 ;
        RECT 372.210 1590.280 420.280 1590.420 ;
        RECT 372.210 1590.220 372.530 1590.280 ;
        RECT 372.210 1545.540 372.530 1545.600 ;
        RECT 372.015 1545.400 372.530 1545.540 ;
        RECT 372.210 1545.340 372.530 1545.400 ;
        RECT 372.210 1497.600 372.530 1497.660 ;
        RECT 372.015 1497.460 372.530 1497.600 ;
        RECT 372.210 1497.400 372.530 1497.460 ;
        RECT 372.210 1490.460 372.530 1490.520 ;
        RECT 372.015 1490.320 372.530 1490.460 ;
        RECT 372.210 1490.260 372.530 1490.320 ;
        RECT 372.210 1401.040 372.530 1401.100 ;
        RECT 372.015 1400.900 372.530 1401.040 ;
        RECT 372.210 1400.840 372.530 1400.900 ;
        RECT 371.290 1345.620 371.610 1345.680 ;
        RECT 372.210 1345.620 372.530 1345.680 ;
        RECT 371.290 1345.480 372.530 1345.620 ;
        RECT 371.290 1345.420 371.610 1345.480 ;
        RECT 372.210 1345.420 372.530 1345.480 ;
        RECT 371.290 1249.060 371.610 1249.120 ;
        RECT 372.210 1249.060 372.530 1249.120 ;
        RECT 371.290 1248.920 372.530 1249.060 ;
        RECT 371.290 1248.860 371.610 1248.920 ;
        RECT 372.210 1248.860 372.530 1248.920 ;
        RECT 371.290 1152.500 371.610 1152.560 ;
        RECT 372.210 1152.500 372.530 1152.560 ;
        RECT 371.290 1152.360 372.530 1152.500 ;
        RECT 371.290 1152.300 371.610 1152.360 ;
        RECT 372.210 1152.300 372.530 1152.360 ;
        RECT 371.290 1007.320 371.610 1007.380 ;
        RECT 372.210 1007.320 372.530 1007.380 ;
        RECT 371.290 1007.180 372.530 1007.320 ;
        RECT 371.290 1007.120 371.610 1007.180 ;
        RECT 372.210 1007.120 372.530 1007.180 ;
        RECT 371.290 910.760 371.610 910.820 ;
        RECT 372.210 910.760 372.530 910.820 ;
        RECT 371.290 910.620 372.530 910.760 ;
        RECT 371.290 910.560 371.610 910.620 ;
        RECT 372.210 910.560 372.530 910.620 ;
        RECT 372.210 814.200 372.530 814.260 ;
        RECT 372.015 814.060 372.530 814.200 ;
        RECT 372.210 814.000 372.530 814.060 ;
        RECT 372.210 766.260 372.530 766.320 ;
        RECT 372.015 766.120 372.530 766.260 ;
        RECT 372.210 766.060 372.530 766.120 ;
        RECT 372.210 717.640 372.530 717.700 ;
        RECT 372.015 717.500 372.530 717.640 ;
        RECT 372.210 717.440 372.530 717.500 ;
        RECT 372.210 669.700 372.530 669.760 ;
        RECT 372.015 669.560 372.530 669.700 ;
        RECT 372.210 669.500 372.530 669.560 ;
        RECT 372.210 524.180 372.530 524.240 ;
        RECT 372.015 524.040 372.530 524.180 ;
        RECT 372.210 523.980 372.530 524.040 ;
        RECT 372.210 476.240 372.530 476.300 ;
        RECT 372.015 476.100 372.530 476.240 ;
        RECT 372.210 476.040 372.530 476.100 ;
        RECT 372.210 331.060 372.530 331.120 ;
        RECT 372.015 330.920 372.530 331.060 ;
        RECT 372.210 330.860 372.530 330.920 ;
        RECT 372.210 283.120 372.530 283.180 ;
        RECT 372.015 282.980 372.530 283.120 ;
        RECT 372.210 282.920 372.530 282.980 ;
        RECT 372.210 234.500 372.530 234.560 ;
        RECT 372.015 234.360 372.530 234.500 ;
        RECT 372.210 234.300 372.530 234.360 ;
        RECT 372.210 186.560 372.530 186.620 ;
        RECT 372.015 186.420 372.530 186.560 ;
        RECT 372.210 186.360 372.530 186.420 ;
        RECT 371.305 137.940 371.595 137.985 ;
        RECT 372.210 137.940 372.530 138.000 ;
        RECT 371.305 137.800 372.530 137.940 ;
        RECT 371.305 137.755 371.595 137.800 ;
        RECT 372.210 137.740 372.530 137.800 ;
        RECT 371.290 48.520 371.610 48.580 ;
        RECT 371.095 48.380 371.610 48.520 ;
        RECT 371.290 48.320 371.610 48.380 ;
      LAYER via ;
        RECT 372.240 1590.220 372.500 1590.480 ;
        RECT 439.860 1590.560 440.120 1590.820 ;
        RECT 372.240 1545.340 372.500 1545.600 ;
        RECT 372.240 1497.400 372.500 1497.660 ;
        RECT 372.240 1490.260 372.500 1490.520 ;
        RECT 372.240 1400.840 372.500 1401.100 ;
        RECT 371.320 1345.420 371.580 1345.680 ;
        RECT 372.240 1345.420 372.500 1345.680 ;
        RECT 371.320 1248.860 371.580 1249.120 ;
        RECT 372.240 1248.860 372.500 1249.120 ;
        RECT 371.320 1152.300 371.580 1152.560 ;
        RECT 372.240 1152.300 372.500 1152.560 ;
        RECT 371.320 1007.120 371.580 1007.380 ;
        RECT 372.240 1007.120 372.500 1007.380 ;
        RECT 371.320 910.560 371.580 910.820 ;
        RECT 372.240 910.560 372.500 910.820 ;
        RECT 372.240 814.000 372.500 814.260 ;
        RECT 372.240 766.060 372.500 766.320 ;
        RECT 372.240 717.440 372.500 717.700 ;
        RECT 372.240 669.500 372.500 669.760 ;
        RECT 372.240 523.980 372.500 524.240 ;
        RECT 372.240 476.040 372.500 476.300 ;
        RECT 372.240 330.860 372.500 331.120 ;
        RECT 372.240 282.920 372.500 283.180 ;
        RECT 372.240 234.300 372.500 234.560 ;
        RECT 372.240 186.360 372.500 186.620 ;
        RECT 372.240 137.740 372.500 138.000 ;
        RECT 371.320 48.320 371.580 48.580 ;
      LAYER met2 ;
        RECT 439.860 1600.000 440.140 1604.000 ;
        RECT 439.920 1590.850 440.060 1600.000 ;
        RECT 439.860 1590.530 440.120 1590.850 ;
        RECT 372.240 1590.190 372.500 1590.510 ;
        RECT 372.300 1545.630 372.440 1590.190 ;
        RECT 372.240 1545.310 372.500 1545.630 ;
        RECT 372.240 1497.370 372.500 1497.690 ;
        RECT 372.300 1490.550 372.440 1497.370 ;
        RECT 372.240 1490.230 372.500 1490.550 ;
        RECT 372.240 1400.810 372.500 1401.130 ;
        RECT 372.300 1393.845 372.440 1400.810 ;
        RECT 371.310 1393.475 371.590 1393.845 ;
        RECT 372.230 1393.475 372.510 1393.845 ;
        RECT 371.380 1345.710 371.520 1393.475 ;
        RECT 371.320 1345.390 371.580 1345.710 ;
        RECT 372.240 1345.390 372.500 1345.710 ;
        RECT 372.300 1297.285 372.440 1345.390 ;
        RECT 371.310 1296.915 371.590 1297.285 ;
        RECT 372.230 1296.915 372.510 1297.285 ;
        RECT 371.380 1249.150 371.520 1296.915 ;
        RECT 371.320 1248.830 371.580 1249.150 ;
        RECT 372.240 1248.830 372.500 1249.150 ;
        RECT 372.300 1200.725 372.440 1248.830 ;
        RECT 371.310 1200.355 371.590 1200.725 ;
        RECT 372.230 1200.355 372.510 1200.725 ;
        RECT 371.380 1152.590 371.520 1200.355 ;
        RECT 371.320 1152.270 371.580 1152.590 ;
        RECT 372.240 1152.270 372.500 1152.590 ;
        RECT 372.300 1104.165 372.440 1152.270 ;
        RECT 371.310 1103.795 371.590 1104.165 ;
        RECT 372.230 1103.795 372.510 1104.165 ;
        RECT 371.380 1055.885 371.520 1103.795 ;
        RECT 371.310 1055.515 371.590 1055.885 ;
        RECT 372.230 1055.515 372.510 1055.885 ;
        RECT 372.300 1007.410 372.440 1055.515 ;
        RECT 371.320 1007.090 371.580 1007.410 ;
        RECT 372.240 1007.090 372.500 1007.410 ;
        RECT 371.380 959.325 371.520 1007.090 ;
        RECT 371.310 958.955 371.590 959.325 ;
        RECT 372.230 958.955 372.510 959.325 ;
        RECT 372.300 910.850 372.440 958.955 ;
        RECT 371.320 910.530 371.580 910.850 ;
        RECT 372.240 910.530 372.500 910.850 ;
        RECT 371.380 862.765 371.520 910.530 ;
        RECT 371.310 862.395 371.590 862.765 ;
        RECT 372.230 862.395 372.510 862.765 ;
        RECT 372.300 814.290 372.440 862.395 ;
        RECT 372.240 813.970 372.500 814.290 ;
        RECT 372.240 766.030 372.500 766.350 ;
        RECT 372.300 725.405 372.440 766.030 ;
        RECT 372.230 725.035 372.510 725.405 ;
        RECT 372.230 724.355 372.510 724.725 ;
        RECT 372.300 717.730 372.440 724.355 ;
        RECT 372.240 717.410 372.500 717.730 ;
        RECT 372.240 669.470 372.500 669.790 ;
        RECT 372.300 628.845 372.440 669.470 ;
        RECT 372.230 628.475 372.510 628.845 ;
        RECT 372.230 627.795 372.510 628.165 ;
        RECT 372.300 524.270 372.440 627.795 ;
        RECT 372.240 523.950 372.500 524.270 ;
        RECT 372.240 476.010 372.500 476.330 ;
        RECT 372.300 331.150 372.440 476.010 ;
        RECT 372.240 330.830 372.500 331.150 ;
        RECT 372.240 282.890 372.500 283.210 ;
        RECT 372.300 234.590 372.440 282.890 ;
        RECT 372.240 234.270 372.500 234.590 ;
        RECT 372.240 186.330 372.500 186.650 ;
        RECT 372.300 138.030 372.440 186.330 ;
        RECT 372.240 137.710 372.500 138.030 ;
        RECT 371.320 48.290 371.580 48.610 ;
        RECT 371.380 2.400 371.520 48.290 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 371.310 1393.520 371.590 1393.800 ;
        RECT 372.230 1393.520 372.510 1393.800 ;
        RECT 371.310 1296.960 371.590 1297.240 ;
        RECT 372.230 1296.960 372.510 1297.240 ;
        RECT 371.310 1200.400 371.590 1200.680 ;
        RECT 372.230 1200.400 372.510 1200.680 ;
        RECT 371.310 1103.840 371.590 1104.120 ;
        RECT 372.230 1103.840 372.510 1104.120 ;
        RECT 371.310 1055.560 371.590 1055.840 ;
        RECT 372.230 1055.560 372.510 1055.840 ;
        RECT 371.310 959.000 371.590 959.280 ;
        RECT 372.230 959.000 372.510 959.280 ;
        RECT 371.310 862.440 371.590 862.720 ;
        RECT 372.230 862.440 372.510 862.720 ;
        RECT 372.230 725.080 372.510 725.360 ;
        RECT 372.230 724.400 372.510 724.680 ;
        RECT 372.230 628.520 372.510 628.800 ;
        RECT 372.230 627.840 372.510 628.120 ;
      LAYER met3 ;
        RECT 371.285 1393.810 371.615 1393.825 ;
        RECT 372.205 1393.810 372.535 1393.825 ;
        RECT 371.285 1393.510 372.535 1393.810 ;
        RECT 371.285 1393.495 371.615 1393.510 ;
        RECT 372.205 1393.495 372.535 1393.510 ;
        RECT 371.285 1297.250 371.615 1297.265 ;
        RECT 372.205 1297.250 372.535 1297.265 ;
        RECT 371.285 1296.950 372.535 1297.250 ;
        RECT 371.285 1296.935 371.615 1296.950 ;
        RECT 372.205 1296.935 372.535 1296.950 ;
        RECT 371.285 1200.690 371.615 1200.705 ;
        RECT 372.205 1200.690 372.535 1200.705 ;
        RECT 371.285 1200.390 372.535 1200.690 ;
        RECT 371.285 1200.375 371.615 1200.390 ;
        RECT 372.205 1200.375 372.535 1200.390 ;
        RECT 371.285 1104.130 371.615 1104.145 ;
        RECT 372.205 1104.130 372.535 1104.145 ;
        RECT 371.285 1103.830 372.535 1104.130 ;
        RECT 371.285 1103.815 371.615 1103.830 ;
        RECT 372.205 1103.815 372.535 1103.830 ;
        RECT 371.285 1055.850 371.615 1055.865 ;
        RECT 372.205 1055.850 372.535 1055.865 ;
        RECT 371.285 1055.550 372.535 1055.850 ;
        RECT 371.285 1055.535 371.615 1055.550 ;
        RECT 372.205 1055.535 372.535 1055.550 ;
        RECT 371.285 959.290 371.615 959.305 ;
        RECT 372.205 959.290 372.535 959.305 ;
        RECT 371.285 958.990 372.535 959.290 ;
        RECT 371.285 958.975 371.615 958.990 ;
        RECT 372.205 958.975 372.535 958.990 ;
        RECT 371.285 862.730 371.615 862.745 ;
        RECT 372.205 862.730 372.535 862.745 ;
        RECT 371.285 862.430 372.535 862.730 ;
        RECT 371.285 862.415 371.615 862.430 ;
        RECT 372.205 862.415 372.535 862.430 ;
        RECT 372.205 725.370 372.535 725.385 ;
        RECT 372.205 725.070 373.210 725.370 ;
        RECT 372.205 725.055 372.535 725.070 ;
        RECT 372.205 724.690 372.535 724.705 ;
        RECT 372.910 724.690 373.210 725.070 ;
        RECT 372.205 724.390 373.210 724.690 ;
        RECT 372.205 724.375 372.535 724.390 ;
        RECT 372.205 628.810 372.535 628.825 ;
        RECT 372.205 628.510 373.210 628.810 ;
        RECT 372.205 628.495 372.535 628.510 ;
        RECT 372.205 628.130 372.535 628.145 ;
        RECT 372.910 628.130 373.210 628.510 ;
        RECT 372.205 627.830 373.210 628.130 ;
        RECT 372.205 627.815 372.535 627.830 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 389.230 16.220 389.550 16.280 ;
        RECT 442.130 16.220 442.450 16.280 ;
        RECT 389.230 16.080 442.450 16.220 ;
        RECT 389.230 16.020 389.550 16.080 ;
        RECT 442.130 16.020 442.450 16.080 ;
      LAYER via ;
        RECT 389.260 16.020 389.520 16.280 ;
        RECT 442.160 16.020 442.420 16.280 ;
      LAYER met2 ;
        RECT 446.760 1601.130 447.040 1604.000 ;
        RECT 444.980 1600.990 447.040 1601.130 ;
        RECT 444.980 1580.050 445.120 1600.990 ;
        RECT 446.760 1600.000 447.040 1600.990 ;
        RECT 442.220 1579.910 445.120 1580.050 ;
        RECT 442.220 16.310 442.360 1579.910 ;
        RECT 389.260 15.990 389.520 16.310 ;
        RECT 442.160 15.990 442.420 16.310 ;
        RECT 389.320 2.400 389.460 15.990 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 413.610 1591.780 413.930 1591.840 ;
        RECT 453.170 1591.780 453.490 1591.840 ;
        RECT 413.610 1591.640 453.490 1591.780 ;
        RECT 413.610 1591.580 413.930 1591.640 ;
        RECT 453.170 1591.580 453.490 1591.640 ;
        RECT 407.170 18.600 407.490 18.660 ;
        RECT 413.610 18.600 413.930 18.660 ;
        RECT 407.170 18.460 413.930 18.600 ;
        RECT 407.170 18.400 407.490 18.460 ;
        RECT 413.610 18.400 413.930 18.460 ;
      LAYER via ;
        RECT 413.640 1591.580 413.900 1591.840 ;
        RECT 453.200 1591.580 453.460 1591.840 ;
        RECT 407.200 18.400 407.460 18.660 ;
        RECT 413.640 18.400 413.900 18.660 ;
      LAYER met2 ;
        RECT 453.200 1600.000 453.480 1604.000 ;
        RECT 453.260 1591.870 453.400 1600.000 ;
        RECT 413.640 1591.550 413.900 1591.870 ;
        RECT 453.200 1591.550 453.460 1591.870 ;
        RECT 413.700 18.690 413.840 1591.550 ;
        RECT 407.200 18.370 407.460 18.690 ;
        RECT 413.640 18.370 413.900 18.690 ;
        RECT 407.260 2.400 407.400 18.370 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.320 1600.000 325.600 1604.000 ;
        RECT 325.380 1591.725 325.520 1600.000 ;
        RECT 68.170 1591.355 68.450 1591.725 ;
        RECT 325.310 1591.355 325.590 1591.725 ;
        RECT 68.240 2.400 68.380 1591.355 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 68.170 1591.400 68.450 1591.680 ;
        RECT 325.310 1591.400 325.590 1591.680 ;
      LAYER met3 ;
        RECT 68.145 1591.690 68.475 1591.705 ;
        RECT 325.285 1591.690 325.615 1591.705 ;
        RECT 68.145 1591.390 325.615 1591.690 ;
        RECT 68.145 1591.375 68.475 1591.390 ;
        RECT 325.285 1591.375 325.615 1591.390 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 1589.740 427.730 1589.800 ;
        RECT 460.070 1589.740 460.390 1589.800 ;
        RECT 427.410 1589.600 460.390 1589.740 ;
        RECT 427.410 1589.540 427.730 1589.600 ;
        RECT 460.070 1589.540 460.390 1589.600 ;
        RECT 424.650 20.640 424.970 20.700 ;
        RECT 427.410 20.640 427.730 20.700 ;
        RECT 424.650 20.500 427.730 20.640 ;
        RECT 424.650 20.440 424.970 20.500 ;
        RECT 427.410 20.440 427.730 20.500 ;
      LAYER via ;
        RECT 427.440 1589.540 427.700 1589.800 ;
        RECT 460.100 1589.540 460.360 1589.800 ;
        RECT 424.680 20.440 424.940 20.700 ;
        RECT 427.440 20.440 427.700 20.700 ;
      LAYER met2 ;
        RECT 460.100 1600.000 460.380 1604.000 ;
        RECT 460.160 1589.830 460.300 1600.000 ;
        RECT 427.440 1589.510 427.700 1589.830 ;
        RECT 460.100 1589.510 460.360 1589.830 ;
        RECT 427.500 20.730 427.640 1589.510 ;
        RECT 424.680 20.410 424.940 20.730 ;
        RECT 427.440 20.410 427.700 20.730 ;
        RECT 424.740 2.400 424.880 20.410 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 1589.400 448.430 1589.460 ;
        RECT 466.970 1589.400 467.290 1589.460 ;
        RECT 448.110 1589.260 467.290 1589.400 ;
        RECT 448.110 1589.200 448.430 1589.260 ;
        RECT 466.970 1589.200 467.290 1589.260 ;
        RECT 442.590 20.640 442.910 20.700 ;
        RECT 448.110 20.640 448.430 20.700 ;
        RECT 442.590 20.500 448.430 20.640 ;
        RECT 442.590 20.440 442.910 20.500 ;
        RECT 448.110 20.440 448.430 20.500 ;
      LAYER via ;
        RECT 448.140 1589.200 448.400 1589.460 ;
        RECT 467.000 1589.200 467.260 1589.460 ;
        RECT 442.620 20.440 442.880 20.700 ;
        RECT 448.140 20.440 448.400 20.700 ;
      LAYER met2 ;
        RECT 467.000 1600.000 467.280 1604.000 ;
        RECT 467.060 1589.490 467.200 1600.000 ;
        RECT 448.140 1589.170 448.400 1589.490 ;
        RECT 467.000 1589.170 467.260 1589.490 ;
        RECT 448.200 20.730 448.340 1589.170 ;
        RECT 442.620 20.410 442.880 20.730 ;
        RECT 448.140 20.410 448.400 20.730 ;
        RECT 442.680 2.400 442.820 20.410 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 1587.700 462.230 1587.760 ;
        RECT 473.410 1587.700 473.730 1587.760 ;
        RECT 461.910 1587.560 473.730 1587.700 ;
        RECT 461.910 1587.500 462.230 1587.560 ;
        RECT 473.410 1587.500 473.730 1587.560 ;
        RECT 460.530 2.960 460.850 3.020 ;
        RECT 461.910 2.960 462.230 3.020 ;
        RECT 460.530 2.820 462.230 2.960 ;
        RECT 460.530 2.760 460.850 2.820 ;
        RECT 461.910 2.760 462.230 2.820 ;
      LAYER via ;
        RECT 461.940 1587.500 462.200 1587.760 ;
        RECT 473.440 1587.500 473.700 1587.760 ;
        RECT 460.560 2.760 460.820 3.020 ;
        RECT 461.940 2.760 462.200 3.020 ;
      LAYER met2 ;
        RECT 473.440 1600.000 473.720 1604.000 ;
        RECT 473.500 1587.790 473.640 1600.000 ;
        RECT 461.940 1587.470 462.200 1587.790 ;
        RECT 473.440 1587.470 473.700 1587.790 ;
        RECT 462.000 3.050 462.140 1587.470 ;
        RECT 460.560 2.730 460.820 3.050 ;
        RECT 461.940 2.730 462.200 3.050 ;
        RECT 460.620 2.400 460.760 2.730 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 477.165 1497.445 477.335 1545.555 ;
        RECT 478.085 1352.605 478.255 1400.715 ;
        RECT 478.085 1256.045 478.255 1304.155 ;
        RECT 477.165 386.325 477.335 434.775 ;
        RECT 477.165 351.305 477.335 385.815 ;
        RECT 478.085 241.485 478.255 289.595 ;
        RECT 478.085 144.925 478.255 193.035 ;
        RECT 478.545 48.365 478.715 96.475 ;
      LAYER mcon ;
        RECT 477.165 1545.385 477.335 1545.555 ;
        RECT 478.085 1400.545 478.255 1400.715 ;
        RECT 478.085 1303.985 478.255 1304.155 ;
        RECT 477.165 434.605 477.335 434.775 ;
        RECT 477.165 385.645 477.335 385.815 ;
        RECT 478.085 289.425 478.255 289.595 ;
        RECT 478.085 192.865 478.255 193.035 ;
        RECT 478.545 96.305 478.715 96.475 ;
      LAYER met1 ;
        RECT 477.090 1545.540 477.410 1545.600 ;
        RECT 476.895 1545.400 477.410 1545.540 ;
        RECT 477.090 1545.340 477.410 1545.400 ;
        RECT 477.105 1497.600 477.395 1497.645 ;
        RECT 478.470 1497.600 478.790 1497.660 ;
        RECT 477.105 1497.460 478.790 1497.600 ;
        RECT 477.105 1497.415 477.395 1497.460 ;
        RECT 478.470 1497.400 478.790 1497.460 ;
        RECT 478.010 1400.700 478.330 1400.760 ;
        RECT 477.815 1400.560 478.330 1400.700 ;
        RECT 478.010 1400.500 478.330 1400.560 ;
        RECT 478.025 1352.760 478.315 1352.805 ;
        RECT 478.470 1352.760 478.790 1352.820 ;
        RECT 478.025 1352.620 478.790 1352.760 ;
        RECT 478.025 1352.575 478.315 1352.620 ;
        RECT 478.470 1352.560 478.790 1352.620 ;
        RECT 478.010 1304.140 478.330 1304.200 ;
        RECT 477.815 1304.000 478.330 1304.140 ;
        RECT 478.010 1303.940 478.330 1304.000 ;
        RECT 478.025 1256.200 478.315 1256.245 ;
        RECT 478.470 1256.200 478.790 1256.260 ;
        RECT 478.025 1256.060 478.790 1256.200 ;
        RECT 478.025 1256.015 478.315 1256.060 ;
        RECT 478.470 1256.000 478.790 1256.060 ;
        RECT 477.090 1159.300 477.410 1159.360 ;
        RECT 478.470 1159.300 478.790 1159.360 ;
        RECT 477.090 1159.160 478.790 1159.300 ;
        RECT 477.090 1159.100 477.410 1159.160 ;
        RECT 478.470 1159.100 478.790 1159.160 ;
        RECT 477.090 1062.740 477.410 1062.800 ;
        RECT 478.470 1062.740 478.790 1062.800 ;
        RECT 477.090 1062.600 478.790 1062.740 ;
        RECT 477.090 1062.540 477.410 1062.600 ;
        RECT 478.470 1062.540 478.790 1062.600 ;
        RECT 477.090 966.180 477.410 966.240 ;
        RECT 478.470 966.180 478.790 966.240 ;
        RECT 477.090 966.040 478.790 966.180 ;
        RECT 477.090 965.980 477.410 966.040 ;
        RECT 478.470 965.980 478.790 966.040 ;
        RECT 477.090 869.620 477.410 869.680 ;
        RECT 478.470 869.620 478.790 869.680 ;
        RECT 477.090 869.480 478.790 869.620 ;
        RECT 477.090 869.420 477.410 869.480 ;
        RECT 478.470 869.420 478.790 869.480 ;
        RECT 477.090 821.000 477.410 821.060 ;
        RECT 478.010 821.000 478.330 821.060 ;
        RECT 477.090 820.860 478.330 821.000 ;
        RECT 477.090 820.800 477.410 820.860 ;
        RECT 478.010 820.800 478.330 820.860 ;
        RECT 477.105 434.760 477.395 434.805 ;
        RECT 477.550 434.760 477.870 434.820 ;
        RECT 477.105 434.620 477.870 434.760 ;
        RECT 477.105 434.575 477.395 434.620 ;
        RECT 477.550 434.560 477.870 434.620 ;
        RECT 477.090 386.480 477.410 386.540 ;
        RECT 476.895 386.340 477.410 386.480 ;
        RECT 477.090 386.280 477.410 386.340 ;
        RECT 477.090 385.800 477.410 385.860 ;
        RECT 476.895 385.660 477.410 385.800 ;
        RECT 477.090 385.600 477.410 385.660 ;
        RECT 477.105 351.460 477.395 351.505 ;
        RECT 477.550 351.460 477.870 351.520 ;
        RECT 477.105 351.320 477.870 351.460 ;
        RECT 477.105 351.275 477.395 351.320 ;
        RECT 477.550 351.260 477.870 351.320 ;
        RECT 477.550 303.520 477.870 303.580 ;
        RECT 478.470 303.520 478.790 303.580 ;
        RECT 477.550 303.380 478.790 303.520 ;
        RECT 477.550 303.320 477.870 303.380 ;
        RECT 478.470 303.320 478.790 303.380 ;
        RECT 478.025 289.580 478.315 289.625 ;
        RECT 478.470 289.580 478.790 289.640 ;
        RECT 478.025 289.440 478.790 289.580 ;
        RECT 478.025 289.395 478.315 289.440 ;
        RECT 478.470 289.380 478.790 289.440 ;
        RECT 478.010 241.640 478.330 241.700 ;
        RECT 477.815 241.500 478.330 241.640 ;
        RECT 478.010 241.440 478.330 241.500 ;
        RECT 477.550 206.960 477.870 207.020 ;
        RECT 478.470 206.960 478.790 207.020 ;
        RECT 477.550 206.820 478.790 206.960 ;
        RECT 477.550 206.760 477.870 206.820 ;
        RECT 478.470 206.760 478.790 206.820 ;
        RECT 478.025 193.020 478.315 193.065 ;
        RECT 478.470 193.020 478.790 193.080 ;
        RECT 478.025 192.880 478.790 193.020 ;
        RECT 478.025 192.835 478.315 192.880 ;
        RECT 478.470 192.820 478.790 192.880 ;
        RECT 478.010 145.080 478.330 145.140 ;
        RECT 477.815 144.940 478.330 145.080 ;
        RECT 478.010 144.880 478.330 144.940 ;
        RECT 477.550 110.400 477.870 110.460 ;
        RECT 478.470 110.400 478.790 110.460 ;
        RECT 477.550 110.260 478.790 110.400 ;
        RECT 477.550 110.200 477.870 110.260 ;
        RECT 478.470 110.200 478.790 110.260 ;
        RECT 478.470 96.460 478.790 96.520 ;
        RECT 478.275 96.320 478.790 96.460 ;
        RECT 478.470 96.260 478.790 96.320 ;
        RECT 478.470 48.520 478.790 48.580 ;
        RECT 478.275 48.380 478.790 48.520 ;
        RECT 478.470 48.320 478.790 48.380 ;
        RECT 477.090 14.180 477.410 14.240 ;
        RECT 478.470 14.180 478.790 14.240 ;
        RECT 477.090 14.040 478.790 14.180 ;
        RECT 477.090 13.980 477.410 14.040 ;
        RECT 478.470 13.980 478.790 14.040 ;
        RECT 477.090 2.960 477.410 3.020 ;
        RECT 478.470 2.960 478.790 3.020 ;
        RECT 477.090 2.820 478.790 2.960 ;
        RECT 477.090 2.760 477.410 2.820 ;
        RECT 478.470 2.760 478.790 2.820 ;
      LAYER via ;
        RECT 477.120 1545.340 477.380 1545.600 ;
        RECT 478.500 1497.400 478.760 1497.660 ;
        RECT 478.040 1400.500 478.300 1400.760 ;
        RECT 478.500 1352.560 478.760 1352.820 ;
        RECT 478.040 1303.940 478.300 1304.200 ;
        RECT 478.500 1256.000 478.760 1256.260 ;
        RECT 477.120 1159.100 477.380 1159.360 ;
        RECT 478.500 1159.100 478.760 1159.360 ;
        RECT 477.120 1062.540 477.380 1062.800 ;
        RECT 478.500 1062.540 478.760 1062.800 ;
        RECT 477.120 965.980 477.380 966.240 ;
        RECT 478.500 965.980 478.760 966.240 ;
        RECT 477.120 869.420 477.380 869.680 ;
        RECT 478.500 869.420 478.760 869.680 ;
        RECT 477.120 820.800 477.380 821.060 ;
        RECT 478.040 820.800 478.300 821.060 ;
        RECT 477.580 434.560 477.840 434.820 ;
        RECT 477.120 386.280 477.380 386.540 ;
        RECT 477.120 385.600 477.380 385.860 ;
        RECT 477.580 351.260 477.840 351.520 ;
        RECT 477.580 303.320 477.840 303.580 ;
        RECT 478.500 303.320 478.760 303.580 ;
        RECT 478.500 289.380 478.760 289.640 ;
        RECT 478.040 241.440 478.300 241.700 ;
        RECT 477.580 206.760 477.840 207.020 ;
        RECT 478.500 206.760 478.760 207.020 ;
        RECT 478.500 192.820 478.760 193.080 ;
        RECT 478.040 144.880 478.300 145.140 ;
        RECT 477.580 110.200 477.840 110.460 ;
        RECT 478.500 110.200 478.760 110.460 ;
        RECT 478.500 96.260 478.760 96.520 ;
        RECT 478.500 48.320 478.760 48.580 ;
        RECT 477.120 13.980 477.380 14.240 ;
        RECT 478.500 13.980 478.760 14.240 ;
        RECT 477.120 2.760 477.380 3.020 ;
        RECT 478.500 2.760 478.760 3.020 ;
      LAYER met2 ;
        RECT 480.340 1600.450 480.620 1604.000 ;
        RECT 479.020 1600.310 480.620 1600.450 ;
        RECT 479.020 1580.050 479.160 1600.310 ;
        RECT 480.340 1600.000 480.620 1600.310 ;
        RECT 477.180 1579.910 479.160 1580.050 ;
        RECT 477.180 1545.630 477.320 1579.910 ;
        RECT 477.120 1545.310 477.380 1545.630 ;
        RECT 478.500 1497.370 478.760 1497.690 ;
        RECT 478.560 1425.010 478.700 1497.370 ;
        RECT 478.100 1424.870 478.700 1425.010 ;
        RECT 478.100 1400.790 478.240 1424.870 ;
        RECT 478.040 1400.470 478.300 1400.790 ;
        RECT 478.500 1352.530 478.760 1352.850 ;
        RECT 478.560 1317.570 478.700 1352.530 ;
        RECT 478.100 1317.430 478.700 1317.570 ;
        RECT 478.100 1304.230 478.240 1317.430 ;
        RECT 478.040 1303.910 478.300 1304.230 ;
        RECT 478.500 1255.970 478.760 1256.290 ;
        RECT 478.560 1221.010 478.700 1255.970 ;
        RECT 478.100 1220.870 478.700 1221.010 ;
        RECT 478.100 1207.525 478.240 1220.870 ;
        RECT 477.110 1207.155 477.390 1207.525 ;
        RECT 478.030 1207.155 478.310 1207.525 ;
        RECT 477.180 1159.390 477.320 1207.155 ;
        RECT 477.120 1159.070 477.380 1159.390 ;
        RECT 478.500 1159.070 478.760 1159.390 ;
        RECT 478.560 1124.450 478.700 1159.070 ;
        RECT 478.100 1124.310 478.700 1124.450 ;
        RECT 478.100 1110.965 478.240 1124.310 ;
        RECT 477.110 1110.595 477.390 1110.965 ;
        RECT 478.030 1110.595 478.310 1110.965 ;
        RECT 477.180 1062.830 477.320 1110.595 ;
        RECT 477.120 1062.510 477.380 1062.830 ;
        RECT 478.500 1062.510 478.760 1062.830 ;
        RECT 478.560 1027.890 478.700 1062.510 ;
        RECT 478.100 1027.750 478.700 1027.890 ;
        RECT 478.100 1014.405 478.240 1027.750 ;
        RECT 477.110 1014.035 477.390 1014.405 ;
        RECT 478.030 1014.035 478.310 1014.405 ;
        RECT 477.180 966.270 477.320 1014.035 ;
        RECT 477.120 965.950 477.380 966.270 ;
        RECT 478.500 965.950 478.760 966.270 ;
        RECT 478.560 931.330 478.700 965.950 ;
        RECT 478.100 931.190 478.700 931.330 ;
        RECT 478.100 917.845 478.240 931.190 ;
        RECT 477.110 917.475 477.390 917.845 ;
        RECT 478.030 917.475 478.310 917.845 ;
        RECT 477.180 869.710 477.320 917.475 ;
        RECT 477.120 869.390 477.380 869.710 ;
        RECT 478.500 869.390 478.760 869.710 ;
        RECT 478.560 834.770 478.700 869.390 ;
        RECT 478.100 834.630 478.700 834.770 ;
        RECT 478.100 821.090 478.240 834.630 ;
        RECT 477.120 820.770 477.380 821.090 ;
        RECT 478.040 820.770 478.300 821.090 ;
        RECT 477.180 773.005 477.320 820.770 ;
        RECT 477.110 772.635 477.390 773.005 ;
        RECT 478.490 772.635 478.770 773.005 ;
        RECT 478.560 738.210 478.700 772.635 ;
        RECT 478.100 738.070 478.700 738.210 ;
        RECT 478.100 700.130 478.240 738.070 ;
        RECT 477.180 699.990 478.240 700.130 ;
        RECT 477.180 676.445 477.320 699.990 ;
        RECT 477.110 676.075 477.390 676.445 ;
        RECT 478.490 676.075 478.770 676.445 ;
        RECT 478.560 641.650 478.700 676.075 ;
        RECT 478.100 641.510 478.700 641.650 ;
        RECT 478.100 603.570 478.240 641.510 ;
        RECT 477.180 603.430 478.240 603.570 ;
        RECT 477.180 579.885 477.320 603.430 ;
        RECT 477.110 579.515 477.390 579.885 ;
        RECT 478.490 579.515 478.770 579.885 ;
        RECT 478.560 545.090 478.700 579.515 ;
        RECT 478.100 544.950 478.700 545.090 ;
        RECT 478.100 507.010 478.240 544.950 ;
        RECT 477.180 506.870 478.240 507.010 ;
        RECT 477.180 483.325 477.320 506.870 ;
        RECT 477.110 482.955 477.390 483.325 ;
        RECT 478.490 482.955 478.770 483.325 ;
        RECT 478.560 448.530 478.700 482.955 ;
        RECT 477.640 448.390 478.700 448.530 ;
        RECT 477.640 434.850 477.780 448.390 ;
        RECT 477.580 434.530 477.840 434.850 ;
        RECT 477.120 386.250 477.380 386.570 ;
        RECT 477.180 385.890 477.320 386.250 ;
        RECT 477.120 385.570 477.380 385.890 ;
        RECT 477.580 351.230 477.840 351.550 ;
        RECT 477.640 303.610 477.780 351.230 ;
        RECT 477.580 303.290 477.840 303.610 ;
        RECT 478.500 303.290 478.760 303.610 ;
        RECT 478.560 289.670 478.700 303.290 ;
        RECT 478.500 289.350 478.760 289.670 ;
        RECT 478.040 241.410 478.300 241.730 ;
        RECT 478.100 207.130 478.240 241.410 ;
        RECT 477.640 207.050 478.240 207.130 ;
        RECT 477.580 206.990 478.240 207.050 ;
        RECT 477.580 206.730 477.840 206.990 ;
        RECT 478.500 206.730 478.760 207.050 ;
        RECT 478.560 193.110 478.700 206.730 ;
        RECT 478.500 192.790 478.760 193.110 ;
        RECT 478.040 144.850 478.300 145.170 ;
        RECT 478.100 110.570 478.240 144.850 ;
        RECT 477.640 110.490 478.240 110.570 ;
        RECT 477.580 110.430 478.240 110.490 ;
        RECT 477.580 110.170 477.840 110.430 ;
        RECT 478.500 110.170 478.760 110.490 ;
        RECT 478.560 96.550 478.700 110.170 ;
        RECT 478.500 96.230 478.760 96.550 ;
        RECT 478.500 48.290 478.760 48.610 ;
        RECT 478.560 14.270 478.700 48.290 ;
        RECT 477.120 13.950 477.380 14.270 ;
        RECT 478.500 13.950 478.760 14.270 ;
        RECT 477.180 3.050 477.320 13.950 ;
        RECT 477.120 2.730 477.380 3.050 ;
        RECT 478.500 2.730 478.760 3.050 ;
        RECT 478.560 2.400 478.700 2.730 ;
        RECT 478.350 -4.800 478.910 2.400 ;
      LAYER via2 ;
        RECT 477.110 1207.200 477.390 1207.480 ;
        RECT 478.030 1207.200 478.310 1207.480 ;
        RECT 477.110 1110.640 477.390 1110.920 ;
        RECT 478.030 1110.640 478.310 1110.920 ;
        RECT 477.110 1014.080 477.390 1014.360 ;
        RECT 478.030 1014.080 478.310 1014.360 ;
        RECT 477.110 917.520 477.390 917.800 ;
        RECT 478.030 917.520 478.310 917.800 ;
        RECT 477.110 772.680 477.390 772.960 ;
        RECT 478.490 772.680 478.770 772.960 ;
        RECT 477.110 676.120 477.390 676.400 ;
        RECT 478.490 676.120 478.770 676.400 ;
        RECT 477.110 579.560 477.390 579.840 ;
        RECT 478.490 579.560 478.770 579.840 ;
        RECT 477.110 483.000 477.390 483.280 ;
        RECT 478.490 483.000 478.770 483.280 ;
      LAYER met3 ;
        RECT 477.085 1207.490 477.415 1207.505 ;
        RECT 478.005 1207.490 478.335 1207.505 ;
        RECT 477.085 1207.190 478.335 1207.490 ;
        RECT 477.085 1207.175 477.415 1207.190 ;
        RECT 478.005 1207.175 478.335 1207.190 ;
        RECT 477.085 1110.930 477.415 1110.945 ;
        RECT 478.005 1110.930 478.335 1110.945 ;
        RECT 477.085 1110.630 478.335 1110.930 ;
        RECT 477.085 1110.615 477.415 1110.630 ;
        RECT 478.005 1110.615 478.335 1110.630 ;
        RECT 477.085 1014.370 477.415 1014.385 ;
        RECT 478.005 1014.370 478.335 1014.385 ;
        RECT 477.085 1014.070 478.335 1014.370 ;
        RECT 477.085 1014.055 477.415 1014.070 ;
        RECT 478.005 1014.055 478.335 1014.070 ;
        RECT 477.085 917.810 477.415 917.825 ;
        RECT 478.005 917.810 478.335 917.825 ;
        RECT 477.085 917.510 478.335 917.810 ;
        RECT 477.085 917.495 477.415 917.510 ;
        RECT 478.005 917.495 478.335 917.510 ;
        RECT 477.085 772.970 477.415 772.985 ;
        RECT 478.465 772.970 478.795 772.985 ;
        RECT 477.085 772.670 478.795 772.970 ;
        RECT 477.085 772.655 477.415 772.670 ;
        RECT 478.465 772.655 478.795 772.670 ;
        RECT 477.085 676.410 477.415 676.425 ;
        RECT 478.465 676.410 478.795 676.425 ;
        RECT 477.085 676.110 478.795 676.410 ;
        RECT 477.085 676.095 477.415 676.110 ;
        RECT 478.465 676.095 478.795 676.110 ;
        RECT 477.085 579.850 477.415 579.865 ;
        RECT 478.465 579.850 478.795 579.865 ;
        RECT 477.085 579.550 478.795 579.850 ;
        RECT 477.085 579.535 477.415 579.550 ;
        RECT 478.465 579.535 478.795 579.550 ;
        RECT 477.085 483.290 477.415 483.305 ;
        RECT 478.465 483.290 478.795 483.305 ;
        RECT 477.085 482.990 478.795 483.290 ;
        RECT 477.085 482.975 477.415 482.990 ;
        RECT 478.465 482.975 478.795 482.990 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 487.210 1587.700 487.530 1587.760 ;
        RECT 489.510 1587.700 489.830 1587.760 ;
        RECT 487.210 1587.560 489.830 1587.700 ;
        RECT 487.210 1587.500 487.530 1587.560 ;
        RECT 489.510 1587.500 489.830 1587.560 ;
        RECT 489.510 20.640 489.830 20.700 ;
        RECT 496.410 20.640 496.730 20.700 ;
        RECT 489.510 20.500 496.730 20.640 ;
        RECT 489.510 20.440 489.830 20.500 ;
        RECT 496.410 20.440 496.730 20.500 ;
      LAYER via ;
        RECT 487.240 1587.500 487.500 1587.760 ;
        RECT 489.540 1587.500 489.800 1587.760 ;
        RECT 489.540 20.440 489.800 20.700 ;
        RECT 496.440 20.440 496.700 20.700 ;
      LAYER met2 ;
        RECT 487.240 1600.000 487.520 1604.000 ;
        RECT 487.300 1587.790 487.440 1600.000 ;
        RECT 487.240 1587.470 487.500 1587.790 ;
        RECT 489.540 1587.470 489.800 1587.790 ;
        RECT 489.600 20.730 489.740 1587.470 ;
        RECT 489.540 20.410 489.800 20.730 ;
        RECT 496.440 20.410 496.700 20.730 ;
        RECT 496.500 2.400 496.640 20.410 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 493.650 1590.420 493.970 1590.480 ;
        RECT 512.050 1590.420 512.370 1590.480 ;
        RECT 493.650 1590.280 512.370 1590.420 ;
        RECT 493.650 1590.220 493.970 1590.280 ;
        RECT 512.050 1590.220 512.370 1590.280 ;
      LAYER via ;
        RECT 493.680 1590.220 493.940 1590.480 ;
        RECT 512.080 1590.220 512.340 1590.480 ;
      LAYER met2 ;
        RECT 493.680 1600.000 493.960 1604.000 ;
        RECT 493.740 1590.510 493.880 1600.000 ;
        RECT 493.680 1590.190 493.940 1590.510 ;
        RECT 512.080 1590.190 512.340 1590.510 ;
        RECT 512.140 16.730 512.280 1590.190 ;
        RECT 512.140 16.590 514.120 16.730 ;
        RECT 513.980 2.400 514.120 16.590 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 503.310 17.920 503.630 17.980 ;
        RECT 531.830 17.920 532.150 17.980 ;
        RECT 503.310 17.780 532.150 17.920 ;
        RECT 503.310 17.720 503.630 17.780 ;
        RECT 531.830 17.720 532.150 17.780 ;
      LAYER via ;
        RECT 503.340 17.720 503.600 17.980 ;
        RECT 531.860 17.720 532.120 17.980 ;
      LAYER met2 ;
        RECT 500.580 1601.130 500.860 1604.000 ;
        RECT 500.580 1600.990 502.620 1601.130 ;
        RECT 500.580 1600.000 500.860 1600.990 ;
        RECT 502.480 1587.700 502.620 1600.990 ;
        RECT 502.480 1587.560 503.540 1587.700 ;
        RECT 503.400 18.010 503.540 1587.560 ;
        RECT 503.340 17.690 503.600 18.010 ;
        RECT 531.860 17.690 532.120 18.010 ;
        RECT 531.920 2.400 532.060 17.690 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 509.750 17.580 510.070 17.640 ;
        RECT 549.770 17.580 550.090 17.640 ;
        RECT 509.750 17.440 550.090 17.580 ;
        RECT 509.750 17.380 510.070 17.440 ;
        RECT 549.770 17.380 550.090 17.440 ;
      LAYER via ;
        RECT 509.780 17.380 510.040 17.640 ;
        RECT 549.800 17.380 550.060 17.640 ;
      LAYER met2 ;
        RECT 507.020 1601.130 507.300 1604.000 ;
        RECT 507.020 1600.990 509.060 1601.130 ;
        RECT 507.020 1600.000 507.300 1600.990 ;
        RECT 508.920 1590.250 509.060 1600.990 ;
        RECT 508.920 1590.110 509.980 1590.250 ;
        RECT 509.840 17.670 509.980 1590.110 ;
        RECT 509.780 17.350 510.040 17.670 ;
        RECT 549.800 17.350 550.060 17.670 ;
        RECT 549.860 2.400 550.000 17.350 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 513.890 1590.420 514.210 1590.480 ;
        RECT 516.650 1590.420 516.970 1590.480 ;
        RECT 513.890 1590.280 516.970 1590.420 ;
        RECT 513.890 1590.220 514.210 1590.280 ;
        RECT 516.650 1590.220 516.970 1590.280 ;
        RECT 516.650 15.880 516.970 15.940 ;
        RECT 567.710 15.880 568.030 15.940 ;
        RECT 516.650 15.740 568.030 15.880 ;
        RECT 516.650 15.680 516.970 15.740 ;
        RECT 567.710 15.680 568.030 15.740 ;
      LAYER via ;
        RECT 513.920 1590.220 514.180 1590.480 ;
        RECT 516.680 1590.220 516.940 1590.480 ;
        RECT 516.680 15.680 516.940 15.940 ;
        RECT 567.740 15.680 568.000 15.940 ;
      LAYER met2 ;
        RECT 513.920 1600.000 514.200 1604.000 ;
        RECT 513.980 1590.510 514.120 1600.000 ;
        RECT 513.920 1590.190 514.180 1590.510 ;
        RECT 516.680 1590.190 516.940 1590.510 ;
        RECT 516.740 15.970 516.880 1590.190 ;
        RECT 516.680 15.650 516.940 15.970 ;
        RECT 567.740 15.650 568.000 15.970 ;
        RECT 567.800 2.400 567.940 15.650 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 523.090 20.640 523.410 20.700 ;
        RECT 585.650 20.640 585.970 20.700 ;
        RECT 523.090 20.500 585.970 20.640 ;
        RECT 523.090 20.440 523.410 20.500 ;
        RECT 585.650 20.440 585.970 20.500 ;
      LAYER via ;
        RECT 523.120 20.440 523.380 20.700 ;
        RECT 585.680 20.440 585.940 20.700 ;
      LAYER met2 ;
        RECT 520.820 1601.130 521.100 1604.000 ;
        RECT 520.820 1600.990 522.860 1601.130 ;
        RECT 520.820 1600.000 521.100 1600.990 ;
        RECT 522.720 1590.250 522.860 1600.990 ;
        RECT 522.720 1590.110 523.320 1590.250 ;
        RECT 523.180 20.730 523.320 1590.110 ;
        RECT 523.120 20.410 523.380 20.730 ;
        RECT 585.680 20.410 585.940 20.730 ;
        RECT 585.740 2.400 585.880 20.410 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 334.105 1497.445 334.275 1545.555 ;
        RECT 332.725 1352.605 332.895 1400.715 ;
        RECT 332.725 1256.045 332.895 1304.155 ;
        RECT 331.805 386.325 331.975 434.775 ;
        RECT 331.805 351.305 331.975 385.815 ;
        RECT 332.725 241.485 332.895 289.595 ;
        RECT 332.725 144.925 332.895 193.035 ;
        RECT 333.185 48.365 333.355 96.475 ;
      LAYER mcon ;
        RECT 334.105 1545.385 334.275 1545.555 ;
        RECT 332.725 1400.545 332.895 1400.715 ;
        RECT 332.725 1303.985 332.895 1304.155 ;
        RECT 331.805 434.605 331.975 434.775 ;
        RECT 331.805 385.645 331.975 385.815 ;
        RECT 332.725 289.425 332.895 289.595 ;
        RECT 332.725 192.865 332.895 193.035 ;
        RECT 333.185 96.305 333.355 96.475 ;
      LAYER met1 ;
        RECT 334.030 1569.680 334.350 1569.740 ;
        RECT 334.950 1569.680 335.270 1569.740 ;
        RECT 334.030 1569.540 335.270 1569.680 ;
        RECT 334.030 1569.480 334.350 1569.540 ;
        RECT 334.950 1569.480 335.270 1569.540 ;
        RECT 334.045 1545.540 334.335 1545.585 ;
        RECT 334.950 1545.540 335.270 1545.600 ;
        RECT 334.045 1545.400 335.270 1545.540 ;
        RECT 334.045 1545.355 334.335 1545.400 ;
        RECT 334.950 1545.340 335.270 1545.400 ;
        RECT 334.030 1497.600 334.350 1497.660 ;
        RECT 333.835 1497.460 334.350 1497.600 ;
        RECT 334.030 1497.400 334.350 1497.460 ;
        RECT 333.110 1473.120 333.430 1473.180 ;
        RECT 334.030 1473.120 334.350 1473.180 ;
        RECT 333.110 1472.980 334.350 1473.120 ;
        RECT 333.110 1472.920 333.430 1472.980 ;
        RECT 334.030 1472.920 334.350 1472.980 ;
        RECT 332.650 1400.700 332.970 1400.760 ;
        RECT 332.455 1400.560 332.970 1400.700 ;
        RECT 332.650 1400.500 332.970 1400.560 ;
        RECT 332.665 1352.760 332.955 1352.805 ;
        RECT 333.110 1352.760 333.430 1352.820 ;
        RECT 332.665 1352.620 333.430 1352.760 ;
        RECT 332.665 1352.575 332.955 1352.620 ;
        RECT 333.110 1352.560 333.430 1352.620 ;
        RECT 332.650 1304.140 332.970 1304.200 ;
        RECT 332.455 1304.000 332.970 1304.140 ;
        RECT 332.650 1303.940 332.970 1304.000 ;
        RECT 332.665 1256.200 332.955 1256.245 ;
        RECT 333.110 1256.200 333.430 1256.260 ;
        RECT 332.665 1256.060 333.430 1256.200 ;
        RECT 332.665 1256.015 332.955 1256.060 ;
        RECT 333.110 1256.000 333.430 1256.060 ;
        RECT 331.730 1159.300 332.050 1159.360 ;
        RECT 333.110 1159.300 333.430 1159.360 ;
        RECT 331.730 1159.160 333.430 1159.300 ;
        RECT 331.730 1159.100 332.050 1159.160 ;
        RECT 333.110 1159.100 333.430 1159.160 ;
        RECT 331.730 1062.740 332.050 1062.800 ;
        RECT 333.110 1062.740 333.430 1062.800 ;
        RECT 331.730 1062.600 333.430 1062.740 ;
        RECT 331.730 1062.540 332.050 1062.600 ;
        RECT 333.110 1062.540 333.430 1062.600 ;
        RECT 331.730 966.180 332.050 966.240 ;
        RECT 333.110 966.180 333.430 966.240 ;
        RECT 331.730 966.040 333.430 966.180 ;
        RECT 331.730 965.980 332.050 966.040 ;
        RECT 333.110 965.980 333.430 966.040 ;
        RECT 331.730 869.620 332.050 869.680 ;
        RECT 333.110 869.620 333.430 869.680 ;
        RECT 331.730 869.480 333.430 869.620 ;
        RECT 331.730 869.420 332.050 869.480 ;
        RECT 333.110 869.420 333.430 869.480 ;
        RECT 331.730 821.000 332.050 821.060 ;
        RECT 332.650 821.000 332.970 821.060 ;
        RECT 331.730 820.860 332.970 821.000 ;
        RECT 331.730 820.800 332.050 820.860 ;
        RECT 332.650 820.800 332.970 820.860 ;
        RECT 331.745 434.760 332.035 434.805 ;
        RECT 332.190 434.760 332.510 434.820 ;
        RECT 331.745 434.620 332.510 434.760 ;
        RECT 331.745 434.575 332.035 434.620 ;
        RECT 332.190 434.560 332.510 434.620 ;
        RECT 331.730 386.480 332.050 386.540 ;
        RECT 331.535 386.340 332.050 386.480 ;
        RECT 331.730 386.280 332.050 386.340 ;
        RECT 331.730 385.800 332.050 385.860 ;
        RECT 331.535 385.660 332.050 385.800 ;
        RECT 331.730 385.600 332.050 385.660 ;
        RECT 331.745 351.460 332.035 351.505 ;
        RECT 332.190 351.460 332.510 351.520 ;
        RECT 331.745 351.320 332.510 351.460 ;
        RECT 331.745 351.275 332.035 351.320 ;
        RECT 332.190 351.260 332.510 351.320 ;
        RECT 332.190 303.520 332.510 303.580 ;
        RECT 333.110 303.520 333.430 303.580 ;
        RECT 332.190 303.380 333.430 303.520 ;
        RECT 332.190 303.320 332.510 303.380 ;
        RECT 333.110 303.320 333.430 303.380 ;
        RECT 332.665 289.580 332.955 289.625 ;
        RECT 333.110 289.580 333.430 289.640 ;
        RECT 332.665 289.440 333.430 289.580 ;
        RECT 332.665 289.395 332.955 289.440 ;
        RECT 333.110 289.380 333.430 289.440 ;
        RECT 332.650 241.640 332.970 241.700 ;
        RECT 332.455 241.500 332.970 241.640 ;
        RECT 332.650 241.440 332.970 241.500 ;
        RECT 332.190 206.960 332.510 207.020 ;
        RECT 333.110 206.960 333.430 207.020 ;
        RECT 332.190 206.820 333.430 206.960 ;
        RECT 332.190 206.760 332.510 206.820 ;
        RECT 333.110 206.760 333.430 206.820 ;
        RECT 332.665 193.020 332.955 193.065 ;
        RECT 333.110 193.020 333.430 193.080 ;
        RECT 332.665 192.880 333.430 193.020 ;
        RECT 332.665 192.835 332.955 192.880 ;
        RECT 333.110 192.820 333.430 192.880 ;
        RECT 332.650 145.080 332.970 145.140 ;
        RECT 332.455 144.940 332.970 145.080 ;
        RECT 332.650 144.880 332.970 144.940 ;
        RECT 332.190 110.400 332.510 110.460 ;
        RECT 333.110 110.400 333.430 110.460 ;
        RECT 332.190 110.260 333.430 110.400 ;
        RECT 332.190 110.200 332.510 110.260 ;
        RECT 333.110 110.200 333.430 110.260 ;
        RECT 333.110 96.460 333.430 96.520 ;
        RECT 332.915 96.320 333.430 96.460 ;
        RECT 333.110 96.260 333.430 96.320 ;
        RECT 333.110 48.520 333.430 48.580 ;
        RECT 332.915 48.380 333.430 48.520 ;
        RECT 333.110 48.320 333.430 48.380 ;
        RECT 91.610 19.620 91.930 19.680 ;
        RECT 333.110 19.620 333.430 19.680 ;
        RECT 91.610 19.480 333.430 19.620 ;
        RECT 91.610 19.420 91.930 19.480 ;
        RECT 333.110 19.420 333.430 19.480 ;
      LAYER via ;
        RECT 334.060 1569.480 334.320 1569.740 ;
        RECT 334.980 1569.480 335.240 1569.740 ;
        RECT 334.980 1545.340 335.240 1545.600 ;
        RECT 334.060 1497.400 334.320 1497.660 ;
        RECT 333.140 1472.920 333.400 1473.180 ;
        RECT 334.060 1472.920 334.320 1473.180 ;
        RECT 332.680 1400.500 332.940 1400.760 ;
        RECT 333.140 1352.560 333.400 1352.820 ;
        RECT 332.680 1303.940 332.940 1304.200 ;
        RECT 333.140 1256.000 333.400 1256.260 ;
        RECT 331.760 1159.100 332.020 1159.360 ;
        RECT 333.140 1159.100 333.400 1159.360 ;
        RECT 331.760 1062.540 332.020 1062.800 ;
        RECT 333.140 1062.540 333.400 1062.800 ;
        RECT 331.760 965.980 332.020 966.240 ;
        RECT 333.140 965.980 333.400 966.240 ;
        RECT 331.760 869.420 332.020 869.680 ;
        RECT 333.140 869.420 333.400 869.680 ;
        RECT 331.760 820.800 332.020 821.060 ;
        RECT 332.680 820.800 332.940 821.060 ;
        RECT 332.220 434.560 332.480 434.820 ;
        RECT 331.760 386.280 332.020 386.540 ;
        RECT 331.760 385.600 332.020 385.860 ;
        RECT 332.220 351.260 332.480 351.520 ;
        RECT 332.220 303.320 332.480 303.580 ;
        RECT 333.140 303.320 333.400 303.580 ;
        RECT 333.140 289.380 333.400 289.640 ;
        RECT 332.680 241.440 332.940 241.700 ;
        RECT 332.220 206.760 332.480 207.020 ;
        RECT 333.140 206.760 333.400 207.020 ;
        RECT 333.140 192.820 333.400 193.080 ;
        RECT 332.680 144.880 332.940 145.140 ;
        RECT 332.220 110.200 332.480 110.460 ;
        RECT 333.140 110.200 333.400 110.460 ;
        RECT 333.140 96.260 333.400 96.520 ;
        RECT 333.140 48.320 333.400 48.580 ;
        RECT 91.640 19.420 91.900 19.680 ;
        RECT 333.140 19.420 333.400 19.680 ;
      LAYER met2 ;
        RECT 334.520 1600.450 334.800 1604.000 ;
        RECT 334.120 1600.310 334.800 1600.450 ;
        RECT 334.120 1569.770 334.260 1600.310 ;
        RECT 334.520 1600.000 334.800 1600.310 ;
        RECT 334.060 1569.450 334.320 1569.770 ;
        RECT 334.980 1569.450 335.240 1569.770 ;
        RECT 335.040 1545.630 335.180 1569.450 ;
        RECT 334.980 1545.310 335.240 1545.630 ;
        RECT 334.060 1497.370 334.320 1497.690 ;
        RECT 334.120 1473.210 334.260 1497.370 ;
        RECT 333.140 1472.890 333.400 1473.210 ;
        RECT 334.060 1472.890 334.320 1473.210 ;
        RECT 333.200 1414.130 333.340 1472.890 ;
        RECT 332.740 1413.990 333.340 1414.130 ;
        RECT 332.740 1400.790 332.880 1413.990 ;
        RECT 332.680 1400.470 332.940 1400.790 ;
        RECT 333.140 1352.530 333.400 1352.850 ;
        RECT 333.200 1317.570 333.340 1352.530 ;
        RECT 332.740 1317.430 333.340 1317.570 ;
        RECT 332.740 1304.230 332.880 1317.430 ;
        RECT 332.680 1303.910 332.940 1304.230 ;
        RECT 333.140 1255.970 333.400 1256.290 ;
        RECT 333.200 1221.010 333.340 1255.970 ;
        RECT 332.740 1220.870 333.340 1221.010 ;
        RECT 332.740 1207.525 332.880 1220.870 ;
        RECT 331.750 1207.155 332.030 1207.525 ;
        RECT 332.670 1207.155 332.950 1207.525 ;
        RECT 331.820 1159.390 331.960 1207.155 ;
        RECT 331.760 1159.070 332.020 1159.390 ;
        RECT 333.140 1159.070 333.400 1159.390 ;
        RECT 333.200 1124.450 333.340 1159.070 ;
        RECT 332.740 1124.310 333.340 1124.450 ;
        RECT 332.740 1110.965 332.880 1124.310 ;
        RECT 331.750 1110.595 332.030 1110.965 ;
        RECT 332.670 1110.595 332.950 1110.965 ;
        RECT 331.820 1062.830 331.960 1110.595 ;
        RECT 331.760 1062.510 332.020 1062.830 ;
        RECT 333.140 1062.510 333.400 1062.830 ;
        RECT 333.200 1027.890 333.340 1062.510 ;
        RECT 332.740 1027.750 333.340 1027.890 ;
        RECT 332.740 1014.405 332.880 1027.750 ;
        RECT 331.750 1014.035 332.030 1014.405 ;
        RECT 332.670 1014.035 332.950 1014.405 ;
        RECT 331.820 966.270 331.960 1014.035 ;
        RECT 331.760 965.950 332.020 966.270 ;
        RECT 333.140 965.950 333.400 966.270 ;
        RECT 333.200 931.330 333.340 965.950 ;
        RECT 332.740 931.190 333.340 931.330 ;
        RECT 332.740 917.845 332.880 931.190 ;
        RECT 331.750 917.475 332.030 917.845 ;
        RECT 332.670 917.475 332.950 917.845 ;
        RECT 331.820 869.710 331.960 917.475 ;
        RECT 331.760 869.390 332.020 869.710 ;
        RECT 333.140 869.390 333.400 869.710 ;
        RECT 333.200 834.770 333.340 869.390 ;
        RECT 332.740 834.630 333.340 834.770 ;
        RECT 332.740 821.090 332.880 834.630 ;
        RECT 331.760 820.770 332.020 821.090 ;
        RECT 332.680 820.770 332.940 821.090 ;
        RECT 331.820 773.005 331.960 820.770 ;
        RECT 331.750 772.635 332.030 773.005 ;
        RECT 333.130 772.635 333.410 773.005 ;
        RECT 333.200 738.210 333.340 772.635 ;
        RECT 332.740 738.070 333.340 738.210 ;
        RECT 332.740 700.130 332.880 738.070 ;
        RECT 331.820 699.990 332.880 700.130 ;
        RECT 331.820 676.445 331.960 699.990 ;
        RECT 331.750 676.075 332.030 676.445 ;
        RECT 333.130 676.075 333.410 676.445 ;
        RECT 333.200 641.650 333.340 676.075 ;
        RECT 332.740 641.510 333.340 641.650 ;
        RECT 332.740 603.570 332.880 641.510 ;
        RECT 331.820 603.430 332.880 603.570 ;
        RECT 331.820 579.885 331.960 603.430 ;
        RECT 331.750 579.515 332.030 579.885 ;
        RECT 333.130 579.515 333.410 579.885 ;
        RECT 333.200 545.090 333.340 579.515 ;
        RECT 332.740 544.950 333.340 545.090 ;
        RECT 332.740 507.010 332.880 544.950 ;
        RECT 331.820 506.870 332.880 507.010 ;
        RECT 331.820 483.325 331.960 506.870 ;
        RECT 331.750 482.955 332.030 483.325 ;
        RECT 333.130 482.955 333.410 483.325 ;
        RECT 333.200 448.530 333.340 482.955 ;
        RECT 332.280 448.390 333.340 448.530 ;
        RECT 332.280 434.850 332.420 448.390 ;
        RECT 332.220 434.530 332.480 434.850 ;
        RECT 331.760 386.250 332.020 386.570 ;
        RECT 331.820 385.890 331.960 386.250 ;
        RECT 331.760 385.570 332.020 385.890 ;
        RECT 332.220 351.230 332.480 351.550 ;
        RECT 332.280 303.610 332.420 351.230 ;
        RECT 332.220 303.290 332.480 303.610 ;
        RECT 333.140 303.290 333.400 303.610 ;
        RECT 333.200 289.670 333.340 303.290 ;
        RECT 333.140 289.350 333.400 289.670 ;
        RECT 332.680 241.410 332.940 241.730 ;
        RECT 332.740 207.130 332.880 241.410 ;
        RECT 332.280 207.050 332.880 207.130 ;
        RECT 332.220 206.990 332.880 207.050 ;
        RECT 332.220 206.730 332.480 206.990 ;
        RECT 333.140 206.730 333.400 207.050 ;
        RECT 333.200 193.110 333.340 206.730 ;
        RECT 333.140 192.790 333.400 193.110 ;
        RECT 332.680 144.850 332.940 145.170 ;
        RECT 332.740 110.570 332.880 144.850 ;
        RECT 332.280 110.490 332.880 110.570 ;
        RECT 332.220 110.430 332.880 110.490 ;
        RECT 332.220 110.170 332.480 110.430 ;
        RECT 333.140 110.170 333.400 110.490 ;
        RECT 333.200 96.550 333.340 110.170 ;
        RECT 333.140 96.230 333.400 96.550 ;
        RECT 333.140 48.290 333.400 48.610 ;
        RECT 333.200 19.710 333.340 48.290 ;
        RECT 91.640 19.390 91.900 19.710 ;
        RECT 333.140 19.390 333.400 19.710 ;
        RECT 91.700 2.400 91.840 19.390 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 331.750 1207.200 332.030 1207.480 ;
        RECT 332.670 1207.200 332.950 1207.480 ;
        RECT 331.750 1110.640 332.030 1110.920 ;
        RECT 332.670 1110.640 332.950 1110.920 ;
        RECT 331.750 1014.080 332.030 1014.360 ;
        RECT 332.670 1014.080 332.950 1014.360 ;
        RECT 331.750 917.520 332.030 917.800 ;
        RECT 332.670 917.520 332.950 917.800 ;
        RECT 331.750 772.680 332.030 772.960 ;
        RECT 333.130 772.680 333.410 772.960 ;
        RECT 331.750 676.120 332.030 676.400 ;
        RECT 333.130 676.120 333.410 676.400 ;
        RECT 331.750 579.560 332.030 579.840 ;
        RECT 333.130 579.560 333.410 579.840 ;
        RECT 331.750 483.000 332.030 483.280 ;
        RECT 333.130 483.000 333.410 483.280 ;
      LAYER met3 ;
        RECT 331.725 1207.490 332.055 1207.505 ;
        RECT 332.645 1207.490 332.975 1207.505 ;
        RECT 331.725 1207.190 332.975 1207.490 ;
        RECT 331.725 1207.175 332.055 1207.190 ;
        RECT 332.645 1207.175 332.975 1207.190 ;
        RECT 331.725 1110.930 332.055 1110.945 ;
        RECT 332.645 1110.930 332.975 1110.945 ;
        RECT 331.725 1110.630 332.975 1110.930 ;
        RECT 331.725 1110.615 332.055 1110.630 ;
        RECT 332.645 1110.615 332.975 1110.630 ;
        RECT 331.725 1014.370 332.055 1014.385 ;
        RECT 332.645 1014.370 332.975 1014.385 ;
        RECT 331.725 1014.070 332.975 1014.370 ;
        RECT 331.725 1014.055 332.055 1014.070 ;
        RECT 332.645 1014.055 332.975 1014.070 ;
        RECT 331.725 917.810 332.055 917.825 ;
        RECT 332.645 917.810 332.975 917.825 ;
        RECT 331.725 917.510 332.975 917.810 ;
        RECT 331.725 917.495 332.055 917.510 ;
        RECT 332.645 917.495 332.975 917.510 ;
        RECT 331.725 772.970 332.055 772.985 ;
        RECT 333.105 772.970 333.435 772.985 ;
        RECT 331.725 772.670 333.435 772.970 ;
        RECT 331.725 772.655 332.055 772.670 ;
        RECT 333.105 772.655 333.435 772.670 ;
        RECT 331.725 676.410 332.055 676.425 ;
        RECT 333.105 676.410 333.435 676.425 ;
        RECT 331.725 676.110 333.435 676.410 ;
        RECT 331.725 676.095 332.055 676.110 ;
        RECT 333.105 676.095 333.435 676.110 ;
        RECT 331.725 579.850 332.055 579.865 ;
        RECT 333.105 579.850 333.435 579.865 ;
        RECT 331.725 579.550 333.435 579.850 ;
        RECT 331.725 579.535 332.055 579.550 ;
        RECT 333.105 579.535 333.435 579.550 ;
        RECT 331.725 483.290 332.055 483.305 ;
        RECT 333.105 483.290 333.435 483.305 ;
        RECT 331.725 482.990 333.435 483.290 ;
        RECT 331.725 482.975 332.055 482.990 ;
        RECT 333.105 482.975 333.435 482.990 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 530.450 19.960 530.770 20.020 ;
        RECT 603.130 19.960 603.450 20.020 ;
        RECT 530.450 19.820 603.450 19.960 ;
        RECT 530.450 19.760 530.770 19.820 ;
        RECT 603.130 19.760 603.450 19.820 ;
      LAYER via ;
        RECT 530.480 19.760 530.740 20.020 ;
        RECT 603.160 19.760 603.420 20.020 ;
      LAYER met2 ;
        RECT 527.260 1600.450 527.540 1604.000 ;
        RECT 527.260 1600.310 529.300 1600.450 ;
        RECT 527.260 1600.000 527.540 1600.310 ;
        RECT 529.160 1582.770 529.300 1600.310 ;
        RECT 529.160 1582.630 530.680 1582.770 ;
        RECT 530.540 20.050 530.680 1582.630 ;
        RECT 530.480 19.730 530.740 20.050 ;
        RECT 603.160 19.730 603.420 20.050 ;
        RECT 603.220 2.400 603.360 19.730 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 534.130 1588.720 534.450 1588.780 ;
        RECT 537.350 1588.720 537.670 1588.780 ;
        RECT 534.130 1588.580 537.670 1588.720 ;
        RECT 534.130 1588.520 534.450 1588.580 ;
        RECT 537.350 1588.520 537.670 1588.580 ;
        RECT 621.070 19.620 621.390 19.680 ;
        RECT 609.660 19.480 621.390 19.620 ;
        RECT 537.350 18.940 537.670 19.000 ;
        RECT 609.660 18.940 609.800 19.480 ;
        RECT 621.070 19.420 621.390 19.480 ;
        RECT 537.350 18.800 609.800 18.940 ;
        RECT 537.350 18.740 537.670 18.800 ;
      LAYER via ;
        RECT 534.160 1588.520 534.420 1588.780 ;
        RECT 537.380 1588.520 537.640 1588.780 ;
        RECT 537.380 18.740 537.640 19.000 ;
        RECT 621.100 19.420 621.360 19.680 ;
      LAYER met2 ;
        RECT 534.160 1600.000 534.440 1604.000 ;
        RECT 534.220 1588.810 534.360 1600.000 ;
        RECT 534.160 1588.490 534.420 1588.810 ;
        RECT 537.380 1588.490 537.640 1588.810 ;
        RECT 537.440 19.030 537.580 1588.490 ;
        RECT 621.100 19.390 621.360 19.710 ;
        RECT 537.380 18.710 537.640 19.030 ;
        RECT 621.160 2.400 621.300 19.390 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 116.910 1592.800 117.230 1592.860 ;
        RECT 116.910 1592.660 304.360 1592.800 ;
        RECT 116.910 1592.600 117.230 1592.660 ;
        RECT 304.220 1592.460 304.360 1592.660 ;
        RECT 343.230 1592.460 343.550 1592.520 ;
        RECT 304.220 1592.320 343.550 1592.460 ;
        RECT 343.230 1592.260 343.550 1592.320 ;
        RECT 115.530 2.960 115.850 3.020 ;
        RECT 116.910 2.960 117.230 3.020 ;
        RECT 115.530 2.820 117.230 2.960 ;
        RECT 115.530 2.760 115.850 2.820 ;
        RECT 116.910 2.760 117.230 2.820 ;
      LAYER via ;
        RECT 116.940 1592.600 117.200 1592.860 ;
        RECT 343.260 1592.260 343.520 1592.520 ;
        RECT 115.560 2.760 115.820 3.020 ;
        RECT 116.940 2.760 117.200 3.020 ;
      LAYER met2 ;
        RECT 343.260 1600.000 343.540 1604.000 ;
        RECT 116.940 1592.570 117.200 1592.890 ;
        RECT 117.000 3.050 117.140 1592.570 ;
        RECT 343.320 1592.550 343.460 1600.000 ;
        RECT 343.260 1592.230 343.520 1592.550 ;
        RECT 115.560 2.730 115.820 3.050 ;
        RECT 116.940 2.730 117.200 3.050 ;
        RECT 115.620 2.400 115.760 2.730 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 151.945 16.745 152.115 20.315 ;
        RECT 179.545 15.385 179.715 20.315 ;
        RECT 227.385 15.385 227.555 20.315 ;
        RECT 276.145 20.145 276.315 20.995 ;
        RECT 333.185 20.485 333.355 21.335 ;
      LAYER mcon ;
        RECT 333.185 21.165 333.355 21.335 ;
        RECT 276.145 20.825 276.315 20.995 ;
        RECT 151.945 20.145 152.115 20.315 ;
        RECT 179.545 20.145 179.715 20.315 ;
        RECT 227.385 20.145 227.555 20.315 ;
      LAYER met1 ;
        RECT 333.125 21.320 333.415 21.365 ;
        RECT 352.890 21.320 353.210 21.380 ;
        RECT 333.125 21.180 353.210 21.320 ;
        RECT 333.125 21.135 333.415 21.180 ;
        RECT 352.890 21.120 353.210 21.180 ;
        RECT 276.085 20.980 276.375 21.025 ;
        RECT 276.085 20.840 304.360 20.980 ;
        RECT 276.085 20.795 276.375 20.840 ;
        RECT 304.220 20.640 304.360 20.840 ;
        RECT 333.125 20.640 333.415 20.685 ;
        RECT 304.220 20.500 333.415 20.640 ;
        RECT 333.125 20.455 333.415 20.500 ;
        RECT 151.885 20.300 152.175 20.345 ;
        RECT 179.485 20.300 179.775 20.345 ;
        RECT 151.885 20.160 179.775 20.300 ;
        RECT 151.885 20.115 152.175 20.160 ;
        RECT 179.485 20.115 179.775 20.160 ;
        RECT 227.325 20.300 227.615 20.345 ;
        RECT 276.085 20.300 276.375 20.345 ;
        RECT 227.325 20.160 276.375 20.300 ;
        RECT 227.325 20.115 227.615 20.160 ;
        RECT 276.085 20.115 276.375 20.160 ;
        RECT 139.450 16.900 139.770 16.960 ;
        RECT 151.885 16.900 152.175 16.945 ;
        RECT 139.450 16.760 152.175 16.900 ;
        RECT 139.450 16.700 139.770 16.760 ;
        RECT 151.885 16.715 152.175 16.760 ;
        RECT 179.485 15.540 179.775 15.585 ;
        RECT 227.325 15.540 227.615 15.585 ;
        RECT 179.485 15.400 227.615 15.540 ;
        RECT 179.485 15.355 179.775 15.400 ;
        RECT 227.325 15.355 227.615 15.400 ;
      LAYER via ;
        RECT 352.920 21.120 353.180 21.380 ;
        RECT 139.480 16.700 139.740 16.960 ;
      LAYER met2 ;
        RECT 352.460 1600.450 352.740 1604.000 ;
        RECT 352.460 1600.310 353.120 1600.450 ;
        RECT 352.460 1600.000 352.740 1600.310 ;
        RECT 352.980 21.410 353.120 1600.310 ;
        RECT 352.920 21.090 353.180 21.410 ;
        RECT 139.480 16.670 139.740 16.990 ;
        RECT 139.540 2.400 139.680 16.670 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 1593.480 158.630 1593.540 ;
        RECT 358.870 1593.480 359.190 1593.540 ;
        RECT 158.310 1593.340 359.190 1593.480 ;
        RECT 158.310 1593.280 158.630 1593.340 ;
        RECT 358.870 1593.280 359.190 1593.340 ;
      LAYER via ;
        RECT 158.340 1593.280 158.600 1593.540 ;
        RECT 358.900 1593.280 359.160 1593.540 ;
      LAYER met2 ;
        RECT 358.900 1600.000 359.180 1604.000 ;
        RECT 358.960 1593.570 359.100 1600.000 ;
        RECT 158.340 1593.250 158.600 1593.570 ;
        RECT 358.900 1593.250 359.160 1593.570 ;
        RECT 158.400 17.410 158.540 1593.250 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.800 1600.450 366.080 1604.000 ;
        RECT 365.800 1600.310 366.460 1600.450 ;
        RECT 365.800 1600.000 366.080 1600.310 ;
        RECT 366.320 18.885 366.460 1600.310 ;
        RECT 174.890 18.515 175.170 18.885 ;
        RECT 366.250 18.515 366.530 18.885 ;
        RECT 174.960 2.400 175.100 18.515 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 174.890 18.560 175.170 18.840 ;
        RECT 366.250 18.560 366.530 18.840 ;
      LAYER met3 ;
        RECT 174.865 18.850 175.195 18.865 ;
        RECT 366.225 18.850 366.555 18.865 ;
        RECT 174.865 18.550 366.555 18.850 ;
        RECT 174.865 18.535 175.195 18.550 ;
        RECT 366.225 18.535 366.555 18.550 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.350 1590.080 192.670 1590.140 ;
        RECT 372.670 1590.080 372.990 1590.140 ;
        RECT 192.350 1589.940 372.990 1590.080 ;
        RECT 192.350 1589.880 192.670 1589.940 ;
        RECT 372.670 1589.880 372.990 1589.940 ;
      LAYER via ;
        RECT 192.380 1589.880 192.640 1590.140 ;
        RECT 372.700 1589.880 372.960 1590.140 ;
      LAYER met2 ;
        RECT 372.700 1600.000 372.980 1604.000 ;
        RECT 372.760 1590.170 372.900 1600.000 ;
        RECT 192.380 1589.850 192.640 1590.170 ;
        RECT 372.700 1589.850 372.960 1590.170 ;
        RECT 192.440 17.410 192.580 1589.850 ;
        RECT 192.440 17.270 193.040 17.410 ;
        RECT 192.900 2.400 193.040 17.270 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 375.045 1497.445 375.215 1511.895 ;
        RECT 374.585 1449.165 374.755 1496.935 ;
        RECT 374.585 1400.885 374.755 1448.655 ;
        RECT 375.045 1256.045 375.215 1304.155 ;
        RECT 375.045 669.545 375.215 717.655 ;
        RECT 375.045 586.245 375.215 613.955 ;
        RECT 375.045 421.345 375.215 469.115 ;
        RECT 375.045 372.725 375.215 420.835 ;
        RECT 374.125 331.245 374.295 355.555 ;
        RECT 374.125 276.165 374.295 324.275 ;
        RECT 375.045 186.065 375.215 227.715 ;
        RECT 374.585 48.365 374.755 137.955 ;
        RECT 328.585 16.575 328.755 16.915 ;
        RECT 327.665 16.405 328.755 16.575 ;
        RECT 352.965 16.065 353.135 16.915 ;
      LAYER mcon ;
        RECT 375.045 1511.725 375.215 1511.895 ;
        RECT 374.585 1496.765 374.755 1496.935 ;
        RECT 374.585 1448.485 374.755 1448.655 ;
        RECT 375.045 1303.985 375.215 1304.155 ;
        RECT 375.045 717.485 375.215 717.655 ;
        RECT 375.045 613.785 375.215 613.955 ;
        RECT 375.045 468.945 375.215 469.115 ;
        RECT 375.045 420.665 375.215 420.835 ;
        RECT 374.125 355.385 374.295 355.555 ;
        RECT 374.125 324.105 374.295 324.275 ;
        RECT 375.045 227.545 375.215 227.715 ;
        RECT 374.585 137.785 374.755 137.955 ;
        RECT 328.585 16.745 328.755 16.915 ;
        RECT 352.965 16.745 353.135 16.915 ;
      LAYER met1 ;
        RECT 374.970 1579.540 375.290 1579.600 ;
        RECT 377.270 1579.540 377.590 1579.600 ;
        RECT 374.970 1579.400 377.590 1579.540 ;
        RECT 374.970 1579.340 375.290 1579.400 ;
        RECT 377.270 1579.340 377.590 1579.400 ;
        RECT 374.970 1511.880 375.290 1511.940 ;
        RECT 374.775 1511.740 375.290 1511.880 ;
        RECT 374.970 1511.680 375.290 1511.740 ;
        RECT 374.970 1497.600 375.290 1497.660 ;
        RECT 374.775 1497.460 375.290 1497.600 ;
        RECT 374.970 1497.400 375.290 1497.460 ;
        RECT 374.525 1496.920 374.815 1496.965 ;
        RECT 374.970 1496.920 375.290 1496.980 ;
        RECT 374.525 1496.780 375.290 1496.920 ;
        RECT 374.525 1496.735 374.815 1496.780 ;
        RECT 374.970 1496.720 375.290 1496.780 ;
        RECT 374.510 1449.320 374.830 1449.380 ;
        RECT 374.315 1449.180 374.830 1449.320 ;
        RECT 374.510 1449.120 374.830 1449.180 ;
        RECT 374.510 1448.640 374.830 1448.700 ;
        RECT 374.315 1448.500 374.830 1448.640 ;
        RECT 374.510 1448.440 374.830 1448.500 ;
        RECT 374.525 1401.040 374.815 1401.085 ;
        RECT 374.970 1401.040 375.290 1401.100 ;
        RECT 374.525 1400.900 375.290 1401.040 ;
        RECT 374.525 1400.855 374.815 1400.900 ;
        RECT 374.970 1400.840 375.290 1400.900 ;
        RECT 374.970 1304.140 375.290 1304.200 ;
        RECT 374.775 1304.000 375.290 1304.140 ;
        RECT 374.970 1303.940 375.290 1304.000 ;
        RECT 374.970 1256.200 375.290 1256.260 ;
        RECT 374.775 1256.060 375.290 1256.200 ;
        RECT 374.970 1256.000 375.290 1256.060 ;
        RECT 374.050 1159.300 374.370 1159.360 ;
        RECT 374.970 1159.300 375.290 1159.360 ;
        RECT 374.050 1159.160 375.290 1159.300 ;
        RECT 374.050 1159.100 374.370 1159.160 ;
        RECT 374.970 1159.100 375.290 1159.160 ;
        RECT 374.050 1062.740 374.370 1062.800 ;
        RECT 374.970 1062.740 375.290 1062.800 ;
        RECT 374.050 1062.600 375.290 1062.740 ;
        RECT 374.050 1062.540 374.370 1062.600 ;
        RECT 374.970 1062.540 375.290 1062.600 ;
        RECT 374.050 966.180 374.370 966.240 ;
        RECT 374.970 966.180 375.290 966.240 ;
        RECT 374.050 966.040 375.290 966.180 ;
        RECT 374.050 965.980 374.370 966.040 ;
        RECT 374.970 965.980 375.290 966.040 ;
        RECT 374.050 869.620 374.370 869.680 ;
        RECT 374.970 869.620 375.290 869.680 ;
        RECT 374.050 869.480 375.290 869.620 ;
        RECT 374.050 869.420 374.370 869.480 ;
        RECT 374.970 869.420 375.290 869.480 ;
        RECT 374.970 717.640 375.290 717.700 ;
        RECT 374.775 717.500 375.290 717.640 ;
        RECT 374.970 717.440 375.290 717.500 ;
        RECT 374.970 669.700 375.290 669.760 ;
        RECT 374.775 669.560 375.290 669.700 ;
        RECT 374.970 669.500 375.290 669.560 ;
        RECT 374.970 613.940 375.290 614.000 ;
        RECT 374.775 613.800 375.290 613.940 ;
        RECT 374.970 613.740 375.290 613.800 ;
        RECT 374.970 586.400 375.290 586.460 ;
        RECT 374.775 586.260 375.290 586.400 ;
        RECT 374.970 586.200 375.290 586.260 ;
        RECT 374.970 469.100 375.290 469.160 ;
        RECT 374.775 468.960 375.290 469.100 ;
        RECT 374.970 468.900 375.290 468.960 ;
        RECT 374.970 421.500 375.290 421.560 ;
        RECT 374.775 421.360 375.290 421.500 ;
        RECT 374.970 421.300 375.290 421.360 ;
        RECT 374.970 420.820 375.290 420.880 ;
        RECT 374.775 420.680 375.290 420.820 ;
        RECT 374.970 420.620 375.290 420.680 ;
        RECT 374.970 372.880 375.290 372.940 ;
        RECT 374.970 372.740 375.485 372.880 ;
        RECT 374.970 372.680 375.290 372.740 ;
        RECT 374.065 355.540 374.355 355.585 ;
        RECT 374.970 355.540 375.290 355.600 ;
        RECT 374.065 355.400 375.290 355.540 ;
        RECT 374.065 355.355 374.355 355.400 ;
        RECT 374.970 355.340 375.290 355.400 ;
        RECT 374.050 331.400 374.370 331.460 ;
        RECT 373.855 331.260 374.370 331.400 ;
        RECT 374.050 331.200 374.370 331.260 ;
        RECT 374.050 324.260 374.370 324.320 ;
        RECT 373.855 324.120 374.370 324.260 ;
        RECT 374.050 324.060 374.370 324.120 ;
        RECT 374.065 276.320 374.355 276.365 ;
        RECT 374.510 276.320 374.830 276.380 ;
        RECT 374.065 276.180 374.830 276.320 ;
        RECT 374.065 276.135 374.355 276.180 ;
        RECT 374.510 276.120 374.830 276.180 ;
        RECT 374.510 234.500 374.830 234.560 ;
        RECT 375.430 234.500 375.750 234.560 ;
        RECT 374.510 234.360 375.750 234.500 ;
        RECT 374.510 234.300 374.830 234.360 ;
        RECT 375.430 234.300 375.750 234.360 ;
        RECT 374.985 227.700 375.275 227.745 ;
        RECT 375.430 227.700 375.750 227.760 ;
        RECT 374.985 227.560 375.750 227.700 ;
        RECT 374.985 227.515 375.275 227.560 ;
        RECT 375.430 227.500 375.750 227.560 ;
        RECT 374.985 186.220 375.275 186.265 ;
        RECT 375.430 186.220 375.750 186.280 ;
        RECT 374.985 186.080 375.750 186.220 ;
        RECT 374.985 186.035 375.275 186.080 ;
        RECT 375.430 186.020 375.750 186.080 ;
        RECT 374.050 148.820 374.370 148.880 ;
        RECT 375.430 148.820 375.750 148.880 ;
        RECT 374.050 148.680 375.750 148.820 ;
        RECT 374.050 148.620 374.370 148.680 ;
        RECT 375.430 148.620 375.750 148.680 ;
        RECT 374.050 137.940 374.370 138.000 ;
        RECT 374.525 137.940 374.815 137.985 ;
        RECT 374.050 137.800 374.815 137.940 ;
        RECT 374.050 137.740 374.370 137.800 ;
        RECT 374.525 137.755 374.815 137.800 ;
        RECT 374.510 48.520 374.830 48.580 ;
        RECT 374.315 48.380 374.830 48.520 ;
        RECT 374.510 48.320 374.830 48.380 ;
        RECT 328.525 16.900 328.815 16.945 ;
        RECT 352.905 16.900 353.195 16.945 ;
        RECT 328.525 16.760 353.195 16.900 ;
        RECT 328.525 16.715 328.815 16.760 ;
        RECT 352.905 16.715 353.195 16.760 ;
        RECT 327.605 16.560 327.895 16.605 ;
        RECT 269.260 16.420 327.895 16.560 ;
        RECT 210.750 16.220 211.070 16.280 ;
        RECT 269.260 16.220 269.400 16.420 ;
        RECT 327.605 16.375 327.895 16.420 ;
        RECT 210.750 16.080 269.400 16.220 ;
        RECT 352.905 16.220 353.195 16.265 ;
        RECT 374.510 16.220 374.830 16.280 ;
        RECT 352.905 16.080 374.830 16.220 ;
        RECT 210.750 16.020 211.070 16.080 ;
        RECT 352.905 16.035 353.195 16.080 ;
        RECT 374.510 16.020 374.830 16.080 ;
      LAYER via ;
        RECT 375.000 1579.340 375.260 1579.600 ;
        RECT 377.300 1579.340 377.560 1579.600 ;
        RECT 375.000 1511.680 375.260 1511.940 ;
        RECT 375.000 1497.400 375.260 1497.660 ;
        RECT 375.000 1496.720 375.260 1496.980 ;
        RECT 374.540 1449.120 374.800 1449.380 ;
        RECT 374.540 1448.440 374.800 1448.700 ;
        RECT 375.000 1400.840 375.260 1401.100 ;
        RECT 375.000 1303.940 375.260 1304.200 ;
        RECT 375.000 1256.000 375.260 1256.260 ;
        RECT 374.080 1159.100 374.340 1159.360 ;
        RECT 375.000 1159.100 375.260 1159.360 ;
        RECT 374.080 1062.540 374.340 1062.800 ;
        RECT 375.000 1062.540 375.260 1062.800 ;
        RECT 374.080 965.980 374.340 966.240 ;
        RECT 375.000 965.980 375.260 966.240 ;
        RECT 374.080 869.420 374.340 869.680 ;
        RECT 375.000 869.420 375.260 869.680 ;
        RECT 375.000 717.440 375.260 717.700 ;
        RECT 375.000 669.500 375.260 669.760 ;
        RECT 375.000 613.740 375.260 614.000 ;
        RECT 375.000 586.200 375.260 586.460 ;
        RECT 375.000 468.900 375.260 469.160 ;
        RECT 375.000 421.300 375.260 421.560 ;
        RECT 375.000 420.620 375.260 420.880 ;
        RECT 375.000 372.680 375.260 372.940 ;
        RECT 375.000 355.340 375.260 355.600 ;
        RECT 374.080 331.200 374.340 331.460 ;
        RECT 374.080 324.060 374.340 324.320 ;
        RECT 374.540 276.120 374.800 276.380 ;
        RECT 374.540 234.300 374.800 234.560 ;
        RECT 375.460 234.300 375.720 234.560 ;
        RECT 375.460 227.500 375.720 227.760 ;
        RECT 375.460 186.020 375.720 186.280 ;
        RECT 374.080 148.620 374.340 148.880 ;
        RECT 375.460 148.620 375.720 148.880 ;
        RECT 374.080 137.740 374.340 138.000 ;
        RECT 374.540 48.320 374.800 48.580 ;
        RECT 210.780 16.020 211.040 16.280 ;
        RECT 374.540 16.020 374.800 16.280 ;
      LAYER met2 ;
        RECT 379.140 1600.450 379.420 1604.000 ;
        RECT 377.360 1600.310 379.420 1600.450 ;
        RECT 377.360 1579.630 377.500 1600.310 ;
        RECT 379.140 1600.000 379.420 1600.310 ;
        RECT 375.000 1579.310 375.260 1579.630 ;
        RECT 377.300 1579.310 377.560 1579.630 ;
        RECT 375.060 1511.970 375.200 1579.310 ;
        RECT 375.000 1511.650 375.260 1511.970 ;
        RECT 375.000 1497.370 375.260 1497.690 ;
        RECT 375.060 1497.010 375.200 1497.370 ;
        RECT 375.000 1496.690 375.260 1497.010 ;
        RECT 374.540 1449.090 374.800 1449.410 ;
        RECT 374.600 1448.730 374.740 1449.090 ;
        RECT 374.540 1448.410 374.800 1448.730 ;
        RECT 375.000 1400.810 375.260 1401.130 ;
        RECT 375.060 1400.530 375.200 1400.810 ;
        RECT 375.060 1400.390 375.660 1400.530 ;
        RECT 375.520 1352.760 375.660 1400.390 ;
        RECT 375.060 1352.620 375.660 1352.760 ;
        RECT 375.060 1304.230 375.200 1352.620 ;
        RECT 375.000 1303.910 375.260 1304.230 ;
        RECT 375.000 1255.970 375.260 1256.290 ;
        RECT 375.060 1207.525 375.200 1255.970 ;
        RECT 374.070 1207.155 374.350 1207.525 ;
        RECT 374.990 1207.155 375.270 1207.525 ;
        RECT 374.140 1159.390 374.280 1207.155 ;
        RECT 374.080 1159.070 374.340 1159.390 ;
        RECT 375.000 1159.070 375.260 1159.390 ;
        RECT 375.060 1110.965 375.200 1159.070 ;
        RECT 374.070 1110.595 374.350 1110.965 ;
        RECT 374.990 1110.595 375.270 1110.965 ;
        RECT 374.140 1062.830 374.280 1110.595 ;
        RECT 374.080 1062.510 374.340 1062.830 ;
        RECT 375.000 1062.510 375.260 1062.830 ;
        RECT 375.060 1014.405 375.200 1062.510 ;
        RECT 374.070 1014.035 374.350 1014.405 ;
        RECT 374.990 1014.035 375.270 1014.405 ;
        RECT 374.140 966.270 374.280 1014.035 ;
        RECT 374.080 965.950 374.340 966.270 ;
        RECT 375.000 965.950 375.260 966.270 ;
        RECT 375.060 917.845 375.200 965.950 ;
        RECT 374.070 917.475 374.350 917.845 ;
        RECT 374.990 917.475 375.270 917.845 ;
        RECT 374.140 869.710 374.280 917.475 ;
        RECT 374.080 869.390 374.340 869.710 ;
        RECT 375.000 869.390 375.260 869.710 ;
        RECT 375.060 787.170 375.200 869.390 ;
        RECT 374.600 787.030 375.200 787.170 ;
        RECT 374.600 786.490 374.740 787.030 ;
        RECT 374.600 786.350 375.200 786.490 ;
        RECT 375.060 725.405 375.200 786.350 ;
        RECT 374.990 725.035 375.270 725.405 ;
        RECT 374.990 724.355 375.270 724.725 ;
        RECT 375.060 717.730 375.200 724.355 ;
        RECT 375.000 717.410 375.260 717.730 ;
        RECT 375.000 669.470 375.260 669.790 ;
        RECT 375.060 628.845 375.200 669.470 ;
        RECT 374.990 628.475 375.270 628.845 ;
        RECT 374.990 627.795 375.270 628.165 ;
        RECT 375.060 614.030 375.200 627.795 ;
        RECT 375.000 613.710 375.260 614.030 ;
        RECT 375.000 586.170 375.260 586.490 ;
        RECT 375.060 477.090 375.200 586.170 ;
        RECT 374.600 476.950 375.200 477.090 ;
        RECT 374.600 469.610 374.740 476.950 ;
        RECT 374.600 469.470 375.200 469.610 ;
        RECT 375.060 469.190 375.200 469.470 ;
        RECT 375.000 468.870 375.260 469.190 ;
        RECT 375.000 421.270 375.260 421.590 ;
        RECT 375.060 420.910 375.200 421.270 ;
        RECT 375.000 420.590 375.260 420.910 ;
        RECT 375.000 372.650 375.260 372.970 ;
        RECT 375.060 355.630 375.200 372.650 ;
        RECT 375.000 355.310 375.260 355.630 ;
        RECT 374.080 331.170 374.340 331.490 ;
        RECT 374.140 324.350 374.280 331.170 ;
        RECT 374.080 324.030 374.340 324.350 ;
        RECT 374.540 276.090 374.800 276.410 ;
        RECT 374.600 234.590 374.740 276.090 ;
        RECT 374.540 234.270 374.800 234.590 ;
        RECT 375.460 234.270 375.720 234.590 ;
        RECT 375.520 227.790 375.660 234.270 ;
        RECT 375.460 227.470 375.720 227.790 ;
        RECT 375.460 185.990 375.720 186.310 ;
        RECT 375.520 148.910 375.660 185.990 ;
        RECT 374.080 148.590 374.340 148.910 ;
        RECT 375.460 148.590 375.720 148.910 ;
        RECT 374.140 138.030 374.280 148.590 ;
        RECT 374.080 137.710 374.340 138.030 ;
        RECT 374.540 48.290 374.800 48.610 ;
        RECT 374.600 16.310 374.740 48.290 ;
        RECT 210.780 15.990 211.040 16.310 ;
        RECT 374.540 15.990 374.800 16.310 ;
        RECT 210.840 2.400 210.980 15.990 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 374.070 1207.200 374.350 1207.480 ;
        RECT 374.990 1207.200 375.270 1207.480 ;
        RECT 374.070 1110.640 374.350 1110.920 ;
        RECT 374.990 1110.640 375.270 1110.920 ;
        RECT 374.070 1014.080 374.350 1014.360 ;
        RECT 374.990 1014.080 375.270 1014.360 ;
        RECT 374.070 917.520 374.350 917.800 ;
        RECT 374.990 917.520 375.270 917.800 ;
        RECT 374.990 725.080 375.270 725.360 ;
        RECT 374.990 724.400 375.270 724.680 ;
        RECT 374.990 628.520 375.270 628.800 ;
        RECT 374.990 627.840 375.270 628.120 ;
      LAYER met3 ;
        RECT 374.045 1207.490 374.375 1207.505 ;
        RECT 374.965 1207.490 375.295 1207.505 ;
        RECT 374.045 1207.190 375.295 1207.490 ;
        RECT 374.045 1207.175 374.375 1207.190 ;
        RECT 374.965 1207.175 375.295 1207.190 ;
        RECT 374.045 1110.930 374.375 1110.945 ;
        RECT 374.965 1110.930 375.295 1110.945 ;
        RECT 374.045 1110.630 375.295 1110.930 ;
        RECT 374.045 1110.615 374.375 1110.630 ;
        RECT 374.965 1110.615 375.295 1110.630 ;
        RECT 374.045 1014.370 374.375 1014.385 ;
        RECT 374.965 1014.370 375.295 1014.385 ;
        RECT 374.045 1014.070 375.295 1014.370 ;
        RECT 374.045 1014.055 374.375 1014.070 ;
        RECT 374.965 1014.055 375.295 1014.070 ;
        RECT 374.045 917.810 374.375 917.825 ;
        RECT 374.965 917.810 375.295 917.825 ;
        RECT 374.045 917.510 375.295 917.810 ;
        RECT 374.045 917.495 374.375 917.510 ;
        RECT 374.965 917.495 375.295 917.510 ;
        RECT 374.965 725.370 375.295 725.385 ;
        RECT 374.965 725.070 375.970 725.370 ;
        RECT 374.965 725.055 375.295 725.070 ;
        RECT 374.965 724.690 375.295 724.705 ;
        RECT 375.670 724.690 375.970 725.070 ;
        RECT 374.965 724.390 375.970 724.690 ;
        RECT 374.965 724.375 375.295 724.390 ;
        RECT 374.965 628.810 375.295 628.825 ;
        RECT 374.965 628.510 375.970 628.810 ;
        RECT 374.965 628.495 375.295 628.510 ;
        RECT 374.965 628.130 375.295 628.145 ;
        RECT 375.670 628.130 375.970 628.510 ;
        RECT 374.965 627.830 375.970 628.130 ;
        RECT 374.965 627.815 375.295 627.830 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 234.210 1588.040 234.530 1588.100 ;
        RECT 386.010 1588.040 386.330 1588.100 ;
        RECT 234.210 1587.900 386.330 1588.040 ;
        RECT 234.210 1587.840 234.530 1587.900 ;
        RECT 386.010 1587.840 386.330 1587.900 ;
        RECT 228.690 16.560 229.010 16.620 ;
        RECT 234.210 16.560 234.530 16.620 ;
        RECT 228.690 16.420 234.530 16.560 ;
        RECT 228.690 16.360 229.010 16.420 ;
        RECT 234.210 16.360 234.530 16.420 ;
      LAYER via ;
        RECT 234.240 1587.840 234.500 1588.100 ;
        RECT 386.040 1587.840 386.300 1588.100 ;
        RECT 228.720 16.360 228.980 16.620 ;
        RECT 234.240 16.360 234.500 16.620 ;
      LAYER met2 ;
        RECT 386.040 1600.000 386.320 1604.000 ;
        RECT 386.100 1588.130 386.240 1600.000 ;
        RECT 234.240 1587.810 234.500 1588.130 ;
        RECT 386.040 1587.810 386.300 1588.130 ;
        RECT 234.300 16.650 234.440 1587.810 ;
        RECT 228.720 16.330 228.980 16.650 ;
        RECT 234.240 16.330 234.500 16.650 ;
        RECT 228.780 2.400 228.920 16.330 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 18.600 50.530 18.660 ;
        RECT 317.930 18.600 318.250 18.660 ;
        RECT 50.210 18.460 318.250 18.600 ;
        RECT 50.210 18.400 50.530 18.460 ;
        RECT 317.930 18.400 318.250 18.460 ;
      LAYER via ;
        RECT 50.240 18.400 50.500 18.660 ;
        RECT 317.960 18.400 318.220 18.660 ;
      LAYER met2 ;
        RECT 318.880 1600.450 319.160 1604.000 ;
        RECT 318.020 1600.310 319.160 1600.450 ;
        RECT 318.020 18.690 318.160 1600.310 ;
        RECT 318.880 1600.000 319.160 1600.310 ;
        RECT 50.240 18.370 50.500 18.690 ;
        RECT 317.960 18.370 318.220 18.690 ;
        RECT 50.300 2.400 50.440 18.370 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 1588.380 255.230 1588.440 ;
        RECT 394.750 1588.380 395.070 1588.440 ;
        RECT 254.910 1588.240 395.070 1588.380 ;
        RECT 254.910 1588.180 255.230 1588.240 ;
        RECT 394.750 1588.180 395.070 1588.240 ;
        RECT 252.610 16.560 252.930 16.620 ;
        RECT 254.910 16.560 255.230 16.620 ;
        RECT 252.610 16.420 255.230 16.560 ;
        RECT 252.610 16.360 252.930 16.420 ;
        RECT 254.910 16.360 255.230 16.420 ;
      LAYER via ;
        RECT 254.940 1588.180 255.200 1588.440 ;
        RECT 394.780 1588.180 395.040 1588.440 ;
        RECT 252.640 16.360 252.900 16.620 ;
        RECT 254.940 16.360 255.200 16.620 ;
      LAYER met2 ;
        RECT 394.780 1600.000 395.060 1604.000 ;
        RECT 394.840 1588.470 394.980 1600.000 ;
        RECT 254.940 1588.150 255.200 1588.470 ;
        RECT 394.780 1588.150 395.040 1588.470 ;
        RECT 255.000 16.650 255.140 1588.150 ;
        RECT 252.640 16.330 252.900 16.650 ;
        RECT 254.940 16.330 255.200 16.650 ;
        RECT 252.700 2.400 252.840 16.330 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 14.860 270.410 14.920 ;
        RECT 400.270 14.860 400.590 14.920 ;
        RECT 270.090 14.720 400.590 14.860 ;
        RECT 270.090 14.660 270.410 14.720 ;
        RECT 400.270 14.660 400.590 14.720 ;
      LAYER via ;
        RECT 270.120 14.660 270.380 14.920 ;
        RECT 400.300 14.660 400.560 14.920 ;
      LAYER met2 ;
        RECT 401.680 1600.450 401.960 1604.000 ;
        RECT 400.360 1600.310 401.960 1600.450 ;
        RECT 400.360 14.950 400.500 1600.310 ;
        RECT 401.680 1600.000 401.960 1600.310 ;
        RECT 270.120 14.630 270.380 14.950 ;
        RECT 400.300 14.630 400.560 14.950 ;
        RECT 270.180 2.400 270.320 14.630 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 1587.360 289.730 1587.420 ;
        RECT 408.550 1587.360 408.870 1587.420 ;
        RECT 289.410 1587.220 408.870 1587.360 ;
        RECT 289.410 1587.160 289.730 1587.220 ;
        RECT 408.550 1587.160 408.870 1587.220 ;
      LAYER via ;
        RECT 289.440 1587.160 289.700 1587.420 ;
        RECT 408.580 1587.160 408.840 1587.420 ;
      LAYER met2 ;
        RECT 408.580 1600.000 408.860 1604.000 ;
        RECT 408.640 1587.450 408.780 1600.000 ;
        RECT 289.440 1587.130 289.700 1587.450 ;
        RECT 408.580 1587.130 408.840 1587.450 ;
        RECT 289.500 3.130 289.640 1587.130 ;
        RECT 288.120 2.990 289.640 3.130 ;
        RECT 288.120 2.400 288.260 2.990 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 375.505 14.025 375.675 17.255 ;
      LAYER mcon ;
        RECT 375.505 17.085 375.675 17.255 ;
      LAYER met1 ;
        RECT 305.970 17.240 306.290 17.300 ;
        RECT 375.445 17.240 375.735 17.285 ;
        RECT 305.970 17.100 375.735 17.240 ;
        RECT 305.970 17.040 306.290 17.100 ;
        RECT 375.445 17.055 375.735 17.100 ;
        RECT 375.445 14.180 375.735 14.225 ;
        RECT 415.450 14.180 415.770 14.240 ;
        RECT 375.445 14.040 415.770 14.180 ;
        RECT 375.445 13.995 375.735 14.040 ;
        RECT 415.450 13.980 415.770 14.040 ;
      LAYER via ;
        RECT 306.000 17.040 306.260 17.300 ;
        RECT 415.480 13.980 415.740 14.240 ;
      LAYER met2 ;
        RECT 415.020 1600.450 415.300 1604.000 ;
        RECT 415.020 1600.310 415.680 1600.450 ;
        RECT 415.020 1600.000 415.300 1600.310 ;
        RECT 306.000 17.010 306.260 17.330 ;
        RECT 306.060 2.400 306.200 17.010 ;
        RECT 415.540 14.270 415.680 1600.310 ;
        RECT 415.480 13.950 415.740 14.270 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 17.920 324.230 17.980 ;
        RECT 421.890 17.920 422.210 17.980 ;
        RECT 323.910 17.780 422.210 17.920 ;
        RECT 323.910 17.720 324.230 17.780 ;
        RECT 421.890 17.720 422.210 17.780 ;
      LAYER via ;
        RECT 323.940 17.720 324.200 17.980 ;
        RECT 421.920 17.720 422.180 17.980 ;
      LAYER met2 ;
        RECT 421.920 1600.000 422.200 1604.000 ;
        RECT 421.980 18.010 422.120 1600.000 ;
        RECT 323.940 17.690 324.200 18.010 ;
        RECT 421.920 17.690 422.180 18.010 ;
        RECT 324.000 2.400 324.140 17.690 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 406.785 18.445 406.955 19.635 ;
      LAYER mcon ;
        RECT 406.785 19.465 406.955 19.635 ;
      LAYER met1 ;
        RECT 406.725 19.620 407.015 19.665 ;
        RECT 428.790 19.620 429.110 19.680 ;
        RECT 406.725 19.480 429.110 19.620 ;
        RECT 406.725 19.435 407.015 19.480 ;
        RECT 428.790 19.420 429.110 19.480 ;
        RECT 341.390 18.940 341.710 19.000 ;
        RECT 341.390 18.800 376.120 18.940 ;
        RECT 341.390 18.740 341.710 18.800 ;
        RECT 375.980 18.600 376.120 18.800 ;
        RECT 406.725 18.600 407.015 18.645 ;
        RECT 375.980 18.460 407.015 18.600 ;
        RECT 406.725 18.415 407.015 18.460 ;
      LAYER via ;
        RECT 428.820 19.420 429.080 19.680 ;
        RECT 341.420 18.740 341.680 19.000 ;
      LAYER met2 ;
        RECT 428.820 1600.000 429.100 1604.000 ;
        RECT 428.880 19.710 429.020 1600.000 ;
        RECT 428.820 19.390 429.080 19.710 ;
        RECT 341.420 18.710 341.680 19.030 ;
        RECT 341.480 2.400 341.620 18.710 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 375.890 1591.440 376.210 1591.500 ;
        RECT 435.230 1591.440 435.550 1591.500 ;
        RECT 375.890 1591.300 435.550 1591.440 ;
        RECT 375.890 1591.240 376.210 1591.300 ;
        RECT 435.230 1591.240 435.550 1591.300 ;
        RECT 360.710 20.640 361.030 20.700 ;
        RECT 375.890 20.640 376.210 20.700 ;
        RECT 360.710 20.500 376.210 20.640 ;
        RECT 360.710 20.440 361.030 20.500 ;
        RECT 375.890 20.440 376.210 20.500 ;
      LAYER via ;
        RECT 375.920 1591.240 376.180 1591.500 ;
        RECT 435.260 1591.240 435.520 1591.500 ;
        RECT 360.740 20.440 361.000 20.700 ;
        RECT 375.920 20.440 376.180 20.700 ;
      LAYER met2 ;
        RECT 435.260 1600.000 435.540 1604.000 ;
        RECT 435.320 1591.530 435.460 1600.000 ;
        RECT 375.920 1591.210 376.180 1591.530 ;
        RECT 435.260 1591.210 435.520 1591.530 ;
        RECT 375.980 20.730 376.120 1591.210 ;
        RECT 360.740 20.410 361.000 20.730 ;
        RECT 375.920 20.410 376.180 20.730 ;
        RECT 360.800 9.930 360.940 20.410 ;
        RECT 359.420 9.790 360.940 9.930 ;
        RECT 359.420 2.400 359.560 9.790 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 406.325 16.745 406.495 19.635 ;
      LAYER mcon ;
        RECT 406.325 19.465 406.495 19.635 ;
      LAYER met1 ;
        RECT 431.090 1587.360 431.410 1587.420 ;
        RECT 442.130 1587.360 442.450 1587.420 ;
        RECT 431.090 1587.220 442.450 1587.360 ;
        RECT 431.090 1587.160 431.410 1587.220 ;
        RECT 442.130 1587.160 442.450 1587.220 ;
        RECT 377.270 19.620 377.590 19.680 ;
        RECT 406.265 19.620 406.555 19.665 ;
        RECT 377.270 19.480 406.555 19.620 ;
        RECT 377.270 19.420 377.590 19.480 ;
        RECT 406.265 19.435 406.555 19.480 ;
        RECT 406.265 16.900 406.555 16.945 ;
        RECT 431.090 16.900 431.410 16.960 ;
        RECT 406.265 16.760 431.410 16.900 ;
        RECT 406.265 16.715 406.555 16.760 ;
        RECT 431.090 16.700 431.410 16.760 ;
      LAYER via ;
        RECT 431.120 1587.160 431.380 1587.420 ;
        RECT 442.160 1587.160 442.420 1587.420 ;
        RECT 377.300 19.420 377.560 19.680 ;
        RECT 431.120 16.700 431.380 16.960 ;
      LAYER met2 ;
        RECT 442.160 1600.000 442.440 1604.000 ;
        RECT 442.220 1587.450 442.360 1600.000 ;
        RECT 431.120 1587.130 431.380 1587.450 ;
        RECT 442.160 1587.130 442.420 1587.450 ;
        RECT 377.300 19.390 377.560 19.710 ;
        RECT 377.360 2.400 377.500 19.390 ;
        RECT 431.180 16.990 431.320 1587.130 ;
        RECT 431.120 16.670 431.380 16.990 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 400.345 19.125 400.515 20.315 ;
      LAYER mcon ;
        RECT 400.345 20.145 400.515 20.315 ;
      LAYER met1 ;
        RECT 437.990 1590.420 438.310 1590.480 ;
        RECT 449.030 1590.420 449.350 1590.480 ;
        RECT 437.990 1590.280 449.350 1590.420 ;
        RECT 437.990 1590.220 438.310 1590.280 ;
        RECT 449.030 1590.220 449.350 1590.280 ;
        RECT 395.210 20.300 395.530 20.360 ;
        RECT 400.285 20.300 400.575 20.345 ;
        RECT 395.210 20.160 400.575 20.300 ;
        RECT 395.210 20.100 395.530 20.160 ;
        RECT 400.285 20.115 400.575 20.160 ;
        RECT 400.285 19.280 400.575 19.325 ;
        RECT 437.990 19.280 438.310 19.340 ;
        RECT 400.285 19.140 438.310 19.280 ;
        RECT 400.285 19.095 400.575 19.140 ;
        RECT 437.990 19.080 438.310 19.140 ;
      LAYER via ;
        RECT 438.020 1590.220 438.280 1590.480 ;
        RECT 449.060 1590.220 449.320 1590.480 ;
        RECT 395.240 20.100 395.500 20.360 ;
        RECT 438.020 19.080 438.280 19.340 ;
      LAYER met2 ;
        RECT 449.060 1600.000 449.340 1604.000 ;
        RECT 449.120 1590.510 449.260 1600.000 ;
        RECT 438.020 1590.190 438.280 1590.510 ;
        RECT 449.060 1590.190 449.320 1590.510 ;
        RECT 395.240 20.070 395.500 20.390 ;
        RECT 395.300 2.400 395.440 20.070 ;
        RECT 438.080 19.370 438.220 1590.190 ;
        RECT 438.020 19.050 438.280 19.370 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 434.845 17.085 435.015 24.055 ;
      LAYER mcon ;
        RECT 434.845 23.885 435.015 24.055 ;
      LAYER met1 ;
        RECT 451.790 1587.360 452.110 1587.420 ;
        RECT 455.470 1587.360 455.790 1587.420 ;
        RECT 451.790 1587.220 455.790 1587.360 ;
        RECT 451.790 1587.160 452.110 1587.220 ;
        RECT 455.470 1587.160 455.790 1587.220 ;
        RECT 434.785 24.040 435.075 24.085 ;
        RECT 451.790 24.040 452.110 24.100 ;
        RECT 434.785 23.900 452.110 24.040 ;
        RECT 434.785 23.855 435.075 23.900 ;
        RECT 451.790 23.840 452.110 23.900 ;
        RECT 413.150 17.240 413.470 17.300 ;
        RECT 434.785 17.240 435.075 17.285 ;
        RECT 413.150 17.100 435.075 17.240 ;
        RECT 413.150 17.040 413.470 17.100 ;
        RECT 434.785 17.055 435.075 17.100 ;
      LAYER via ;
        RECT 451.820 1587.160 452.080 1587.420 ;
        RECT 455.500 1587.160 455.760 1587.420 ;
        RECT 451.820 23.840 452.080 24.100 ;
        RECT 413.180 17.040 413.440 17.300 ;
      LAYER met2 ;
        RECT 455.500 1600.000 455.780 1604.000 ;
        RECT 455.560 1587.450 455.700 1600.000 ;
        RECT 451.820 1587.130 452.080 1587.450 ;
        RECT 455.500 1587.130 455.760 1587.450 ;
        RECT 451.880 24.130 452.020 1587.130 ;
        RECT 451.820 23.810 452.080 24.130 ;
        RECT 413.180 17.010 413.440 17.330 ;
        RECT 413.240 2.400 413.380 17.010 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 74.130 18.940 74.450 19.000 ;
        RECT 324.830 18.940 325.150 19.000 ;
        RECT 74.130 18.800 325.150 18.940 ;
        RECT 74.130 18.740 74.450 18.800 ;
        RECT 324.830 18.740 325.150 18.800 ;
      LAYER via ;
        RECT 74.160 18.740 74.420 19.000 ;
        RECT 324.860 18.740 325.120 19.000 ;
      LAYER met2 ;
        RECT 327.620 1600.450 327.900 1604.000 ;
        RECT 326.300 1600.310 327.900 1600.450 ;
        RECT 326.300 1580.050 326.440 1600.310 ;
        RECT 327.620 1600.000 327.900 1600.310 ;
        RECT 324.920 1579.910 326.440 1580.050 ;
        RECT 324.920 19.030 325.060 1579.910 ;
        RECT 74.160 18.710 74.420 19.030 ;
        RECT 324.860 18.710 325.120 19.030 ;
        RECT 74.220 2.400 74.360 18.710 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 430.630 15.200 430.950 15.260 ;
        RECT 463.290 15.200 463.610 15.260 ;
        RECT 430.630 15.060 463.610 15.200 ;
        RECT 430.630 15.000 430.950 15.060 ;
        RECT 463.290 15.000 463.610 15.060 ;
      LAYER via ;
        RECT 430.660 15.000 430.920 15.260 ;
        RECT 463.320 15.000 463.580 15.260 ;
      LAYER met2 ;
        RECT 462.400 1600.450 462.680 1604.000 ;
        RECT 462.400 1600.310 463.520 1600.450 ;
        RECT 462.400 1600.000 462.680 1600.310 ;
        RECT 463.380 15.290 463.520 1600.310 ;
        RECT 430.660 14.970 430.920 15.290 ;
        RECT 463.320 14.970 463.580 15.290 ;
        RECT 430.720 2.400 430.860 14.970 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 462.830 1579.880 463.150 1579.940 ;
        RECT 467.430 1579.880 467.750 1579.940 ;
        RECT 462.830 1579.740 467.750 1579.880 ;
        RECT 462.830 1579.680 463.150 1579.740 ;
        RECT 467.430 1579.680 467.750 1579.740 ;
        RECT 448.570 19.280 448.890 19.340 ;
        RECT 462.830 19.280 463.150 19.340 ;
        RECT 448.570 19.140 463.150 19.280 ;
        RECT 448.570 19.080 448.890 19.140 ;
        RECT 462.830 19.080 463.150 19.140 ;
      LAYER via ;
        RECT 462.860 1579.680 463.120 1579.940 ;
        RECT 467.460 1579.680 467.720 1579.940 ;
        RECT 448.600 19.080 448.860 19.340 ;
        RECT 462.860 19.080 463.120 19.340 ;
      LAYER met2 ;
        RECT 468.840 1600.450 469.120 1604.000 ;
        RECT 467.520 1600.310 469.120 1600.450 ;
        RECT 467.520 1579.970 467.660 1600.310 ;
        RECT 468.840 1600.000 469.120 1600.310 ;
        RECT 462.860 1579.650 463.120 1579.970 ;
        RECT 467.460 1579.650 467.720 1579.970 ;
        RECT 462.920 19.370 463.060 1579.650 ;
        RECT 448.600 19.050 448.860 19.370 ;
        RECT 462.860 19.050 463.120 19.370 ;
        RECT 448.660 2.400 448.800 19.050 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.810 1587.360 469.130 1587.420 ;
        RECT 475.710 1587.360 476.030 1587.420 ;
        RECT 468.810 1587.220 476.030 1587.360 ;
        RECT 468.810 1587.160 469.130 1587.220 ;
        RECT 475.710 1587.160 476.030 1587.220 ;
        RECT 466.510 20.640 466.830 20.700 ;
        RECT 468.810 20.640 469.130 20.700 ;
        RECT 466.510 20.500 469.130 20.640 ;
        RECT 466.510 20.440 466.830 20.500 ;
        RECT 468.810 20.440 469.130 20.500 ;
      LAYER via ;
        RECT 468.840 1587.160 469.100 1587.420 ;
        RECT 475.740 1587.160 476.000 1587.420 ;
        RECT 466.540 20.440 466.800 20.700 ;
        RECT 468.840 20.440 469.100 20.700 ;
      LAYER met2 ;
        RECT 475.740 1600.000 476.020 1604.000 ;
        RECT 475.800 1587.450 475.940 1600.000 ;
        RECT 468.840 1587.130 469.100 1587.450 ;
        RECT 475.740 1587.130 476.000 1587.450 ;
        RECT 468.900 20.730 469.040 1587.130 ;
        RECT 466.540 20.410 466.800 20.730 ;
        RECT 468.840 20.410 469.100 20.730 ;
        RECT 466.600 2.400 466.740 20.410 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 482.610 20.640 482.930 20.700 ;
        RECT 484.450 20.640 484.770 20.700 ;
        RECT 482.610 20.500 484.770 20.640 ;
        RECT 482.610 20.440 482.930 20.500 ;
        RECT 484.450 20.440 484.770 20.500 ;
      LAYER via ;
        RECT 482.640 20.440 482.900 20.700 ;
        RECT 484.480 20.440 484.740 20.700 ;
      LAYER met2 ;
        RECT 482.640 1600.000 482.920 1604.000 ;
        RECT 482.700 20.730 482.840 1600.000 ;
        RECT 482.640 20.410 482.900 20.730 ;
        RECT 484.480 20.410 484.740 20.730 ;
        RECT 484.540 2.400 484.680 20.410 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 489.050 17.240 489.370 17.300 ;
        RECT 502.390 17.240 502.710 17.300 ;
        RECT 489.050 17.100 502.710 17.240 ;
        RECT 489.050 17.040 489.370 17.100 ;
        RECT 502.390 17.040 502.710 17.100 ;
      LAYER via ;
        RECT 489.080 17.040 489.340 17.300 ;
        RECT 502.420 17.040 502.680 17.300 ;
      LAYER met2 ;
        RECT 489.080 1600.000 489.360 1604.000 ;
        RECT 489.140 17.330 489.280 1600.000 ;
        RECT 489.080 17.010 489.340 17.330 ;
        RECT 502.420 17.010 502.680 17.330 ;
        RECT 502.480 2.400 502.620 17.010 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 495.950 1588.720 496.270 1588.780 ;
        RECT 500.090 1588.720 500.410 1588.780 ;
        RECT 495.950 1588.580 500.410 1588.720 ;
        RECT 495.950 1588.520 496.270 1588.580 ;
        RECT 500.090 1588.520 500.410 1588.580 ;
        RECT 500.090 20.640 500.410 20.700 ;
        RECT 519.870 20.640 520.190 20.700 ;
        RECT 500.090 20.500 520.190 20.640 ;
        RECT 500.090 20.440 500.410 20.500 ;
        RECT 519.870 20.440 520.190 20.500 ;
      LAYER via ;
        RECT 495.980 1588.520 496.240 1588.780 ;
        RECT 500.120 1588.520 500.380 1588.780 ;
        RECT 500.120 20.440 500.380 20.700 ;
        RECT 519.900 20.440 520.160 20.700 ;
      LAYER met2 ;
        RECT 495.980 1600.000 496.260 1604.000 ;
        RECT 496.040 1588.810 496.180 1600.000 ;
        RECT 495.980 1588.490 496.240 1588.810 ;
        RECT 500.120 1588.490 500.380 1588.810 ;
        RECT 500.180 20.730 500.320 1588.490 ;
        RECT 500.120 20.410 500.380 20.730 ;
        RECT 519.900 20.410 520.160 20.730 ;
        RECT 519.960 2.400 520.100 20.410 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 502.850 1588.380 503.170 1588.440 ;
        RECT 520.790 1588.380 521.110 1588.440 ;
        RECT 502.850 1588.240 521.110 1588.380 ;
        RECT 502.850 1588.180 503.170 1588.240 ;
        RECT 520.790 1588.180 521.110 1588.240 ;
        RECT 520.790 15.540 521.110 15.600 ;
        RECT 537.810 15.540 538.130 15.600 ;
        RECT 520.790 15.400 538.130 15.540 ;
        RECT 520.790 15.340 521.110 15.400 ;
        RECT 537.810 15.340 538.130 15.400 ;
      LAYER via ;
        RECT 502.880 1588.180 503.140 1588.440 ;
        RECT 520.820 1588.180 521.080 1588.440 ;
        RECT 520.820 15.340 521.080 15.600 ;
        RECT 537.840 15.340 538.100 15.600 ;
      LAYER met2 ;
        RECT 502.880 1600.000 503.160 1604.000 ;
        RECT 502.940 1588.470 503.080 1600.000 ;
        RECT 502.880 1588.150 503.140 1588.470 ;
        RECT 520.820 1588.150 521.080 1588.470 ;
        RECT 520.880 15.630 521.020 1588.150 ;
        RECT 520.820 15.310 521.080 15.630 ;
        RECT 537.840 15.310 538.100 15.630 ;
        RECT 537.900 2.400 538.040 15.310 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 510.210 17.240 510.530 17.300 ;
        RECT 555.750 17.240 556.070 17.300 ;
        RECT 510.210 17.100 556.070 17.240 ;
        RECT 510.210 17.040 510.530 17.100 ;
        RECT 555.750 17.040 556.070 17.100 ;
      LAYER via ;
        RECT 510.240 17.040 510.500 17.300 ;
        RECT 555.780 17.040 556.040 17.300 ;
      LAYER met2 ;
        RECT 509.320 1600.450 509.600 1604.000 ;
        RECT 509.320 1600.310 510.440 1600.450 ;
        RECT 509.320 1600.000 509.600 1600.310 ;
        RECT 510.300 17.330 510.440 1600.310 ;
        RECT 510.240 17.010 510.500 17.330 ;
        RECT 555.780 17.010 556.040 17.330 ;
        RECT 555.840 2.400 555.980 17.010 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 517.110 16.220 517.430 16.280 ;
        RECT 573.690 16.220 574.010 16.280 ;
        RECT 517.110 16.080 574.010 16.220 ;
        RECT 517.110 16.020 517.430 16.080 ;
        RECT 573.690 16.020 574.010 16.080 ;
      LAYER via ;
        RECT 517.140 16.020 517.400 16.280 ;
        RECT 573.720 16.020 573.980 16.280 ;
      LAYER met2 ;
        RECT 516.220 1600.450 516.500 1604.000 ;
        RECT 516.220 1600.310 517.340 1600.450 ;
        RECT 516.220 1600.000 516.500 1600.310 ;
        RECT 517.200 16.310 517.340 1600.310 ;
        RECT 517.140 15.990 517.400 16.310 ;
        RECT 573.720 15.990 573.980 16.310 ;
        RECT 573.780 2.400 573.920 15.990 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 524.010 20.300 524.330 20.360 ;
        RECT 591.170 20.300 591.490 20.360 ;
        RECT 524.010 20.160 591.490 20.300 ;
        RECT 524.010 20.100 524.330 20.160 ;
        RECT 591.170 20.100 591.490 20.160 ;
      LAYER via ;
        RECT 524.040 20.100 524.300 20.360 ;
        RECT 591.200 20.100 591.460 20.360 ;
      LAYER met2 ;
        RECT 523.120 1600.450 523.400 1604.000 ;
        RECT 523.120 1600.310 524.240 1600.450 ;
        RECT 523.120 1600.000 523.400 1600.310 ;
        RECT 524.100 20.390 524.240 1600.310 ;
        RECT 524.040 20.070 524.300 20.390 ;
        RECT 591.200 20.070 591.460 20.390 ;
        RECT 591.260 2.400 591.400 20.070 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 103.110 1591.780 103.430 1591.840 ;
        RECT 336.790 1591.780 337.110 1591.840 ;
        RECT 103.110 1591.640 337.110 1591.780 ;
        RECT 103.110 1591.580 103.430 1591.640 ;
        RECT 336.790 1591.580 337.110 1591.640 ;
        RECT 97.590 16.900 97.910 16.960 ;
        RECT 103.110 16.900 103.430 16.960 ;
        RECT 97.590 16.760 103.430 16.900 ;
        RECT 97.590 16.700 97.910 16.760 ;
        RECT 103.110 16.700 103.430 16.760 ;
      LAYER via ;
        RECT 103.140 1591.580 103.400 1591.840 ;
        RECT 336.820 1591.580 337.080 1591.840 ;
        RECT 97.620 16.700 97.880 16.960 ;
        RECT 103.140 16.700 103.400 16.960 ;
      LAYER met2 ;
        RECT 336.820 1600.000 337.100 1604.000 ;
        RECT 336.880 1591.870 337.020 1600.000 ;
        RECT 103.140 1591.550 103.400 1591.870 ;
        RECT 336.820 1591.550 337.080 1591.870 ;
        RECT 103.200 16.990 103.340 1591.550 ;
        RECT 97.620 16.670 97.880 16.990 ;
        RECT 103.140 16.670 103.400 16.990 ;
        RECT 97.680 2.400 97.820 16.670 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 530.910 19.280 531.230 19.340 ;
        RECT 609.110 19.280 609.430 19.340 ;
        RECT 530.910 19.140 609.430 19.280 ;
        RECT 530.910 19.080 531.230 19.140 ;
        RECT 609.110 19.080 609.430 19.140 ;
      LAYER via ;
        RECT 530.940 19.080 531.200 19.340 ;
        RECT 609.140 19.080 609.400 19.340 ;
      LAYER met2 ;
        RECT 529.560 1600.450 529.840 1604.000 ;
        RECT 529.560 1600.310 531.140 1600.450 ;
        RECT 529.560 1600.000 529.840 1600.310 ;
        RECT 531.000 19.370 531.140 1600.310 ;
        RECT 530.940 19.050 531.200 19.370 ;
        RECT 609.140 19.050 609.400 19.370 ;
        RECT 609.200 2.400 609.340 19.050 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 622.065 1539.265 622.235 1591.455 ;
        RECT 621.145 1490.985 621.315 1538.755 ;
        RECT 622.065 1462.085 622.235 1490.475 ;
        RECT 622.065 1369.605 622.235 1400.715 ;
        RECT 621.605 1297.185 621.775 1318.095 ;
        RECT 621.605 1110.865 621.775 1124.975 ;
        RECT 621.605 1014.305 621.775 1028.415 ;
        RECT 621.605 917.745 621.775 931.855 ;
        RECT 621.605 821.185 621.775 835.295 ;
        RECT 622.065 234.685 622.235 282.795 ;
      LAYER mcon ;
        RECT 622.065 1591.285 622.235 1591.455 ;
        RECT 621.145 1538.585 621.315 1538.755 ;
        RECT 622.065 1490.305 622.235 1490.475 ;
        RECT 622.065 1400.545 622.235 1400.715 ;
        RECT 621.605 1317.925 621.775 1318.095 ;
        RECT 621.605 1124.805 621.775 1124.975 ;
        RECT 621.605 1028.245 621.775 1028.415 ;
        RECT 621.605 931.685 621.775 931.855 ;
        RECT 621.605 835.125 621.775 835.295 ;
        RECT 622.065 282.625 622.235 282.795 ;
      LAYER met1 ;
        RECT 536.430 1591.440 536.750 1591.500 ;
        RECT 622.005 1591.440 622.295 1591.485 ;
        RECT 536.430 1591.300 622.295 1591.440 ;
        RECT 536.430 1591.240 536.750 1591.300 ;
        RECT 622.005 1591.255 622.295 1591.300 ;
        RECT 622.005 1539.420 622.295 1539.465 ;
        RECT 622.450 1539.420 622.770 1539.480 ;
        RECT 622.005 1539.280 622.770 1539.420 ;
        RECT 622.005 1539.235 622.295 1539.280 ;
        RECT 622.450 1539.220 622.770 1539.280 ;
        RECT 621.085 1538.740 621.375 1538.785 ;
        RECT 621.990 1538.740 622.310 1538.800 ;
        RECT 621.085 1538.600 622.310 1538.740 ;
        RECT 621.085 1538.555 621.375 1538.600 ;
        RECT 621.990 1538.540 622.310 1538.600 ;
        RECT 621.070 1491.140 621.390 1491.200 ;
        RECT 621.070 1491.000 621.585 1491.140 ;
        RECT 621.070 1490.940 621.390 1491.000 ;
        RECT 621.070 1490.460 621.390 1490.520 ;
        RECT 622.005 1490.460 622.295 1490.505 ;
        RECT 621.070 1490.320 622.295 1490.460 ;
        RECT 621.070 1490.260 621.390 1490.320 ;
        RECT 622.005 1490.275 622.295 1490.320 ;
        RECT 621.990 1462.240 622.310 1462.300 ;
        RECT 621.795 1462.100 622.310 1462.240 ;
        RECT 621.990 1462.040 622.310 1462.100 ;
        RECT 621.990 1414.780 622.310 1415.040 ;
        RECT 622.080 1414.360 622.220 1414.780 ;
        RECT 621.990 1414.100 622.310 1414.360 ;
        RECT 621.990 1400.700 622.310 1400.760 ;
        RECT 621.795 1400.560 622.310 1400.700 ;
        RECT 621.990 1400.500 622.310 1400.560 ;
        RECT 621.990 1369.760 622.310 1369.820 ;
        RECT 621.795 1369.620 622.310 1369.760 ;
        RECT 621.990 1369.560 622.310 1369.620 ;
        RECT 621.530 1318.080 621.850 1318.140 ;
        RECT 621.335 1317.940 621.850 1318.080 ;
        RECT 621.530 1317.880 621.850 1317.940 ;
        RECT 621.530 1297.340 621.850 1297.400 ;
        RECT 621.335 1297.200 621.850 1297.340 ;
        RECT 621.530 1297.140 621.850 1297.200 ;
        RECT 621.530 1269.600 621.850 1269.860 ;
        RECT 621.620 1269.120 621.760 1269.600 ;
        RECT 621.990 1269.120 622.310 1269.180 ;
        RECT 621.620 1268.980 622.310 1269.120 ;
        RECT 621.990 1268.920 622.310 1268.980 ;
        RECT 621.990 1221.860 622.310 1221.920 ;
        RECT 621.620 1221.720 622.310 1221.860 ;
        RECT 621.620 1221.240 621.760 1221.720 ;
        RECT 621.990 1221.660 622.310 1221.720 ;
        RECT 621.530 1220.980 621.850 1221.240 ;
        RECT 621.530 1173.040 621.850 1173.300 ;
        RECT 621.620 1172.560 621.760 1173.040 ;
        RECT 621.990 1172.560 622.310 1172.620 ;
        RECT 621.620 1172.420 622.310 1172.560 ;
        RECT 621.990 1172.360 622.310 1172.420 ;
        RECT 621.530 1124.960 621.850 1125.020 ;
        RECT 621.335 1124.820 621.850 1124.960 ;
        RECT 621.530 1124.760 621.850 1124.820 ;
        RECT 621.530 1111.020 621.850 1111.080 ;
        RECT 621.335 1110.880 621.850 1111.020 ;
        RECT 621.530 1110.820 621.850 1110.880 ;
        RECT 621.530 1076.480 621.850 1076.740 ;
        RECT 621.620 1076.000 621.760 1076.480 ;
        RECT 621.990 1076.000 622.310 1076.060 ;
        RECT 621.620 1075.860 622.310 1076.000 ;
        RECT 621.990 1075.800 622.310 1075.860 ;
        RECT 621.530 1028.400 621.850 1028.460 ;
        RECT 621.335 1028.260 621.850 1028.400 ;
        RECT 621.530 1028.200 621.850 1028.260 ;
        RECT 621.530 1014.460 621.850 1014.520 ;
        RECT 621.335 1014.320 621.850 1014.460 ;
        RECT 621.530 1014.260 621.850 1014.320 ;
        RECT 621.530 979.920 621.850 980.180 ;
        RECT 621.620 979.440 621.760 979.920 ;
        RECT 621.990 979.440 622.310 979.500 ;
        RECT 621.620 979.300 622.310 979.440 ;
        RECT 621.990 979.240 622.310 979.300 ;
        RECT 621.530 931.840 621.850 931.900 ;
        RECT 621.335 931.700 621.850 931.840 ;
        RECT 621.530 931.640 621.850 931.700 ;
        RECT 621.530 917.900 621.850 917.960 ;
        RECT 621.335 917.760 621.850 917.900 ;
        RECT 621.530 917.700 621.850 917.760 ;
        RECT 621.530 883.360 621.850 883.620 ;
        RECT 621.620 882.880 621.760 883.360 ;
        RECT 621.990 882.880 622.310 882.940 ;
        RECT 621.620 882.740 622.310 882.880 ;
        RECT 621.990 882.680 622.310 882.740 ;
        RECT 621.530 835.280 621.850 835.340 ;
        RECT 621.335 835.140 621.850 835.280 ;
        RECT 621.530 835.080 621.850 835.140 ;
        RECT 621.530 821.340 621.850 821.400 ;
        RECT 621.335 821.200 621.850 821.340 ;
        RECT 621.530 821.140 621.850 821.200 ;
        RECT 621.530 786.800 621.850 787.060 ;
        RECT 621.620 786.320 621.760 786.800 ;
        RECT 621.990 786.320 622.310 786.380 ;
        RECT 621.620 786.180 622.310 786.320 ;
        RECT 621.990 786.120 622.310 786.180 ;
        RECT 621.990 772.720 622.310 772.780 ;
        RECT 622.910 772.720 623.230 772.780 ;
        RECT 621.990 772.580 623.230 772.720 ;
        RECT 621.990 772.520 622.310 772.580 ;
        RECT 622.910 772.520 623.230 772.580 ;
        RECT 621.530 689.900 621.850 690.160 ;
        RECT 621.620 689.760 621.760 689.900 ;
        RECT 621.990 689.760 622.310 689.820 ;
        RECT 621.620 689.620 622.310 689.760 ;
        RECT 621.990 689.560 622.310 689.620 ;
        RECT 621.990 676.160 622.310 676.220 ;
        RECT 622.910 676.160 623.230 676.220 ;
        RECT 621.990 676.020 623.230 676.160 ;
        RECT 621.990 675.960 622.310 676.020 ;
        RECT 622.910 675.960 623.230 676.020 ;
        RECT 621.530 593.340 621.850 593.600 ;
        RECT 621.620 593.200 621.760 593.340 ;
        RECT 621.990 593.200 622.310 593.260 ;
        RECT 621.620 593.060 622.310 593.200 ;
        RECT 621.990 593.000 622.310 593.060 ;
        RECT 621.990 579.600 622.310 579.660 ;
        RECT 622.910 579.600 623.230 579.660 ;
        RECT 621.990 579.460 623.230 579.600 ;
        RECT 621.990 579.400 622.310 579.460 ;
        RECT 622.910 579.400 623.230 579.460 ;
        RECT 621.530 496.780 621.850 497.040 ;
        RECT 621.620 496.640 621.760 496.780 ;
        RECT 621.990 496.640 622.310 496.700 ;
        RECT 621.620 496.500 622.310 496.640 ;
        RECT 621.990 496.440 622.310 496.500 ;
        RECT 621.990 483.040 622.310 483.100 ;
        RECT 622.910 483.040 623.230 483.100 ;
        RECT 621.990 482.900 623.230 483.040 ;
        RECT 621.990 482.840 622.310 482.900 ;
        RECT 622.910 482.840 623.230 482.900 ;
        RECT 621.530 400.220 621.850 400.480 ;
        RECT 621.620 399.740 621.760 400.220 ;
        RECT 621.990 399.740 622.310 399.800 ;
        RECT 621.620 399.600 622.310 399.740 ;
        RECT 621.990 399.540 622.310 399.600 ;
        RECT 621.990 331.400 622.310 331.460 ;
        RECT 622.910 331.400 623.230 331.460 ;
        RECT 621.990 331.260 623.230 331.400 ;
        RECT 621.990 331.200 622.310 331.260 ;
        RECT 622.910 331.200 623.230 331.260 ;
        RECT 621.990 303.180 622.310 303.240 ;
        RECT 622.910 303.180 623.230 303.240 ;
        RECT 621.990 303.040 623.230 303.180 ;
        RECT 621.990 302.980 622.310 303.040 ;
        RECT 622.910 302.980 623.230 303.040 ;
        RECT 621.990 282.780 622.310 282.840 ;
        RECT 621.795 282.640 622.310 282.780 ;
        RECT 621.990 282.580 622.310 282.640 ;
        RECT 622.005 234.840 622.295 234.885 ;
        RECT 622.450 234.840 622.770 234.900 ;
        RECT 622.005 234.700 622.770 234.840 ;
        RECT 622.005 234.655 622.295 234.700 ;
        RECT 622.450 234.640 622.770 234.700 ;
        RECT 621.990 138.280 622.310 138.340 ;
        RECT 622.910 138.280 623.230 138.340 ;
        RECT 621.990 138.140 623.230 138.280 ;
        RECT 621.990 138.080 622.310 138.140 ;
        RECT 622.910 138.080 623.230 138.140 ;
        RECT 621.990 90.000 622.310 90.060 ;
        RECT 622.910 90.000 623.230 90.060 ;
        RECT 621.990 89.860 623.230 90.000 ;
        RECT 621.990 89.800 622.310 89.860 ;
        RECT 622.910 89.800 623.230 89.860 ;
        RECT 621.990 65.520 622.310 65.580 ;
        RECT 626.590 65.520 626.910 65.580 ;
        RECT 621.990 65.380 626.910 65.520 ;
        RECT 621.990 65.320 622.310 65.380 ;
        RECT 626.590 65.320 626.910 65.380 ;
      LAYER via ;
        RECT 536.460 1591.240 536.720 1591.500 ;
        RECT 622.480 1539.220 622.740 1539.480 ;
        RECT 622.020 1538.540 622.280 1538.800 ;
        RECT 621.100 1490.940 621.360 1491.200 ;
        RECT 621.100 1490.260 621.360 1490.520 ;
        RECT 622.020 1462.040 622.280 1462.300 ;
        RECT 622.020 1414.780 622.280 1415.040 ;
        RECT 622.020 1414.100 622.280 1414.360 ;
        RECT 622.020 1400.500 622.280 1400.760 ;
        RECT 622.020 1369.560 622.280 1369.820 ;
        RECT 621.560 1317.880 621.820 1318.140 ;
        RECT 621.560 1297.140 621.820 1297.400 ;
        RECT 621.560 1269.600 621.820 1269.860 ;
        RECT 622.020 1268.920 622.280 1269.180 ;
        RECT 622.020 1221.660 622.280 1221.920 ;
        RECT 621.560 1220.980 621.820 1221.240 ;
        RECT 621.560 1173.040 621.820 1173.300 ;
        RECT 622.020 1172.360 622.280 1172.620 ;
        RECT 621.560 1124.760 621.820 1125.020 ;
        RECT 621.560 1110.820 621.820 1111.080 ;
        RECT 621.560 1076.480 621.820 1076.740 ;
        RECT 622.020 1075.800 622.280 1076.060 ;
        RECT 621.560 1028.200 621.820 1028.460 ;
        RECT 621.560 1014.260 621.820 1014.520 ;
        RECT 621.560 979.920 621.820 980.180 ;
        RECT 622.020 979.240 622.280 979.500 ;
        RECT 621.560 931.640 621.820 931.900 ;
        RECT 621.560 917.700 621.820 917.960 ;
        RECT 621.560 883.360 621.820 883.620 ;
        RECT 622.020 882.680 622.280 882.940 ;
        RECT 621.560 835.080 621.820 835.340 ;
        RECT 621.560 821.140 621.820 821.400 ;
        RECT 621.560 786.800 621.820 787.060 ;
        RECT 622.020 786.120 622.280 786.380 ;
        RECT 622.020 772.520 622.280 772.780 ;
        RECT 622.940 772.520 623.200 772.780 ;
        RECT 621.560 689.900 621.820 690.160 ;
        RECT 622.020 689.560 622.280 689.820 ;
        RECT 622.020 675.960 622.280 676.220 ;
        RECT 622.940 675.960 623.200 676.220 ;
        RECT 621.560 593.340 621.820 593.600 ;
        RECT 622.020 593.000 622.280 593.260 ;
        RECT 622.020 579.400 622.280 579.660 ;
        RECT 622.940 579.400 623.200 579.660 ;
        RECT 621.560 496.780 621.820 497.040 ;
        RECT 622.020 496.440 622.280 496.700 ;
        RECT 622.020 482.840 622.280 483.100 ;
        RECT 622.940 482.840 623.200 483.100 ;
        RECT 621.560 400.220 621.820 400.480 ;
        RECT 622.020 399.540 622.280 399.800 ;
        RECT 622.020 331.200 622.280 331.460 ;
        RECT 622.940 331.200 623.200 331.460 ;
        RECT 622.020 302.980 622.280 303.240 ;
        RECT 622.940 302.980 623.200 303.240 ;
        RECT 622.020 282.580 622.280 282.840 ;
        RECT 622.480 234.640 622.740 234.900 ;
        RECT 622.020 138.080 622.280 138.340 ;
        RECT 622.940 138.080 623.200 138.340 ;
        RECT 622.020 89.800 622.280 90.060 ;
        RECT 622.940 89.800 623.200 90.060 ;
        RECT 622.020 65.320 622.280 65.580 ;
        RECT 626.620 65.320 626.880 65.580 ;
      LAYER met2 ;
        RECT 536.460 1600.000 536.740 1604.000 ;
        RECT 536.520 1591.530 536.660 1600.000 ;
        RECT 536.460 1591.210 536.720 1591.530 ;
        RECT 622.480 1539.250 622.740 1539.510 ;
        RECT 622.080 1539.190 622.740 1539.250 ;
        RECT 622.080 1539.110 622.680 1539.190 ;
        RECT 622.080 1538.830 622.220 1539.110 ;
        RECT 622.020 1538.510 622.280 1538.830 ;
        RECT 621.100 1490.910 621.360 1491.230 ;
        RECT 621.160 1490.550 621.300 1490.910 ;
        RECT 621.100 1490.230 621.360 1490.550 ;
        RECT 622.020 1462.010 622.280 1462.330 ;
        RECT 622.080 1415.070 622.220 1462.010 ;
        RECT 622.020 1414.750 622.280 1415.070 ;
        RECT 622.020 1414.070 622.280 1414.390 ;
        RECT 622.080 1400.790 622.220 1414.070 ;
        RECT 622.020 1400.470 622.280 1400.790 ;
        RECT 622.020 1369.530 622.280 1369.850 ;
        RECT 622.080 1345.450 622.220 1369.530 ;
        RECT 621.620 1345.310 622.220 1345.450 ;
        RECT 621.620 1318.170 621.760 1345.310 ;
        RECT 621.560 1317.850 621.820 1318.170 ;
        RECT 621.560 1297.110 621.820 1297.430 ;
        RECT 621.620 1269.890 621.760 1297.110 ;
        RECT 621.560 1269.570 621.820 1269.890 ;
        RECT 622.020 1268.890 622.280 1269.210 ;
        RECT 622.080 1221.950 622.220 1268.890 ;
        RECT 622.020 1221.630 622.280 1221.950 ;
        RECT 621.560 1220.950 621.820 1221.270 ;
        RECT 621.620 1173.330 621.760 1220.950 ;
        RECT 621.560 1173.010 621.820 1173.330 ;
        RECT 622.020 1172.330 622.280 1172.650 ;
        RECT 622.080 1159.130 622.220 1172.330 ;
        RECT 621.620 1158.990 622.220 1159.130 ;
        RECT 621.620 1125.050 621.760 1158.990 ;
        RECT 621.560 1124.730 621.820 1125.050 ;
        RECT 621.560 1110.790 621.820 1111.110 ;
        RECT 621.620 1076.770 621.760 1110.790 ;
        RECT 621.560 1076.450 621.820 1076.770 ;
        RECT 622.020 1075.770 622.280 1076.090 ;
        RECT 622.080 1062.570 622.220 1075.770 ;
        RECT 621.620 1062.430 622.220 1062.570 ;
        RECT 621.620 1028.490 621.760 1062.430 ;
        RECT 621.560 1028.170 621.820 1028.490 ;
        RECT 621.560 1014.230 621.820 1014.550 ;
        RECT 621.620 980.210 621.760 1014.230 ;
        RECT 621.560 979.890 621.820 980.210 ;
        RECT 622.020 979.210 622.280 979.530 ;
        RECT 622.080 966.010 622.220 979.210 ;
        RECT 621.620 965.870 622.220 966.010 ;
        RECT 621.620 931.930 621.760 965.870 ;
        RECT 621.560 931.610 621.820 931.930 ;
        RECT 621.560 917.670 621.820 917.990 ;
        RECT 621.620 883.650 621.760 917.670 ;
        RECT 621.560 883.330 621.820 883.650 ;
        RECT 622.020 882.650 622.280 882.970 ;
        RECT 622.080 869.450 622.220 882.650 ;
        RECT 621.620 869.310 622.220 869.450 ;
        RECT 621.620 835.370 621.760 869.310 ;
        RECT 621.560 835.050 621.820 835.370 ;
        RECT 621.560 821.110 621.820 821.430 ;
        RECT 621.620 787.090 621.760 821.110 ;
        RECT 621.560 786.770 621.820 787.090 ;
        RECT 622.020 786.090 622.280 786.410 ;
        RECT 622.080 772.810 622.220 786.090 ;
        RECT 622.020 772.490 622.280 772.810 ;
        RECT 622.940 772.490 623.200 772.810 ;
        RECT 623.000 724.725 623.140 772.490 ;
        RECT 621.550 724.355 621.830 724.725 ;
        RECT 622.930 724.355 623.210 724.725 ;
        RECT 621.620 690.190 621.760 724.355 ;
        RECT 621.560 689.870 621.820 690.190 ;
        RECT 622.020 689.530 622.280 689.850 ;
        RECT 622.080 676.250 622.220 689.530 ;
        RECT 622.020 675.930 622.280 676.250 ;
        RECT 622.940 675.930 623.200 676.250 ;
        RECT 623.000 628.165 623.140 675.930 ;
        RECT 621.550 627.795 621.830 628.165 ;
        RECT 622.930 627.795 623.210 628.165 ;
        RECT 621.620 593.630 621.760 627.795 ;
        RECT 621.560 593.310 621.820 593.630 ;
        RECT 622.020 592.970 622.280 593.290 ;
        RECT 622.080 579.690 622.220 592.970 ;
        RECT 622.020 579.370 622.280 579.690 ;
        RECT 622.940 579.370 623.200 579.690 ;
        RECT 623.000 531.605 623.140 579.370 ;
        RECT 621.550 531.235 621.830 531.605 ;
        RECT 622.930 531.235 623.210 531.605 ;
        RECT 621.620 497.070 621.760 531.235 ;
        RECT 621.560 496.750 621.820 497.070 ;
        RECT 622.020 496.410 622.280 496.730 ;
        RECT 622.080 483.130 622.220 496.410 ;
        RECT 622.020 482.810 622.280 483.130 ;
        RECT 622.940 482.810 623.200 483.130 ;
        RECT 623.000 435.045 623.140 482.810 ;
        RECT 621.550 434.675 621.830 435.045 ;
        RECT 622.930 434.675 623.210 435.045 ;
        RECT 621.620 400.510 621.760 434.675 ;
        RECT 621.560 400.190 621.820 400.510 ;
        RECT 622.020 399.510 622.280 399.830 ;
        RECT 622.080 331.490 622.220 399.510 ;
        RECT 622.020 331.170 622.280 331.490 ;
        RECT 622.940 331.170 623.200 331.490 ;
        RECT 623.000 303.270 623.140 331.170 ;
        RECT 622.020 302.950 622.280 303.270 ;
        RECT 622.940 302.950 623.200 303.270 ;
        RECT 622.080 282.870 622.220 302.950 ;
        RECT 622.020 282.550 622.280 282.870 ;
        RECT 622.480 234.610 622.740 234.930 ;
        RECT 622.540 210.645 622.680 234.610 ;
        RECT 622.470 210.275 622.750 210.645 ;
        RECT 622.010 161.995 622.290 162.365 ;
        RECT 622.080 138.370 622.220 161.995 ;
        RECT 622.020 138.050 622.280 138.370 ;
        RECT 622.940 138.050 623.200 138.370 ;
        RECT 623.000 90.090 623.140 138.050 ;
        RECT 622.020 89.770 622.280 90.090 ;
        RECT 622.940 89.770 623.200 90.090 ;
        RECT 622.080 65.610 622.220 89.770 ;
        RECT 622.020 65.290 622.280 65.610 ;
        RECT 626.620 65.290 626.880 65.610 ;
        RECT 626.680 33.730 626.820 65.290 ;
        RECT 626.680 33.590 627.280 33.730 ;
        RECT 627.140 2.400 627.280 33.590 ;
        RECT 626.930 -4.800 627.490 2.400 ;
      LAYER via2 ;
        RECT 621.550 724.400 621.830 724.680 ;
        RECT 622.930 724.400 623.210 724.680 ;
        RECT 621.550 627.840 621.830 628.120 ;
        RECT 622.930 627.840 623.210 628.120 ;
        RECT 621.550 531.280 621.830 531.560 ;
        RECT 622.930 531.280 623.210 531.560 ;
        RECT 621.550 434.720 621.830 435.000 ;
        RECT 622.930 434.720 623.210 435.000 ;
        RECT 622.470 210.320 622.750 210.600 ;
        RECT 622.010 162.040 622.290 162.320 ;
      LAYER met3 ;
        RECT 621.525 724.690 621.855 724.705 ;
        RECT 622.905 724.690 623.235 724.705 ;
        RECT 621.525 724.390 623.235 724.690 ;
        RECT 621.525 724.375 621.855 724.390 ;
        RECT 622.905 724.375 623.235 724.390 ;
        RECT 621.525 628.130 621.855 628.145 ;
        RECT 622.905 628.130 623.235 628.145 ;
        RECT 621.525 627.830 623.235 628.130 ;
        RECT 621.525 627.815 621.855 627.830 ;
        RECT 622.905 627.815 623.235 627.830 ;
        RECT 621.525 531.570 621.855 531.585 ;
        RECT 622.905 531.570 623.235 531.585 ;
        RECT 621.525 531.270 623.235 531.570 ;
        RECT 621.525 531.255 621.855 531.270 ;
        RECT 622.905 531.255 623.235 531.270 ;
        RECT 621.525 435.010 621.855 435.025 ;
        RECT 622.905 435.010 623.235 435.025 ;
        RECT 621.525 434.710 623.235 435.010 ;
        RECT 621.525 434.695 621.855 434.710 ;
        RECT 622.905 434.695 623.235 434.710 ;
        RECT 622.445 210.620 622.775 210.625 ;
        RECT 622.190 210.610 622.775 210.620 ;
        RECT 622.190 210.310 623.000 210.610 ;
        RECT 622.190 210.300 622.775 210.310 ;
        RECT 622.445 210.295 622.775 210.300 ;
        RECT 621.985 162.340 622.315 162.345 ;
        RECT 621.985 162.330 622.570 162.340 ;
        RECT 621.985 162.030 622.770 162.330 ;
        RECT 621.985 162.020 622.570 162.030 ;
        RECT 621.985 162.015 622.315 162.020 ;
      LAYER via3 ;
        RECT 622.220 210.300 622.540 210.620 ;
        RECT 622.220 162.020 622.540 162.340 ;
      LAYER met4 ;
        RECT 622.215 210.295 622.545 210.625 ;
        RECT 622.230 162.345 622.530 210.295 ;
        RECT 622.215 162.015 622.545 162.345 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 345.560 1600.450 345.840 1604.000 ;
        RECT 345.560 1600.310 346.680 1600.450 ;
        RECT 345.560 1600.000 345.840 1600.310 ;
        RECT 346.540 18.205 346.680 1600.310 ;
        RECT 121.530 17.835 121.810 18.205 ;
        RECT 346.470 17.835 346.750 18.205 ;
        RECT 121.600 2.400 121.740 17.835 ;
        RECT 121.390 -4.800 121.950 2.400 ;
      LAYER via2 ;
        RECT 121.530 17.880 121.810 18.160 ;
        RECT 346.470 17.880 346.750 18.160 ;
      LAYER met3 ;
        RECT 121.505 18.170 121.835 18.185 ;
        RECT 346.445 18.170 346.775 18.185 ;
        RECT 121.505 17.870 346.775 18.170 ;
        RECT 121.505 17.855 121.835 17.870 ;
        RECT 346.445 17.855 346.775 17.870 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 151.410 1593.820 151.730 1593.880 ;
        RECT 354.730 1593.820 355.050 1593.880 ;
        RECT 151.410 1593.680 355.050 1593.820 ;
        RECT 151.410 1593.620 151.730 1593.680 ;
        RECT 354.730 1593.620 355.050 1593.680 ;
        RECT 145.430 20.300 145.750 20.360 ;
        RECT 151.410 20.300 151.730 20.360 ;
        RECT 145.430 20.160 151.730 20.300 ;
        RECT 145.430 20.100 145.750 20.160 ;
        RECT 151.410 20.100 151.730 20.160 ;
      LAYER via ;
        RECT 151.440 1593.620 151.700 1593.880 ;
        RECT 354.760 1593.620 355.020 1593.880 ;
        RECT 145.460 20.100 145.720 20.360 ;
        RECT 151.440 20.100 151.700 20.360 ;
      LAYER met2 ;
        RECT 354.760 1600.000 355.040 1604.000 ;
        RECT 354.820 1593.910 354.960 1600.000 ;
        RECT 151.440 1593.590 151.700 1593.910 ;
        RECT 354.760 1593.590 355.020 1593.910 ;
        RECT 151.500 20.390 151.640 1593.590 ;
        RECT 145.460 20.070 145.720 20.390 ;
        RECT 151.440 20.070 151.700 20.390 ;
        RECT 145.520 2.400 145.660 20.070 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 304.665 20.655 304.835 20.995 ;
        RECT 331.345 20.825 331.515 26.095 ;
        RECT 203.465 15.725 203.635 20.655 ;
        RECT 303.745 20.485 304.835 20.655 ;
      LAYER mcon ;
        RECT 331.345 25.925 331.515 26.095 ;
        RECT 304.665 20.825 304.835 20.995 ;
        RECT 203.465 20.485 203.635 20.655 ;
      LAYER met1 ;
        RECT 331.285 26.080 331.575 26.125 ;
        RECT 359.330 26.080 359.650 26.140 ;
        RECT 331.285 25.940 359.650 26.080 ;
        RECT 331.285 25.895 331.575 25.940 ;
        RECT 359.330 25.880 359.650 25.940 ;
        RECT 304.605 20.980 304.895 21.025 ;
        RECT 331.285 20.980 331.575 21.025 ;
        RECT 304.605 20.840 331.575 20.980 ;
        RECT 304.605 20.795 304.895 20.840 ;
        RECT 331.285 20.795 331.575 20.840 ;
        RECT 203.405 20.640 203.695 20.685 ;
        RECT 303.685 20.640 303.975 20.685 ;
        RECT 203.405 20.500 303.975 20.640 ;
        RECT 203.405 20.455 203.695 20.500 ;
        RECT 303.685 20.455 303.975 20.500 ;
        RECT 163.370 16.560 163.690 16.620 ;
        RECT 163.370 16.420 180.620 16.560 ;
        RECT 163.370 16.360 163.690 16.420 ;
        RECT 180.480 15.880 180.620 16.420 ;
        RECT 203.405 15.880 203.695 15.925 ;
        RECT 180.480 15.740 203.695 15.880 ;
        RECT 203.405 15.695 203.695 15.740 ;
      LAYER via ;
        RECT 359.360 25.880 359.620 26.140 ;
        RECT 163.400 16.360 163.660 16.620 ;
      LAYER met2 ;
        RECT 361.200 1600.450 361.480 1604.000 ;
        RECT 359.420 1600.310 361.480 1600.450 ;
        RECT 359.420 26.170 359.560 1600.310 ;
        RECT 361.200 1600.000 361.480 1600.310 ;
        RECT 359.360 25.850 359.620 26.170 ;
        RECT 163.400 16.330 163.660 16.650 ;
        RECT 163.460 2.400 163.600 16.330 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 185.910 1589.740 186.230 1589.800 ;
        RECT 368.070 1589.740 368.390 1589.800 ;
        RECT 185.910 1589.600 368.390 1589.740 ;
        RECT 185.910 1589.540 186.230 1589.600 ;
        RECT 368.070 1589.540 368.390 1589.600 ;
        RECT 180.850 16.560 181.170 16.620 ;
        RECT 185.910 16.560 186.230 16.620 ;
        RECT 180.850 16.420 186.230 16.560 ;
        RECT 180.850 16.360 181.170 16.420 ;
        RECT 185.910 16.360 186.230 16.420 ;
      LAYER via ;
        RECT 185.940 1589.540 186.200 1589.800 ;
        RECT 368.100 1589.540 368.360 1589.800 ;
        RECT 180.880 16.360 181.140 16.620 ;
        RECT 185.940 16.360 186.200 16.620 ;
      LAYER met2 ;
        RECT 368.100 1600.000 368.380 1604.000 ;
        RECT 368.160 1589.830 368.300 1600.000 ;
        RECT 185.940 1589.510 186.200 1589.830 ;
        RECT 368.100 1589.510 368.360 1589.830 ;
        RECT 186.000 16.650 186.140 1589.510 ;
        RECT 180.880 16.330 181.140 16.650 ;
        RECT 185.940 16.330 186.200 16.650 ;
        RECT 180.940 2.400 181.080 16.330 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 375.000 1600.450 375.280 1604.000 ;
        RECT 373.220 1600.310 375.280 1600.450 ;
        RECT 373.220 19.565 373.360 1600.310 ;
        RECT 375.000 1600.000 375.280 1600.310 ;
        RECT 198.810 19.195 199.090 19.565 ;
        RECT 373.150 19.195 373.430 19.565 ;
        RECT 198.880 2.400 199.020 19.195 ;
        RECT 198.670 -4.800 199.230 2.400 ;
      LAYER via2 ;
        RECT 198.810 19.240 199.090 19.520 ;
        RECT 373.150 19.240 373.430 19.520 ;
      LAYER met3 ;
        RECT 198.785 19.530 199.115 19.545 ;
        RECT 373.125 19.530 373.455 19.545 ;
        RECT 198.785 19.230 373.455 19.530 ;
        RECT 198.785 19.215 199.115 19.230 ;
        RECT 373.125 19.215 373.455 19.230 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 220.410 1589.400 220.730 1589.460 ;
        RECT 381.410 1589.400 381.730 1589.460 ;
        RECT 220.410 1589.260 381.730 1589.400 ;
        RECT 220.410 1589.200 220.730 1589.260 ;
        RECT 381.410 1589.200 381.730 1589.260 ;
        RECT 216.730 16.560 217.050 16.620 ;
        RECT 220.410 16.560 220.730 16.620 ;
        RECT 216.730 16.420 220.730 16.560 ;
        RECT 216.730 16.360 217.050 16.420 ;
        RECT 220.410 16.360 220.730 16.420 ;
      LAYER via ;
        RECT 220.440 1589.200 220.700 1589.460 ;
        RECT 381.440 1589.200 381.700 1589.460 ;
        RECT 216.760 16.360 217.020 16.620 ;
        RECT 220.440 16.360 220.700 16.620 ;
      LAYER met2 ;
        RECT 381.440 1600.000 381.720 1604.000 ;
        RECT 381.500 1589.490 381.640 1600.000 ;
        RECT 220.440 1589.170 220.700 1589.490 ;
        RECT 381.440 1589.170 381.700 1589.490 ;
        RECT 220.500 16.650 220.640 1589.170 ;
        RECT 216.760 16.330 217.020 16.650 ;
        RECT 220.440 16.330 220.700 16.650 ;
        RECT 216.820 2.400 216.960 16.330 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 270.625 14.365 270.795 15.895 ;
      LAYER mcon ;
        RECT 270.625 15.725 270.795 15.895 ;
      LAYER met1 ;
        RECT 270.565 15.880 270.855 15.925 ;
        RECT 386.470 15.880 386.790 15.940 ;
        RECT 270.565 15.740 386.790 15.880 ;
        RECT 270.565 15.695 270.855 15.740 ;
        RECT 386.470 15.680 386.790 15.740 ;
        RECT 234.670 14.520 234.990 14.580 ;
        RECT 270.565 14.520 270.855 14.565 ;
        RECT 234.670 14.380 270.855 14.520 ;
        RECT 234.670 14.320 234.990 14.380 ;
        RECT 270.565 14.335 270.855 14.380 ;
      LAYER via ;
        RECT 386.500 15.680 386.760 15.940 ;
        RECT 234.700 14.320 234.960 14.580 ;
      LAYER met2 ;
        RECT 388.340 1600.450 388.620 1604.000 ;
        RECT 386.560 1600.310 388.620 1600.450 ;
        RECT 386.560 15.970 386.700 1600.310 ;
        RECT 388.340 1600.000 388.620 1600.310 ;
        RECT 386.500 15.650 386.760 15.970 ;
        RECT 234.700 14.290 234.960 14.610 ;
        RECT 234.760 2.400 234.900 14.290 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 56.190 16.900 56.510 16.960 ;
        RECT 61.710 16.900 62.030 16.960 ;
        RECT 56.190 16.760 62.030 16.900 ;
        RECT 56.190 16.700 56.510 16.760 ;
        RECT 61.710 16.700 62.030 16.760 ;
      LAYER via ;
        RECT 56.220 16.700 56.480 16.960 ;
        RECT 61.740 16.700 62.000 16.960 ;
      LAYER met2 ;
        RECT 320.720 1600.000 321.000 1604.000 ;
        RECT 320.780 1592.405 320.920 1600.000 ;
        RECT 61.730 1592.035 62.010 1592.405 ;
        RECT 320.710 1592.035 320.990 1592.405 ;
        RECT 61.800 16.990 61.940 1592.035 ;
        RECT 56.220 16.670 56.480 16.990 ;
        RECT 61.740 16.670 62.000 16.990 ;
        RECT 56.280 2.400 56.420 16.670 ;
        RECT 56.070 -4.800 56.630 2.400 ;
      LAYER via2 ;
        RECT 61.730 1592.080 62.010 1592.360 ;
        RECT 320.710 1592.080 320.990 1592.360 ;
      LAYER met3 ;
        RECT 61.705 1592.370 62.035 1592.385 ;
        RECT 320.685 1592.370 321.015 1592.385 ;
        RECT 61.705 1592.070 321.015 1592.370 ;
        RECT 61.705 1592.055 62.035 1592.070 ;
        RECT 320.685 1592.055 321.015 1592.070 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 324.370 1579.880 324.690 1579.940 ;
        RECT 328.510 1579.880 328.830 1579.940 ;
        RECT 324.370 1579.740 328.830 1579.880 ;
        RECT 324.370 1579.680 324.690 1579.740 ;
        RECT 328.510 1579.680 328.830 1579.740 ;
        RECT 80.110 19.280 80.430 19.340 ;
        RECT 324.370 19.280 324.690 19.340 ;
        RECT 80.110 19.140 324.690 19.280 ;
        RECT 80.110 19.080 80.430 19.140 ;
        RECT 324.370 19.080 324.690 19.140 ;
      LAYER via ;
        RECT 324.400 1579.680 324.660 1579.940 ;
        RECT 328.540 1579.680 328.800 1579.940 ;
        RECT 80.140 19.080 80.400 19.340 ;
        RECT 324.400 19.080 324.660 19.340 ;
      LAYER met2 ;
        RECT 329.920 1600.450 330.200 1604.000 ;
        RECT 328.600 1600.310 330.200 1600.450 ;
        RECT 328.600 1579.970 328.740 1600.310 ;
        RECT 329.920 1600.000 330.200 1600.310 ;
        RECT 324.400 1579.650 324.660 1579.970 ;
        RECT 328.540 1579.650 328.800 1579.970 ;
        RECT 324.460 19.370 324.600 1579.650 ;
        RECT 80.140 19.050 80.400 19.370 ;
        RECT 324.400 19.050 324.660 19.370 ;
        RECT 80.200 2.400 80.340 19.050 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 1592.120 110.330 1592.180 ;
        RECT 338.630 1592.120 338.950 1592.180 ;
        RECT 110.010 1591.980 338.950 1592.120 ;
        RECT 110.010 1591.920 110.330 1591.980 ;
        RECT 338.630 1591.920 338.950 1591.980 ;
        RECT 103.570 14.860 103.890 14.920 ;
        RECT 110.010 14.860 110.330 14.920 ;
        RECT 103.570 14.720 110.330 14.860 ;
        RECT 103.570 14.660 103.890 14.720 ;
        RECT 110.010 14.660 110.330 14.720 ;
      LAYER via ;
        RECT 110.040 1591.920 110.300 1592.180 ;
        RECT 338.660 1591.920 338.920 1592.180 ;
        RECT 103.600 14.660 103.860 14.920 ;
        RECT 110.040 14.660 110.300 14.920 ;
      LAYER met2 ;
        RECT 338.660 1600.000 338.940 1604.000 ;
        RECT 338.720 1592.210 338.860 1600.000 ;
        RECT 110.040 1591.890 110.300 1592.210 ;
        RECT 338.660 1591.890 338.920 1592.210 ;
        RECT 110.100 14.950 110.240 1591.890 ;
        RECT 103.600 14.630 103.860 14.950 ;
        RECT 110.040 14.630 110.300 14.950 ;
        RECT 103.660 2.400 103.800 14.630 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 345.530 1579.880 345.850 1579.940 ;
        RECT 346.910 1579.880 347.230 1579.940 ;
        RECT 345.530 1579.740 347.230 1579.880 ;
        RECT 345.530 1579.680 345.850 1579.740 ;
        RECT 346.910 1579.680 347.230 1579.740 ;
        RECT 127.490 19.960 127.810 20.020 ;
        RECT 345.530 19.960 345.850 20.020 ;
        RECT 127.490 19.820 345.850 19.960 ;
        RECT 127.490 19.760 127.810 19.820 ;
        RECT 345.530 19.760 345.850 19.820 ;
      LAYER via ;
        RECT 345.560 1579.680 345.820 1579.940 ;
        RECT 346.940 1579.680 347.200 1579.940 ;
        RECT 127.520 19.760 127.780 20.020 ;
        RECT 345.560 19.760 345.820 20.020 ;
      LAYER met2 ;
        RECT 347.860 1600.450 348.140 1604.000 ;
        RECT 347.000 1600.310 348.140 1600.450 ;
        RECT 347.000 1579.970 347.140 1600.310 ;
        RECT 347.860 1600.000 348.140 1600.310 ;
        RECT 345.560 1579.650 345.820 1579.970 ;
        RECT 346.940 1579.650 347.200 1579.970 ;
        RECT 345.620 20.050 345.760 1579.650 ;
        RECT 127.520 19.730 127.780 20.050 ;
        RECT 345.560 19.730 345.820 20.050 ;
        RECT 127.580 2.400 127.720 19.730 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 2.960 26.610 3.020 ;
        RECT 27.210 2.960 27.530 3.020 ;
        RECT 26.290 2.820 27.530 2.960 ;
        RECT 26.290 2.760 26.610 2.820 ;
        RECT 27.210 2.760 27.530 2.820 ;
      LAYER via ;
        RECT 26.320 2.760 26.580 3.020 ;
        RECT 27.240 2.760 27.500 3.020 ;
      LAYER met2 ;
        RECT 309.680 1600.000 309.960 1604.000 ;
        RECT 309.740 1590.365 309.880 1600.000 ;
        RECT 27.230 1589.995 27.510 1590.365 ;
        RECT 309.670 1589.995 309.950 1590.365 ;
        RECT 27.300 3.050 27.440 1589.995 ;
        RECT 26.320 2.730 26.580 3.050 ;
        RECT 27.240 2.730 27.500 3.050 ;
        RECT 26.380 2.400 26.520 2.730 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 27.230 1590.040 27.510 1590.320 ;
        RECT 309.670 1590.040 309.950 1590.320 ;
      LAYER met3 ;
        RECT 27.205 1590.330 27.535 1590.345 ;
        RECT 309.645 1590.330 309.975 1590.345 ;
        RECT 27.205 1590.030 309.975 1590.330 ;
        RECT 27.205 1590.015 27.535 1590.030 ;
        RECT 309.645 1590.015 309.975 1590.030 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 17.920 32.590 17.980 ;
        RECT 310.570 17.920 310.890 17.980 ;
        RECT 32.270 17.780 310.890 17.920 ;
        RECT 32.270 17.720 32.590 17.780 ;
        RECT 310.570 17.720 310.890 17.780 ;
      LAYER via ;
        RECT 32.300 17.720 32.560 17.980 ;
        RECT 310.600 17.720 310.860 17.980 ;
      LAYER met2 ;
        RECT 311.980 1600.450 312.260 1604.000 ;
        RECT 310.660 1600.310 312.260 1600.450 ;
        RECT 310.660 18.010 310.800 1600.310 ;
        RECT 311.980 1600.000 312.260 1600.310 ;
        RECT 32.300 17.690 32.560 18.010 ;
        RECT 310.600 17.690 310.860 18.010 ;
        RECT 32.360 2.400 32.500 17.690 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.480 3243.600 684.050 3244.660 ;
        RECT 1331.480 3243.600 1334.050 3244.660 ;
        RECT 1931.480 3243.600 1934.050 3244.660 ;
        RECT 2581.480 3243.600 2584.050 3244.660 ;
        RECT 2581.480 2043.600 2584.050 2044.660 ;
        RECT 1552.430 1611.575 1555.000 1612.635 ;
      LAYER via3 ;
        RECT 682.500 3243.620 684.020 3244.630 ;
        RECT 1332.500 3243.620 1334.020 3244.630 ;
        RECT 1932.500 3243.620 1934.020 3244.630 ;
        RECT 2582.500 3243.620 2584.020 3244.630 ;
        RECT 2582.500 2043.620 2584.020 2044.630 ;
        RECT 1552.460 1611.605 1553.980 1612.615 ;
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 364.020 3271.235 367.020 3529.000 ;
        RECT 382.020 3271.235 385.020 3538.400 ;
        RECT 400.020 3271.235 403.020 3547.800 ;
        RECT 418.020 3271.235 421.020 3557.200 ;
        RECT 544.020 3271.235 547.020 3529.000 ;
        RECT 562.020 3271.235 565.020 3538.400 ;
        RECT 580.020 3271.235 583.020 3547.800 ;
        RECT 598.020 3271.235 601.020 3557.200 ;
        RECT 682.470 2803.670 684.070 3244.680 ;
        RECT 382.020 2715.000 385.020 2785.000 ;
        RECT 400.020 2715.000 403.020 2785.000 ;
        RECT 418.020 2715.000 421.020 2785.000 ;
        RECT 562.020 2715.000 565.020 2785.000 ;
        RECT 580.020 2715.000 583.020 2785.000 ;
        RECT 598.020 2715.000 601.020 2785.000 ;
        RECT 724.020 2715.000 727.020 3529.000 ;
        RECT 742.020 2715.000 745.020 3538.400 ;
        RECT 760.020 2715.000 763.020 3547.800 ;
        RECT 778.020 2715.000 781.020 3557.200 ;
        RECT 904.020 2715.000 907.020 3529.000 ;
        RECT 922.020 2715.000 925.020 3538.400 ;
        RECT 940.020 3271.235 943.020 3547.800 ;
        RECT 958.020 3271.235 961.020 3557.200 ;
        RECT 1084.020 3271.235 1087.020 3529.000 ;
        RECT 1102.020 3271.235 1105.020 3538.400 ;
        RECT 1120.020 3271.235 1123.020 3547.800 ;
        RECT 1138.020 3271.235 1141.020 3557.200 ;
        RECT 1264.020 3271.235 1267.020 3529.000 ;
        RECT 1282.020 3271.235 1285.020 3538.400 ;
        RECT 1300.020 3271.235 1303.020 3547.800 ;
        RECT 1318.020 3271.235 1321.020 3557.200 ;
        RECT 1332.470 2803.670 1334.070 3244.680 ;
        RECT 940.020 2715.000 943.020 2785.000 ;
        RECT 958.020 2715.000 961.020 2785.000 ;
        RECT 1102.020 2715.000 1105.020 2785.000 ;
        RECT 1120.020 2715.000 1123.020 2785.000 ;
        RECT 1138.020 2715.000 1141.020 2785.000 ;
        RECT 1282.020 2715.000 1285.020 2785.000 ;
        RECT 1300.020 2715.000 1303.020 2785.000 ;
        RECT 1318.020 2715.000 1321.020 2785.000 ;
        RECT 320.970 1610.640 322.570 2688.240 ;
        RECT 364.020 -9.320 367.020 1585.000 ;
        RECT 382.020 -18.720 385.020 1585.000 ;
        RECT 400.020 -28.120 403.020 1585.000 ;
        RECT 418.020 -37.520 421.020 1585.000 ;
        RECT 544.020 -9.320 547.020 1585.000 ;
        RECT 562.020 -18.720 565.020 1585.000 ;
        RECT 580.020 -28.120 583.020 1585.000 ;
        RECT 598.020 -37.520 601.020 1585.000 ;
        RECT 724.020 -9.320 727.020 1585.000 ;
        RECT 742.020 -18.720 745.020 1585.000 ;
        RECT 760.020 -28.120 763.020 1585.000 ;
        RECT 778.020 -37.520 781.020 1585.000 ;
        RECT 904.020 -9.320 907.020 1585.000 ;
        RECT 922.020 -18.720 925.020 1585.000 ;
        RECT 940.020 -28.120 943.020 1585.000 ;
        RECT 958.020 -37.520 961.020 1585.000 ;
        RECT 1084.020 -9.320 1087.020 1585.000 ;
        RECT 1102.020 -18.720 1105.020 1585.000 ;
        RECT 1120.020 -28.120 1123.020 1585.000 ;
        RECT 1138.020 -37.520 1141.020 1585.000 ;
        RECT 1264.020 -9.320 1267.020 1585.000 ;
        RECT 1282.020 -18.720 1285.020 1585.000 ;
        RECT 1300.020 -28.120 1303.020 1585.000 ;
        RECT 1318.020 -37.520 1321.020 1585.000 ;
        RECT 1444.020 -9.320 1447.020 3529.000 ;
        RECT 1462.020 -18.720 1465.020 3538.400 ;
        RECT 1480.020 -28.120 1483.020 3547.800 ;
        RECT 1498.020 -37.520 1501.020 3557.200 ;
        RECT 1624.020 3271.235 1627.020 3529.000 ;
        RECT 1642.020 3271.235 1645.020 3538.400 ;
        RECT 1660.020 3271.235 1663.020 3547.800 ;
        RECT 1678.020 3271.235 1681.020 3557.200 ;
        RECT 1804.020 3271.235 1807.020 3529.000 ;
        RECT 1822.020 3271.235 1825.020 3538.400 ;
        RECT 1840.020 3271.235 1843.020 3547.800 ;
        RECT 1858.020 3271.235 1861.020 3557.200 ;
        RECT 1932.470 2803.670 1934.070 3244.680 ;
        RECT 1624.020 2071.235 1627.020 2785.000 ;
        RECT 1642.020 2071.235 1645.020 2785.000 ;
        RECT 1660.020 2071.235 1663.020 2785.000 ;
        RECT 1678.020 2071.235 1681.020 2785.000 ;
        RECT 1804.020 2071.235 1807.020 2785.000 ;
        RECT 1822.020 2071.235 1825.020 2785.000 ;
        RECT 1840.020 2071.235 1843.020 2785.000 ;
        RECT 1858.020 2071.235 1861.020 2785.000 ;
        RECT 1552.410 1611.555 1554.010 2052.565 ;
        RECT 1984.020 1515.000 1987.020 3529.000 ;
        RECT 2002.020 1515.000 2005.020 3538.400 ;
        RECT 2020.020 1515.000 2023.020 3547.800 ;
        RECT 2038.020 1515.000 2041.020 3557.200 ;
        RECT 2164.020 1515.000 2167.020 3529.000 ;
        RECT 2182.020 3271.235 2185.020 3538.400 ;
        RECT 2200.020 3271.235 2203.020 3547.800 ;
        RECT 2218.020 3271.235 2221.020 3557.200 ;
        RECT 2344.020 3271.235 2347.020 3529.000 ;
        RECT 2362.020 3271.235 2365.020 3538.400 ;
        RECT 2380.020 3271.235 2383.020 3547.800 ;
        RECT 2398.020 3271.235 2401.020 3557.200 ;
        RECT 2524.020 3271.235 2527.020 3529.000 ;
        RECT 2542.020 3271.235 2545.020 3538.400 ;
        RECT 2560.020 3271.235 2563.020 3547.800 ;
        RECT 2578.020 3271.235 2581.020 3557.200 ;
        RECT 2582.470 2803.670 2584.070 3244.680 ;
        RECT 2182.020 2071.235 2185.020 2785.000 ;
        RECT 2200.020 2071.235 2203.020 2785.000 ;
        RECT 2218.020 2071.235 2221.020 2785.000 ;
        RECT 2344.020 2071.235 2347.020 2785.000 ;
        RECT 2362.020 2071.235 2365.020 2785.000 ;
        RECT 2380.020 2071.235 2383.020 2785.000 ;
        RECT 2398.020 2071.235 2401.020 2785.000 ;
        RECT 2524.020 2071.235 2527.020 2785.000 ;
        RECT 2542.020 2071.235 2545.020 2785.000 ;
        RECT 2560.020 2071.235 2563.020 2785.000 ;
        RECT 2578.020 2071.235 2581.020 2785.000 ;
        RECT 2582.470 1603.670 2584.070 2044.680 ;
        RECT 1570.970 410.640 1572.570 1488.240 ;
        RECT 1624.020 -9.320 1627.020 385.000 ;
        RECT 1642.020 -18.720 1645.020 385.000 ;
        RECT 1660.020 -28.120 1663.020 385.000 ;
        RECT 1678.020 -37.520 1681.020 385.000 ;
        RECT 1804.020 -9.320 1807.020 385.000 ;
        RECT 1822.020 -18.720 1825.020 385.000 ;
        RECT 1840.020 -28.120 1843.020 385.000 ;
        RECT 1858.020 -37.520 1861.020 385.000 ;
        RECT 1984.020 -9.320 1987.020 385.000 ;
        RECT 2002.020 -18.720 2005.020 385.000 ;
        RECT 2020.020 -28.120 2023.020 385.000 ;
        RECT 2038.020 -37.520 2041.020 385.000 ;
        RECT 2164.020 -9.320 2167.020 385.000 ;
        RECT 2182.020 -18.720 2185.020 385.000 ;
        RECT 2200.020 -28.120 2203.020 385.000 ;
        RECT 2218.020 -37.520 2221.020 385.000 ;
        RECT 2344.020 -9.320 2347.020 385.000 ;
        RECT 2362.020 -18.720 2365.020 385.000 ;
        RECT 2380.020 -28.120 2383.020 385.000 ;
        RECT 2398.020 -37.520 2401.020 385.000 ;
        RECT 2524.020 -9.320 2527.020 385.000 ;
        RECT 2542.020 -18.720 2545.020 385.000 ;
        RECT 2560.020 -28.120 2563.020 385.000 ;
        RECT 2578.020 -37.520 2581.020 385.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 682.680 3125.090 683.860 3126.270 ;
        RECT 682.680 3123.490 683.860 3124.670 ;
        RECT 682.680 3107.090 683.860 3108.270 ;
        RECT 682.680 3105.490 683.860 3106.670 ;
        RECT 682.680 3089.090 683.860 3090.270 ;
        RECT 682.680 3087.490 683.860 3088.670 ;
        RECT 682.680 3071.090 683.860 3072.270 ;
        RECT 682.680 3069.490 683.860 3070.670 ;
        RECT 682.680 2945.090 683.860 2946.270 ;
        RECT 682.680 2943.490 683.860 2944.670 ;
        RECT 682.680 2927.090 683.860 2928.270 ;
        RECT 682.680 2925.490 683.860 2926.670 ;
        RECT 682.680 2909.090 683.860 2910.270 ;
        RECT 682.680 2907.490 683.860 2908.670 ;
        RECT 682.680 2891.090 683.860 2892.270 ;
        RECT 682.680 2889.490 683.860 2890.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 1332.680 3125.090 1333.860 3126.270 ;
        RECT 1332.680 3123.490 1333.860 3124.670 ;
        RECT 1332.680 3107.090 1333.860 3108.270 ;
        RECT 1332.680 3105.490 1333.860 3106.670 ;
        RECT 1332.680 3089.090 1333.860 3090.270 ;
        RECT 1332.680 3087.490 1333.860 3088.670 ;
        RECT 1332.680 3071.090 1333.860 3072.270 ;
        RECT 1332.680 3069.490 1333.860 3070.670 ;
        RECT 1332.680 2945.090 1333.860 2946.270 ;
        RECT 1332.680 2943.490 1333.860 2944.670 ;
        RECT 1332.680 2927.090 1333.860 2928.270 ;
        RECT 1332.680 2925.490 1333.860 2926.670 ;
        RECT 1332.680 2909.090 1333.860 2910.270 ;
        RECT 1332.680 2907.490 1333.860 2908.670 ;
        RECT 1332.680 2891.090 1333.860 2892.270 ;
        RECT 1332.680 2889.490 1333.860 2890.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 321.180 2585.090 322.360 2586.270 ;
        RECT 321.180 2583.490 322.360 2584.670 ;
        RECT 321.180 2567.090 322.360 2568.270 ;
        RECT 321.180 2565.490 322.360 2566.670 ;
        RECT 321.180 2549.090 322.360 2550.270 ;
        RECT 321.180 2547.490 322.360 2548.670 ;
        RECT 321.180 2531.090 322.360 2532.270 ;
        RECT 321.180 2529.490 322.360 2530.670 ;
        RECT 321.180 2405.090 322.360 2406.270 ;
        RECT 321.180 2403.490 322.360 2404.670 ;
        RECT 321.180 2387.090 322.360 2388.270 ;
        RECT 321.180 2385.490 322.360 2386.670 ;
        RECT 321.180 2369.090 322.360 2370.270 ;
        RECT 321.180 2367.490 322.360 2368.670 ;
        RECT 321.180 2351.090 322.360 2352.270 ;
        RECT 321.180 2349.490 322.360 2350.670 ;
        RECT 321.180 2225.090 322.360 2226.270 ;
        RECT 321.180 2223.490 322.360 2224.670 ;
        RECT 321.180 2207.090 322.360 2208.270 ;
        RECT 321.180 2205.490 322.360 2206.670 ;
        RECT 321.180 2189.090 322.360 2190.270 ;
        RECT 321.180 2187.490 322.360 2188.670 ;
        RECT 321.180 2171.090 322.360 2172.270 ;
        RECT 321.180 2169.490 322.360 2170.670 ;
        RECT 321.180 2045.090 322.360 2046.270 ;
        RECT 321.180 2043.490 322.360 2044.670 ;
        RECT 321.180 2027.090 322.360 2028.270 ;
        RECT 321.180 2025.490 322.360 2026.670 ;
        RECT 321.180 2009.090 322.360 2010.270 ;
        RECT 321.180 2007.490 322.360 2008.670 ;
        RECT 321.180 1991.090 322.360 1992.270 ;
        RECT 321.180 1989.490 322.360 1990.670 ;
        RECT 321.180 1865.090 322.360 1866.270 ;
        RECT 321.180 1863.490 322.360 1864.670 ;
        RECT 321.180 1847.090 322.360 1848.270 ;
        RECT 321.180 1845.490 322.360 1846.670 ;
        RECT 321.180 1829.090 322.360 1830.270 ;
        RECT 321.180 1827.490 322.360 1828.670 ;
        RECT 321.180 1811.090 322.360 1812.270 ;
        RECT 321.180 1809.490 322.360 1810.670 ;
        RECT 321.180 1685.090 322.360 1686.270 ;
        RECT 321.180 1683.490 322.360 1684.670 ;
        RECT 321.180 1667.090 322.360 1668.270 ;
        RECT 321.180 1665.490 322.360 1666.670 ;
        RECT 321.180 1649.090 322.360 1650.270 ;
        RECT 321.180 1647.490 322.360 1648.670 ;
        RECT 321.180 1631.090 322.360 1632.270 ;
        RECT 321.180 1629.490 322.360 1630.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1932.680 3125.090 1933.860 3126.270 ;
        RECT 1932.680 3123.490 1933.860 3124.670 ;
        RECT 1932.680 3107.090 1933.860 3108.270 ;
        RECT 1932.680 3105.490 1933.860 3106.670 ;
        RECT 1932.680 3089.090 1933.860 3090.270 ;
        RECT 1932.680 3087.490 1933.860 3088.670 ;
        RECT 1932.680 3071.090 1933.860 3072.270 ;
        RECT 1932.680 3069.490 1933.860 3070.670 ;
        RECT 1932.680 2945.090 1933.860 2946.270 ;
        RECT 1932.680 2943.490 1933.860 2944.670 ;
        RECT 1932.680 2927.090 1933.860 2928.270 ;
        RECT 1932.680 2925.490 1933.860 2926.670 ;
        RECT 1932.680 2909.090 1933.860 2910.270 ;
        RECT 1932.680 2907.490 1933.860 2908.670 ;
        RECT 1932.680 2891.090 1933.860 2892.270 ;
        RECT 1932.680 2889.490 1933.860 2890.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1552.620 2045.090 1553.800 2046.270 ;
        RECT 1552.620 2043.490 1553.800 2044.670 ;
        RECT 1552.620 2027.090 1553.800 2028.270 ;
        RECT 1552.620 2025.490 1553.800 2026.670 ;
        RECT 1552.620 2009.090 1553.800 2010.270 ;
        RECT 1552.620 2007.490 1553.800 2008.670 ;
        RECT 1552.620 1991.090 1553.800 1992.270 ;
        RECT 1552.620 1989.490 1553.800 1990.670 ;
        RECT 1552.620 1865.090 1553.800 1866.270 ;
        RECT 1552.620 1863.490 1553.800 1864.670 ;
        RECT 1552.620 1847.090 1553.800 1848.270 ;
        RECT 1552.620 1845.490 1553.800 1846.670 ;
        RECT 1552.620 1829.090 1553.800 1830.270 ;
        RECT 1552.620 1827.490 1553.800 1828.670 ;
        RECT 1552.620 1811.090 1553.800 1812.270 ;
        RECT 1552.620 1809.490 1553.800 1810.670 ;
        RECT 1552.620 1685.090 1553.800 1686.270 ;
        RECT 1552.620 1683.490 1553.800 1684.670 ;
        RECT 1552.620 1667.090 1553.800 1668.270 ;
        RECT 1552.620 1665.490 1553.800 1666.670 ;
        RECT 1552.620 1649.090 1553.800 1650.270 ;
        RECT 1552.620 1647.490 1553.800 1648.670 ;
        RECT 1552.620 1631.090 1553.800 1632.270 ;
        RECT 1552.620 1629.490 1553.800 1630.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2582.680 3125.090 2583.860 3126.270 ;
        RECT 2582.680 3123.490 2583.860 3124.670 ;
        RECT 2582.680 3107.090 2583.860 3108.270 ;
        RECT 2582.680 3105.490 2583.860 3106.670 ;
        RECT 2582.680 3089.090 2583.860 3090.270 ;
        RECT 2582.680 3087.490 2583.860 3088.670 ;
        RECT 2582.680 3071.090 2583.860 3072.270 ;
        RECT 2582.680 3069.490 2583.860 3070.670 ;
        RECT 2582.680 2945.090 2583.860 2946.270 ;
        RECT 2582.680 2943.490 2583.860 2944.670 ;
        RECT 2582.680 2927.090 2583.860 2928.270 ;
        RECT 2582.680 2925.490 2583.860 2926.670 ;
        RECT 2582.680 2909.090 2583.860 2910.270 ;
        RECT 2582.680 2907.490 2583.860 2908.670 ;
        RECT 2582.680 2891.090 2583.860 2892.270 ;
        RECT 2582.680 2889.490 2583.860 2890.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2582.680 2027.090 2583.860 2028.270 ;
        RECT 2582.680 2025.490 2583.860 2026.670 ;
        RECT 2582.680 2009.090 2583.860 2010.270 ;
        RECT 2582.680 2007.490 2583.860 2008.670 ;
        RECT 2582.680 1991.090 2583.860 1992.270 ;
        RECT 2582.680 1989.490 2583.860 1990.670 ;
        RECT 2582.680 1865.090 2583.860 1866.270 ;
        RECT 2582.680 1863.490 2583.860 1864.670 ;
        RECT 2582.680 1847.090 2583.860 1848.270 ;
        RECT 2582.680 1845.490 2583.860 1846.670 ;
        RECT 2582.680 1829.090 2583.860 1830.270 ;
        RECT 2582.680 1827.490 2583.860 1828.670 ;
        RECT 2582.680 1811.090 2583.860 1812.270 ;
        RECT 2582.680 1809.490 2583.860 1810.670 ;
        RECT 2582.680 1685.090 2583.860 1686.270 ;
        RECT 2582.680 1683.490 2583.860 1684.670 ;
        RECT 2582.680 1667.090 2583.860 1668.270 ;
        RECT 2582.680 1665.490 2583.860 1666.670 ;
        RECT 2582.680 1649.090 2583.860 1650.270 ;
        RECT 2582.680 1647.490 2583.860 1648.670 ;
        RECT 2582.680 1631.090 2583.860 1632.270 ;
        RECT 2582.680 1629.490 2583.860 1630.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1571.180 1469.090 1572.360 1470.270 ;
        RECT 1571.180 1467.490 1572.360 1468.670 ;
        RECT 1571.180 1451.090 1572.360 1452.270 ;
        RECT 1571.180 1449.490 1572.360 1450.670 ;
        RECT 1571.180 1325.090 1572.360 1326.270 ;
        RECT 1571.180 1323.490 1572.360 1324.670 ;
        RECT 1571.180 1307.090 1572.360 1308.270 ;
        RECT 1571.180 1305.490 1572.360 1306.670 ;
        RECT 1571.180 1289.090 1572.360 1290.270 ;
        RECT 1571.180 1287.490 1572.360 1288.670 ;
        RECT 1571.180 1271.090 1572.360 1272.270 ;
        RECT 1571.180 1269.490 1572.360 1270.670 ;
        RECT 1571.180 1145.090 1572.360 1146.270 ;
        RECT 1571.180 1143.490 1572.360 1144.670 ;
        RECT 1571.180 1127.090 1572.360 1128.270 ;
        RECT 1571.180 1125.490 1572.360 1126.670 ;
        RECT 1571.180 1109.090 1572.360 1110.270 ;
        RECT 1571.180 1107.490 1572.360 1108.670 ;
        RECT 1571.180 1091.090 1572.360 1092.270 ;
        RECT 1571.180 1089.490 1572.360 1090.670 ;
        RECT 1571.180 965.090 1572.360 966.270 ;
        RECT 1571.180 963.490 1572.360 964.670 ;
        RECT 1571.180 947.090 1572.360 948.270 ;
        RECT 1571.180 945.490 1572.360 946.670 ;
        RECT 1571.180 929.090 1572.360 930.270 ;
        RECT 1571.180 927.490 1572.360 928.670 ;
        RECT 1571.180 911.090 1572.360 912.270 ;
        RECT 1571.180 909.490 1572.360 910.670 ;
        RECT 1571.180 785.090 1572.360 786.270 ;
        RECT 1571.180 783.490 1572.360 784.670 ;
        RECT 1571.180 767.090 1572.360 768.270 ;
        RECT 1571.180 765.490 1572.360 766.670 ;
        RECT 1571.180 749.090 1572.360 750.270 ;
        RECT 1571.180 747.490 1572.360 748.670 ;
        RECT 1571.180 731.090 1572.360 732.270 ;
        RECT 1571.180 729.490 1572.360 730.670 ;
        RECT 1571.180 605.090 1572.360 606.270 ;
        RECT 1571.180 603.490 1572.360 604.670 ;
        RECT 1571.180 587.090 1572.360 588.270 ;
        RECT 1571.180 585.490 1572.360 586.670 ;
        RECT 1571.180 569.090 1572.360 570.270 ;
        RECT 1571.180 567.490 1572.360 568.670 ;
        RECT 1571.180 551.090 1572.360 552.270 ;
        RECT 1571.180 549.490 1572.360 550.670 ;
        RECT 1571.180 425.090 1572.360 426.270 ;
        RECT 1571.180 423.490 1572.360 424.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 682.470 3126.380 684.070 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 1332.470 3126.380 1334.070 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1932.470 3126.380 1934.070 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2582.470 3126.380 2584.070 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 682.470 3123.370 684.070 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 1332.470 3123.370 1334.070 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1932.470 3123.370 1934.070 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2582.470 3123.370 2584.070 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 682.470 3108.380 684.070 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 1332.470 3108.380 1334.070 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1932.470 3108.380 1934.070 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2582.470 3108.380 2584.070 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 682.470 3105.370 684.070 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 1332.470 3105.370 1334.070 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1932.470 3105.370 1934.070 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2582.470 3105.370 2584.070 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 682.470 3090.380 684.070 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1332.470 3090.380 1334.070 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1932.470 3090.380 1934.070 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2582.470 3090.380 2584.070 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 682.470 3087.370 684.070 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1332.470 3087.370 1334.070 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1932.470 3087.370 1934.070 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2582.470 3087.370 2584.070 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 682.470 3072.380 684.070 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1332.470 3072.380 1334.070 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1932.470 3072.380 1934.070 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2582.470 3072.380 2584.070 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 682.470 3069.370 684.070 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1332.470 3069.370 1334.070 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1932.470 3069.370 1934.070 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2582.470 3069.370 2584.070 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 682.470 2946.380 684.070 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 1332.470 2946.380 1334.070 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1932.470 2946.380 1934.070 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2582.470 2946.380 2584.070 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 682.470 2943.370 684.070 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 1332.470 2943.370 1334.070 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1932.470 2943.370 1934.070 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2582.470 2943.370 2584.070 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 682.470 2928.380 684.070 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 1332.470 2928.380 1334.070 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1932.470 2928.380 1934.070 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2582.470 2928.380 2584.070 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 682.470 2925.370 684.070 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 1332.470 2925.370 1334.070 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1932.470 2925.370 1934.070 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2582.470 2925.370 2584.070 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 682.470 2910.380 684.070 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1332.470 2910.380 1334.070 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1932.470 2910.380 1934.070 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2582.470 2910.380 2584.070 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 682.470 2907.370 684.070 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1332.470 2907.370 1334.070 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1932.470 2907.370 1934.070 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2582.470 2907.370 2584.070 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 682.470 2892.380 684.070 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1332.470 2892.380 1334.070 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1932.470 2892.380 1934.070 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2582.470 2892.380 2584.070 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 682.470 2889.370 684.070 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1332.470 2889.370 1334.070 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1932.470 2889.370 1934.070 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2582.470 2889.370 2584.070 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 320.970 2586.380 322.570 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 320.970 2583.370 322.570 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 320.970 2568.380 322.570 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 320.970 2565.370 322.570 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 320.970 2550.380 322.570 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 320.970 2547.370 322.570 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 320.970 2532.380 322.570 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 320.970 2529.370 322.570 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 320.970 2406.380 322.570 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 320.970 2403.370 322.570 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 320.970 2388.380 322.570 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 320.970 2385.370 322.570 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 320.970 2370.380 322.570 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 320.970 2367.370 322.570 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 320.970 2352.380 322.570 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 320.970 2349.370 322.570 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 320.970 2226.380 322.570 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 320.970 2223.370 322.570 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 320.970 2208.380 322.570 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 320.970 2205.370 322.570 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 320.970 2190.380 322.570 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 320.970 2187.370 322.570 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 320.970 2172.380 322.570 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 320.970 2169.370 322.570 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 320.970 2046.380 322.570 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1552.410 2046.380 1554.010 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 320.970 2043.370 322.570 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1552.410 2043.370 1554.010 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 320.970 2028.380 322.570 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1552.410 2028.380 1554.010 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2582.470 2028.380 2584.070 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 320.970 2025.370 322.570 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1552.410 2025.370 1554.010 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2582.470 2025.370 2584.070 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 320.970 2010.380 322.570 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1552.410 2010.380 1554.010 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2582.470 2010.380 2584.070 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 320.970 2007.370 322.570 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1552.410 2007.370 1554.010 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2582.470 2007.370 2584.070 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 320.970 1992.380 322.570 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1552.410 1992.380 1554.010 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2582.470 1992.380 2584.070 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 320.970 1989.370 322.570 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1552.410 1989.370 1554.010 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2582.470 1989.370 2584.070 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 320.970 1866.380 322.570 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1552.410 1866.380 1554.010 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2582.470 1866.380 2584.070 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 320.970 1863.370 322.570 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1552.410 1863.370 1554.010 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2582.470 1863.370 2584.070 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 320.970 1848.380 322.570 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1552.410 1848.380 1554.010 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2582.470 1848.380 2584.070 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 320.970 1845.370 322.570 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1552.410 1845.370 1554.010 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2582.470 1845.370 2584.070 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 320.970 1830.380 322.570 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1552.410 1830.380 1554.010 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2582.470 1830.380 2584.070 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 320.970 1827.370 322.570 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1552.410 1827.370 1554.010 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2582.470 1827.370 2584.070 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 320.970 1812.380 322.570 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1552.410 1812.380 1554.010 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2582.470 1812.380 2584.070 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 320.970 1809.370 322.570 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1552.410 1809.370 1554.010 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2582.470 1809.370 2584.070 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 320.970 1686.380 322.570 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1552.410 1686.380 1554.010 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2582.470 1686.380 2584.070 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 320.970 1683.370 322.570 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1552.410 1683.370 1554.010 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2582.470 1683.370 2584.070 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 320.970 1668.380 322.570 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1552.410 1668.380 1554.010 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2582.470 1668.380 2584.070 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 320.970 1665.370 322.570 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1552.410 1665.370 1554.010 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2582.470 1665.370 2584.070 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 320.970 1650.380 322.570 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1552.410 1650.380 1554.010 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2582.470 1650.380 2584.070 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 320.970 1647.370 322.570 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1552.410 1647.370 1554.010 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2582.470 1647.370 2584.070 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 320.970 1632.380 322.570 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1552.410 1632.380 1554.010 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2582.470 1632.380 2584.070 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 320.970 1629.370 322.570 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1552.410 1629.370 1554.010 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2582.470 1629.370 2584.070 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1570.970 1470.380 1572.570 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1570.970 1467.370 1572.570 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1570.970 1452.380 1572.570 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1570.970 1449.370 1572.570 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1570.970 1326.380 1572.570 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1570.970 1323.370 1572.570 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1570.970 1308.380 1572.570 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1570.970 1305.370 1572.570 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1570.970 1290.380 1572.570 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1570.970 1287.370 1572.570 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1570.970 1272.380 1572.570 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1570.970 1269.370 1572.570 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1570.970 1146.380 1572.570 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1570.970 1143.370 1572.570 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1570.970 1128.380 1572.570 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1570.970 1125.370 1572.570 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1570.970 1110.380 1572.570 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1570.970 1107.370 1572.570 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1570.970 1092.380 1572.570 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1570.970 1089.370 1572.570 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1570.970 966.380 1572.570 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1570.970 963.370 1572.570 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1570.970 948.380 1572.570 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1570.970 945.370 1572.570 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1570.970 930.380 1572.570 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1570.970 927.370 1572.570 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1570.970 912.380 1572.570 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1570.970 909.370 1572.570 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1570.970 786.380 1572.570 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1570.970 783.370 1572.570 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1570.970 768.380 1572.570 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1570.970 765.370 1572.570 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1570.970 750.380 1572.570 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1570.970 747.370 1572.570 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1570.970 732.380 1572.570 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1570.970 729.370 1572.570 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1570.970 606.380 1572.570 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1570.970 603.370 1572.570 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1570.970 588.380 1572.570 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1570.970 585.370 1572.570 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1570.970 570.380 1572.570 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1570.970 567.370 1572.570 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1570.970 552.380 1572.570 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1570.970 549.370 1572.570 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1570.970 426.380 1572.570 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1570.970 423.370 1572.570 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.040 3251.235 686.300 3252.140 ;
        RECT 1331.040 3251.235 1336.300 3252.140 ;
        RECT 1931.040 3251.235 1936.300 3252.140 ;
        RECT 2581.040 3251.235 2586.300 3252.140 ;
        RECT 681.480 3250.400 686.300 3251.235 ;
        RECT 1331.480 3250.400 1336.300 3251.235 ;
        RECT 1931.480 3250.400 1936.300 3251.235 ;
        RECT 2581.480 3250.400 2586.300 3251.235 ;
        RECT 2581.040 2051.235 2586.300 2052.140 ;
        RECT 2581.480 2050.400 2586.300 2051.235 ;
        RECT 1550.180 1605.000 1555.000 1605.835 ;
        RECT 1550.180 1604.095 1555.440 1605.000 ;
      LAYER via3 ;
        RECT 684.720 3250.440 686.240 3252.050 ;
        RECT 1334.720 3250.440 1336.240 3252.050 ;
        RECT 1934.720 3250.440 1936.240 3252.050 ;
        RECT 2584.720 3250.440 2586.240 3252.050 ;
        RECT 2584.720 2050.440 2586.240 2052.050 ;
        RECT 1550.240 1604.185 1551.760 1605.795 ;
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 292.020 3271.235 295.020 3538.400 ;
        RECT 310.020 3271.235 313.020 3547.800 ;
        RECT 328.020 3271.235 331.020 3557.200 ;
        RECT 454.020 3271.235 457.020 3529.000 ;
        RECT 472.020 3271.235 475.020 3538.400 ;
        RECT 490.020 3271.235 493.020 3547.800 ;
        RECT 508.020 3271.235 511.020 3557.200 ;
        RECT 634.020 3271.235 637.020 3529.000 ;
        RECT 652.020 3271.235 655.020 3538.400 ;
        RECT 670.020 3271.235 673.020 3547.800 ;
        RECT 688.020 3271.235 691.020 3557.200 ;
        RECT 684.690 2804.060 686.310 3252.140 ;
        RECT 814.020 2715.000 817.020 3529.000 ;
        RECT 832.020 2715.000 835.020 3538.400 ;
        RECT 850.020 2715.000 853.020 3547.800 ;
        RECT 868.020 2715.000 871.020 3557.200 ;
        RECT 994.020 3271.235 997.020 3529.000 ;
        RECT 1012.020 3271.235 1015.020 3538.400 ;
        RECT 1030.020 3271.235 1033.020 3547.800 ;
        RECT 1048.020 3271.235 1051.020 3557.200 ;
        RECT 1174.020 3271.235 1177.020 3529.000 ;
        RECT 1192.020 3271.235 1195.020 3538.400 ;
        RECT 1210.020 3271.235 1213.020 3547.800 ;
        RECT 1228.020 3271.235 1231.020 3557.200 ;
        RECT 1334.690 2804.060 1336.310 3252.140 ;
        RECT 1354.020 2715.000 1357.020 3529.000 ;
        RECT 1372.020 2715.000 1375.020 3538.400 ;
        RECT 1390.020 2715.000 1393.020 3547.800 ;
        RECT 1408.020 2715.000 1411.020 3557.200 ;
        RECT 1534.020 3271.235 1537.020 3529.000 ;
        RECT 1552.020 3271.235 1555.020 3538.400 ;
        RECT 1570.020 3271.235 1573.020 3547.800 ;
        RECT 1588.020 3271.235 1591.020 3557.200 ;
        RECT 1714.020 3271.235 1717.020 3529.000 ;
        RECT 1732.020 3271.235 1735.020 3538.400 ;
        RECT 1750.020 3271.235 1753.020 3547.800 ;
        RECT 1768.020 3271.235 1771.020 3557.200 ;
        RECT 1894.020 3271.235 1897.020 3529.000 ;
        RECT 1912.020 3271.235 1915.020 3538.400 ;
        RECT 1930.020 3271.235 1933.020 3547.800 ;
        RECT 1948.020 3271.235 1951.020 3557.200 ;
        RECT 1934.690 2804.060 1936.310 3252.140 ;
        RECT 397.770 1610.640 399.370 2688.240 ;
        RECT 1534.020 2071.235 1537.020 2785.000 ;
        RECT 1552.020 2071.235 1555.020 2785.000 ;
        RECT 1570.020 2071.235 1573.020 2785.000 ;
        RECT 1588.020 2071.235 1591.020 2785.000 ;
        RECT 1714.020 2071.235 1717.020 2785.000 ;
        RECT 1732.020 2071.235 1735.020 2785.000 ;
        RECT 1750.020 2071.235 1753.020 2785.000 ;
        RECT 1768.020 2071.235 1771.020 2785.000 ;
        RECT 1894.020 2071.235 1897.020 2785.000 ;
        RECT 1912.020 2071.235 1915.020 2785.000 ;
        RECT 1930.020 2071.235 1933.020 2785.000 ;
        RECT 1948.020 2071.235 1951.020 2785.000 ;
        RECT 1550.170 1604.095 1551.790 2052.175 ;
        RECT 292.020 -18.720 295.020 1585.000 ;
        RECT 310.020 -28.120 313.020 1585.000 ;
        RECT 328.020 -37.520 331.020 1585.000 ;
        RECT 454.020 -9.320 457.020 1585.000 ;
        RECT 472.020 -18.720 475.020 1585.000 ;
        RECT 490.020 -28.120 493.020 1585.000 ;
        RECT 508.020 -37.520 511.020 1585.000 ;
        RECT 634.020 -9.320 637.020 1585.000 ;
        RECT 652.020 -18.720 655.020 1585.000 ;
        RECT 670.020 -28.120 673.020 1585.000 ;
        RECT 688.020 -37.520 691.020 1585.000 ;
        RECT 814.020 -9.320 817.020 1585.000 ;
        RECT 832.020 -18.720 835.020 1585.000 ;
        RECT 850.020 -28.120 853.020 1585.000 ;
        RECT 868.020 -37.520 871.020 1585.000 ;
        RECT 994.020 -9.320 997.020 1585.000 ;
        RECT 1012.020 -18.720 1015.020 1585.000 ;
        RECT 1030.020 -28.120 1033.020 1585.000 ;
        RECT 1048.020 -37.520 1051.020 1585.000 ;
        RECT 1174.020 -9.320 1177.020 1585.000 ;
        RECT 1192.020 -18.720 1195.020 1585.000 ;
        RECT 1210.020 -28.120 1213.020 1585.000 ;
        RECT 1228.020 -37.520 1231.020 1585.000 ;
        RECT 1354.020 -9.320 1357.020 1585.000 ;
        RECT 1372.020 -18.720 1375.020 1585.000 ;
        RECT 1390.020 -28.120 1393.020 1585.000 ;
        RECT 1408.020 -37.520 1411.020 1585.000 ;
        RECT 1534.020 1515.000 1537.020 1585.000 ;
        RECT 1552.020 1515.000 1555.020 1585.000 ;
        RECT 1570.020 1515.000 1573.020 1585.000 ;
        RECT 1714.020 1515.000 1717.020 1585.000 ;
        RECT 1732.020 1515.000 1735.020 1585.000 ;
        RECT 1750.020 1515.000 1753.020 1585.000 ;
        RECT 1894.020 1515.000 1897.020 1585.000 ;
        RECT 1912.020 1515.000 1915.020 1585.000 ;
        RECT 1930.020 1515.000 1933.020 1585.000 ;
        RECT 2074.020 1515.000 2077.020 3529.000 ;
        RECT 2092.020 1515.000 2095.020 3538.400 ;
        RECT 2110.020 1515.000 2113.020 3547.800 ;
        RECT 2128.020 1515.000 2131.020 3557.200 ;
        RECT 2254.020 3271.235 2257.020 3529.000 ;
        RECT 2272.020 3271.235 2275.020 3538.400 ;
        RECT 2290.020 3271.235 2293.020 3547.800 ;
        RECT 2308.020 3271.235 2311.020 3557.200 ;
        RECT 2434.020 3271.235 2437.020 3529.000 ;
        RECT 2452.020 3271.235 2455.020 3538.400 ;
        RECT 2470.020 3271.235 2473.020 3547.800 ;
        RECT 2488.020 3271.235 2491.020 3557.200 ;
        RECT 2584.690 2804.060 2586.310 3252.140 ;
        RECT 2254.020 2071.235 2257.020 2785.000 ;
        RECT 2272.020 2071.235 2275.020 2785.000 ;
        RECT 2290.020 2071.235 2293.020 2785.000 ;
        RECT 2308.020 2071.235 2311.020 2785.000 ;
        RECT 2434.020 2071.235 2437.020 2785.000 ;
        RECT 2452.020 2071.235 2455.020 2785.000 ;
        RECT 2470.020 2071.235 2473.020 2785.000 ;
        RECT 2488.020 2071.235 2491.020 2785.000 ;
        RECT 2584.690 1604.060 2586.310 2052.140 ;
        RECT 2254.020 1515.000 2257.020 1585.000 ;
        RECT 2272.020 1515.000 2275.020 1585.000 ;
        RECT 2290.020 1515.000 2293.020 1585.000 ;
        RECT 2434.020 1515.000 2437.020 1585.000 ;
        RECT 2452.020 1515.000 2455.020 1585.000 ;
        RECT 2470.020 1515.000 2473.020 1585.000 ;
        RECT 2614.020 1515.000 2617.020 3529.000 ;
        RECT 2632.020 1515.000 2635.020 3538.400 ;
        RECT 2650.020 1515.000 2653.020 3547.800 ;
        RECT 1647.770 410.640 1649.370 1488.240 ;
        RECT 1534.020 -9.320 1537.020 385.000 ;
        RECT 1552.020 -18.720 1555.020 385.000 ;
        RECT 1570.020 -28.120 1573.020 385.000 ;
        RECT 1588.020 -37.520 1591.020 385.000 ;
        RECT 1714.020 -9.320 1717.020 385.000 ;
        RECT 1732.020 -18.720 1735.020 385.000 ;
        RECT 1750.020 -28.120 1753.020 385.000 ;
        RECT 1768.020 -37.520 1771.020 385.000 ;
        RECT 1894.020 -9.320 1897.020 385.000 ;
        RECT 1912.020 -18.720 1915.020 385.000 ;
        RECT 1930.020 -28.120 1933.020 385.000 ;
        RECT 1948.020 -37.520 1951.020 385.000 ;
        RECT 2074.020 -9.320 2077.020 385.000 ;
        RECT 2092.020 -18.720 2095.020 385.000 ;
        RECT 2110.020 -28.120 2113.020 385.000 ;
        RECT 2128.020 -37.520 2131.020 385.000 ;
        RECT 2254.020 -9.320 2257.020 385.000 ;
        RECT 2272.020 -18.720 2275.020 385.000 ;
        RECT 2290.020 -28.120 2293.020 385.000 ;
        RECT 2308.020 -37.520 2311.020 385.000 ;
        RECT 2434.020 -9.320 2437.020 385.000 ;
        RECT 2452.020 -18.720 2455.020 385.000 ;
        RECT 2470.020 -28.120 2473.020 385.000 ;
        RECT 2488.020 -37.520 2491.020 385.000 ;
        RECT 2614.020 -9.320 2617.020 385.000 ;
        RECT 2632.020 -18.720 2635.020 385.000 ;
        RECT 2650.020 -28.120 2653.020 385.000 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 684.910 3215.090 686.090 3216.270 ;
        RECT 684.910 3213.490 686.090 3214.670 ;
        RECT 684.910 3197.090 686.090 3198.270 ;
        RECT 684.910 3195.490 686.090 3196.670 ;
        RECT 684.910 3179.090 686.090 3180.270 ;
        RECT 684.910 3177.490 686.090 3178.670 ;
        RECT 684.910 3161.090 686.090 3162.270 ;
        RECT 684.910 3159.490 686.090 3160.670 ;
        RECT 684.910 3035.090 686.090 3036.270 ;
        RECT 684.910 3033.490 686.090 3034.670 ;
        RECT 684.910 3017.090 686.090 3018.270 ;
        RECT 684.910 3015.490 686.090 3016.670 ;
        RECT 684.910 2999.090 686.090 3000.270 ;
        RECT 684.910 2997.490 686.090 2998.670 ;
        RECT 684.910 2981.090 686.090 2982.270 ;
        RECT 684.910 2979.490 686.090 2980.670 ;
        RECT 684.910 2855.090 686.090 2856.270 ;
        RECT 684.910 2853.490 686.090 2854.670 ;
        RECT 684.910 2837.090 686.090 2838.270 ;
        RECT 684.910 2835.490 686.090 2836.670 ;
        RECT 684.910 2819.090 686.090 2820.270 ;
        RECT 684.910 2817.490 686.090 2818.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 1334.910 3215.090 1336.090 3216.270 ;
        RECT 1334.910 3213.490 1336.090 3214.670 ;
        RECT 1334.910 3197.090 1336.090 3198.270 ;
        RECT 1334.910 3195.490 1336.090 3196.670 ;
        RECT 1334.910 3179.090 1336.090 3180.270 ;
        RECT 1334.910 3177.490 1336.090 3178.670 ;
        RECT 1334.910 3161.090 1336.090 3162.270 ;
        RECT 1334.910 3159.490 1336.090 3160.670 ;
        RECT 1334.910 3035.090 1336.090 3036.270 ;
        RECT 1334.910 3033.490 1336.090 3034.670 ;
        RECT 1334.910 3017.090 1336.090 3018.270 ;
        RECT 1334.910 3015.490 1336.090 3016.670 ;
        RECT 1334.910 2999.090 1336.090 3000.270 ;
        RECT 1334.910 2997.490 1336.090 2998.670 ;
        RECT 1334.910 2981.090 1336.090 2982.270 ;
        RECT 1334.910 2979.490 1336.090 2980.670 ;
        RECT 1334.910 2855.090 1336.090 2856.270 ;
        RECT 1334.910 2853.490 1336.090 2854.670 ;
        RECT 1334.910 2837.090 1336.090 2838.270 ;
        RECT 1334.910 2835.490 1336.090 2836.670 ;
        RECT 1334.910 2819.090 1336.090 2820.270 ;
        RECT 1334.910 2817.490 1336.090 2818.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1934.910 3215.090 1936.090 3216.270 ;
        RECT 1934.910 3213.490 1936.090 3214.670 ;
        RECT 1934.910 3197.090 1936.090 3198.270 ;
        RECT 1934.910 3195.490 1936.090 3196.670 ;
        RECT 1934.910 3179.090 1936.090 3180.270 ;
        RECT 1934.910 3177.490 1936.090 3178.670 ;
        RECT 1934.910 3161.090 1936.090 3162.270 ;
        RECT 1934.910 3159.490 1936.090 3160.670 ;
        RECT 1934.910 3035.090 1936.090 3036.270 ;
        RECT 1934.910 3033.490 1936.090 3034.670 ;
        RECT 1934.910 3017.090 1936.090 3018.270 ;
        RECT 1934.910 3015.490 1936.090 3016.670 ;
        RECT 1934.910 2999.090 1936.090 3000.270 ;
        RECT 1934.910 2997.490 1936.090 2998.670 ;
        RECT 1934.910 2981.090 1936.090 2982.270 ;
        RECT 1934.910 2979.490 1936.090 2980.670 ;
        RECT 1934.910 2855.090 1936.090 2856.270 ;
        RECT 1934.910 2853.490 1936.090 2854.670 ;
        RECT 1934.910 2837.090 1936.090 2838.270 ;
        RECT 1934.910 2835.490 1936.090 2836.670 ;
        RECT 1934.910 2819.090 1936.090 2820.270 ;
        RECT 1934.910 2817.490 1936.090 2818.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 397.980 2675.090 399.160 2676.270 ;
        RECT 397.980 2673.490 399.160 2674.670 ;
        RECT 397.980 2657.090 399.160 2658.270 ;
        RECT 397.980 2655.490 399.160 2656.670 ;
        RECT 397.980 2639.090 399.160 2640.270 ;
        RECT 397.980 2637.490 399.160 2638.670 ;
        RECT 397.980 2621.090 399.160 2622.270 ;
        RECT 397.980 2619.490 399.160 2620.670 ;
        RECT 397.980 2495.090 399.160 2496.270 ;
        RECT 397.980 2493.490 399.160 2494.670 ;
        RECT 397.980 2477.090 399.160 2478.270 ;
        RECT 397.980 2475.490 399.160 2476.670 ;
        RECT 397.980 2459.090 399.160 2460.270 ;
        RECT 397.980 2457.490 399.160 2458.670 ;
        RECT 397.980 2441.090 399.160 2442.270 ;
        RECT 397.980 2439.490 399.160 2440.670 ;
        RECT 397.980 2315.090 399.160 2316.270 ;
        RECT 397.980 2313.490 399.160 2314.670 ;
        RECT 397.980 2297.090 399.160 2298.270 ;
        RECT 397.980 2295.490 399.160 2296.670 ;
        RECT 397.980 2279.090 399.160 2280.270 ;
        RECT 397.980 2277.490 399.160 2278.670 ;
        RECT 397.980 2261.090 399.160 2262.270 ;
        RECT 397.980 2259.490 399.160 2260.670 ;
        RECT 397.980 2135.090 399.160 2136.270 ;
        RECT 397.980 2133.490 399.160 2134.670 ;
        RECT 397.980 2117.090 399.160 2118.270 ;
        RECT 397.980 2115.490 399.160 2116.670 ;
        RECT 397.980 2099.090 399.160 2100.270 ;
        RECT 397.980 2097.490 399.160 2098.670 ;
        RECT 397.980 2081.090 399.160 2082.270 ;
        RECT 397.980 2079.490 399.160 2080.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 397.980 1955.090 399.160 1956.270 ;
        RECT 397.980 1953.490 399.160 1954.670 ;
        RECT 397.980 1937.090 399.160 1938.270 ;
        RECT 397.980 1935.490 399.160 1936.670 ;
        RECT 397.980 1919.090 399.160 1920.270 ;
        RECT 397.980 1917.490 399.160 1918.670 ;
        RECT 397.980 1901.090 399.160 1902.270 ;
        RECT 397.980 1899.490 399.160 1900.670 ;
        RECT 397.980 1775.090 399.160 1776.270 ;
        RECT 397.980 1773.490 399.160 1774.670 ;
        RECT 397.980 1757.090 399.160 1758.270 ;
        RECT 397.980 1755.490 399.160 1756.670 ;
        RECT 397.980 1739.090 399.160 1740.270 ;
        RECT 397.980 1737.490 399.160 1738.670 ;
        RECT 397.980 1721.090 399.160 1722.270 ;
        RECT 397.980 1719.490 399.160 1720.670 ;
        RECT 1550.390 1955.090 1551.570 1956.270 ;
        RECT 1550.390 1953.490 1551.570 1954.670 ;
        RECT 1550.390 1937.090 1551.570 1938.270 ;
        RECT 1550.390 1935.490 1551.570 1936.670 ;
        RECT 1550.390 1919.090 1551.570 1920.270 ;
        RECT 1550.390 1917.490 1551.570 1918.670 ;
        RECT 1550.390 1901.090 1551.570 1902.270 ;
        RECT 1550.390 1899.490 1551.570 1900.670 ;
        RECT 1550.390 1775.090 1551.570 1776.270 ;
        RECT 1550.390 1773.490 1551.570 1774.670 ;
        RECT 1550.390 1757.090 1551.570 1758.270 ;
        RECT 1550.390 1755.490 1551.570 1756.670 ;
        RECT 1550.390 1739.090 1551.570 1740.270 ;
        RECT 1550.390 1737.490 1551.570 1738.670 ;
        RECT 1550.390 1721.090 1551.570 1722.270 ;
        RECT 1550.390 1719.490 1551.570 1720.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2584.910 3215.090 2586.090 3216.270 ;
        RECT 2584.910 3213.490 2586.090 3214.670 ;
        RECT 2584.910 3197.090 2586.090 3198.270 ;
        RECT 2584.910 3195.490 2586.090 3196.670 ;
        RECT 2584.910 3179.090 2586.090 3180.270 ;
        RECT 2584.910 3177.490 2586.090 3178.670 ;
        RECT 2584.910 3161.090 2586.090 3162.270 ;
        RECT 2584.910 3159.490 2586.090 3160.670 ;
        RECT 2584.910 3035.090 2586.090 3036.270 ;
        RECT 2584.910 3033.490 2586.090 3034.670 ;
        RECT 2584.910 3017.090 2586.090 3018.270 ;
        RECT 2584.910 3015.490 2586.090 3016.670 ;
        RECT 2584.910 2999.090 2586.090 3000.270 ;
        RECT 2584.910 2997.490 2586.090 2998.670 ;
        RECT 2584.910 2981.090 2586.090 2982.270 ;
        RECT 2584.910 2979.490 2586.090 2980.670 ;
        RECT 2584.910 2855.090 2586.090 2856.270 ;
        RECT 2584.910 2853.490 2586.090 2854.670 ;
        RECT 2584.910 2837.090 2586.090 2838.270 ;
        RECT 2584.910 2835.490 2586.090 2836.670 ;
        RECT 2584.910 2819.090 2586.090 2820.270 ;
        RECT 2584.910 2817.490 2586.090 2818.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2584.910 1955.090 2586.090 1956.270 ;
        RECT 2584.910 1953.490 2586.090 1954.670 ;
        RECT 2584.910 1937.090 2586.090 1938.270 ;
        RECT 2584.910 1935.490 2586.090 1936.670 ;
        RECT 2584.910 1919.090 2586.090 1920.270 ;
        RECT 2584.910 1917.490 2586.090 1918.670 ;
        RECT 2584.910 1901.090 2586.090 1902.270 ;
        RECT 2584.910 1899.490 2586.090 1900.670 ;
        RECT 2584.910 1775.090 2586.090 1776.270 ;
        RECT 2584.910 1773.490 2586.090 1774.670 ;
        RECT 2584.910 1757.090 2586.090 1758.270 ;
        RECT 2584.910 1755.490 2586.090 1756.670 ;
        RECT 2584.910 1739.090 2586.090 1740.270 ;
        RECT 2584.910 1737.490 2586.090 1738.670 ;
        RECT 2584.910 1721.090 2586.090 1722.270 ;
        RECT 2584.910 1719.490 2586.090 1720.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1647.980 1415.090 1649.160 1416.270 ;
        RECT 1647.980 1413.490 1649.160 1414.670 ;
        RECT 1647.980 1397.090 1649.160 1398.270 ;
        RECT 1647.980 1395.490 1649.160 1396.670 ;
        RECT 1647.980 1379.090 1649.160 1380.270 ;
        RECT 1647.980 1377.490 1649.160 1378.670 ;
        RECT 1647.980 1361.090 1649.160 1362.270 ;
        RECT 1647.980 1359.490 1649.160 1360.670 ;
        RECT 1647.980 1235.090 1649.160 1236.270 ;
        RECT 1647.980 1233.490 1649.160 1234.670 ;
        RECT 1647.980 1217.090 1649.160 1218.270 ;
        RECT 1647.980 1215.490 1649.160 1216.670 ;
        RECT 1647.980 1199.090 1649.160 1200.270 ;
        RECT 1647.980 1197.490 1649.160 1198.670 ;
        RECT 1647.980 1181.090 1649.160 1182.270 ;
        RECT 1647.980 1179.490 1649.160 1180.670 ;
        RECT 1647.980 1055.090 1649.160 1056.270 ;
        RECT 1647.980 1053.490 1649.160 1054.670 ;
        RECT 1647.980 1037.090 1649.160 1038.270 ;
        RECT 1647.980 1035.490 1649.160 1036.670 ;
        RECT 1647.980 1019.090 1649.160 1020.270 ;
        RECT 1647.980 1017.490 1649.160 1018.670 ;
        RECT 1647.980 1001.090 1649.160 1002.270 ;
        RECT 1647.980 999.490 1649.160 1000.670 ;
        RECT 1647.980 875.090 1649.160 876.270 ;
        RECT 1647.980 873.490 1649.160 874.670 ;
        RECT 1647.980 857.090 1649.160 858.270 ;
        RECT 1647.980 855.490 1649.160 856.670 ;
        RECT 1647.980 839.090 1649.160 840.270 ;
        RECT 1647.980 837.490 1649.160 838.670 ;
        RECT 1647.980 821.090 1649.160 822.270 ;
        RECT 1647.980 819.490 1649.160 820.670 ;
        RECT 1647.980 695.090 1649.160 696.270 ;
        RECT 1647.980 693.490 1649.160 694.670 ;
        RECT 1647.980 677.090 1649.160 678.270 ;
        RECT 1647.980 675.490 1649.160 676.670 ;
        RECT 1647.980 659.090 1649.160 660.270 ;
        RECT 1647.980 657.490 1649.160 658.670 ;
        RECT 1647.980 641.090 1649.160 642.270 ;
        RECT 1647.980 639.490 1649.160 640.670 ;
        RECT 1647.980 515.090 1649.160 516.270 ;
        RECT 1647.980 513.490 1649.160 514.670 ;
        RECT 1647.980 497.090 1649.160 498.270 ;
        RECT 1647.980 495.490 1649.160 496.670 ;
        RECT 1647.980 479.090 1649.160 480.270 ;
        RECT 1647.980 477.490 1649.160 478.670 ;
        RECT 1647.980 461.090 1649.160 462.270 ;
        RECT 1647.980 459.490 1649.160 460.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 684.690 3216.380 686.310 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1334.690 3216.380 1336.310 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1934.690 3216.380 1936.310 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2584.690 3216.380 2586.310 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 684.690 3213.370 686.310 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1334.690 3213.370 1336.310 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1934.690 3213.370 1936.310 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2584.690 3213.370 2586.310 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 684.690 3198.380 686.310 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1334.690 3198.380 1336.310 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1934.690 3198.380 1936.310 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2584.690 3198.380 2586.310 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 684.690 3195.370 686.310 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1334.690 3195.370 1336.310 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1934.690 3195.370 1936.310 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2584.690 3195.370 2586.310 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 684.690 3180.380 686.310 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1334.690 3180.380 1336.310 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1934.690 3180.380 1936.310 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2584.690 3180.380 2586.310 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 684.690 3177.370 686.310 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1334.690 3177.370 1336.310 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1934.690 3177.370 1936.310 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2584.690 3177.370 2586.310 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 684.690 3162.380 686.310 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 1334.690 3162.380 1336.310 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1934.690 3162.380 1936.310 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2584.690 3162.380 2586.310 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 684.690 3159.370 686.310 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 1334.690 3159.370 1336.310 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1934.690 3159.370 1936.310 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2584.690 3159.370 2586.310 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 684.690 3036.380 686.310 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1334.690 3036.380 1336.310 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1934.690 3036.380 1936.310 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2584.690 3036.380 2586.310 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 684.690 3033.370 686.310 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1334.690 3033.370 1336.310 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1934.690 3033.370 1936.310 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2584.690 3033.370 2586.310 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 684.690 3018.380 686.310 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1334.690 3018.380 1336.310 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1934.690 3018.380 1936.310 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2584.690 3018.380 2586.310 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 684.690 3015.370 686.310 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1334.690 3015.370 1336.310 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1934.690 3015.370 1936.310 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2584.690 3015.370 2586.310 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 684.690 3000.380 686.310 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1334.690 3000.380 1336.310 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1934.690 3000.380 1936.310 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2584.690 3000.380 2586.310 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 684.690 2997.370 686.310 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1334.690 2997.370 1336.310 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1934.690 2997.370 1936.310 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2584.690 2997.370 2586.310 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 684.690 2982.380 686.310 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 1334.690 2982.380 1336.310 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1934.690 2982.380 1936.310 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2584.690 2982.380 2586.310 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 684.690 2979.370 686.310 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 1334.690 2979.370 1336.310 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1934.690 2979.370 1936.310 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2584.690 2979.370 2586.310 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 684.690 2856.380 686.310 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1334.690 2856.380 1336.310 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1934.690 2856.380 1936.310 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2584.690 2856.380 2586.310 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 684.690 2853.370 686.310 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1334.690 2853.370 1336.310 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1934.690 2853.370 1936.310 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2584.690 2853.370 2586.310 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 684.690 2838.380 686.310 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1334.690 2838.380 1336.310 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1934.690 2838.380 1936.310 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2584.690 2838.380 2586.310 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 684.690 2835.370 686.310 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1334.690 2835.370 1336.310 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1934.690 2835.370 1936.310 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2584.690 2835.370 2586.310 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 684.690 2820.380 686.310 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1334.690 2820.380 1336.310 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1934.690 2820.380 1936.310 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2584.690 2820.380 2586.310 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 684.690 2817.370 686.310 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1334.690 2817.370 1336.310 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1934.690 2817.370 1936.310 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2584.690 2817.370 2586.310 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 397.770 2676.380 399.370 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 397.770 2673.370 399.370 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 397.770 2658.380 399.370 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 397.770 2655.370 399.370 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 397.770 2640.380 399.370 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 397.770 2637.370 399.370 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 397.770 2622.380 399.370 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 397.770 2619.370 399.370 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 397.770 2496.380 399.370 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 397.770 2493.370 399.370 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 397.770 2478.380 399.370 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 397.770 2475.370 399.370 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 397.770 2460.380 399.370 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 397.770 2457.370 399.370 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 397.770 2442.380 399.370 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 397.770 2439.370 399.370 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 397.770 2316.380 399.370 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 397.770 2313.370 399.370 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 397.770 2298.380 399.370 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 397.770 2295.370 399.370 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 397.770 2280.380 399.370 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 397.770 2277.370 399.370 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 397.770 2262.380 399.370 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 397.770 2259.370 399.370 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 397.770 2136.380 399.370 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 397.770 2133.370 399.370 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 397.770 2118.380 399.370 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 397.770 2115.370 399.370 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 397.770 2100.380 399.370 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 397.770 2097.370 399.370 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 397.770 2082.380 399.370 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 397.770 2079.370 399.370 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 397.770 1956.380 399.370 1956.390 ;
        RECT 1550.170 1956.380 1551.790 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2584.690 1956.380 2586.310 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 397.770 1953.370 399.370 1953.380 ;
        RECT 1550.170 1953.370 1551.790 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2584.690 1953.370 2586.310 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 397.770 1938.380 399.370 1938.390 ;
        RECT 1550.170 1938.380 1551.790 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2584.690 1938.380 2586.310 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 397.770 1935.370 399.370 1935.380 ;
        RECT 1550.170 1935.370 1551.790 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2584.690 1935.370 2586.310 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 397.770 1920.380 399.370 1920.390 ;
        RECT 1550.170 1920.380 1551.790 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2584.690 1920.380 2586.310 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 397.770 1917.370 399.370 1917.380 ;
        RECT 1550.170 1917.370 1551.790 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2584.690 1917.370 2586.310 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 397.770 1902.380 399.370 1902.390 ;
        RECT 1550.170 1902.380 1551.790 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2584.690 1902.380 2586.310 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 397.770 1899.370 399.370 1899.380 ;
        RECT 1550.170 1899.370 1551.790 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2584.690 1899.370 2586.310 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 397.770 1776.380 399.370 1776.390 ;
        RECT 1550.170 1776.380 1551.790 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2584.690 1776.380 2586.310 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 397.770 1773.370 399.370 1773.380 ;
        RECT 1550.170 1773.370 1551.790 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2584.690 1773.370 2586.310 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 397.770 1758.380 399.370 1758.390 ;
        RECT 1550.170 1758.380 1551.790 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2584.690 1758.380 2586.310 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 397.770 1755.370 399.370 1755.380 ;
        RECT 1550.170 1755.370 1551.790 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2584.690 1755.370 2586.310 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 397.770 1740.380 399.370 1740.390 ;
        RECT 1550.170 1740.380 1551.790 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2584.690 1740.380 2586.310 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 397.770 1737.370 399.370 1737.380 ;
        RECT 1550.170 1737.370 1551.790 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2584.690 1737.370 2586.310 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 397.770 1722.380 399.370 1722.390 ;
        RECT 1550.170 1722.380 1551.790 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2584.690 1722.380 2586.310 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 397.770 1719.370 399.370 1719.380 ;
        RECT 1550.170 1719.370 1551.790 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2584.690 1719.370 2586.310 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1647.770 1416.380 1649.370 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1647.770 1413.370 1649.370 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1647.770 1398.380 1649.370 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1647.770 1395.370 1649.370 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1647.770 1380.380 1649.370 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1647.770 1377.370 1649.370 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1647.770 1362.380 1649.370 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1647.770 1359.370 1649.370 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1647.770 1236.380 1649.370 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1647.770 1233.370 1649.370 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1647.770 1218.380 1649.370 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1647.770 1215.370 1649.370 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1647.770 1200.380 1649.370 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1647.770 1197.370 1649.370 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1647.770 1182.380 1649.370 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1647.770 1179.370 1649.370 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1647.770 1056.380 1649.370 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1647.770 1053.370 1649.370 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1647.770 1038.380 1649.370 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1647.770 1035.370 1649.370 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1647.770 1020.380 1649.370 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1647.770 1017.370 1649.370 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1647.770 1002.380 1649.370 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1647.770 999.370 1649.370 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1647.770 876.380 1649.370 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1647.770 873.370 1649.370 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1647.770 858.380 1649.370 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1647.770 855.370 1649.370 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1647.770 840.380 1649.370 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1647.770 837.370 1649.370 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1647.770 822.380 1649.370 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1647.770 819.370 1649.370 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1647.770 696.380 1649.370 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1647.770 693.370 1649.370 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1647.770 678.380 1649.370 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1647.770 675.370 1649.370 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1647.770 660.380 1649.370 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1647.770 657.370 1649.370 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1647.770 642.380 1649.370 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1647.770 639.370 1649.370 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1647.770 516.380 1649.370 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1647.770 513.370 1649.370 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1647.770 498.380 1649.370 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1647.770 495.370 1649.370 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1647.770 480.380 1649.370 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1647.770 477.370 1649.370 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1647.770 462.380 1649.370 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1647.770 459.370 1649.370 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 724.645 3252.185 724.815 3253.035 ;
        RECT 772.485 3251.845 772.655 3253.035 ;
        RECT 786.285 3251.845 786.915 3252.015 ;
      LAYER li1 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER li1 ;
        RECT 821.245 3250.825 821.415 3251.675 ;
        RECT 869.085 3250.825 869.255 3252.015 ;
        RECT 884.265 3251.845 884.435 3252.695 ;
        RECT 917.845 3252.525 918.015 3253.375 ;
        RECT 965.685 3252.185 965.855 3253.375 ;
        RECT 1014.445 3252.525 1014.615 3253.375 ;
        RECT 979.485 3252.185 980.115 3252.355 ;
        RECT 1062.285 3252.185 1062.455 3253.375 ;
        RECT 1111.045 3252.525 1111.215 3253.375 ;
        RECT 1076.085 3252.185 1076.715 3252.355 ;
        RECT 1158.885 3252.185 1159.055 3253.375 ;
        RECT 1207.645 3252.525 1207.815 3253.375 ;
        RECT 1172.685 3252.185 1173.315 3252.355 ;
        RECT 1255.485 3252.185 1255.655 3253.375 ;
        RECT 1594.045 3253.205 1594.215 3254.055 ;
        RECT 1559.085 3252.865 1559.715 3253.035 ;
        RECT 1641.885 3252.865 1642.055 3254.055 ;
        RECT 1690.645 3253.205 1690.815 3254.055 ;
        RECT 1655.685 3252.865 1656.315 3253.035 ;
        RECT 1738.485 3252.865 1738.655 3254.055 ;
        RECT 1787.245 3253.205 1787.415 3254.055 ;
        RECT 1752.285 3252.865 1752.915 3253.035 ;
        RECT 1835.085 3252.865 1835.255 3254.055 ;
        RECT 2270.245 3253.205 2270.415 3254.055 ;
        RECT 1849.345 3252.865 1849.975 3253.035 ;
        RECT 2235.285 3252.865 2235.915 3253.035 ;
        RECT 2318.085 3252.865 2318.255 3254.055 ;
        RECT 2366.845 3253.205 2367.015 3254.055 ;
        RECT 2331.885 3252.865 2332.515 3253.035 ;
        RECT 2414.685 3252.865 2414.855 3254.055 ;
        RECT 2463.445 3253.205 2463.615 3254.055 ;
        RECT 2428.485 3252.865 2429.115 3253.035 ;
        RECT 2511.285 3252.865 2511.455 3254.055 ;
        RECT 2525.545 3252.865 2526.175 3253.035 ;
        RECT 1269.285 3252.185 1270.375 3252.355 ;
        RECT 1270.205 3251.505 1270.375 3252.185 ;
        RECT 1304.245 3251.845 1304.415 3252.695 ;
      LAYER li1 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER li1 ;
        RECT 1352.545 3251.165 1352.715 3252.015 ;
        RECT 1400.385 3250.825 1400.555 3252.015 ;
        RECT 1449.145 3251.505 1449.315 3252.355 ;
        RECT 1496.985 3251.505 1497.155 3252.695 ;
      LAYER li1 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER li1 ;
        RECT 1932.145 3251.165 1932.315 3252.355 ;
        RECT 1948.245 3251.165 1948.415 3252.695 ;
        RECT 1980.445 3251.505 1980.615 3252.695 ;
        RECT 2028.745 3250.825 2028.915 3251.675 ;
        RECT 2076.585 3250.825 2076.755 3252.015 ;
        RECT 2125.345 3251.505 2125.515 3252.355 ;
        RECT 2173.185 3251.505 2173.355 3252.695 ;
      LAYER li1 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER li1 ;
        RECT 432.085 2789.445 432.255 2792.335 ;
        RECT 432.545 2788.085 432.715 2791.995 ;
        RECT 484.525 2787.745 484.695 2791.995 ;
        RECT 487.745 2791.825 487.915 2793.355 ;
        RECT 507.065 2789.105 507.235 2793.695 ;
        RECT 507.525 2792.505 507.695 2793.695 ;
        RECT 484.985 2787.745 485.155 2788.935 ;
        RECT 613.785 2788.085 613.955 2789.275 ;
        RECT 625.745 2788.085 625.915 2789.275 ;
        RECT 648.285 2789.105 648.455 2793.695 ;
        RECT 1103.685 2793.185 1103.855 2794.375 ;
        RECT 1111.045 2793.185 1111.215 2794.375 ;
        RECT 1153.825 2791.825 1153.995 2794.035 ;
        RECT 1111.045 2789.785 1111.215 2790.635 ;
        RECT 1158.885 2789.785 1159.055 2790.975 ;
        RECT 647.365 2787.745 649.375 2787.915 ;
        RECT 1462.485 2787.405 1462.655 2793.015 ;
        RECT 1510.325 2792.505 1510.495 2795.055 ;
        RECT 1510.785 2793.185 1510.955 2794.715 ;
        RECT 1511.245 2793.185 1511.415 2794.715 ;
        RECT 1511.245 2792.335 1511.415 2792.675 ;
        RECT 1511.705 2792.505 1511.875 2795.055 ;
        RECT 1512.165 2792.335 1512.335 2794.715 ;
        RECT 1559.085 2792.845 1559.255 2794.715 ;
        RECT 1670.865 2793.185 1671.035 2794.375 ;
        RECT 1729.285 2793.355 1729.455 2793.695 ;
        RECT 1727.905 2793.185 1729.455 2793.355 ;
        RECT 1511.245 2792.165 1512.335 2792.335 ;
        RECT 1723.305 2791.145 1723.475 2792.335 ;
        RECT 1727.905 2792.165 1728.075 2793.185 ;
        RECT 1728.365 2792.165 1728.535 2793.015 ;
        RECT 2114.765 2790.805 2114.935 2793.015 ;
        RECT 2163.065 2790.805 2163.235 2793.015 ;
        RECT 2090.845 2790.465 2091.935 2790.635 ;
        RECT 2090.845 2788.765 2091.015 2790.465 ;
        RECT 2091.305 2790.125 2092.395 2790.295 ;
        RECT 2091.305 2788.425 2091.475 2790.125 ;
        RECT 2092.225 2787.915 2092.395 2788.935 ;
        RECT 2162.605 2788.425 2162.775 2790.295 ;
        RECT 2091.305 2787.745 2092.395 2787.915 ;
        RECT 2163.065 2787.745 2163.235 2788.935 ;
        RECT 2163.525 2788.765 2163.695 2790.635 ;
        RECT 2163.985 2790.465 2164.155 2793.355 ;
        RECT 2208.145 2788.765 2208.315 2793.015 ;
        RECT 2208.605 2788.425 2208.775 2793.355 ;
        RECT 2217.805 2789.785 2217.975 2793.695 ;
        RECT 2235.745 2788.085 2235.915 2792.675 ;
        RECT 2259.205 2792.505 2259.375 2794.035 ;
        RECT 2259.665 2792.845 2259.835 2794.035 ;
        RECT 2261.045 2789.785 2261.215 2793.355 ;
        RECT 2245.405 2787.745 2245.575 2789.615 ;
        RECT 2261.505 2789.105 2261.675 2792.675 ;
        RECT 2266.565 2788.085 2266.735 2793.015 ;
        RECT 2283.585 2787.745 2283.755 2792.335 ;
        RECT 2290.945 2789.275 2291.115 2789.615 ;
        RECT 2290.945 2789.105 2292.035 2789.275 ;
        RECT 2312.565 2787.745 2312.735 2793.355 ;
        RECT 2401.345 2793.185 2401.515 2794.035 ;
        RECT 2344.305 2789.955 2344.475 2792.335 ;
        RECT 2343.385 2789.785 2344.475 2789.955 ;
        RECT 2376.045 2787.745 2376.215 2789.955 ;
        RECT 2376.505 2789.785 2376.675 2792.335 ;
        RECT 2376.965 2792.165 2377.135 2793.015 ;
        RECT 727.405 2712.265 727.575 2718.555 ;
        RECT 761.905 2711.925 762.075 2717.875 ;
        RECT 762.365 2712.605 762.535 2718.555 ;
      LAYER li1 ;
        RECT 305.450 1610.795 1394.270 2688.085 ;
      LAYER li1 ;
        RECT 1410.045 2052.665 1410.215 2061.335 ;
      LAYER li1 ;
        RECT 1555.000 1605.000 1931.480 2051.235 ;
        RECT 2205.000 1605.000 2581.480 2051.235 ;
        RECT 1555.450 410.795 2644.270 1488.085 ;
      LAYER mcon ;
        RECT 1594.045 3253.885 1594.215 3254.055 ;
        RECT 917.845 3253.205 918.015 3253.375 ;
        RECT 724.645 3252.865 724.815 3253.035 ;
        RECT 772.485 3252.865 772.655 3253.035 ;
        RECT 884.265 3252.525 884.435 3252.695 ;
        RECT 965.685 3253.205 965.855 3253.375 ;
        RECT 1014.445 3253.205 1014.615 3253.375 ;
        RECT 1062.285 3253.205 1062.455 3253.375 ;
        RECT 1111.045 3253.205 1111.215 3253.375 ;
        RECT 1158.885 3253.205 1159.055 3253.375 ;
        RECT 1207.645 3253.205 1207.815 3253.375 ;
        RECT 1255.485 3253.205 1255.655 3253.375 ;
        RECT 1641.885 3253.885 1642.055 3254.055 ;
        RECT 1690.645 3253.885 1690.815 3254.055 ;
        RECT 1738.485 3253.885 1738.655 3254.055 ;
        RECT 1787.245 3253.885 1787.415 3254.055 ;
        RECT 1835.085 3253.885 1835.255 3254.055 ;
        RECT 2270.245 3253.885 2270.415 3254.055 ;
        RECT 2318.085 3253.885 2318.255 3254.055 ;
        RECT 2366.845 3253.885 2367.015 3254.055 ;
        RECT 2414.685 3253.885 2414.855 3254.055 ;
        RECT 2463.445 3253.885 2463.615 3254.055 ;
        RECT 2511.285 3253.885 2511.455 3254.055 ;
        RECT 1559.545 3252.865 1559.715 3253.035 ;
        RECT 1656.145 3252.865 1656.315 3253.035 ;
        RECT 1752.745 3252.865 1752.915 3253.035 ;
        RECT 1849.805 3252.865 1849.975 3253.035 ;
        RECT 2235.745 3252.865 2235.915 3253.035 ;
        RECT 2332.345 3252.865 2332.515 3253.035 ;
        RECT 2428.945 3252.865 2429.115 3253.035 ;
        RECT 2526.005 3252.865 2526.175 3253.035 ;
        RECT 1304.245 3252.525 1304.415 3252.695 ;
        RECT 979.945 3252.185 980.115 3252.355 ;
        RECT 1076.545 3252.185 1076.715 3252.355 ;
        RECT 1173.145 3252.185 1173.315 3252.355 ;
        RECT 786.745 3251.845 786.915 3252.015 ;
        RECT 869.085 3251.845 869.255 3252.015 ;
        RECT 821.245 3251.505 821.415 3251.675 ;
        RECT 1496.985 3252.525 1497.155 3252.695 ;
        RECT 1449.145 3252.185 1449.315 3252.355 ;
        RECT 1352.545 3251.845 1352.715 3252.015 ;
        RECT 1400.385 3251.845 1400.555 3252.015 ;
        RECT 1948.245 3252.525 1948.415 3252.695 ;
        RECT 1932.145 3252.185 1932.315 3252.355 ;
        RECT 1980.445 3252.525 1980.615 3252.695 ;
        RECT 2173.185 3252.525 2173.355 3252.695 ;
        RECT 2125.345 3252.185 2125.515 3252.355 ;
        RECT 2076.585 3251.845 2076.755 3252.015 ;
        RECT 2028.745 3251.505 2028.915 3251.675 ;
        RECT 1510.325 2794.885 1510.495 2795.055 ;
        RECT 1103.685 2794.205 1103.855 2794.375 ;
        RECT 507.065 2793.525 507.235 2793.695 ;
        RECT 487.745 2793.185 487.915 2793.355 ;
        RECT 432.085 2792.165 432.255 2792.335 ;
        RECT 432.545 2791.825 432.715 2791.995 ;
        RECT 484.525 2791.825 484.695 2791.995 ;
        RECT 507.525 2793.525 507.695 2793.695 ;
        RECT 648.285 2793.525 648.455 2793.695 ;
        RECT 1111.045 2794.205 1111.215 2794.375 ;
        RECT 1153.825 2793.865 1153.995 2794.035 ;
        RECT 1462.485 2792.845 1462.655 2793.015 ;
        RECT 1158.885 2790.805 1159.055 2790.975 ;
        RECT 1111.045 2790.465 1111.215 2790.635 ;
        RECT 613.785 2789.105 613.955 2789.275 ;
        RECT 484.985 2788.765 485.155 2788.935 ;
        RECT 625.745 2789.105 625.915 2789.275 ;
        RECT 649.205 2787.745 649.375 2787.915 ;
        RECT 1511.705 2794.885 1511.875 2795.055 ;
        RECT 1510.785 2794.545 1510.955 2794.715 ;
        RECT 1511.245 2794.545 1511.415 2794.715 ;
        RECT 1511.245 2792.505 1511.415 2792.675 ;
        RECT 1512.165 2794.545 1512.335 2794.715 ;
        RECT 1559.085 2794.545 1559.255 2794.715 ;
        RECT 1670.865 2794.205 1671.035 2794.375 ;
        RECT 2259.205 2793.865 2259.375 2794.035 ;
        RECT 1729.285 2793.525 1729.455 2793.695 ;
        RECT 2217.805 2793.525 2217.975 2793.695 ;
        RECT 2163.985 2793.185 2164.155 2793.355 ;
        RECT 1723.305 2792.165 1723.475 2792.335 ;
        RECT 1728.365 2792.845 1728.535 2793.015 ;
        RECT 2114.765 2792.845 2114.935 2793.015 ;
        RECT 2163.065 2792.845 2163.235 2793.015 ;
        RECT 2208.605 2793.185 2208.775 2793.355 ;
        RECT 2091.765 2790.465 2091.935 2790.635 ;
        RECT 2163.525 2790.465 2163.695 2790.635 ;
        RECT 2208.145 2792.845 2208.315 2793.015 ;
        RECT 2092.225 2790.125 2092.395 2790.295 ;
        RECT 2162.605 2790.125 2162.775 2790.295 ;
        RECT 2092.225 2788.765 2092.395 2788.935 ;
        RECT 2163.065 2788.765 2163.235 2788.935 ;
        RECT 2259.665 2793.865 2259.835 2794.035 ;
        RECT 2401.345 2793.865 2401.515 2794.035 ;
        RECT 2261.045 2793.185 2261.215 2793.355 ;
        RECT 2235.745 2792.505 2235.915 2792.675 ;
        RECT 2312.565 2793.185 2312.735 2793.355 ;
        RECT 2266.565 2792.845 2266.735 2793.015 ;
        RECT 2261.505 2792.505 2261.675 2792.675 ;
        RECT 2245.405 2789.445 2245.575 2789.615 ;
        RECT 2283.585 2792.165 2283.755 2792.335 ;
        RECT 2290.945 2789.445 2291.115 2789.615 ;
        RECT 2291.865 2789.105 2292.035 2789.275 ;
        RECT 2376.965 2792.845 2377.135 2793.015 ;
        RECT 2344.305 2792.165 2344.475 2792.335 ;
        RECT 2376.505 2792.165 2376.675 2792.335 ;
        RECT 2376.045 2789.785 2376.215 2789.955 ;
        RECT 727.405 2718.385 727.575 2718.555 ;
        RECT 762.365 2718.385 762.535 2718.555 ;
        RECT 761.905 2717.705 762.075 2717.875 ;
        RECT 1410.045 2061.165 1410.215 2061.335 ;
      LAYER met1 ;
        RECT 1324.410 3266.960 1324.730 3267.020 ;
        RECT 1890.670 3266.960 1890.990 3267.020 ;
        RECT 1324.410 3266.820 1890.990 3266.960 ;
        RECT 1324.410 3266.760 1324.730 3266.820 ;
        RECT 1890.670 3266.760 1890.990 3266.820 ;
        RECT 1917.810 3266.960 1918.130 3267.020 ;
        RECT 2542.030 3266.960 2542.350 3267.020 ;
        RECT 1917.810 3266.820 2542.350 3266.960 ;
        RECT 1917.810 3266.760 1918.130 3266.820 ;
        RECT 2542.030 3266.760 2542.350 3266.820 ;
        RECT 1295.890 3264.580 1296.210 3264.640 ;
        RECT 1317.970 3264.580 1318.290 3264.640 ;
        RECT 1324.410 3264.580 1324.730 3264.640 ;
        RECT 1295.890 3264.440 1324.730 3264.580 ;
        RECT 1295.890 3264.380 1296.210 3264.440 ;
        RECT 1317.970 3264.380 1318.290 3264.440 ;
        RECT 1324.410 3264.380 1324.730 3264.440 ;
        RECT 1890.670 3264.580 1890.990 3264.640 ;
        RECT 1917.810 3264.580 1918.130 3264.640 ;
        RECT 1890.670 3264.440 1918.130 3264.580 ;
        RECT 1890.670 3264.380 1890.990 3264.440 ;
        RECT 1917.810 3264.380 1918.130 3264.440 ;
        RECT 2542.030 3264.240 2542.350 3264.300 ;
        RECT 2566.870 3264.240 2567.190 3264.300 ;
        RECT 2542.030 3264.100 2567.190 3264.240 ;
        RECT 2542.030 3264.040 2542.350 3264.100 ;
        RECT 2566.870 3264.040 2567.190 3264.100 ;
        RECT 646.370 3263.900 646.690 3263.960 ;
        RECT 668.450 3263.900 668.770 3263.960 ;
        RECT 696.970 3263.900 697.290 3263.960 ;
        RECT 646.370 3263.760 697.290 3263.900 ;
        RECT 2566.960 3263.900 2567.100 3264.040 ;
        RECT 2594.470 3263.900 2594.790 3263.960 ;
        RECT 2566.960 3263.760 2594.790 3263.900 ;
        RECT 646.370 3263.700 646.690 3263.760 ;
        RECT 668.450 3263.700 668.770 3263.760 ;
        RECT 696.970 3263.700 697.290 3263.760 ;
        RECT 2594.470 3263.700 2594.790 3263.760 ;
        RECT 1593.985 3254.040 1594.275 3254.085 ;
        RECT 1641.825 3254.040 1642.115 3254.085 ;
        RECT 1593.985 3253.900 1642.115 3254.040 ;
        RECT 1593.985 3253.855 1594.275 3253.900 ;
        RECT 1641.825 3253.855 1642.115 3253.900 ;
        RECT 1690.585 3254.040 1690.875 3254.085 ;
        RECT 1738.425 3254.040 1738.715 3254.085 ;
        RECT 1690.585 3253.900 1738.715 3254.040 ;
        RECT 1690.585 3253.855 1690.875 3253.900 ;
        RECT 1738.425 3253.855 1738.715 3253.900 ;
        RECT 1787.185 3254.040 1787.475 3254.085 ;
        RECT 1835.025 3254.040 1835.315 3254.085 ;
        RECT 1787.185 3253.900 1835.315 3254.040 ;
        RECT 1787.185 3253.855 1787.475 3253.900 ;
        RECT 1835.025 3253.855 1835.315 3253.900 ;
        RECT 2270.185 3254.040 2270.475 3254.085 ;
        RECT 2318.025 3254.040 2318.315 3254.085 ;
        RECT 2270.185 3253.900 2318.315 3254.040 ;
        RECT 2270.185 3253.855 2270.475 3253.900 ;
        RECT 2318.025 3253.855 2318.315 3253.900 ;
        RECT 2366.785 3254.040 2367.075 3254.085 ;
        RECT 2414.625 3254.040 2414.915 3254.085 ;
        RECT 2366.785 3253.900 2414.915 3254.040 ;
        RECT 2366.785 3253.855 2367.075 3253.900 ;
        RECT 2414.625 3253.855 2414.915 3253.900 ;
        RECT 2463.385 3254.040 2463.675 3254.085 ;
        RECT 2511.225 3254.040 2511.515 3254.085 ;
        RECT 2463.385 3253.900 2511.515 3254.040 ;
        RECT 2463.385 3253.855 2463.675 3253.900 ;
        RECT 2511.225 3253.855 2511.515 3253.900 ;
        RECT 917.785 3253.360 918.075 3253.405 ;
        RECT 965.625 3253.360 965.915 3253.405 ;
        RECT 917.785 3253.220 965.915 3253.360 ;
        RECT 917.785 3253.175 918.075 3253.220 ;
        RECT 965.625 3253.175 965.915 3253.220 ;
        RECT 1014.385 3253.360 1014.675 3253.405 ;
        RECT 1062.225 3253.360 1062.515 3253.405 ;
        RECT 1014.385 3253.220 1062.515 3253.360 ;
        RECT 1014.385 3253.175 1014.675 3253.220 ;
        RECT 1062.225 3253.175 1062.515 3253.220 ;
        RECT 1110.985 3253.360 1111.275 3253.405 ;
        RECT 1158.825 3253.360 1159.115 3253.405 ;
        RECT 1110.985 3253.220 1159.115 3253.360 ;
        RECT 1110.985 3253.175 1111.275 3253.220 ;
        RECT 1158.825 3253.175 1159.115 3253.220 ;
        RECT 1207.585 3253.360 1207.875 3253.405 ;
        RECT 1255.425 3253.360 1255.715 3253.405 ;
        RECT 1593.985 3253.360 1594.275 3253.405 ;
        RECT 1690.585 3253.360 1690.875 3253.405 ;
        RECT 1787.185 3253.360 1787.475 3253.405 ;
        RECT 2270.185 3253.360 2270.475 3253.405 ;
        RECT 2366.785 3253.360 2367.075 3253.405 ;
        RECT 2463.385 3253.360 2463.675 3253.405 ;
        RECT 1207.585 3253.220 1255.715 3253.360 ;
        RECT 1207.585 3253.175 1207.875 3253.220 ;
        RECT 1255.425 3253.175 1255.715 3253.220 ;
        RECT 1565.540 3253.220 1594.275 3253.360 ;
        RECT 724.585 3253.020 724.875 3253.065 ;
        RECT 772.425 3253.020 772.715 3253.065 ;
        RECT 1559.025 3253.020 1559.315 3253.065 ;
        RECT 724.585 3252.880 772.715 3253.020 ;
        RECT 724.585 3252.835 724.875 3252.880 ;
        RECT 772.425 3252.835 772.715 3252.880 ;
        RECT 1510.800 3252.880 1559.315 3253.020 ;
        RECT 884.205 3252.680 884.495 3252.725 ;
        RECT 917.785 3252.680 918.075 3252.725 ;
        RECT 1014.385 3252.680 1014.675 3252.725 ;
        RECT 1110.985 3252.680 1111.275 3252.725 ;
        RECT 1207.585 3252.680 1207.875 3252.725 ;
        RECT 884.205 3252.540 918.075 3252.680 ;
        RECT 884.205 3252.495 884.495 3252.540 ;
        RECT 917.785 3252.495 918.075 3252.540 ;
        RECT 985.940 3252.540 1014.675 3252.680 ;
        RECT 688.230 3252.340 688.550 3252.400 ;
        RECT 724.585 3252.340 724.875 3252.385 ;
        RECT 688.230 3252.200 724.875 3252.340 ;
        RECT 688.230 3252.140 688.550 3252.200 ;
        RECT 724.585 3252.155 724.875 3252.200 ;
        RECT 965.625 3252.340 965.915 3252.385 ;
        RECT 979.425 3252.340 979.715 3252.385 ;
        RECT 965.625 3252.200 979.715 3252.340 ;
        RECT 965.625 3252.155 965.915 3252.200 ;
        RECT 979.425 3252.155 979.715 3252.200 ;
        RECT 979.885 3252.340 980.175 3252.385 ;
        RECT 985.940 3252.340 986.080 3252.540 ;
        RECT 1014.385 3252.495 1014.675 3252.540 ;
        RECT 1082.540 3252.540 1111.275 3252.680 ;
        RECT 979.885 3252.200 986.080 3252.340 ;
        RECT 1062.225 3252.340 1062.515 3252.385 ;
        RECT 1076.025 3252.340 1076.315 3252.385 ;
        RECT 1062.225 3252.200 1076.315 3252.340 ;
        RECT 979.885 3252.155 980.175 3252.200 ;
        RECT 1062.225 3252.155 1062.515 3252.200 ;
        RECT 1076.025 3252.155 1076.315 3252.200 ;
        RECT 1076.485 3252.340 1076.775 3252.385 ;
        RECT 1082.540 3252.340 1082.680 3252.540 ;
        RECT 1110.985 3252.495 1111.275 3252.540 ;
        RECT 1179.140 3252.540 1207.875 3252.680 ;
        RECT 1076.485 3252.200 1082.680 3252.340 ;
        RECT 1158.825 3252.340 1159.115 3252.385 ;
        RECT 1172.625 3252.340 1172.915 3252.385 ;
        RECT 1158.825 3252.200 1172.915 3252.340 ;
        RECT 1076.485 3252.155 1076.775 3252.200 ;
        RECT 1158.825 3252.155 1159.115 3252.200 ;
        RECT 1172.625 3252.155 1172.915 3252.200 ;
        RECT 1173.085 3252.340 1173.375 3252.385 ;
        RECT 1179.140 3252.340 1179.280 3252.540 ;
        RECT 1207.585 3252.495 1207.875 3252.540 ;
        RECT 1304.185 3252.680 1304.475 3252.725 ;
        RECT 1332.230 3252.680 1332.550 3252.740 ;
        RECT 1304.185 3252.540 1332.550 3252.680 ;
        RECT 1304.185 3252.495 1304.475 3252.540 ;
        RECT 1332.230 3252.480 1332.550 3252.540 ;
        RECT 1496.925 3252.680 1497.215 3252.725 ;
        RECT 1510.800 3252.680 1510.940 3252.880 ;
        RECT 1559.025 3252.835 1559.315 3252.880 ;
        RECT 1559.485 3253.020 1559.775 3253.065 ;
        RECT 1565.540 3253.020 1565.680 3253.220 ;
        RECT 1593.985 3253.175 1594.275 3253.220 ;
        RECT 1662.140 3253.220 1690.875 3253.360 ;
        RECT 1559.485 3252.880 1565.680 3253.020 ;
        RECT 1641.825 3253.020 1642.115 3253.065 ;
        RECT 1655.625 3253.020 1655.915 3253.065 ;
        RECT 1641.825 3252.880 1655.915 3253.020 ;
        RECT 1559.485 3252.835 1559.775 3252.880 ;
        RECT 1641.825 3252.835 1642.115 3252.880 ;
        RECT 1655.625 3252.835 1655.915 3252.880 ;
        RECT 1656.085 3253.020 1656.375 3253.065 ;
        RECT 1662.140 3253.020 1662.280 3253.220 ;
        RECT 1690.585 3253.175 1690.875 3253.220 ;
        RECT 1758.740 3253.220 1787.475 3253.360 ;
        RECT 1656.085 3252.880 1662.280 3253.020 ;
        RECT 1738.425 3253.020 1738.715 3253.065 ;
        RECT 1752.225 3253.020 1752.515 3253.065 ;
        RECT 1738.425 3252.880 1752.515 3253.020 ;
        RECT 1656.085 3252.835 1656.375 3252.880 ;
        RECT 1738.425 3252.835 1738.715 3252.880 ;
        RECT 1752.225 3252.835 1752.515 3252.880 ;
        RECT 1752.685 3253.020 1752.975 3253.065 ;
        RECT 1758.740 3253.020 1758.880 3253.220 ;
        RECT 1787.185 3253.175 1787.475 3253.220 ;
        RECT 2241.740 3253.220 2270.475 3253.360 ;
        RECT 1752.685 3252.880 1758.880 3253.020 ;
        RECT 1835.025 3253.020 1835.315 3253.065 ;
        RECT 1849.285 3253.020 1849.575 3253.065 ;
        RECT 1835.025 3252.880 1849.575 3253.020 ;
        RECT 1752.685 3252.835 1752.975 3252.880 ;
        RECT 1835.025 3252.835 1835.315 3252.880 ;
        RECT 1849.285 3252.835 1849.575 3252.880 ;
        RECT 1849.745 3253.020 1850.035 3253.065 ;
        RECT 2235.225 3253.020 2235.515 3253.065 ;
        RECT 1849.745 3252.880 1883.540 3253.020 ;
        RECT 1849.745 3252.835 1850.035 3252.880 ;
        RECT 1496.925 3252.540 1510.940 3252.680 ;
        RECT 1883.400 3252.680 1883.540 3252.880 ;
        RECT 2187.000 3252.880 2235.515 3253.020 ;
        RECT 1948.185 3252.680 1948.475 3252.725 ;
        RECT 1980.385 3252.680 1980.675 3252.725 ;
        RECT 1883.400 3252.540 1897.340 3252.680 ;
        RECT 1496.925 3252.495 1497.215 3252.540 ;
        RECT 1173.085 3252.200 1179.280 3252.340 ;
        RECT 1255.425 3252.340 1255.715 3252.385 ;
        RECT 1269.225 3252.340 1269.515 3252.385 ;
        RECT 1255.425 3252.200 1269.515 3252.340 ;
        RECT 1173.085 3252.155 1173.375 3252.200 ;
        RECT 1255.425 3252.155 1255.715 3252.200 ;
        RECT 1269.225 3252.155 1269.515 3252.200 ;
        RECT 1414.110 3252.340 1414.430 3252.400 ;
        RECT 1449.085 3252.340 1449.375 3252.385 ;
        RECT 1414.110 3252.200 1449.375 3252.340 ;
        RECT 1897.200 3252.340 1897.340 3252.540 ;
        RECT 1948.185 3252.540 1980.675 3252.680 ;
        RECT 1948.185 3252.495 1948.475 3252.540 ;
        RECT 1980.385 3252.495 1980.675 3252.540 ;
        RECT 2173.125 3252.680 2173.415 3252.725 ;
        RECT 2187.000 3252.680 2187.140 3252.880 ;
        RECT 2235.225 3252.835 2235.515 3252.880 ;
        RECT 2235.685 3253.020 2235.975 3253.065 ;
        RECT 2241.740 3253.020 2241.880 3253.220 ;
        RECT 2270.185 3253.175 2270.475 3253.220 ;
        RECT 2338.340 3253.220 2367.075 3253.360 ;
        RECT 2235.685 3252.880 2241.880 3253.020 ;
        RECT 2318.025 3253.020 2318.315 3253.065 ;
        RECT 2331.825 3253.020 2332.115 3253.065 ;
        RECT 2318.025 3252.880 2332.115 3253.020 ;
        RECT 2235.685 3252.835 2235.975 3252.880 ;
        RECT 2318.025 3252.835 2318.315 3252.880 ;
        RECT 2331.825 3252.835 2332.115 3252.880 ;
        RECT 2332.285 3253.020 2332.575 3253.065 ;
        RECT 2338.340 3253.020 2338.480 3253.220 ;
        RECT 2366.785 3253.175 2367.075 3253.220 ;
        RECT 2434.940 3253.220 2463.675 3253.360 ;
        RECT 2332.285 3252.880 2338.480 3253.020 ;
        RECT 2414.625 3253.020 2414.915 3253.065 ;
        RECT 2428.425 3253.020 2428.715 3253.065 ;
        RECT 2414.625 3252.880 2428.715 3253.020 ;
        RECT 2332.285 3252.835 2332.575 3252.880 ;
        RECT 2414.625 3252.835 2414.915 3252.880 ;
        RECT 2428.425 3252.835 2428.715 3252.880 ;
        RECT 2428.885 3253.020 2429.175 3253.065 ;
        RECT 2434.940 3253.020 2435.080 3253.220 ;
        RECT 2463.385 3253.175 2463.675 3253.220 ;
        RECT 2428.885 3252.880 2435.080 3253.020 ;
        RECT 2511.225 3253.020 2511.515 3253.065 ;
        RECT 2525.485 3253.020 2525.775 3253.065 ;
        RECT 2511.225 3252.880 2525.775 3253.020 ;
        RECT 2428.885 3252.835 2429.175 3252.880 ;
        RECT 2511.225 3252.835 2511.515 3252.880 ;
        RECT 2525.485 3252.835 2525.775 3252.880 ;
        RECT 2525.945 3253.020 2526.235 3253.065 ;
        RECT 2525.945 3252.880 2559.740 3253.020 ;
        RECT 2525.945 3252.835 2526.235 3252.880 ;
        RECT 2173.125 3252.540 2187.140 3252.680 ;
        RECT 2559.600 3252.680 2559.740 3252.880 ;
        RECT 2559.600 3252.540 2573.540 3252.680 ;
        RECT 2173.125 3252.495 2173.415 3252.540 ;
        RECT 1932.085 3252.340 1932.375 3252.385 ;
        RECT 2125.285 3252.340 2125.575 3252.385 ;
        RECT 1897.200 3252.200 1932.375 3252.340 ;
        RECT 1414.110 3252.140 1414.430 3252.200 ;
        RECT 1449.085 3252.155 1449.375 3252.200 ;
        RECT 1932.085 3252.155 1932.375 3252.200 ;
        RECT 2090.400 3252.200 2125.575 3252.340 ;
        RECT 2573.400 3252.340 2573.540 3252.540 ;
        RECT 2582.050 3252.340 2582.370 3252.400 ;
        RECT 2573.400 3252.200 2582.370 3252.340 ;
        RECT 772.425 3252.000 772.715 3252.045 ;
        RECT 786.225 3252.000 786.515 3252.045 ;
        RECT 772.425 3251.860 786.515 3252.000 ;
        RECT 772.425 3251.815 772.715 3251.860 ;
        RECT 786.225 3251.815 786.515 3251.860 ;
        RECT 786.685 3252.000 786.975 3252.045 ;
        RECT 869.025 3252.000 869.315 3252.045 ;
        RECT 884.205 3252.000 884.495 3252.045 ;
        RECT 786.685 3251.860 792.880 3252.000 ;
        RECT 786.685 3251.815 786.975 3251.860 ;
        RECT 792.740 3251.660 792.880 3251.860 ;
        RECT 869.025 3251.860 884.495 3252.000 ;
        RECT 869.025 3251.815 869.315 3251.860 ;
        RECT 884.205 3251.815 884.495 3251.860 ;
        RECT 1304.185 3251.815 1304.475 3252.045 ;
        RECT 1352.485 3252.000 1352.775 3252.045 ;
        RECT 1400.325 3252.000 1400.615 3252.045 ;
        RECT 1352.485 3251.860 1400.615 3252.000 ;
        RECT 1352.485 3251.815 1352.775 3251.860 ;
        RECT 1400.325 3251.815 1400.615 3251.860 ;
        RECT 2076.525 3252.000 2076.815 3252.045 ;
        RECT 2090.400 3252.000 2090.540 3252.200 ;
        RECT 2125.285 3252.155 2125.575 3252.200 ;
        RECT 2582.050 3252.140 2582.370 3252.200 ;
        RECT 2076.525 3251.860 2090.540 3252.000 ;
        RECT 2076.525 3251.815 2076.815 3251.860 ;
        RECT 821.185 3251.660 821.475 3251.705 ;
        RECT 792.740 3251.520 821.475 3251.660 ;
        RECT 821.185 3251.475 821.475 3251.520 ;
        RECT 1270.145 3251.660 1270.435 3251.705 ;
        RECT 1304.260 3251.660 1304.400 3251.815 ;
        RECT 1270.145 3251.520 1304.400 3251.660 ;
        RECT 1449.085 3251.660 1449.375 3251.705 ;
        RECT 1496.925 3251.660 1497.215 3251.705 ;
        RECT 1449.085 3251.520 1497.215 3251.660 ;
        RECT 1270.145 3251.475 1270.435 3251.520 ;
        RECT 1449.085 3251.475 1449.375 3251.520 ;
        RECT 1496.925 3251.475 1497.215 3251.520 ;
        RECT 1980.385 3251.660 1980.675 3251.705 ;
        RECT 2028.685 3251.660 2028.975 3251.705 ;
        RECT 1980.385 3251.520 2028.975 3251.660 ;
        RECT 1980.385 3251.475 1980.675 3251.520 ;
        RECT 2028.685 3251.475 2028.975 3251.520 ;
        RECT 2125.285 3251.660 2125.575 3251.705 ;
        RECT 2173.125 3251.660 2173.415 3251.705 ;
        RECT 2125.285 3251.520 2173.415 3251.660 ;
        RECT 2125.285 3251.475 2125.575 3251.520 ;
        RECT 2173.125 3251.475 2173.415 3251.520 ;
        RECT 1332.230 3251.320 1332.550 3251.380 ;
        RECT 1352.485 3251.320 1352.775 3251.365 ;
      LAYER met1 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met1 ;
        RECT 821.185 3250.980 821.475 3251.025 ;
        RECT 869.025 3250.980 869.315 3251.025 ;
        RECT 821.185 3250.840 869.315 3250.980 ;
        RECT 821.185 3250.795 821.475 3250.840 ;
        RECT 869.025 3250.795 869.315 3250.840 ;
        RECT 696.970 2898.060 697.290 2898.120 ;
        RECT 938.470 2898.060 938.790 2898.120 ;
        RECT 696.970 2897.920 938.790 2898.060 ;
        RECT 696.970 2897.860 697.290 2897.920 ;
        RECT 938.470 2897.860 938.790 2897.920 ;
      LAYER met1 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met1 ;
        RECT 1332.230 3251.180 1352.775 3251.320 ;
        RECT 1932.085 3251.320 1932.375 3251.365 ;
        RECT 1935.750 3251.320 1936.070 3251.380 ;
        RECT 1948.185 3251.320 1948.475 3251.365 ;
        RECT 1332.230 3251.120 1332.550 3251.180 ;
        RECT 1352.485 3251.135 1352.775 3251.180 ;
        RECT 1400.325 3250.980 1400.615 3251.025 ;
        RECT 1411.350 3250.980 1411.670 3251.040 ;
        RECT 1414.110 3250.980 1414.430 3251.040 ;
        RECT 1400.325 3250.840 1414.430 3250.980 ;
        RECT 1400.325 3250.795 1400.615 3250.840 ;
        RECT 1411.350 3250.780 1411.670 3250.840 ;
        RECT 1414.110 3250.780 1414.430 3250.840 ;
        RECT 1473.450 3229.560 1473.770 3229.620 ;
        RECT 1536.930 3229.560 1537.250 3229.620 ;
        RECT 1473.450 3229.420 1537.250 3229.560 ;
        RECT 1473.450 3229.360 1473.770 3229.420 ;
        RECT 1536.930 3229.360 1537.250 3229.420 ;
        RECT 1459.190 3222.420 1459.510 3222.480 ;
        RECT 1535.550 3222.420 1535.870 3222.480 ;
        RECT 1459.190 3222.280 1535.870 3222.420 ;
        RECT 1459.190 3222.220 1459.510 3222.280 ;
        RECT 1535.550 3222.220 1535.870 3222.280 ;
        RECT 1452.290 3215.620 1452.610 3215.680 ;
        RECT 1535.550 3215.620 1535.870 3215.680 ;
        RECT 1452.290 3215.480 1535.870 3215.620 ;
        RECT 1452.290 3215.420 1452.610 3215.480 ;
        RECT 1535.550 3215.420 1535.870 3215.480 ;
        RECT 1438.490 3208.820 1438.810 3208.880 ;
        RECT 1538.310 3208.820 1538.630 3208.880 ;
        RECT 1438.490 3208.680 1538.630 3208.820 ;
        RECT 1438.490 3208.620 1438.810 3208.680 ;
        RECT 1538.310 3208.620 1538.630 3208.680 ;
        RECT 1431.590 3201.680 1431.910 3201.740 ;
        RECT 1538.310 3201.680 1538.630 3201.740 ;
        RECT 1431.590 3201.540 1538.630 3201.680 ;
        RECT 1431.590 3201.480 1431.910 3201.540 ;
        RECT 1538.310 3201.480 1538.630 3201.540 ;
        RECT 1424.690 3194.880 1425.010 3194.940 ;
        RECT 1533.250 3194.880 1533.570 3194.940 ;
        RECT 1424.690 3194.740 1533.570 3194.880 ;
        RECT 1424.690 3194.680 1425.010 3194.740 ;
        RECT 1533.250 3194.680 1533.570 3194.740 ;
        RECT 1472.990 3188.080 1473.310 3188.140 ;
        RECT 1534.170 3188.080 1534.490 3188.140 ;
        RECT 1472.990 3187.940 1534.490 3188.080 ;
        RECT 1472.990 3187.880 1473.310 3187.940 ;
        RECT 1534.170 3187.880 1534.490 3187.940 ;
        RECT 1514.390 2898.400 1514.710 2898.460 ;
        RECT 1534.630 2898.400 1534.950 2898.460 ;
        RECT 1514.390 2898.260 1534.950 2898.400 ;
        RECT 1514.390 2898.200 1514.710 2898.260 ;
        RECT 1534.630 2898.200 1534.950 2898.260 ;
        RECT 1410.890 2894.660 1411.210 2894.720 ;
        RECT 1538.310 2894.660 1538.630 2894.720 ;
        RECT 1410.890 2894.520 1538.630 2894.660 ;
        RECT 1410.890 2894.460 1411.210 2894.520 ;
        RECT 1538.310 2894.460 1538.630 2894.520 ;
      LAYER met1 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met1 ;
        RECT 1932.085 3251.180 1948.475 3251.320 ;
        RECT 1932.085 3251.135 1932.375 3251.180 ;
        RECT 1935.750 3251.120 1936.070 3251.180 ;
        RECT 1948.185 3251.135 1948.475 3251.180 ;
        RECT 2028.685 3250.980 2028.975 3251.025 ;
        RECT 2076.525 3250.980 2076.815 3251.025 ;
        RECT 2028.685 3250.840 2076.815 3250.980 ;
        RECT 2028.685 3250.795 2028.975 3250.840 ;
        RECT 2076.525 3250.795 2076.815 3250.840 ;
        RECT 1945.870 2901.460 1946.190 2901.520 ;
        RECT 2189.210 2901.460 2189.530 2901.520 ;
        RECT 1945.870 2901.320 2189.530 2901.460 ;
        RECT 1945.870 2901.260 1946.190 2901.320 ;
        RECT 2189.210 2901.260 2189.530 2901.320 ;
      LAYER met1 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met1 ;
        RECT 1510.265 2795.040 1510.555 2795.085 ;
        RECT 1511.645 2795.040 1511.935 2795.085 ;
        RECT 1510.265 2794.900 1511.935 2795.040 ;
        RECT 1510.265 2794.855 1510.555 2794.900 ;
        RECT 1511.645 2794.855 1511.935 2794.900 ;
        RECT 1510.725 2794.700 1511.015 2794.745 ;
        RECT 1511.185 2794.700 1511.475 2794.745 ;
        RECT 1510.725 2794.560 1511.475 2794.700 ;
        RECT 1510.725 2794.515 1511.015 2794.560 ;
        RECT 1511.185 2794.515 1511.475 2794.560 ;
        RECT 1512.105 2794.700 1512.395 2794.745 ;
        RECT 1559.025 2794.700 1559.315 2794.745 ;
        RECT 1512.105 2794.560 1559.315 2794.700 ;
        RECT 1512.105 2794.515 1512.395 2794.560 ;
        RECT 1559.025 2794.515 1559.315 2794.560 ;
        RECT 330.810 2794.360 331.130 2794.420 ;
        RECT 1001.030 2794.360 1001.350 2794.420 ;
        RECT 330.810 2794.220 1001.350 2794.360 ;
        RECT 330.810 2794.160 331.130 2794.220 ;
        RECT 1001.030 2794.160 1001.350 2794.220 ;
        RECT 1103.625 2794.360 1103.915 2794.405 ;
        RECT 1110.985 2794.360 1111.275 2794.405 ;
        RECT 1103.625 2794.220 1111.275 2794.360 ;
        RECT 1103.625 2794.175 1103.915 2794.220 ;
        RECT 1110.985 2794.175 1111.275 2794.220 ;
        RECT 1410.430 2794.360 1410.750 2794.420 ;
        RECT 1419.630 2794.360 1419.950 2794.420 ;
        RECT 1587.070 2794.360 1587.390 2794.420 ;
        RECT 1410.430 2794.220 1419.400 2794.360 ;
        RECT 1410.430 2794.160 1410.750 2794.220 ;
        RECT 337.250 2794.020 337.570 2794.080 ;
        RECT 1007.470 2794.020 1007.790 2794.080 ;
        RECT 337.250 2793.880 1007.790 2794.020 ;
        RECT 337.250 2793.820 337.570 2793.880 ;
        RECT 1007.470 2793.820 1007.790 2793.880 ;
        RECT 1100.390 2794.020 1100.710 2794.080 ;
        RECT 1146.850 2794.020 1147.170 2794.080 ;
        RECT 1153.765 2794.020 1154.055 2794.065 ;
        RECT 1100.390 2793.880 1154.055 2794.020 ;
        RECT 1100.390 2793.820 1100.710 2793.880 ;
        RECT 1146.850 2793.820 1147.170 2793.880 ;
        RECT 1153.765 2793.835 1154.055 2793.880 ;
        RECT 397.510 2793.680 397.830 2793.740 ;
        RECT 444.430 2793.680 444.750 2793.740 ;
        RECT 492.730 2793.680 493.050 2793.740 ;
        RECT 507.005 2793.680 507.295 2793.725 ;
        RECT 397.510 2793.540 507.295 2793.680 ;
        RECT 397.510 2793.480 397.830 2793.540 ;
        RECT 444.430 2793.480 444.750 2793.540 ;
        RECT 492.730 2793.480 493.050 2793.540 ;
        RECT 507.005 2793.495 507.295 2793.540 ;
        RECT 507.465 2793.680 507.755 2793.725 ;
        RECT 524.470 2793.680 524.790 2793.740 ;
        RECT 507.465 2793.540 524.790 2793.680 ;
        RECT 507.465 2793.495 507.755 2793.540 ;
        RECT 524.470 2793.480 524.790 2793.540 ;
        RECT 627.510 2793.680 627.830 2793.740 ;
        RECT 648.225 2793.680 648.515 2793.725 ;
        RECT 627.510 2793.540 648.515 2793.680 ;
        RECT 627.510 2793.480 627.830 2793.540 ;
        RECT 648.225 2793.495 648.515 2793.540 ;
        RECT 1042.430 2793.680 1042.750 2793.740 ;
        RECT 1055.770 2793.680 1056.090 2793.740 ;
        RECT 1042.430 2793.540 1056.090 2793.680 ;
        RECT 1042.430 2793.480 1042.750 2793.540 ;
        RECT 1055.770 2793.480 1056.090 2793.540 ;
        RECT 1089.810 2793.680 1090.130 2793.740 ;
        RECT 1129.830 2793.680 1130.150 2793.740 ;
        RECT 1173.070 2793.680 1173.390 2793.740 ;
        RECT 1089.810 2793.540 1173.390 2793.680 ;
        RECT 1089.810 2793.480 1090.130 2793.540 ;
        RECT 1129.830 2793.480 1130.150 2793.540 ;
        RECT 1173.070 2793.480 1173.390 2793.540 ;
        RECT 392.450 2793.340 392.770 2793.400 ;
        RECT 439.370 2793.340 439.690 2793.400 ;
        RECT 485.370 2793.340 485.690 2793.400 ;
        RECT 392.450 2793.200 485.690 2793.340 ;
        RECT 392.450 2793.140 392.770 2793.200 ;
        RECT 439.370 2793.140 439.690 2793.200 ;
        RECT 485.370 2793.140 485.690 2793.200 ;
        RECT 487.685 2793.340 487.975 2793.385 ;
        RECT 510.210 2793.340 510.530 2793.400 ;
        RECT 700.190 2793.340 700.510 2793.400 ;
        RECT 1103.610 2793.340 1103.930 2793.400 ;
        RECT 487.685 2793.200 508.600 2793.340 ;
        RECT 487.685 2793.155 487.975 2793.200 ;
        RECT 386.930 2793.000 387.250 2793.060 ;
        RECT 433.390 2793.000 433.710 2793.060 ;
        RECT 474.330 2793.000 474.650 2793.060 ;
        RECT 508.460 2793.000 508.600 2793.200 ;
        RECT 510.210 2793.200 700.510 2793.340 ;
        RECT 1103.415 2793.200 1103.930 2793.340 ;
        RECT 510.210 2793.140 510.530 2793.200 ;
        RECT 700.190 2793.140 700.510 2793.200 ;
        RECT 1103.610 2793.140 1103.930 2793.200 ;
        RECT 1110.985 2793.340 1111.275 2793.385 ;
        RECT 1136.270 2793.340 1136.590 2793.400 ;
        RECT 1179.970 2793.340 1180.290 2793.400 ;
        RECT 1110.985 2793.200 1180.290 2793.340 ;
        RECT 1419.260 2793.340 1419.400 2794.220 ;
        RECT 1419.630 2794.220 1587.390 2794.360 ;
        RECT 1419.630 2794.160 1419.950 2794.220 ;
        RECT 1587.070 2794.160 1587.390 2794.220 ;
        RECT 1631.690 2794.360 1632.010 2794.420 ;
        RECT 1670.805 2794.360 1671.095 2794.405 ;
        RECT 1631.690 2794.220 1671.095 2794.360 ;
        RECT 1631.690 2794.160 1632.010 2794.220 ;
        RECT 1670.805 2794.175 1671.095 2794.220 ;
        RECT 1671.250 2794.360 1671.570 2794.420 ;
        RECT 1718.170 2794.360 1718.490 2794.420 ;
        RECT 1723.690 2794.360 1724.010 2794.420 ;
        RECT 1671.250 2794.220 1724.010 2794.360 ;
        RECT 1671.250 2794.160 1671.570 2794.220 ;
        RECT 1718.170 2794.160 1718.490 2794.220 ;
        RECT 1723.690 2794.160 1724.010 2794.220 ;
        RECT 1724.150 2794.360 1724.470 2794.420 ;
        RECT 1766.470 2794.360 1766.790 2794.420 ;
        RECT 1724.150 2794.220 1766.790 2794.360 ;
        RECT 1724.150 2794.160 1724.470 2794.220 ;
        RECT 1766.470 2794.160 1766.790 2794.220 ;
        RECT 2231.990 2794.360 2232.310 2794.420 ;
        RECT 2402.650 2794.360 2402.970 2794.420 ;
        RECT 2231.990 2794.220 2402.970 2794.360 ;
        RECT 2231.990 2794.160 2232.310 2794.220 ;
        RECT 2402.650 2794.160 2402.970 2794.220 ;
        RECT 1421.010 2794.020 1421.330 2794.080 ;
        RECT 1601.330 2794.020 1601.650 2794.080 ;
        RECT 1421.010 2793.880 1601.650 2794.020 ;
        RECT 1421.010 2793.820 1421.330 2793.880 ;
        RECT 1601.330 2793.820 1601.650 2793.880 ;
        RECT 1662.510 2794.020 1662.830 2794.080 ;
        RECT 1706.210 2794.020 1706.530 2794.080 ;
        RECT 1752.670 2794.020 1752.990 2794.080 ;
        RECT 1662.510 2793.880 1752.990 2794.020 ;
        RECT 1662.510 2793.820 1662.830 2793.880 ;
        RECT 1706.210 2793.820 1706.530 2793.880 ;
        RECT 1752.670 2793.820 1752.990 2793.880 ;
        RECT 2208.070 2794.020 2208.390 2794.080 ;
        RECT 2259.145 2794.020 2259.435 2794.065 ;
        RECT 2208.070 2793.880 2259.435 2794.020 ;
        RECT 2208.070 2793.820 2208.390 2793.880 ;
        RECT 2259.145 2793.835 2259.435 2793.880 ;
        RECT 2259.605 2794.020 2259.895 2794.065 ;
        RECT 2286.730 2794.020 2287.050 2794.080 ;
        RECT 2332.730 2794.020 2333.050 2794.080 ;
        RECT 2377.350 2794.020 2377.670 2794.080 ;
        RECT 2259.605 2793.880 2377.670 2794.020 ;
        RECT 2259.605 2793.835 2259.895 2793.880 ;
        RECT 2286.730 2793.820 2287.050 2793.880 ;
        RECT 2332.730 2793.820 2333.050 2793.880 ;
        RECT 2377.350 2793.820 2377.670 2793.880 ;
        RECT 2401.285 2794.020 2401.575 2794.065 ;
        RECT 2415.070 2794.020 2415.390 2794.080 ;
        RECT 2401.285 2793.880 2415.390 2794.020 ;
        RECT 2401.285 2793.835 2401.575 2793.880 ;
        RECT 2415.070 2793.820 2415.390 2793.880 ;
        RECT 1420.550 2793.680 1420.870 2793.740 ;
        RECT 1600.870 2793.680 1601.190 2793.740 ;
        RECT 1420.550 2793.540 1601.190 2793.680 ;
        RECT 1420.550 2793.480 1420.870 2793.540 ;
        RECT 1600.870 2793.480 1601.190 2793.540 ;
        RECT 1624.790 2793.680 1625.110 2793.740 ;
        RECT 1671.250 2793.680 1671.570 2793.740 ;
        RECT 1624.790 2793.540 1671.570 2793.680 ;
        RECT 1624.790 2793.480 1625.110 2793.540 ;
        RECT 1671.250 2793.480 1671.570 2793.540 ;
        RECT 1681.370 2793.680 1681.690 2793.740 ;
        RECT 1728.750 2793.680 1729.070 2793.740 ;
        RECT 1681.370 2793.540 1729.070 2793.680 ;
        RECT 1681.370 2793.480 1681.690 2793.540 ;
        RECT 1728.750 2793.480 1729.070 2793.540 ;
        RECT 1729.225 2793.680 1729.515 2793.725 ;
        RECT 1746.690 2793.680 1747.010 2793.740 ;
        RECT 1729.225 2793.540 1747.010 2793.680 ;
        RECT 1729.225 2793.495 1729.515 2793.540 ;
        RECT 1746.690 2793.480 1747.010 2793.540 ;
        RECT 2217.745 2793.680 2218.035 2793.725 ;
        RECT 2268.330 2793.680 2268.650 2793.740 ;
        RECT 2312.950 2793.680 2313.270 2793.740 ;
        RECT 2360.790 2793.680 2361.110 2793.740 ;
        RECT 2408.170 2793.680 2408.490 2793.740 ;
        RECT 2217.745 2793.540 2408.490 2793.680 ;
        RECT 2217.745 2793.495 2218.035 2793.540 ;
        RECT 2268.330 2793.480 2268.650 2793.540 ;
        RECT 2312.950 2793.480 2313.270 2793.540 ;
        RECT 2360.790 2793.480 2361.110 2793.540 ;
        RECT 2408.170 2793.480 2408.490 2793.540 ;
        RECT 1510.725 2793.340 1511.015 2793.385 ;
        RECT 1419.260 2793.200 1511.015 2793.340 ;
        RECT 1110.985 2793.155 1111.275 2793.200 ;
        RECT 1136.270 2793.140 1136.590 2793.200 ;
        RECT 1179.970 2793.140 1180.290 2793.200 ;
        RECT 1510.725 2793.155 1511.015 2793.200 ;
        RECT 1511.185 2793.340 1511.475 2793.385 ;
        RECT 1614.210 2793.340 1614.530 2793.400 ;
        RECT 1511.185 2793.200 1614.530 2793.340 ;
        RECT 1511.185 2793.155 1511.475 2793.200 ;
        RECT 1614.210 2793.140 1614.530 2793.200 ;
        RECT 1638.590 2793.340 1638.910 2793.400 ;
        RECT 1670.805 2793.340 1671.095 2793.385 ;
        RECT 1679.530 2793.340 1679.850 2793.400 ;
        RECT 1724.150 2793.340 1724.470 2793.400 ;
        RECT 1638.590 2793.200 1670.560 2793.340 ;
        RECT 1638.590 2793.140 1638.910 2793.200 ;
        RECT 513.890 2793.000 514.210 2793.060 ;
        RECT 386.930 2792.860 433.710 2793.000 ;
        RECT 386.930 2792.800 387.250 2792.860 ;
        RECT 433.390 2792.800 433.710 2792.860 ;
        RECT 439.000 2792.860 508.140 2793.000 ;
        RECT 508.460 2792.860 514.210 2793.000 ;
        RECT 379.570 2792.660 379.890 2792.720 ;
        RECT 426.950 2792.660 427.270 2792.720 ;
        RECT 439.000 2792.660 439.140 2792.860 ;
        RECT 474.330 2792.800 474.650 2792.860 ;
        RECT 478.470 2792.660 478.790 2792.720 ;
        RECT 507.465 2792.660 507.755 2792.705 ;
        RECT 379.570 2792.520 439.140 2792.660 ;
        RECT 439.460 2792.520 507.755 2792.660 ;
        RECT 508.000 2792.660 508.140 2792.860 ;
        RECT 513.890 2792.800 514.210 2792.860 ;
        RECT 524.010 2793.000 524.330 2793.060 ;
        RECT 720.890 2793.000 721.210 2793.060 ;
        RECT 524.010 2792.860 721.210 2793.000 ;
        RECT 524.010 2792.800 524.330 2792.860 ;
        RECT 720.890 2792.800 721.210 2792.860 ;
        RECT 1062.670 2793.000 1062.990 2793.060 ;
        RECT 1065.430 2793.000 1065.750 2793.060 ;
        RECT 1111.430 2793.000 1111.750 2793.060 ;
        RECT 1159.270 2793.000 1159.590 2793.060 ;
        RECT 1062.670 2792.860 1159.590 2793.000 ;
        RECT 1062.670 2792.800 1062.990 2792.860 ;
        RECT 1065.430 2792.800 1065.750 2792.860 ;
        RECT 1111.430 2792.800 1111.750 2792.860 ;
        RECT 1159.270 2792.800 1159.590 2792.860 ;
        RECT 1462.425 2793.000 1462.715 2793.045 ;
        RECT 1462.870 2793.000 1463.190 2793.060 ;
        RECT 1462.425 2792.860 1463.190 2793.000 ;
        RECT 1462.425 2792.815 1462.715 2792.860 ;
        RECT 1462.870 2792.800 1463.190 2792.860 ;
        RECT 1559.025 2793.000 1559.315 2793.045 ;
        RECT 1617.430 2793.000 1617.750 2793.060 ;
        RECT 1665.730 2793.000 1666.050 2793.060 ;
        RECT 1669.410 2793.000 1669.730 2793.060 ;
        RECT 1559.025 2792.860 1669.730 2793.000 ;
        RECT 1670.420 2793.000 1670.560 2793.200 ;
        RECT 1670.805 2793.200 1724.470 2793.340 ;
        RECT 1670.805 2793.155 1671.095 2793.200 ;
        RECT 1679.530 2793.140 1679.850 2793.200 ;
        RECT 1724.150 2793.140 1724.470 2793.200 ;
        RECT 1681.370 2793.000 1681.690 2793.060 ;
        RECT 1670.420 2792.860 1681.690 2793.000 ;
        RECT 1559.025 2792.815 1559.315 2792.860 ;
        RECT 1617.430 2792.800 1617.750 2792.860 ;
        RECT 1665.730 2792.800 1666.050 2792.860 ;
        RECT 1669.410 2792.800 1669.730 2792.860 ;
        RECT 1681.370 2792.800 1681.690 2792.860 ;
        RECT 1683.670 2793.000 1683.990 2793.060 ;
        RECT 1688.730 2793.000 1689.050 2793.060 ;
        RECT 1728.305 2793.000 1728.595 2793.045 ;
        RECT 1683.670 2792.860 1728.595 2793.000 ;
        RECT 1728.840 2793.000 1728.980 2793.480 ;
        RECT 1732.430 2793.340 1732.750 2793.400 ;
        RECT 1780.270 2793.340 1780.590 2793.400 ;
        RECT 1732.430 2793.200 1780.590 2793.340 ;
        RECT 1732.430 2793.140 1732.750 2793.200 ;
        RECT 1780.270 2793.140 1780.590 2793.200 ;
        RECT 2091.230 2793.340 2091.550 2793.400 ;
        RECT 2163.925 2793.340 2164.215 2793.385 ;
        RECT 2091.230 2793.200 2164.215 2793.340 ;
        RECT 2091.230 2793.140 2091.550 2793.200 ;
        RECT 2163.925 2793.155 2164.215 2793.200 ;
        RECT 2208.545 2793.340 2208.835 2793.385 ;
        RECT 2260.985 2793.340 2261.275 2793.385 ;
        RECT 2208.545 2793.200 2261.275 2793.340 ;
        RECT 2208.545 2793.155 2208.835 2793.200 ;
        RECT 2260.985 2793.155 2261.275 2793.200 ;
        RECT 2270.170 2793.340 2270.490 2793.400 ;
        RECT 2273.390 2793.340 2273.710 2793.400 ;
        RECT 2312.505 2793.340 2312.795 2793.385 ;
        RECT 2326.290 2793.340 2326.610 2793.400 ;
        RECT 2374.130 2793.340 2374.450 2793.400 ;
        RECT 2401.285 2793.340 2401.575 2793.385 ;
        RECT 2270.170 2793.200 2312.795 2793.340 ;
        RECT 2270.170 2793.140 2270.490 2793.200 ;
        RECT 2273.390 2793.140 2273.710 2793.200 ;
        RECT 2312.505 2793.155 2312.795 2793.200 ;
        RECT 2314.420 2793.200 2401.575 2793.340 ;
        RECT 1773.370 2793.000 1773.690 2793.060 ;
        RECT 1728.840 2792.860 1773.690 2793.000 ;
        RECT 1683.670 2792.800 1683.990 2792.860 ;
        RECT 1688.730 2792.800 1689.050 2792.860 ;
        RECT 1728.305 2792.815 1728.595 2792.860 ;
        RECT 1773.370 2792.800 1773.690 2792.860 ;
        RECT 2114.705 2793.000 2114.995 2793.045 ;
        RECT 2163.005 2793.000 2163.295 2793.045 ;
        RECT 2114.705 2792.860 2163.295 2793.000 ;
        RECT 2114.705 2792.815 2114.995 2792.860 ;
        RECT 2163.005 2792.815 2163.295 2792.860 ;
        RECT 2208.085 2793.000 2208.375 2793.045 ;
        RECT 2259.605 2793.000 2259.895 2793.045 ;
        RECT 2208.085 2792.860 2259.895 2793.000 ;
        RECT 2208.085 2792.815 2208.375 2792.860 ;
        RECT 2259.605 2792.815 2259.895 2792.860 ;
        RECT 2266.505 2793.000 2266.795 2793.045 ;
        RECT 2279.830 2793.000 2280.150 2793.060 ;
        RECT 2314.420 2793.000 2314.560 2793.200 ;
        RECT 2326.290 2793.140 2326.610 2793.200 ;
        RECT 2374.130 2793.140 2374.450 2793.200 ;
        RECT 2401.285 2793.155 2401.575 2793.200 ;
        RECT 2266.505 2792.860 2314.560 2793.000 ;
        RECT 2314.790 2793.000 2315.110 2793.060 ;
        RECT 2343.310 2793.000 2343.630 2793.060 ;
        RECT 2376.905 2793.000 2377.195 2793.045 ;
        RECT 2314.790 2792.860 2377.195 2793.000 ;
        RECT 2266.505 2792.815 2266.795 2792.860 ;
        RECT 2279.830 2792.800 2280.150 2792.860 ;
        RECT 2314.790 2792.800 2315.110 2792.860 ;
        RECT 2343.310 2792.800 2343.630 2792.860 ;
        RECT 2376.905 2792.815 2377.195 2792.860 ;
        RECT 2377.350 2793.000 2377.670 2793.060 ;
        RECT 2421.970 2793.000 2422.290 2793.060 ;
        RECT 2377.350 2792.860 2422.290 2793.000 ;
        RECT 2377.350 2792.800 2377.670 2792.860 ;
        RECT 2421.970 2792.800 2422.290 2792.860 ;
        RECT 520.790 2792.660 521.110 2792.720 ;
        RECT 508.000 2792.520 521.110 2792.660 ;
        RECT 379.570 2792.460 379.890 2792.520 ;
        RECT 426.950 2792.460 427.270 2792.520 ;
        RECT 403.950 2792.320 404.270 2792.380 ;
        RECT 432.025 2792.320 432.315 2792.365 ;
        RECT 403.950 2792.180 432.315 2792.320 ;
        RECT 403.950 2792.120 404.270 2792.180 ;
        RECT 432.025 2792.135 432.315 2792.180 ;
        RECT 433.390 2792.320 433.710 2792.380 ;
        RECT 439.460 2792.320 439.600 2792.520 ;
        RECT 478.470 2792.460 478.790 2792.520 ;
        RECT 507.465 2792.475 507.755 2792.520 ;
        RECT 520.790 2792.460 521.110 2792.520 ;
        RECT 542.410 2792.660 542.730 2792.720 ;
        RECT 741.590 2792.660 741.910 2792.720 ;
        RECT 542.410 2792.520 741.910 2792.660 ;
        RECT 542.410 2792.460 542.730 2792.520 ;
        RECT 741.590 2792.460 741.910 2792.520 ;
        RECT 1093.950 2792.660 1094.270 2792.720 ;
        RECT 1140.410 2792.660 1140.730 2792.720 ;
        RECT 1186.870 2792.660 1187.190 2792.720 ;
        RECT 1093.950 2792.520 1187.190 2792.660 ;
        RECT 1093.950 2792.460 1094.270 2792.520 ;
        RECT 1140.410 2792.460 1140.730 2792.520 ;
        RECT 1186.870 2792.460 1187.190 2792.520 ;
        RECT 1420.090 2792.660 1420.410 2792.720 ;
        RECT 1510.265 2792.660 1510.555 2792.705 ;
        RECT 1420.090 2792.520 1510.555 2792.660 ;
        RECT 1420.090 2792.460 1420.410 2792.520 ;
        RECT 1510.265 2792.475 1510.555 2792.520 ;
        RECT 1510.710 2792.660 1511.030 2792.720 ;
        RECT 1511.185 2792.660 1511.475 2792.705 ;
        RECT 1510.710 2792.520 1511.475 2792.660 ;
        RECT 1510.710 2792.460 1511.030 2792.520 ;
        RECT 1511.185 2792.475 1511.475 2792.520 ;
        RECT 1511.645 2792.660 1511.935 2792.705 ;
        RECT 1593.970 2792.660 1594.290 2792.720 ;
        RECT 1511.645 2792.520 1594.290 2792.660 ;
        RECT 1511.645 2792.475 1511.935 2792.520 ;
        RECT 1593.970 2792.460 1594.290 2792.520 ;
        RECT 2235.685 2792.660 2235.975 2792.705 ;
        RECT 2258.670 2792.660 2258.990 2792.720 ;
        RECT 2235.685 2792.520 2258.990 2792.660 ;
        RECT 2235.685 2792.475 2235.975 2792.520 ;
        RECT 2258.670 2792.460 2258.990 2792.520 ;
        RECT 2259.145 2792.660 2259.435 2792.705 ;
        RECT 2261.445 2792.660 2261.735 2792.705 ;
        RECT 2259.145 2792.520 2261.735 2792.660 ;
        RECT 2259.145 2792.475 2259.435 2792.520 ;
        RECT 2261.445 2792.475 2261.735 2792.520 ;
        RECT 2261.890 2792.660 2262.210 2792.720 ;
        RECT 2269.710 2792.660 2270.030 2792.720 ;
        RECT 2308.350 2792.660 2308.670 2792.720 ;
        RECT 2356.650 2792.660 2356.970 2792.720 ;
        RECT 2401.730 2792.660 2402.050 2792.720 ;
        RECT 2261.890 2792.520 2263.960 2792.660 ;
        RECT 2261.890 2792.460 2262.210 2792.520 ;
        RECT 433.390 2792.180 439.600 2792.320 ;
        RECT 449.030 2792.320 449.350 2792.380 ;
        RECT 496.870 2792.320 497.190 2792.380 ;
        RECT 500.550 2792.320 500.870 2792.380 ;
        RECT 449.030 2792.180 500.870 2792.320 ;
        RECT 433.390 2792.120 433.710 2792.180 ;
        RECT 449.030 2792.120 449.350 2792.180 ;
        RECT 496.870 2792.120 497.190 2792.180 ;
        RECT 500.550 2792.120 500.870 2792.180 ;
        RECT 502.850 2792.320 503.170 2792.380 ;
        RECT 700.650 2792.320 700.970 2792.380 ;
        RECT 502.850 2792.180 700.970 2792.320 ;
        RECT 502.850 2792.120 503.170 2792.180 ;
        RECT 700.650 2792.120 700.970 2792.180 ;
        RECT 1409.510 2792.320 1409.830 2792.380 ;
        RECT 1647.790 2792.320 1648.110 2792.380 ;
        RECT 1695.170 2792.320 1695.490 2792.380 ;
        RECT 1723.245 2792.320 1723.535 2792.365 ;
        RECT 1727.845 2792.320 1728.135 2792.365 ;
        RECT 1409.510 2792.180 1723.000 2792.320 ;
        RECT 1409.510 2792.120 1409.830 2792.180 ;
        RECT 1647.790 2792.120 1648.110 2792.180 ;
        RECT 1695.170 2792.120 1695.490 2792.180 ;
        RECT 368.530 2791.980 368.850 2792.040 ;
        RECT 414.530 2791.980 414.850 2792.040 ;
        RECT 432.485 2791.980 432.775 2792.025 ;
        RECT 368.530 2791.840 432.775 2791.980 ;
        RECT 368.530 2791.780 368.850 2791.840 ;
        RECT 414.530 2791.780 414.850 2791.840 ;
        RECT 432.485 2791.795 432.775 2791.840 ;
        RECT 484.465 2791.980 484.755 2792.025 ;
        RECT 487.685 2791.980 487.975 2792.025 ;
        RECT 484.465 2791.840 487.975 2791.980 ;
        RECT 484.465 2791.795 484.755 2791.840 ;
        RECT 487.685 2791.795 487.975 2791.840 ;
        RECT 488.130 2791.980 488.450 2792.040 ;
        RECT 693.290 2791.980 693.610 2792.040 ;
        RECT 488.130 2791.840 693.610 2791.980 ;
        RECT 488.130 2791.780 488.450 2791.840 ;
        RECT 693.290 2791.780 693.610 2791.840 ;
        RECT 1055.770 2791.980 1056.090 2792.040 ;
        RECT 1059.450 2791.980 1059.770 2792.040 ;
        RECT 1105.450 2791.980 1105.770 2792.040 ;
        RECT 1152.370 2791.980 1152.690 2792.040 ;
        RECT 1055.770 2791.840 1152.690 2791.980 ;
        RECT 1055.770 2791.780 1056.090 2791.840 ;
        RECT 1059.450 2791.780 1059.770 2791.840 ;
        RECT 1105.450 2791.780 1105.770 2791.840 ;
        RECT 1152.370 2791.780 1152.690 2791.840 ;
        RECT 1153.765 2791.980 1154.055 2792.025 ;
        RECT 1409.970 2791.980 1410.290 2792.040 ;
        RECT 1642.730 2791.980 1643.050 2792.040 ;
        RECT 1683.670 2791.980 1683.990 2792.040 ;
        RECT 1153.765 2791.840 1166.860 2791.980 ;
        RECT 1153.765 2791.795 1154.055 2791.840 ;
        RECT 407.170 2791.640 407.490 2791.700 ;
        RECT 409.930 2791.640 410.250 2791.700 ;
        RECT 455.470 2791.640 455.790 2791.700 ;
        RECT 407.170 2791.500 455.790 2791.640 ;
        RECT 407.170 2791.440 407.490 2791.500 ;
        RECT 409.930 2791.440 410.250 2791.500 ;
        RECT 455.470 2791.440 455.790 2791.500 ;
        RECT 461.450 2791.640 461.770 2791.700 ;
        RECT 687.310 2791.640 687.630 2791.700 ;
        RECT 461.450 2791.500 687.630 2791.640 ;
        RECT 461.450 2791.440 461.770 2791.500 ;
        RECT 687.310 2791.440 687.630 2791.500 ;
        RECT 1031.850 2791.640 1032.170 2791.700 ;
        RECT 1076.470 2791.640 1076.790 2791.700 ;
        RECT 1119.710 2791.640 1120.030 2791.700 ;
        RECT 1166.170 2791.640 1166.490 2791.700 ;
        RECT 1031.850 2791.500 1166.490 2791.640 ;
        RECT 1166.720 2791.640 1166.860 2791.840 ;
        RECT 1409.970 2791.840 1683.990 2791.980 ;
        RECT 1722.860 2791.980 1723.000 2792.180 ;
        RECT 1723.245 2792.180 1728.135 2792.320 ;
        RECT 1723.245 2792.135 1723.535 2792.180 ;
        RECT 1727.845 2792.135 1728.135 2792.180 ;
        RECT 1728.305 2792.320 1728.595 2792.365 ;
        RECT 1732.430 2792.320 1732.750 2792.380 ;
        RECT 1741.170 2792.320 1741.490 2792.380 ;
        RECT 1787.170 2792.320 1787.490 2792.380 ;
        RECT 1728.305 2792.180 1732.750 2792.320 ;
        RECT 1728.305 2792.135 1728.595 2792.180 ;
        RECT 1732.430 2792.120 1732.750 2792.180 ;
        RECT 1732.980 2792.180 1787.490 2792.320 ;
        RECT 1732.980 2791.980 1733.120 2792.180 ;
        RECT 1741.170 2792.120 1741.490 2792.180 ;
        RECT 1787.170 2792.120 1787.490 2792.180 ;
        RECT 1790.390 2792.320 1790.710 2792.380 ;
        RECT 2263.270 2792.320 2263.590 2792.380 ;
        RECT 1790.390 2792.180 2263.590 2792.320 ;
        RECT 2263.820 2792.320 2263.960 2792.520 ;
        RECT 2269.710 2792.520 2402.050 2792.660 ;
        RECT 2269.710 2792.460 2270.030 2792.520 ;
        RECT 2308.350 2792.460 2308.670 2792.520 ;
        RECT 2356.650 2792.460 2356.970 2792.520 ;
        RECT 2401.730 2792.460 2402.050 2792.520 ;
        RECT 2283.525 2792.320 2283.815 2792.365 ;
        RECT 2263.820 2792.180 2283.815 2792.320 ;
        RECT 1790.390 2792.120 1790.710 2792.180 ;
        RECT 2263.270 2792.120 2263.590 2792.180 ;
        RECT 2283.525 2792.135 2283.815 2792.180 ;
        RECT 2297.310 2792.320 2297.630 2792.380 ;
        RECT 2340.090 2792.320 2340.410 2792.380 ;
        RECT 2343.770 2792.320 2344.090 2792.380 ;
        RECT 2297.310 2792.180 2344.090 2792.320 ;
        RECT 2297.310 2792.120 2297.630 2792.180 ;
        RECT 2340.090 2792.120 2340.410 2792.180 ;
        RECT 2343.770 2792.120 2344.090 2792.180 ;
        RECT 2344.245 2792.320 2344.535 2792.365 ;
        RECT 2350.210 2792.320 2350.530 2792.380 ;
        RECT 2376.445 2792.320 2376.735 2792.365 ;
        RECT 2344.245 2792.180 2376.735 2792.320 ;
        RECT 2344.245 2792.135 2344.535 2792.180 ;
        RECT 2350.210 2792.120 2350.530 2792.180 ;
        RECT 2376.445 2792.135 2376.735 2792.180 ;
        RECT 2376.905 2792.320 2377.195 2792.365 ;
        RECT 2387.930 2792.320 2388.250 2792.380 ;
        RECT 2376.905 2792.180 2388.250 2792.320 ;
        RECT 2376.905 2792.135 2377.195 2792.180 ;
        RECT 2387.930 2792.120 2388.250 2792.180 ;
        RECT 1742.090 2791.980 1742.410 2792.040 ;
        RECT 1722.860 2791.840 1733.120 2791.980 ;
        RECT 1733.440 2791.840 1742.410 2791.980 ;
        RECT 1409.970 2791.780 1410.290 2791.840 ;
        RECT 1642.730 2791.780 1643.050 2791.840 ;
        RECT 1683.670 2791.780 1683.990 2791.840 ;
        RECT 1193.770 2791.640 1194.090 2791.700 ;
        RECT 1166.720 2791.500 1194.090 2791.640 ;
        RECT 1031.850 2791.440 1032.170 2791.500 ;
        RECT 1076.470 2791.440 1076.790 2791.500 ;
        RECT 1119.710 2791.440 1120.030 2791.500 ;
        RECT 1166.170 2791.440 1166.490 2791.500 ;
        RECT 1193.770 2791.440 1194.090 2791.500 ;
        RECT 1409.050 2791.640 1409.370 2791.700 ;
        RECT 1652.390 2791.640 1652.710 2791.700 ;
        RECT 1669.410 2791.640 1669.730 2791.700 ;
        RECT 1712.650 2791.640 1712.970 2791.700 ;
        RECT 1733.440 2791.640 1733.580 2791.840 ;
        RECT 1742.090 2791.780 1742.410 2791.840 ;
        RECT 1797.290 2791.980 1797.610 2792.040 ;
        RECT 2380.570 2791.980 2380.890 2792.040 ;
        RECT 1797.290 2791.840 2380.890 2791.980 ;
        RECT 1797.290 2791.780 1797.610 2791.840 ;
        RECT 2380.570 2791.780 2380.890 2791.840 ;
        RECT 2381.490 2791.980 2381.810 2792.040 ;
        RECT 2385.630 2791.980 2385.950 2792.040 ;
        RECT 2428.870 2791.980 2429.190 2792.040 ;
        RECT 2381.490 2791.840 2429.190 2791.980 ;
        RECT 2381.490 2791.780 2381.810 2791.840 ;
        RECT 2385.630 2791.780 2385.950 2791.840 ;
        RECT 2428.870 2791.780 2429.190 2791.840 ;
        RECT 1409.050 2791.500 1669.180 2791.640 ;
        RECT 1409.050 2791.440 1409.370 2791.500 ;
        RECT 1652.390 2791.440 1652.710 2791.500 ;
        RECT 371.290 2791.300 371.610 2791.360 ;
        RECT 686.850 2791.300 687.170 2791.360 ;
        RECT 371.290 2791.160 687.170 2791.300 ;
        RECT 371.290 2791.100 371.610 2791.160 ;
        RECT 686.850 2791.100 687.170 2791.160 ;
        RECT 1614.210 2791.300 1614.530 2791.360 ;
        RECT 1662.510 2791.300 1662.830 2791.360 ;
        RECT 1614.210 2791.160 1662.830 2791.300 ;
        RECT 1669.040 2791.300 1669.180 2791.500 ;
        RECT 1669.410 2791.500 1733.580 2791.640 ;
        RECT 1746.690 2791.640 1747.010 2791.700 ;
        RECT 1788.550 2791.640 1788.870 2791.700 ;
        RECT 1746.690 2791.500 1788.870 2791.640 ;
        RECT 1669.410 2791.440 1669.730 2791.500 ;
        RECT 1712.650 2791.440 1712.970 2791.500 ;
        RECT 1746.690 2791.440 1747.010 2791.500 ;
        RECT 1788.550 2791.440 1788.870 2791.500 ;
        RECT 1797.750 2791.640 1798.070 2791.700 ;
        RECT 2387.470 2791.640 2387.790 2791.700 ;
        RECT 1797.750 2791.500 2387.790 2791.640 ;
        RECT 1797.750 2791.440 1798.070 2791.500 ;
        RECT 2387.470 2791.440 2387.790 2791.500 ;
        RECT 1699.310 2791.300 1699.630 2791.360 ;
        RECT 1723.245 2791.300 1723.535 2791.345 ;
        RECT 1669.040 2791.160 1723.535 2791.300 ;
        RECT 1614.210 2791.100 1614.530 2791.160 ;
        RECT 1662.510 2791.100 1662.830 2791.160 ;
        RECT 1699.310 2791.100 1699.630 2791.160 ;
        RECT 1723.245 2791.115 1723.535 2791.160 ;
        RECT 1723.690 2791.300 1724.010 2791.360 ;
        RECT 1760.030 2791.300 1760.350 2791.360 ;
        RECT 1723.690 2791.160 1760.350 2791.300 ;
        RECT 1723.690 2791.100 1724.010 2791.160 ;
        RECT 1760.030 2791.100 1760.350 2791.160 ;
        RECT 1790.850 2791.300 1791.170 2791.360 ;
        RECT 2381.030 2791.300 2381.350 2791.360 ;
        RECT 1790.850 2791.160 2381.350 2791.300 ;
        RECT 1790.850 2791.100 1791.170 2791.160 ;
        RECT 2381.030 2791.100 2381.350 2791.160 ;
        RECT 2387.930 2791.300 2388.250 2791.360 ;
        RECT 2391.150 2791.300 2391.470 2791.360 ;
        RECT 2435.770 2791.300 2436.090 2791.360 ;
        RECT 2387.930 2791.160 2436.090 2791.300 ;
        RECT 2387.930 2791.100 2388.250 2791.160 ;
        RECT 2391.150 2791.100 2391.470 2791.160 ;
        RECT 2435.770 2791.100 2436.090 2791.160 ;
        RECT 362.550 2790.960 362.870 2791.020 ;
        RECT 407.170 2790.960 407.490 2791.020 ;
        RECT 362.550 2790.820 407.490 2790.960 ;
        RECT 362.550 2790.760 362.870 2790.820 ;
        RECT 407.170 2790.760 407.490 2790.820 ;
        RECT 419.130 2790.960 419.450 2791.020 ;
        RECT 748.490 2790.960 748.810 2791.020 ;
        RECT 419.130 2790.820 748.810 2790.960 ;
        RECT 419.130 2790.760 419.450 2790.820 ;
        RECT 748.490 2790.760 748.810 2790.820 ;
        RECT 1018.970 2790.960 1019.290 2791.020 ;
        RECT 1062.670 2790.960 1062.990 2791.020 ;
        RECT 1018.970 2790.820 1062.990 2790.960 ;
        RECT 1018.970 2790.760 1019.290 2790.820 ;
        RECT 1062.670 2790.760 1062.990 2790.820 ;
        RECT 1158.825 2790.960 1159.115 2791.005 ;
        RECT 1159.730 2790.960 1160.050 2791.020 ;
        RECT 1158.825 2790.820 1160.050 2790.960 ;
        RECT 1158.825 2790.775 1159.115 2790.820 ;
        RECT 1159.730 2790.760 1160.050 2790.820 ;
        RECT 1417.790 2790.960 1418.110 2791.020 ;
        RECT 2114.705 2790.960 2114.995 2791.005 ;
        RECT 1417.790 2790.820 2114.995 2790.960 ;
        RECT 1417.790 2790.760 1418.110 2790.820 ;
        RECT 2114.705 2790.775 2114.995 2790.820 ;
        RECT 2163.005 2790.960 2163.295 2791.005 ;
        RECT 2237.970 2790.960 2238.290 2791.020 ;
        RECT 2394.370 2790.960 2394.690 2791.020 ;
        RECT 2163.005 2790.820 2238.290 2790.960 ;
        RECT 2163.005 2790.775 2163.295 2790.820 ;
        RECT 2237.970 2790.760 2238.290 2790.820 ;
        RECT 2259.680 2790.820 2394.690 2790.960 ;
        RECT 384.170 2790.620 384.490 2790.680 ;
        RECT 727.790 2790.620 728.110 2790.680 ;
        RECT 384.170 2790.480 728.110 2790.620 ;
        RECT 384.170 2790.420 384.490 2790.480 ;
        RECT 727.790 2790.420 728.110 2790.480 ;
        RECT 1069.570 2790.620 1069.890 2790.680 ;
        RECT 1110.985 2790.620 1111.275 2790.665 ;
        RECT 1069.570 2790.480 1111.275 2790.620 ;
        RECT 1069.570 2790.420 1069.890 2790.480 ;
        RECT 1110.985 2790.435 1111.275 2790.480 ;
        RECT 1418.710 2790.620 1419.030 2790.680 ;
        RECT 2091.230 2790.620 2091.550 2790.680 ;
        RECT 1418.710 2790.480 2091.550 2790.620 ;
        RECT 1418.710 2790.420 1419.030 2790.480 ;
        RECT 2091.230 2790.420 2091.550 2790.480 ;
        RECT 2091.705 2790.620 2091.995 2790.665 ;
        RECT 2163.465 2790.620 2163.755 2790.665 ;
        RECT 2091.705 2790.480 2163.755 2790.620 ;
        RECT 2091.705 2790.435 2091.995 2790.480 ;
        RECT 2163.465 2790.435 2163.755 2790.480 ;
        RECT 2163.925 2790.620 2164.215 2790.665 ;
        RECT 2249.470 2790.620 2249.790 2790.680 ;
        RECT 2163.925 2790.480 2249.790 2790.620 ;
        RECT 2163.925 2790.435 2164.215 2790.480 ;
        RECT 2249.470 2790.420 2249.790 2790.480 ;
        RECT 406.250 2790.280 406.570 2790.340 ;
        RECT 762.750 2790.280 763.070 2790.340 ;
        RECT 406.250 2790.140 763.070 2790.280 ;
        RECT 406.250 2790.080 406.570 2790.140 ;
        RECT 762.750 2790.080 763.070 2790.140 ;
        RECT 1419.170 2790.280 1419.490 2790.340 ;
        RECT 2090.770 2790.280 2091.090 2790.340 ;
        RECT 1419.170 2790.140 2091.090 2790.280 ;
        RECT 1419.170 2790.080 1419.490 2790.140 ;
        RECT 2090.770 2790.080 2091.090 2790.140 ;
        RECT 2092.165 2790.280 2092.455 2790.325 ;
        RECT 2162.545 2790.280 2162.835 2790.325 ;
        RECT 2092.165 2790.140 2162.835 2790.280 ;
        RECT 2092.165 2790.095 2092.455 2790.140 ;
        RECT 2162.545 2790.095 2162.835 2790.140 ;
        RECT 2162.990 2790.280 2163.310 2790.340 ;
        RECT 2256.370 2790.280 2256.690 2790.340 ;
        RECT 2162.990 2790.140 2256.690 2790.280 ;
        RECT 2162.990 2790.080 2163.310 2790.140 ;
        RECT 2256.370 2790.080 2256.690 2790.140 ;
        RECT 396.590 2789.940 396.910 2790.000 ;
        RECT 762.290 2789.940 762.610 2790.000 ;
        RECT 396.590 2789.800 762.610 2789.940 ;
        RECT 396.590 2789.740 396.910 2789.800 ;
        RECT 762.290 2789.740 762.610 2789.800 ;
        RECT 1110.985 2789.940 1111.275 2789.985 ;
        RECT 1117.870 2789.940 1118.190 2790.000 ;
        RECT 1158.825 2789.940 1159.115 2789.985 ;
        RECT 1110.985 2789.800 1159.115 2789.940 ;
        RECT 1110.985 2789.755 1111.275 2789.800 ;
        RECT 1117.870 2789.740 1118.190 2789.800 ;
        RECT 1158.825 2789.755 1159.115 2789.800 ;
        RECT 1411.350 2789.940 1411.670 2790.000 ;
        RECT 2217.745 2789.940 2218.035 2789.985 ;
        RECT 1411.350 2789.800 2218.035 2789.940 ;
        RECT 1411.350 2789.740 1411.670 2789.800 ;
        RECT 2217.745 2789.755 2218.035 2789.800 ;
        RECT 2218.190 2789.940 2218.510 2790.000 ;
        RECT 2259.680 2789.940 2259.820 2790.820 ;
        RECT 2394.370 2790.760 2394.690 2790.820 ;
        RECT 2394.830 2790.960 2395.150 2791.020 ;
        RECT 2442.670 2790.960 2442.990 2791.020 ;
        RECT 2394.830 2790.820 2442.990 2790.960 ;
        RECT 2394.830 2790.760 2395.150 2790.820 ;
        RECT 2442.670 2790.760 2442.990 2790.820 ;
        RECT 2415.070 2790.620 2415.390 2790.680 ;
        RECT 2218.190 2789.800 2259.820 2789.940 ;
        RECT 2260.140 2790.480 2415.390 2790.620 ;
        RECT 2218.190 2789.740 2218.510 2789.800 ;
        RECT 374.970 2789.600 375.290 2789.660 ;
        RECT 420.970 2789.600 421.290 2789.660 ;
        RECT 374.970 2789.460 421.290 2789.600 ;
        RECT 374.970 2789.400 375.290 2789.460 ;
        RECT 420.970 2789.400 421.290 2789.460 ;
        RECT 432.025 2789.600 432.315 2789.645 ;
        RECT 449.030 2789.600 449.350 2789.660 ;
        RECT 432.025 2789.460 449.350 2789.600 ;
        RECT 432.025 2789.415 432.315 2789.460 ;
        RECT 449.030 2789.400 449.350 2789.460 ;
        RECT 468.810 2789.600 469.130 2789.660 ;
        RECT 686.390 2789.600 686.710 2789.660 ;
        RECT 468.810 2789.460 686.710 2789.600 ;
        RECT 468.810 2789.400 469.130 2789.460 ;
        RECT 686.390 2789.400 686.710 2789.460 ;
        RECT 1010.690 2789.600 1011.010 2789.660 ;
        RECT 1055.770 2789.600 1056.090 2789.660 ;
        RECT 1010.690 2789.460 1056.090 2789.600 ;
        RECT 1010.690 2789.400 1011.010 2789.460 ;
        RECT 1055.770 2789.400 1056.090 2789.460 ;
        RECT 1411.810 2789.600 1412.130 2789.660 ;
        RECT 2245.345 2789.600 2245.635 2789.645 ;
        RECT 1411.810 2789.460 2245.635 2789.600 ;
        RECT 1411.810 2789.400 1412.130 2789.460 ;
        RECT 2245.345 2789.415 2245.635 2789.460 ;
        RECT 2245.790 2789.600 2246.110 2789.660 ;
        RECT 2260.140 2789.600 2260.280 2790.480 ;
        RECT 2415.070 2790.420 2415.390 2790.480 ;
        RECT 2408.170 2790.280 2408.490 2790.340 ;
        RECT 2245.790 2789.460 2260.280 2789.600 ;
        RECT 2260.600 2790.140 2408.490 2790.280 ;
        RECT 2245.790 2789.400 2246.110 2789.460 ;
        RECT 507.005 2789.260 507.295 2789.305 ;
        RECT 538.270 2789.260 538.590 2789.320 ;
        RECT 507.005 2789.120 538.590 2789.260 ;
        RECT 507.005 2789.075 507.295 2789.120 ;
        RECT 538.270 2789.060 538.590 2789.120 ;
        RECT 613.725 2789.260 614.015 2789.305 ;
        RECT 625.685 2789.260 625.975 2789.305 ;
        RECT 613.725 2789.120 625.975 2789.260 ;
        RECT 613.725 2789.075 614.015 2789.120 ;
        RECT 625.685 2789.075 625.975 2789.120 ;
        RECT 648.225 2789.260 648.515 2789.305 ;
        RECT 1042.430 2789.260 1042.750 2789.320 ;
        RECT 648.225 2789.120 1042.750 2789.260 ;
        RECT 648.225 2789.075 648.515 2789.120 ;
        RECT 1042.430 2789.060 1042.750 2789.120 ;
        RECT 1412.270 2789.260 1412.590 2789.320 ;
        RECT 2238.890 2789.260 2239.210 2789.320 ;
        RECT 2260.600 2789.260 2260.740 2790.140 ;
        RECT 2408.170 2790.080 2408.490 2790.140 ;
        RECT 2260.985 2789.940 2261.275 2789.985 ;
        RECT 2291.330 2789.940 2291.650 2790.000 ;
        RECT 2297.310 2789.940 2297.630 2790.000 ;
        RECT 2260.985 2789.800 2297.630 2789.940 ;
        RECT 2260.985 2789.755 2261.275 2789.800 ;
        RECT 2291.330 2789.740 2291.650 2789.800 ;
        RECT 2297.310 2789.740 2297.630 2789.800 ;
        RECT 2304.210 2789.940 2304.530 2790.000 ;
        RECT 2343.325 2789.940 2343.615 2789.985 ;
        RECT 2304.210 2789.800 2343.615 2789.940 ;
        RECT 2304.210 2789.740 2304.530 2789.800 ;
        RECT 2343.325 2789.755 2343.615 2789.800 ;
        RECT 2343.770 2789.940 2344.090 2790.000 ;
        RECT 2375.985 2789.940 2376.275 2789.985 ;
        RECT 2343.770 2789.800 2376.275 2789.940 ;
        RECT 2343.770 2789.740 2344.090 2789.800 ;
        RECT 2375.985 2789.755 2376.275 2789.800 ;
        RECT 2376.445 2789.940 2376.735 2789.985 ;
        RECT 2394.830 2789.940 2395.150 2790.000 ;
        RECT 2376.445 2789.800 2395.150 2789.940 ;
        RECT 2376.445 2789.755 2376.735 2789.800 ;
        RECT 2394.830 2789.740 2395.150 2789.800 ;
        RECT 2273.390 2789.600 2273.710 2789.660 ;
        RECT 2290.885 2789.600 2291.175 2789.645 ;
        RECT 2304.300 2789.600 2304.440 2789.740 ;
        RECT 2273.390 2789.460 2291.175 2789.600 ;
        RECT 2273.390 2789.400 2273.710 2789.460 ;
        RECT 2290.885 2789.415 2291.175 2789.460 ;
        RECT 2291.420 2789.460 2304.440 2789.600 ;
        RECT 2321.690 2789.600 2322.010 2789.660 ;
        RECT 2442.670 2789.600 2442.990 2789.660 ;
        RECT 2321.690 2789.460 2442.990 2789.600 ;
        RECT 1412.270 2789.120 2238.200 2789.260 ;
        RECT 1412.270 2789.060 1412.590 2789.120 ;
        RECT 446.730 2788.920 447.050 2788.980 ;
        RECT 484.925 2788.920 485.215 2788.965 ;
        RECT 446.730 2788.780 485.215 2788.920 ;
        RECT 446.730 2788.720 447.050 2788.780 ;
        RECT 484.925 2788.735 485.215 2788.780 ;
        RECT 485.370 2788.920 485.690 2788.980 ;
        RECT 531.370 2788.920 531.690 2788.980 ;
        RECT 485.370 2788.780 531.690 2788.920 ;
        RECT 485.370 2788.720 485.690 2788.780 ;
        RECT 531.370 2788.720 531.690 2788.780 ;
        RECT 606.810 2788.920 607.130 2788.980 ;
        RECT 1031.850 2788.920 1032.170 2788.980 ;
        RECT 606.810 2788.780 1032.170 2788.920 ;
        RECT 606.810 2788.720 607.130 2788.780 ;
        RECT 1031.850 2788.720 1032.170 2788.780 ;
        RECT 1038.290 2788.920 1038.610 2788.980 ;
        RECT 1089.810 2788.920 1090.130 2788.980 ;
        RECT 1038.290 2788.780 1090.130 2788.920 ;
        RECT 1038.290 2788.720 1038.610 2788.780 ;
        RECT 1089.810 2788.720 1090.130 2788.780 ;
        RECT 1412.730 2788.920 1413.050 2788.980 ;
        RECT 2090.785 2788.920 2091.075 2788.965 ;
        RECT 1412.730 2788.780 2091.075 2788.920 ;
        RECT 1412.730 2788.720 1413.050 2788.780 ;
        RECT 2090.785 2788.735 2091.075 2788.780 ;
        RECT 2092.165 2788.920 2092.455 2788.965 ;
        RECT 2163.005 2788.920 2163.295 2788.965 ;
        RECT 2092.165 2788.780 2163.295 2788.920 ;
        RECT 2092.165 2788.735 2092.455 2788.780 ;
        RECT 2163.005 2788.735 2163.295 2788.780 ;
        RECT 2163.465 2788.920 2163.755 2788.965 ;
        RECT 2208.085 2788.920 2208.375 2788.965 ;
        RECT 2163.465 2788.780 2208.375 2788.920 ;
        RECT 2163.465 2788.735 2163.755 2788.780 ;
        RECT 2208.085 2788.735 2208.375 2788.780 ;
        RECT 455.470 2788.580 455.790 2788.640 ;
        RECT 500.090 2788.580 500.410 2788.640 ;
        RECT 455.470 2788.440 500.410 2788.580 ;
        RECT 455.470 2788.380 455.790 2788.440 ;
        RECT 500.090 2788.380 500.410 2788.440 ;
        RECT 500.550 2788.580 500.870 2788.640 ;
        RECT 541.490 2788.580 541.810 2788.640 ;
        RECT 500.550 2788.440 541.810 2788.580 ;
        RECT 500.550 2788.380 500.870 2788.440 ;
        RECT 541.490 2788.380 541.810 2788.440 ;
        RECT 586.110 2788.580 586.430 2788.640 ;
        RECT 1018.970 2788.580 1019.290 2788.640 ;
        RECT 586.110 2788.440 1019.290 2788.580 ;
        RECT 586.110 2788.380 586.430 2788.440 ;
        RECT 1018.970 2788.380 1019.290 2788.440 ;
        RECT 1024.490 2788.580 1024.810 2788.640 ;
        RECT 1069.570 2788.580 1069.890 2788.640 ;
        RECT 1024.490 2788.440 1069.890 2788.580 ;
        RECT 1024.490 2788.380 1024.810 2788.440 ;
        RECT 1069.570 2788.380 1069.890 2788.440 ;
        RECT 1413.190 2788.580 1413.510 2788.640 ;
        RECT 2091.245 2788.580 2091.535 2788.625 ;
        RECT 1413.190 2788.440 2091.535 2788.580 ;
        RECT 1413.190 2788.380 1413.510 2788.440 ;
        RECT 2091.245 2788.395 2091.535 2788.440 ;
        RECT 2162.545 2788.580 2162.835 2788.625 ;
        RECT 2208.545 2788.580 2208.835 2788.625 ;
        RECT 2162.545 2788.440 2208.835 2788.580 ;
        RECT 2162.545 2788.395 2162.835 2788.440 ;
        RECT 2208.545 2788.395 2208.835 2788.440 ;
        RECT 432.485 2788.240 432.775 2788.285 ;
        RECT 462.370 2788.240 462.690 2788.300 ;
        RECT 504.230 2788.240 504.550 2788.300 ;
        RECT 613.725 2788.240 614.015 2788.285 ;
        RECT 432.485 2788.100 504.550 2788.240 ;
        RECT 432.485 2788.055 432.775 2788.100 ;
        RECT 462.370 2788.040 462.690 2788.100 ;
        RECT 504.230 2788.040 504.550 2788.100 ;
        RECT 513.060 2788.100 614.015 2788.240 ;
        RECT 420.970 2787.900 421.290 2787.960 ;
        RECT 467.890 2787.900 468.210 2787.960 ;
        RECT 484.465 2787.900 484.755 2787.945 ;
        RECT 420.970 2787.760 484.755 2787.900 ;
        RECT 420.970 2787.700 421.290 2787.760 ;
        RECT 467.890 2787.700 468.210 2787.760 ;
        RECT 484.465 2787.715 484.755 2787.760 ;
        RECT 484.925 2787.900 485.215 2787.945 ;
        RECT 513.060 2787.900 513.200 2788.100 ;
        RECT 613.725 2788.055 614.015 2788.100 ;
        RECT 625.685 2788.240 625.975 2788.285 ;
        RECT 648.670 2788.240 648.990 2788.300 ;
        RECT 1052.550 2788.240 1052.870 2788.300 ;
        RECT 1100.390 2788.240 1100.710 2788.300 ;
        RECT 625.685 2788.100 647.980 2788.240 ;
        RECT 625.685 2788.055 625.975 2788.100 ;
        RECT 484.925 2787.760 513.200 2787.900 ;
        RECT 537.350 2787.900 537.670 2787.960 ;
        RECT 647.305 2787.900 647.595 2787.945 ;
        RECT 537.350 2787.760 647.595 2787.900 ;
        RECT 484.925 2787.715 485.215 2787.760 ;
        RECT 537.350 2787.700 537.670 2787.760 ;
        RECT 647.305 2787.715 647.595 2787.760 ;
        RECT 647.840 2787.560 647.980 2788.100 ;
        RECT 648.670 2788.100 1100.710 2788.240 ;
        RECT 648.670 2788.040 648.990 2788.100 ;
        RECT 1052.550 2788.040 1052.870 2788.100 ;
        RECT 1100.390 2788.040 1100.710 2788.100 ;
        RECT 1413.650 2788.240 1413.970 2788.300 ;
        RECT 2235.685 2788.240 2235.975 2788.285 ;
        RECT 1413.650 2788.100 2235.975 2788.240 ;
        RECT 2238.060 2788.240 2238.200 2789.120 ;
        RECT 2238.890 2789.120 2260.740 2789.260 ;
        RECT 2261.445 2789.260 2261.735 2789.305 ;
        RECT 2291.420 2789.260 2291.560 2789.460 ;
        RECT 2321.690 2789.400 2322.010 2789.460 ;
        RECT 2442.670 2789.400 2442.990 2789.460 ;
        RECT 2261.445 2789.120 2291.560 2789.260 ;
        RECT 2291.805 2789.260 2292.095 2789.305 ;
        RECT 2435.770 2789.260 2436.090 2789.320 ;
        RECT 2291.805 2789.120 2436.090 2789.260 ;
        RECT 2238.890 2789.060 2239.210 2789.120 ;
        RECT 2261.445 2789.075 2261.735 2789.120 ;
        RECT 2291.805 2789.075 2292.095 2789.120 ;
        RECT 2435.770 2789.060 2436.090 2789.120 ;
        RECT 2259.590 2788.920 2259.910 2788.980 ;
        RECT 2421.970 2788.920 2422.290 2788.980 ;
        RECT 2259.590 2788.780 2422.290 2788.920 ;
        RECT 2259.590 2788.720 2259.910 2788.780 ;
        RECT 2421.970 2788.720 2422.290 2788.780 ;
        RECT 2252.690 2788.580 2253.010 2788.640 ;
        RECT 2415.530 2788.580 2415.850 2788.640 ;
        RECT 2252.690 2788.440 2415.850 2788.580 ;
        RECT 2252.690 2788.380 2253.010 2788.440 ;
        RECT 2415.530 2788.380 2415.850 2788.440 ;
        RECT 2266.505 2788.240 2266.795 2788.285 ;
        RECT 2238.060 2788.100 2266.795 2788.240 ;
        RECT 1413.650 2788.040 1413.970 2788.100 ;
        RECT 2235.685 2788.055 2235.975 2788.100 ;
        RECT 2266.505 2788.055 2266.795 2788.100 ;
        RECT 2267.410 2788.240 2267.730 2788.300 ;
        RECT 2428.870 2788.240 2429.190 2788.300 ;
        RECT 2267.410 2788.100 2429.190 2788.240 ;
        RECT 2267.410 2788.040 2267.730 2788.100 ;
        RECT 2428.870 2788.040 2429.190 2788.100 ;
        RECT 649.145 2787.900 649.435 2787.945 ;
        RECT 707.090 2787.900 707.410 2787.960 ;
        RECT 649.145 2787.760 707.410 2787.900 ;
        RECT 649.145 2787.715 649.435 2787.760 ;
        RECT 707.090 2787.700 707.410 2787.760 ;
        RECT 1045.190 2787.900 1045.510 2787.960 ;
        RECT 1093.950 2787.900 1094.270 2787.960 ;
        RECT 1045.190 2787.760 1094.270 2787.900 ;
        RECT 1045.190 2787.700 1045.510 2787.760 ;
        RECT 1093.950 2787.700 1094.270 2787.760 ;
        RECT 1414.110 2787.900 1414.430 2787.960 ;
        RECT 2091.245 2787.900 2091.535 2787.945 ;
        RECT 1414.110 2787.760 2091.535 2787.900 ;
        RECT 1414.110 2787.700 1414.430 2787.760 ;
        RECT 2091.245 2787.715 2091.535 2787.760 ;
        RECT 2091.690 2787.900 2092.010 2787.960 ;
        RECT 2162.530 2787.900 2162.850 2787.960 ;
        RECT 2091.690 2787.760 2162.850 2787.900 ;
        RECT 2091.690 2787.700 2092.010 2787.760 ;
        RECT 2162.530 2787.700 2162.850 2787.760 ;
        RECT 2163.005 2787.900 2163.295 2787.945 ;
        RECT 2208.070 2787.900 2208.390 2787.960 ;
        RECT 2163.005 2787.760 2208.390 2787.900 ;
        RECT 2163.005 2787.715 2163.295 2787.760 ;
        RECT 2208.070 2787.700 2208.390 2787.760 ;
        RECT 2245.345 2787.900 2245.635 2787.945 ;
        RECT 2270.170 2787.900 2270.490 2787.960 ;
        RECT 2245.345 2787.760 2270.490 2787.900 ;
        RECT 2245.345 2787.715 2245.635 2787.760 ;
        RECT 2270.170 2787.700 2270.490 2787.760 ;
        RECT 2283.525 2787.900 2283.815 2787.945 ;
        RECT 2298.230 2787.900 2298.550 2787.960 ;
        RECT 2283.525 2787.760 2298.550 2787.900 ;
        RECT 2283.525 2787.715 2283.815 2787.760 ;
        RECT 2298.230 2787.700 2298.550 2787.760 ;
        RECT 2312.505 2787.900 2312.795 2787.945 ;
        RECT 2321.230 2787.900 2321.550 2787.960 ;
        RECT 2367.230 2787.900 2367.550 2787.960 ;
        RECT 2373.210 2787.900 2373.530 2787.960 ;
        RECT 2312.505 2787.760 2373.530 2787.900 ;
        RECT 2312.505 2787.715 2312.795 2787.760 ;
        RECT 2321.230 2787.700 2321.550 2787.760 ;
        RECT 2367.230 2787.700 2367.550 2787.760 ;
        RECT 2373.210 2787.700 2373.530 2787.760 ;
        RECT 2375.985 2787.900 2376.275 2787.945 ;
        RECT 2381.490 2787.900 2381.810 2787.960 ;
        RECT 2375.985 2787.760 2381.810 2787.900 ;
        RECT 2375.985 2787.715 2376.275 2787.760 ;
        RECT 2381.490 2787.700 2381.810 2787.760 ;
        RECT 2381.950 2787.900 2382.270 2787.960 ;
        RECT 2415.070 2787.900 2415.390 2787.960 ;
        RECT 2381.950 2787.760 2415.390 2787.900 ;
        RECT 2381.950 2787.700 2382.270 2787.760 ;
        RECT 2415.070 2787.700 2415.390 2787.760 ;
        RECT 658.790 2787.560 659.110 2787.620 ;
        RECT 647.840 2787.420 659.110 2787.560 ;
        RECT 658.790 2787.360 659.110 2787.420 ;
        RECT 1417.330 2787.560 1417.650 2787.620 ;
        RECT 1462.425 2787.560 1462.715 2787.605 ;
        RECT 1417.330 2787.420 1462.715 2787.560 ;
        RECT 1417.330 2787.360 1417.650 2787.420 ;
        RECT 1462.425 2787.375 1462.715 2787.420 ;
        RECT 482.610 2725.340 482.930 2725.400 ;
        RECT 948.130 2725.340 948.450 2725.400 ;
        RECT 482.610 2725.200 948.450 2725.340 ;
        RECT 482.610 2725.140 482.930 2725.200 ;
        RECT 948.130 2725.140 948.450 2725.200 ;
        RECT 470.650 2725.000 470.970 2725.060 ;
        RECT 942.150 2725.000 942.470 2725.060 ;
        RECT 470.650 2724.860 942.470 2725.000 ;
        RECT 470.650 2724.800 470.970 2724.860 ;
        RECT 942.150 2724.800 942.470 2724.860 ;
        RECT 510.210 2724.660 510.530 2724.720 ;
        RECT 989.530 2724.660 989.850 2724.720 ;
        RECT 510.210 2724.520 989.850 2724.660 ;
        RECT 510.210 2724.460 510.530 2724.520 ;
        RECT 989.530 2724.460 989.850 2724.520 ;
        RECT 460.530 2724.320 460.850 2724.380 ;
        RECT 942.610 2724.320 942.930 2724.380 ;
        RECT 460.530 2724.180 942.930 2724.320 ;
        RECT 460.530 2724.120 460.850 2724.180 ;
        RECT 942.610 2724.120 942.930 2724.180 ;
        RECT 449.950 2723.980 450.270 2724.040 ;
        RECT 943.070 2723.980 943.390 2724.040 ;
        RECT 449.950 2723.840 943.390 2723.980 ;
        RECT 449.950 2723.780 450.270 2723.840 ;
        RECT 943.070 2723.780 943.390 2723.840 ;
        RECT 530.910 2723.640 531.230 2723.700 ;
        RECT 1030.930 2723.640 1031.250 2723.700 ;
        RECT 530.910 2723.500 1031.250 2723.640 ;
        RECT 530.910 2723.440 531.230 2723.500 ;
        RECT 1030.930 2723.440 1031.250 2723.500 ;
        RECT 439.830 2723.300 440.150 2723.360 ;
        RECT 943.530 2723.300 943.850 2723.360 ;
        RECT 439.830 2723.160 943.850 2723.300 ;
        RECT 439.830 2723.100 440.150 2723.160 ;
        RECT 943.530 2723.100 943.850 2723.160 ;
        RECT 551.610 2722.960 551.930 2723.020 ;
        RECT 1062.210 2722.960 1062.530 2723.020 ;
        RECT 551.610 2722.820 1062.530 2722.960 ;
        RECT 551.610 2722.760 551.930 2722.820 ;
        RECT 1062.210 2722.760 1062.530 2722.820 ;
        RECT 429.250 2722.620 429.570 2722.680 ;
        RECT 943.990 2722.620 944.310 2722.680 ;
        RECT 429.250 2722.480 944.310 2722.620 ;
        RECT 429.250 2722.420 429.570 2722.480 ;
        RECT 943.990 2722.420 944.310 2722.480 ;
        RECT 419.130 2722.280 419.450 2722.340 ;
        RECT 944.450 2722.280 944.770 2722.340 ;
        RECT 419.130 2722.140 944.770 2722.280 ;
        RECT 419.130 2722.080 419.450 2722.140 ;
        RECT 944.450 2722.080 944.770 2722.140 ;
        RECT 408.550 2721.940 408.870 2722.000 ;
        RECT 979.870 2721.940 980.190 2722.000 ;
        RECT 408.550 2721.800 980.190 2721.940 ;
        RECT 408.550 2721.740 408.870 2721.800 ;
        RECT 979.870 2721.740 980.190 2721.800 ;
        RECT 433.850 2721.600 434.170 2721.660 ;
        RECT 865.330 2721.600 865.650 2721.660 ;
        RECT 433.850 2721.460 865.650 2721.600 ;
        RECT 433.850 2721.400 434.170 2721.460 ;
        RECT 865.330 2721.400 865.650 2721.460 ;
        RECT 441.210 2721.260 441.530 2721.320 ;
        RECT 875.450 2721.260 875.770 2721.320 ;
        RECT 441.210 2721.120 875.770 2721.260 ;
        RECT 441.210 2721.060 441.530 2721.120 ;
        RECT 875.450 2721.060 875.770 2721.120 ;
        RECT 434.310 2720.920 434.630 2720.980 ;
        RECT 854.750 2720.920 855.070 2720.980 ;
        RECT 434.310 2720.780 855.070 2720.920 ;
        RECT 434.310 2720.720 434.630 2720.780 ;
        RECT 854.750 2720.720 855.070 2720.780 ;
        RECT 427.410 2720.580 427.730 2720.640 ;
        RECT 844.170 2720.580 844.490 2720.640 ;
        RECT 427.410 2720.440 844.490 2720.580 ;
        RECT 427.410 2720.380 427.730 2720.440 ;
        RECT 844.170 2720.380 844.490 2720.440 ;
        RECT 413.610 2720.240 413.930 2720.300 ;
        RECT 823.470 2720.240 823.790 2720.300 ;
        RECT 413.610 2720.100 823.790 2720.240 ;
        RECT 413.610 2720.040 413.930 2720.100 ;
        RECT 823.470 2720.040 823.790 2720.100 ;
        RECT 365.310 2719.900 365.630 2719.960 ;
        RECT 740.670 2719.900 740.990 2719.960 ;
        RECT 365.310 2719.760 740.990 2719.900 ;
        RECT 365.310 2719.700 365.630 2719.760 ;
        RECT 740.670 2719.700 740.990 2719.760 ;
        RECT 289.410 2719.560 289.730 2719.620 ;
        RECT 564.030 2719.560 564.350 2719.620 ;
        RECT 289.410 2719.420 564.350 2719.560 ;
        RECT 289.410 2719.360 289.730 2719.420 ;
        RECT 564.030 2719.360 564.350 2719.420 ;
        RECT 288.950 2719.220 289.270 2719.280 ;
        RECT 553.910 2719.220 554.230 2719.280 ;
        RECT 288.950 2719.080 554.230 2719.220 ;
        RECT 288.950 2719.020 289.270 2719.080 ;
        RECT 553.910 2719.020 554.230 2719.080 ;
        RECT 1103.610 2718.680 1103.930 2718.940 ;
        RECT 358.410 2718.540 358.730 2718.600 ;
        RECT 377.270 2718.540 377.590 2718.600 ;
        RECT 358.410 2718.400 377.590 2718.540 ;
        RECT 358.410 2718.340 358.730 2718.400 ;
        RECT 377.270 2718.340 377.590 2718.400 ;
        RECT 379.110 2718.540 379.430 2718.600 ;
        RECT 727.345 2718.540 727.635 2718.585 ;
        RECT 379.110 2718.400 727.635 2718.540 ;
        RECT 379.110 2718.340 379.430 2718.400 ;
        RECT 727.345 2718.355 727.635 2718.400 ;
        RECT 727.790 2718.540 728.110 2718.600 ;
        RECT 762.305 2718.540 762.595 2718.585 ;
        RECT 727.790 2718.400 762.595 2718.540 ;
        RECT 727.790 2718.340 728.110 2718.400 ;
        RECT 762.305 2718.355 762.595 2718.400 ;
        RECT 762.750 2718.540 763.070 2718.600 ;
        RECT 813.350 2718.540 813.670 2718.600 ;
        RECT 762.750 2718.400 813.670 2718.540 ;
        RECT 762.750 2718.340 763.070 2718.400 ;
        RECT 813.350 2718.340 813.670 2718.400 ;
        RECT 1027.710 2718.540 1028.030 2718.600 ;
        RECT 1093.490 2718.540 1093.810 2718.600 ;
        RECT 1027.710 2718.400 1093.810 2718.540 ;
        RECT 1027.710 2718.340 1028.030 2718.400 ;
        RECT 1093.490 2718.340 1093.810 2718.400 ;
        RECT 1102.690 2718.540 1103.010 2718.600 ;
        RECT 1103.700 2718.540 1103.840 2718.680 ;
        RECT 1102.690 2718.400 1103.840 2718.540 ;
        RECT 1138.110 2718.540 1138.430 2718.600 ;
        RECT 1290.370 2718.540 1290.690 2718.600 ;
        RECT 1138.110 2718.400 1290.690 2718.540 ;
        RECT 1102.690 2718.340 1103.010 2718.400 ;
        RECT 1138.110 2718.340 1138.430 2718.400 ;
        RECT 1290.370 2718.340 1290.690 2718.400 ;
        RECT 392.910 2718.200 393.230 2718.260 ;
        RECT 782.070 2718.200 782.390 2718.260 ;
        RECT 392.910 2718.060 782.390 2718.200 ;
        RECT 392.910 2718.000 393.230 2718.060 ;
        RECT 782.070 2718.000 782.390 2718.060 ;
        RECT 1034.610 2718.200 1034.930 2718.260 ;
        RECT 1103.610 2718.200 1103.930 2718.260 ;
        RECT 1034.610 2718.060 1103.930 2718.200 ;
        RECT 1034.610 2718.000 1034.930 2718.060 ;
        RECT 1103.610 2718.000 1103.930 2718.060 ;
        RECT 1145.010 2718.200 1145.330 2718.260 ;
        RECT 1300.950 2718.200 1301.270 2718.260 ;
        RECT 1145.010 2718.060 1301.270 2718.200 ;
        RECT 1145.010 2718.000 1145.330 2718.060 ;
        RECT 1300.950 2718.000 1301.270 2718.060 ;
        RECT 305.050 2717.860 305.370 2717.920 ;
        RECT 310.110 2717.860 310.430 2717.920 ;
        RECT 305.050 2717.720 310.430 2717.860 ;
        RECT 305.050 2717.660 305.370 2717.720 ;
        RECT 310.110 2717.660 310.430 2717.720 ;
        RECT 325.750 2717.860 326.070 2717.920 ;
        RECT 330.810 2717.860 331.130 2717.920 ;
        RECT 325.750 2717.720 331.130 2717.860 ;
        RECT 325.750 2717.660 326.070 2717.720 ;
        RECT 330.810 2717.660 331.130 2717.720 ;
        RECT 351.510 2717.860 351.830 2717.920 ;
        RECT 356.570 2717.860 356.890 2717.920 ;
        RECT 351.510 2717.720 356.890 2717.860 ;
        RECT 351.510 2717.660 351.830 2717.720 ;
        RECT 356.570 2717.660 356.890 2717.720 ;
        RECT 399.810 2717.860 400.130 2717.920 ;
        RECT 761.845 2717.860 762.135 2717.905 ;
        RECT 399.810 2717.720 762.135 2717.860 ;
        RECT 399.810 2717.660 400.130 2717.720 ;
        RECT 761.845 2717.675 762.135 2717.720 ;
        RECT 762.290 2717.860 762.610 2717.920 ;
        RECT 792.650 2717.860 792.970 2717.920 ;
        RECT 762.290 2717.720 792.970 2717.860 ;
        RECT 762.290 2717.660 762.610 2717.720 ;
        RECT 792.650 2717.660 792.970 2717.720 ;
        RECT 1041.510 2717.860 1041.830 2717.920 ;
        RECT 1114.190 2717.860 1114.510 2717.920 ;
        RECT 1041.510 2717.720 1114.510 2717.860 ;
        RECT 1041.510 2717.660 1041.830 2717.720 ;
        RECT 1114.190 2717.660 1114.510 2717.720 ;
        RECT 1151.910 2717.860 1152.230 2717.920 ;
        RECT 1311.070 2717.860 1311.390 2717.920 ;
        RECT 1151.910 2717.720 1311.390 2717.860 ;
        RECT 1151.910 2717.660 1152.230 2717.720 ;
        RECT 1311.070 2717.660 1311.390 2717.720 ;
        RECT 287.110 2717.520 287.430 2717.580 ;
        RECT 512.510 2717.520 512.830 2717.580 ;
        RECT 287.110 2717.380 512.830 2717.520 ;
        RECT 287.110 2717.320 287.430 2717.380 ;
        RECT 512.510 2717.320 512.830 2717.380 ;
        RECT 636.710 2717.520 637.030 2717.580 ;
        RECT 1045.190 2717.520 1045.510 2717.580 ;
        RECT 636.710 2717.380 1045.510 2717.520 ;
        RECT 636.710 2717.320 637.030 2717.380 ;
        RECT 1045.190 2717.320 1045.510 2717.380 ;
        RECT 1048.410 2717.520 1048.730 2717.580 ;
        RECT 1124.310 2717.520 1124.630 2717.580 ;
        RECT 1048.410 2717.380 1124.630 2717.520 ;
        RECT 1048.410 2717.320 1048.730 2717.380 ;
        RECT 1124.310 2717.320 1124.630 2717.380 ;
        RECT 1158.810 2717.520 1159.130 2717.580 ;
        RECT 1321.650 2717.520 1321.970 2717.580 ;
        RECT 1158.810 2717.380 1321.970 2717.520 ;
        RECT 1158.810 2717.320 1159.130 2717.380 ;
        RECT 1321.650 2717.320 1321.970 2717.380 ;
        RECT 287.570 2717.180 287.890 2717.240 ;
        RECT 522.630 2717.180 522.950 2717.240 ;
        RECT 287.570 2717.040 522.950 2717.180 ;
        RECT 287.570 2716.980 287.890 2717.040 ;
        RECT 522.630 2716.980 522.950 2717.040 ;
        RECT 616.010 2717.180 616.330 2717.240 ;
        RECT 1038.290 2717.180 1038.610 2717.240 ;
        RECT 616.010 2717.040 1038.610 2717.180 ;
        RECT 616.010 2716.980 616.330 2717.040 ;
        RECT 1038.290 2716.980 1038.610 2717.040 ;
        RECT 1054.850 2717.180 1055.170 2717.240 ;
        RECT 1134.890 2717.180 1135.210 2717.240 ;
        RECT 1054.850 2717.040 1135.210 2717.180 ;
        RECT 1054.850 2716.980 1055.170 2717.040 ;
        RECT 1134.890 2716.980 1135.210 2717.040 ;
        RECT 1165.710 2717.180 1166.030 2717.240 ;
        RECT 1332.230 2717.180 1332.550 2717.240 ;
        RECT 1165.710 2717.040 1332.550 2717.180 ;
        RECT 1165.710 2716.980 1166.030 2717.040 ;
        RECT 1332.230 2716.980 1332.550 2717.040 ;
        RECT 288.030 2716.840 288.350 2716.900 ;
        RECT 533.210 2716.840 533.530 2716.900 ;
        RECT 288.030 2716.700 533.530 2716.840 ;
        RECT 288.030 2716.640 288.350 2716.700 ;
        RECT 533.210 2716.640 533.530 2716.700 ;
        RECT 595.310 2716.840 595.630 2716.900 ;
        RECT 1024.490 2716.840 1024.810 2716.900 ;
        RECT 595.310 2716.700 1024.810 2716.840 ;
        RECT 595.310 2716.640 595.630 2716.700 ;
        RECT 1024.490 2716.640 1024.810 2716.700 ;
        RECT 1061.750 2716.840 1062.070 2716.900 ;
        RECT 1155.590 2716.840 1155.910 2716.900 ;
        RECT 1061.750 2716.700 1155.910 2716.840 ;
        RECT 1061.750 2716.640 1062.070 2716.700 ;
        RECT 1155.590 2716.640 1155.910 2716.700 ;
        RECT 1165.250 2716.840 1165.570 2716.900 ;
        RECT 1342.350 2716.840 1342.670 2716.900 ;
        RECT 1165.250 2716.700 1342.670 2716.840 ;
        RECT 1165.250 2716.640 1165.570 2716.700 ;
        RECT 1342.350 2716.640 1342.670 2716.700 ;
        RECT 455.010 2716.500 455.330 2716.560 ;
        RECT 896.150 2716.500 896.470 2716.560 ;
        RECT 455.010 2716.360 896.470 2716.500 ;
        RECT 455.010 2716.300 455.330 2716.360 ;
        RECT 896.150 2716.300 896.470 2716.360 ;
        RECT 1076.010 2716.500 1076.330 2716.560 ;
        RECT 1176.290 2716.500 1176.610 2716.560 ;
        RECT 1076.010 2716.360 1176.610 2716.500 ;
        RECT 1076.010 2716.300 1076.330 2716.360 ;
        RECT 1176.290 2716.300 1176.610 2716.360 ;
        RECT 1179.510 2716.500 1179.830 2716.560 ;
        RECT 1363.050 2716.500 1363.370 2716.560 ;
        RECT 1179.510 2716.360 1363.370 2716.500 ;
        RECT 1179.510 2716.300 1179.830 2716.360 ;
        RECT 1363.050 2716.300 1363.370 2716.360 ;
        RECT 288.490 2716.160 288.810 2716.220 ;
        RECT 543.330 2716.160 543.650 2716.220 ;
        RECT 288.490 2716.020 543.650 2716.160 ;
        RECT 288.490 2715.960 288.810 2716.020 ;
        RECT 543.330 2715.960 543.650 2716.020 ;
        RECT 574.610 2716.160 574.930 2716.220 ;
        RECT 1010.690 2716.160 1011.010 2716.220 ;
        RECT 574.610 2716.020 1011.010 2716.160 ;
        RECT 574.610 2715.960 574.930 2716.020 ;
        RECT 1010.690 2715.960 1011.010 2716.020 ;
        RECT 1055.310 2716.160 1055.630 2716.220 ;
        RECT 1145.470 2716.160 1145.790 2716.220 ;
        RECT 1055.310 2716.020 1145.790 2716.160 ;
        RECT 1055.310 2715.960 1055.630 2716.020 ;
        RECT 1145.470 2715.960 1145.790 2716.020 ;
        RECT 1172.610 2716.160 1172.930 2716.220 ;
        RECT 1352.930 2716.160 1353.250 2716.220 ;
        RECT 1172.610 2716.020 1353.250 2716.160 ;
        RECT 1172.610 2715.960 1172.930 2716.020 ;
        RECT 1352.930 2715.960 1353.250 2716.020 ;
        RECT 468.350 2715.820 468.670 2715.880 ;
        RECT 916.850 2715.820 917.170 2715.880 ;
        RECT 468.350 2715.680 917.170 2715.820 ;
        RECT 468.350 2715.620 468.670 2715.680 ;
        RECT 916.850 2715.620 917.170 2715.680 ;
        RECT 1013.910 2715.820 1014.230 2715.880 ;
        RECT 1072.790 2715.820 1073.110 2715.880 ;
        RECT 1013.910 2715.680 1073.110 2715.820 ;
        RECT 1013.910 2715.620 1014.230 2715.680 ;
        RECT 1072.790 2715.620 1073.110 2715.680 ;
        RECT 1082.910 2715.820 1083.230 2715.880 ;
        RECT 1186.870 2715.820 1187.190 2715.880 ;
        RECT 1082.910 2715.680 1187.190 2715.820 ;
        RECT 1082.910 2715.620 1083.230 2715.680 ;
        RECT 1186.870 2715.620 1187.190 2715.680 ;
        RECT 1193.310 2715.820 1193.630 2715.880 ;
        RECT 1383.750 2715.820 1384.070 2715.880 ;
        RECT 1193.310 2715.680 1384.070 2715.820 ;
        RECT 1193.310 2715.620 1193.630 2715.680 ;
        RECT 1383.750 2715.620 1384.070 2715.680 ;
        RECT 286.190 2715.480 286.510 2715.540 ;
        RECT 398.430 2715.480 398.750 2715.540 ;
        RECT 286.190 2715.340 398.750 2715.480 ;
        RECT 286.190 2715.280 286.510 2715.340 ;
        RECT 398.430 2715.280 398.750 2715.340 ;
        RECT 475.250 2715.480 475.570 2715.540 ;
        RECT 937.550 2715.480 937.870 2715.540 ;
        RECT 475.250 2715.340 937.870 2715.480 ;
        RECT 475.250 2715.280 475.570 2715.340 ;
        RECT 937.550 2715.280 937.870 2715.340 ;
        RECT 1020.810 2715.280 1021.130 2715.540 ;
        RECT 1069.110 2715.480 1069.430 2715.540 ;
        RECT 1166.170 2715.480 1166.490 2715.540 ;
        RECT 1069.110 2715.340 1166.490 2715.480 ;
        RECT 1069.110 2715.280 1069.430 2715.340 ;
        RECT 1166.170 2715.280 1166.490 2715.340 ;
        RECT 1186.410 2715.480 1186.730 2715.540 ;
        RECT 1373.630 2715.480 1373.950 2715.540 ;
        RECT 1186.410 2715.340 1373.950 2715.480 ;
        RECT 1186.410 2715.280 1186.730 2715.340 ;
        RECT 1373.630 2715.280 1373.950 2715.340 ;
        RECT 337.710 2715.140 338.030 2715.200 ;
        RECT 491.810 2715.140 492.130 2715.200 ;
        RECT 337.710 2715.000 492.130 2715.140 ;
        RECT 337.710 2714.940 338.030 2715.000 ;
        RECT 491.810 2714.940 492.130 2715.000 ;
        RECT 496.410 2715.140 496.730 2715.200 ;
        RECT 968.830 2715.140 969.150 2715.200 ;
        RECT 496.410 2715.000 969.150 2715.140 ;
        RECT 1020.900 2715.140 1021.040 2715.280 ;
        RECT 1082.910 2715.140 1083.230 2715.200 ;
        RECT 1020.900 2715.000 1083.230 2715.140 ;
        RECT 496.410 2714.940 496.730 2715.000 ;
        RECT 968.830 2714.940 969.150 2715.000 ;
        RECT 1082.910 2714.940 1083.230 2715.000 ;
        RECT 1089.350 2715.140 1089.670 2715.200 ;
        RECT 1196.990 2715.140 1197.310 2715.200 ;
        RECT 1089.350 2715.000 1197.310 2715.140 ;
        RECT 1089.350 2714.940 1089.670 2715.000 ;
        RECT 1196.990 2714.940 1197.310 2715.000 ;
        RECT 1200.210 2715.140 1200.530 2715.200 ;
        RECT 1394.330 2715.140 1394.650 2715.200 ;
        RECT 1200.210 2715.000 1394.650 2715.140 ;
        RECT 1200.210 2714.940 1200.530 2715.000 ;
        RECT 1394.330 2714.940 1394.650 2715.000 ;
        RECT 286.650 2714.800 286.970 2714.860 ;
        RECT 501.930 2714.800 502.250 2714.860 ;
        RECT 286.650 2714.660 502.250 2714.800 ;
        RECT 286.650 2714.600 286.970 2714.660 ;
        RECT 501.930 2714.600 502.250 2714.660 ;
        RECT 542.870 2714.800 543.190 2714.860 ;
        RECT 719.970 2714.800 720.290 2714.860 ;
        RECT 542.870 2714.660 720.290 2714.800 ;
        RECT 542.870 2714.600 543.190 2714.660 ;
        RECT 719.970 2714.600 720.290 2714.660 ;
        RECT 720.890 2714.800 721.210 2714.860 ;
        RECT 1020.810 2714.800 1021.130 2714.860 ;
        RECT 720.890 2714.660 1021.130 2714.800 ;
        RECT 720.890 2714.600 721.210 2714.660 ;
        RECT 1020.810 2714.600 1021.130 2714.660 ;
        RECT 1130.750 2714.800 1131.070 2714.860 ;
        RECT 1280.250 2714.800 1280.570 2714.860 ;
        RECT 1130.750 2714.660 1280.570 2714.800 ;
        RECT 1130.750 2714.600 1131.070 2714.660 ;
        RECT 1280.250 2714.600 1280.570 2714.660 ;
        RECT 527.690 2714.460 528.010 2714.520 ;
        RECT 699.270 2714.460 699.590 2714.520 ;
        RECT 527.690 2714.320 699.590 2714.460 ;
        RECT 527.690 2714.260 528.010 2714.320 ;
        RECT 699.270 2714.260 699.590 2714.320 ;
        RECT 700.650 2714.460 700.970 2714.520 ;
        RECT 979.410 2714.460 979.730 2714.520 ;
        RECT 700.650 2714.320 979.730 2714.460 ;
        RECT 700.650 2714.260 700.970 2714.320 ;
        RECT 979.410 2714.260 979.730 2714.320 ;
        RECT 1131.210 2714.460 1131.530 2714.520 ;
        RECT 1269.670 2714.460 1269.990 2714.520 ;
        RECT 1131.210 2714.320 1269.990 2714.460 ;
        RECT 1131.210 2714.260 1131.530 2714.320 ;
        RECT 1269.670 2714.260 1269.990 2714.320 ;
        RECT 520.790 2714.120 521.110 2714.180 ;
        RECT 688.690 2714.120 689.010 2714.180 ;
        RECT 520.790 2713.980 689.010 2714.120 ;
        RECT 520.790 2713.920 521.110 2713.980 ;
        RECT 688.690 2713.920 689.010 2713.980 ;
        RECT 693.290 2714.120 693.610 2714.180 ;
        RECT 958.710 2714.120 959.030 2714.180 ;
        RECT 693.290 2713.980 959.030 2714.120 ;
        RECT 693.290 2713.920 693.610 2713.980 ;
        RECT 958.710 2713.920 959.030 2713.980 ;
        RECT 1117.410 2714.120 1117.730 2714.180 ;
        RECT 1248.970 2714.120 1249.290 2714.180 ;
        RECT 1117.410 2713.980 1249.290 2714.120 ;
        RECT 1117.410 2713.920 1117.730 2713.980 ;
        RECT 1248.970 2713.920 1249.290 2713.980 ;
        RECT 513.890 2713.780 514.210 2713.840 ;
        RECT 678.570 2713.780 678.890 2713.840 ;
        RECT 513.890 2713.640 678.890 2713.780 ;
        RECT 513.890 2713.580 514.210 2713.640 ;
        RECT 678.570 2713.580 678.890 2713.640 ;
        RECT 686.390 2713.780 686.710 2713.840 ;
        RECT 927.430 2713.780 927.750 2713.840 ;
        RECT 686.390 2713.640 927.750 2713.780 ;
        RECT 686.390 2713.580 686.710 2713.640 ;
        RECT 927.430 2713.580 927.750 2713.640 ;
        RECT 1123.390 2713.780 1123.710 2713.840 ;
        RECT 1259.550 2713.780 1259.870 2713.840 ;
        RECT 1123.390 2713.640 1259.870 2713.780 ;
        RECT 1123.390 2713.580 1123.710 2713.640 ;
        RECT 1259.550 2713.580 1259.870 2713.640 ;
        RECT 351.050 2713.440 351.370 2713.500 ;
        RECT 367.150 2713.440 367.470 2713.500 ;
        RECT 351.050 2713.300 367.470 2713.440 ;
        RECT 351.050 2713.240 351.370 2713.300 ;
        RECT 367.150 2713.240 367.470 2713.300 ;
        RECT 500.090 2713.440 500.410 2713.500 ;
        RECT 657.410 2713.440 657.730 2713.500 ;
        RECT 500.090 2713.300 657.730 2713.440 ;
        RECT 500.090 2713.240 500.410 2713.300 ;
        RECT 657.410 2713.240 657.730 2713.300 ;
        RECT 658.790 2713.440 659.110 2713.500 ;
        RECT 886.030 2713.440 886.350 2713.500 ;
        RECT 658.790 2713.300 886.350 2713.440 ;
        RECT 658.790 2713.240 659.110 2713.300 ;
        RECT 886.030 2713.240 886.350 2713.300 ;
        RECT 1110.510 2713.440 1110.830 2713.500 ;
        RECT 1238.850 2713.440 1239.170 2713.500 ;
        RECT 1110.510 2713.300 1239.170 2713.440 ;
        RECT 1110.510 2713.240 1110.830 2713.300 ;
        RECT 1238.850 2713.240 1239.170 2713.300 ;
        RECT 506.990 2713.100 507.310 2713.160 ;
        RECT 667.990 2713.100 668.310 2713.160 ;
        RECT 506.990 2712.960 668.310 2713.100 ;
        RECT 506.990 2712.900 507.310 2712.960 ;
        RECT 667.990 2712.900 668.310 2712.960 ;
        RECT 687.310 2713.100 687.630 2713.160 ;
        RECT 906.730 2713.100 907.050 2713.160 ;
        RECT 687.310 2712.960 907.050 2713.100 ;
        RECT 687.310 2712.900 687.630 2712.960 ;
        RECT 906.730 2712.900 907.050 2712.960 ;
        RECT 1102.690 2713.100 1103.010 2713.160 ;
        RECT 1228.270 2713.100 1228.590 2713.160 ;
        RECT 1102.690 2712.960 1228.590 2713.100 ;
        RECT 1102.690 2712.900 1103.010 2712.960 ;
        RECT 1228.270 2712.900 1228.590 2712.960 ;
        RECT 541.490 2712.760 541.810 2712.820 ;
        RECT 730.090 2712.760 730.410 2712.820 ;
        RECT 761.370 2712.760 761.690 2712.820 ;
        RECT 541.490 2712.620 730.410 2712.760 ;
        RECT 541.490 2712.560 541.810 2712.620 ;
        RECT 730.090 2712.560 730.410 2712.620 ;
        RECT 734.780 2712.620 761.690 2712.760 ;
        RECT 534.590 2712.420 534.910 2712.480 ;
        RECT 709.390 2712.420 709.710 2712.480 ;
        RECT 534.590 2712.280 709.710 2712.420 ;
        RECT 534.590 2712.220 534.910 2712.280 ;
        RECT 709.390 2712.220 709.710 2712.280 ;
        RECT 727.345 2712.420 727.635 2712.465 ;
        RECT 734.780 2712.420 734.920 2712.620 ;
        RECT 761.370 2712.560 761.690 2712.620 ;
        RECT 762.305 2712.760 762.595 2712.805 ;
        RECT 771.950 2712.760 772.270 2712.820 ;
        RECT 834.050 2712.760 834.370 2712.820 ;
        RECT 762.305 2712.620 772.270 2712.760 ;
        RECT 762.305 2712.575 762.595 2712.620 ;
        RECT 771.950 2712.560 772.270 2712.620 ;
        RECT 783.080 2712.620 834.370 2712.760 ;
        RECT 727.345 2712.280 734.920 2712.420 ;
        RECT 748.490 2712.420 748.810 2712.480 ;
        RECT 783.080 2712.420 783.220 2712.620 ;
        RECT 834.050 2712.560 834.370 2712.620 ;
        RECT 1089.810 2712.760 1090.130 2712.820 ;
        RECT 1207.570 2712.760 1207.890 2712.820 ;
        RECT 1089.810 2712.620 1207.890 2712.760 ;
        RECT 1089.810 2712.560 1090.130 2712.620 ;
        RECT 1207.570 2712.560 1207.890 2712.620 ;
        RECT 748.490 2712.280 783.220 2712.420 ;
        RECT 1096.710 2712.420 1097.030 2712.480 ;
        RECT 1217.690 2712.420 1218.010 2712.480 ;
        RECT 1096.710 2712.280 1218.010 2712.420 ;
        RECT 727.345 2712.235 727.635 2712.280 ;
        RECT 748.490 2712.220 748.810 2712.280 ;
        RECT 1096.710 2712.220 1097.030 2712.280 ;
        RECT 1217.690 2712.220 1218.010 2712.280 ;
        RECT 686.850 2712.080 687.170 2712.140 ;
        RECT 750.790 2712.080 751.110 2712.140 ;
        RECT 686.850 2711.940 751.110 2712.080 ;
        RECT 686.850 2711.880 687.170 2711.940 ;
        RECT 750.790 2711.880 751.110 2711.940 ;
        RECT 761.845 2712.080 762.135 2712.125 ;
        RECT 802.770 2712.080 803.090 2712.140 ;
        RECT 761.845 2711.940 803.090 2712.080 ;
        RECT 761.845 2711.895 762.135 2711.940 ;
        RECT 802.770 2711.880 803.090 2711.940 ;
        RECT 1408.590 2697.800 1408.910 2697.860 ;
        RECT 2321.690 2697.800 2322.010 2697.860 ;
        RECT 1408.590 2697.660 2322.010 2697.800 ;
        RECT 1408.590 2697.600 1408.910 2697.660 ;
        RECT 2321.690 2697.600 2322.010 2697.660 ;
      LAYER met1 ;
        RECT 300.000 1610.640 1396.500 2695.780 ;
      LAYER met1 ;
        RECT 1408.590 2691.000 1408.910 2691.060 ;
        RECT 2273.390 2691.000 2273.710 2691.060 ;
        RECT 1408.590 2690.860 2273.710 2691.000 ;
        RECT 1408.590 2690.800 1408.910 2690.860 ;
        RECT 2273.390 2690.800 2273.710 2690.860 ;
        RECT 1408.590 2677.060 1408.910 2677.120 ;
        RECT 2267.410 2677.060 2267.730 2677.120 ;
        RECT 1408.590 2676.920 2267.730 2677.060 ;
        RECT 1408.590 2676.860 1408.910 2676.920 ;
        RECT 2267.410 2676.860 2267.730 2676.920 ;
        RECT 1408.590 2670.260 1408.910 2670.320 ;
        RECT 2259.590 2670.260 2259.910 2670.320 ;
        RECT 1408.590 2670.120 2259.910 2670.260 ;
        RECT 1408.590 2670.060 1408.910 2670.120 ;
        RECT 2259.590 2670.060 2259.910 2670.120 ;
        RECT 1408.590 2656.320 1408.910 2656.380 ;
        RECT 2252.690 2656.320 2253.010 2656.380 ;
        RECT 1408.590 2656.180 2253.010 2656.320 ;
        RECT 1408.590 2656.120 1408.910 2656.180 ;
        RECT 2252.690 2656.120 2253.010 2656.180 ;
        RECT 1408.590 2649.520 1408.910 2649.580 ;
        RECT 2245.790 2649.520 2246.110 2649.580 ;
        RECT 1408.590 2649.380 2246.110 2649.520 ;
        RECT 1408.590 2649.320 1408.910 2649.380 ;
        RECT 2245.790 2649.320 2246.110 2649.380 ;
        RECT 1408.590 2635.580 1408.910 2635.640 ;
        RECT 2238.890 2635.580 2239.210 2635.640 ;
        RECT 1408.590 2635.440 2239.210 2635.580 ;
        RECT 1408.590 2635.380 1408.910 2635.440 ;
        RECT 2238.890 2635.380 2239.210 2635.440 ;
        RECT 1408.590 2628.780 1408.910 2628.840 ;
        RECT 2231.990 2628.780 2232.310 2628.840 ;
        RECT 1408.590 2628.640 2232.310 2628.780 ;
        RECT 1408.590 2628.580 1408.910 2628.640 ;
        RECT 2231.990 2628.580 2232.310 2628.640 ;
        RECT 1408.590 2614.840 1408.910 2614.900 ;
        RECT 2218.190 2614.840 2218.510 2614.900 ;
        RECT 1408.590 2614.700 2218.510 2614.840 ;
        RECT 1408.590 2614.640 1408.910 2614.700 ;
        RECT 2218.190 2614.640 2218.510 2614.700 ;
        RECT 1408.590 2608.040 1408.910 2608.100 ;
        RECT 1797.750 2608.040 1798.070 2608.100 ;
        RECT 1408.590 2607.900 1798.070 2608.040 ;
        RECT 1408.590 2607.840 1408.910 2607.900 ;
        RECT 1797.750 2607.840 1798.070 2607.900 ;
        RECT 1408.590 2594.440 1408.910 2594.500 ;
        RECT 1797.290 2594.440 1797.610 2594.500 ;
        RECT 1408.590 2594.300 1797.610 2594.440 ;
        RECT 1408.590 2594.240 1408.910 2594.300 ;
        RECT 1797.290 2594.240 1797.610 2594.300 ;
        RECT 1408.590 2587.300 1408.910 2587.360 ;
        RECT 1790.850 2587.300 1791.170 2587.360 ;
        RECT 1408.590 2587.160 1791.170 2587.300 ;
        RECT 1408.590 2587.100 1408.910 2587.160 ;
        RECT 1790.850 2587.100 1791.170 2587.160 ;
        RECT 1408.590 2573.700 1408.910 2573.760 ;
        RECT 1783.490 2573.700 1783.810 2573.760 ;
        RECT 1408.590 2573.560 1783.810 2573.700 ;
        RECT 1408.590 2573.500 1408.910 2573.560 ;
        RECT 1783.490 2573.500 1783.810 2573.560 ;
        RECT 1408.590 2566.560 1408.910 2566.620 ;
        RECT 2366.770 2566.560 2367.090 2566.620 ;
        RECT 1408.590 2566.420 2367.090 2566.560 ;
        RECT 1408.590 2566.360 1408.910 2566.420 ;
        RECT 2366.770 2566.360 2367.090 2566.420 ;
        RECT 1408.590 2552.960 1408.910 2553.020 ;
        RECT 2359.870 2552.960 2360.190 2553.020 ;
        RECT 1408.590 2552.820 2360.190 2552.960 ;
        RECT 1408.590 2552.760 1408.910 2552.820 ;
        RECT 2359.870 2552.760 2360.190 2552.820 ;
        RECT 1408.590 2546.160 1408.910 2546.220 ;
        RECT 2352.970 2546.160 2353.290 2546.220 ;
        RECT 1408.590 2546.020 2353.290 2546.160 ;
        RECT 1408.590 2545.960 1408.910 2546.020 ;
        RECT 2352.970 2545.960 2353.290 2546.020 ;
        RECT 1408.590 2532.220 1408.910 2532.280 ;
        RECT 2346.070 2532.220 2346.390 2532.280 ;
        RECT 1408.590 2532.080 2346.390 2532.220 ;
        RECT 1408.590 2532.020 1408.910 2532.080 ;
        RECT 2346.070 2532.020 2346.390 2532.080 ;
        RECT 1408.590 2525.420 1408.910 2525.480 ;
        RECT 2339.630 2525.420 2339.950 2525.480 ;
        RECT 1408.590 2525.280 2339.950 2525.420 ;
        RECT 1408.590 2525.220 1408.910 2525.280 ;
        RECT 2339.630 2525.220 2339.950 2525.280 ;
        RECT 1408.590 2511.480 1408.910 2511.540 ;
        RECT 2339.170 2511.480 2339.490 2511.540 ;
        RECT 1408.590 2511.340 2339.490 2511.480 ;
        RECT 1408.590 2511.280 1408.910 2511.340 ;
        RECT 2339.170 2511.280 2339.490 2511.340 ;
        RECT 1408.590 2504.680 1408.910 2504.740 ;
        RECT 2332.270 2504.680 2332.590 2504.740 ;
        RECT 1408.590 2504.540 2332.590 2504.680 ;
        RECT 1408.590 2504.480 1408.910 2504.540 ;
        RECT 2332.270 2504.480 2332.590 2504.540 ;
        RECT 1408.590 2497.540 1408.910 2497.600 ;
        RECT 2325.370 2497.540 2325.690 2497.600 ;
        RECT 1408.590 2497.400 2325.690 2497.540 ;
        RECT 1408.590 2497.340 1408.910 2497.400 ;
        RECT 2325.370 2497.340 2325.690 2497.400 ;
        RECT 1408.590 2483.940 1408.910 2484.000 ;
        RECT 2318.470 2483.940 2318.790 2484.000 ;
        RECT 1408.590 2483.800 2318.790 2483.940 ;
        RECT 1408.590 2483.740 1408.910 2483.800 ;
        RECT 2318.470 2483.740 2318.790 2483.800 ;
        RECT 1408.590 2477.140 1408.910 2477.200 ;
        RECT 2311.570 2477.140 2311.890 2477.200 ;
        RECT 1408.590 2477.000 2311.890 2477.140 ;
        RECT 1408.590 2476.940 1408.910 2477.000 ;
        RECT 2311.570 2476.940 2311.890 2477.000 ;
        RECT 1408.590 2463.200 1408.910 2463.260 ;
        RECT 2305.130 2463.200 2305.450 2463.260 ;
        RECT 1408.590 2463.060 2305.450 2463.200 ;
        RECT 1408.590 2463.000 1408.910 2463.060 ;
        RECT 2305.130 2463.000 2305.450 2463.060 ;
        RECT 1408.590 2456.400 1408.910 2456.460 ;
        RECT 2304.670 2456.400 2304.990 2456.460 ;
        RECT 1408.590 2456.260 2304.990 2456.400 ;
        RECT 1408.590 2456.200 1408.910 2456.260 ;
        RECT 2304.670 2456.200 2304.990 2456.260 ;
        RECT 1408.590 2442.460 1408.910 2442.520 ;
        RECT 2297.770 2442.460 2298.090 2442.520 ;
        RECT 1408.590 2442.320 2298.090 2442.460 ;
        RECT 1408.590 2442.260 1408.910 2442.320 ;
        RECT 2297.770 2442.260 2298.090 2442.320 ;
        RECT 1408.590 2435.660 1408.910 2435.720 ;
        RECT 2290.870 2435.660 2291.190 2435.720 ;
        RECT 1408.590 2435.520 2291.190 2435.660 ;
        RECT 1408.590 2435.460 1408.910 2435.520 ;
        RECT 2290.870 2435.460 2291.190 2435.520 ;
        RECT 1408.590 2421.720 1408.910 2421.780 ;
        RECT 2283.970 2421.720 2284.290 2421.780 ;
        RECT 1408.590 2421.580 2284.290 2421.720 ;
        RECT 1408.590 2421.520 1408.910 2421.580 ;
        RECT 2283.970 2421.520 2284.290 2421.580 ;
        RECT 1408.590 2414.920 1408.910 2414.980 ;
        RECT 2277.070 2414.920 2277.390 2414.980 ;
        RECT 1408.590 2414.780 2277.390 2414.920 ;
        RECT 1408.590 2414.720 1408.910 2414.780 ;
        RECT 2277.070 2414.720 2277.390 2414.780 ;
        RECT 1408.590 2400.980 1408.910 2401.040 ;
        RECT 2266.950 2400.980 2267.270 2401.040 ;
        RECT 1408.590 2400.840 2267.270 2400.980 ;
        RECT 1408.590 2400.780 1408.910 2400.840 ;
        RECT 2266.950 2400.780 2267.270 2400.840 ;
        RECT 1408.590 2394.180 1408.910 2394.240 ;
        RECT 1790.390 2394.180 1790.710 2394.240 ;
        RECT 1408.590 2394.040 1790.710 2394.180 ;
        RECT 1408.590 2393.980 1408.910 2394.040 ;
        RECT 1790.390 2393.980 1790.710 2394.040 ;
        RECT 1408.590 2380.240 1408.910 2380.300 ;
        RECT 2263.270 2380.240 2263.590 2380.300 ;
        RECT 1408.590 2380.100 2263.590 2380.240 ;
        RECT 1408.590 2380.040 1408.910 2380.100 ;
        RECT 2263.270 2380.040 2263.590 2380.100 ;
        RECT 1408.590 2373.440 1408.910 2373.500 ;
        RECT 1794.530 2373.440 1794.850 2373.500 ;
        RECT 1408.590 2373.300 1794.850 2373.440 ;
        RECT 1408.590 2373.240 1408.910 2373.300 ;
        RECT 1794.530 2373.240 1794.850 2373.300 ;
        RECT 1408.590 2359.840 1408.910 2359.900 ;
        RECT 1787.630 2359.840 1787.950 2359.900 ;
        RECT 1408.590 2359.700 1787.950 2359.840 ;
        RECT 1408.590 2359.640 1408.910 2359.700 ;
        RECT 1787.630 2359.640 1787.950 2359.700 ;
        RECT 1408.590 2352.700 1408.910 2352.760 ;
        RECT 1780.270 2352.700 1780.590 2352.760 ;
        RECT 1408.590 2352.560 1780.590 2352.700 ;
        RECT 1408.590 2352.500 1408.910 2352.560 ;
        RECT 1780.270 2352.500 1780.590 2352.560 ;
        RECT 1408.590 2339.100 1408.910 2339.160 ;
        RECT 1773.370 2339.100 1773.690 2339.160 ;
        RECT 1408.590 2338.960 1773.690 2339.100 ;
        RECT 1408.590 2338.900 1408.910 2338.960 ;
        RECT 1773.370 2338.900 1773.690 2338.960 ;
        RECT 1408.590 2331.960 1408.910 2332.020 ;
        RECT 1766.470 2331.960 1766.790 2332.020 ;
        RECT 1408.590 2331.820 1766.790 2331.960 ;
        RECT 1408.590 2331.760 1408.910 2331.820 ;
        RECT 1766.470 2331.760 1766.790 2331.820 ;
        RECT 1408.590 2318.360 1408.910 2318.420 ;
        RECT 1760.030 2318.360 1760.350 2318.420 ;
        RECT 1408.590 2318.220 1760.350 2318.360 ;
        RECT 1408.590 2318.160 1408.910 2318.220 ;
        RECT 1760.030 2318.160 1760.350 2318.220 ;
        RECT 1408.590 2311.560 1408.910 2311.620 ;
        RECT 1760.950 2311.560 1761.270 2311.620 ;
        RECT 1408.590 2311.420 1761.270 2311.560 ;
        RECT 1408.590 2311.360 1408.910 2311.420 ;
        RECT 1760.950 2311.360 1761.270 2311.420 ;
        RECT 1408.590 2297.620 1408.910 2297.680 ;
        RECT 1752.670 2297.620 1752.990 2297.680 ;
        RECT 1408.590 2297.480 1752.990 2297.620 ;
        RECT 1408.590 2297.420 1408.910 2297.480 ;
        RECT 1752.670 2297.420 1752.990 2297.480 ;
        RECT 1408.590 2290.820 1408.910 2290.880 ;
        RECT 1745.770 2290.820 1746.090 2290.880 ;
        RECT 1408.590 2290.680 1746.090 2290.820 ;
        RECT 1408.590 2290.620 1408.910 2290.680 ;
        RECT 1745.770 2290.620 1746.090 2290.680 ;
        RECT 1408.590 2276.880 1408.910 2276.940 ;
        RECT 1738.870 2276.880 1739.190 2276.940 ;
        RECT 1408.590 2276.740 1739.190 2276.880 ;
        RECT 1408.590 2276.680 1408.910 2276.740 ;
        RECT 1738.870 2276.680 1739.190 2276.740 ;
        RECT 1408.590 2270.080 1408.910 2270.140 ;
        RECT 1731.970 2270.080 1732.290 2270.140 ;
        RECT 1408.590 2269.940 1732.290 2270.080 ;
        RECT 1408.590 2269.880 1408.910 2269.940 ;
        RECT 1731.970 2269.880 1732.290 2269.940 ;
        RECT 1408.590 2262.940 1408.910 2263.000 ;
        RECT 1725.070 2262.940 1725.390 2263.000 ;
        RECT 1408.590 2262.800 1725.390 2262.940 ;
        RECT 1408.590 2262.740 1408.910 2262.800 ;
        RECT 1725.070 2262.740 1725.390 2262.800 ;
        RECT 1408.590 2249.340 1408.910 2249.400 ;
        RECT 1718.630 2249.340 1718.950 2249.400 ;
        RECT 1408.590 2249.200 1718.950 2249.340 ;
        RECT 1408.590 2249.140 1408.910 2249.200 ;
        RECT 1718.630 2249.140 1718.950 2249.200 ;
        RECT 1408.590 2242.540 1408.910 2242.600 ;
        RECT 1718.170 2242.540 1718.490 2242.600 ;
        RECT 1408.590 2242.400 1718.490 2242.540 ;
        RECT 1408.590 2242.340 1408.910 2242.400 ;
        RECT 1718.170 2242.340 1718.490 2242.400 ;
        RECT 1408.590 2228.600 1408.910 2228.660 ;
        RECT 1711.270 2228.600 1711.590 2228.660 ;
        RECT 1408.590 2228.460 1711.590 2228.600 ;
        RECT 1408.590 2228.400 1408.910 2228.460 ;
        RECT 1711.270 2228.400 1711.590 2228.460 ;
        RECT 1408.590 2221.800 1408.910 2221.860 ;
        RECT 1704.370 2221.800 1704.690 2221.860 ;
        RECT 1408.590 2221.660 1704.690 2221.800 ;
        RECT 1408.590 2221.600 1408.910 2221.660 ;
        RECT 1704.370 2221.600 1704.690 2221.660 ;
        RECT 1408.590 2207.860 1408.910 2207.920 ;
        RECT 1697.470 2207.860 1697.790 2207.920 ;
        RECT 1408.590 2207.720 1697.790 2207.860 ;
        RECT 1408.590 2207.660 1408.910 2207.720 ;
        RECT 1697.470 2207.660 1697.790 2207.720 ;
        RECT 1408.590 2201.060 1408.910 2201.120 ;
        RECT 1690.570 2201.060 1690.890 2201.120 ;
        RECT 1408.590 2200.920 1690.890 2201.060 ;
        RECT 1408.590 2200.860 1408.910 2200.920 ;
        RECT 1690.570 2200.860 1690.890 2200.920 ;
        RECT 1408.590 2187.120 1408.910 2187.180 ;
        RECT 1684.130 2187.120 1684.450 2187.180 ;
        RECT 1408.590 2186.980 1684.450 2187.120 ;
        RECT 1408.590 2186.920 1408.910 2186.980 ;
        RECT 1684.130 2186.920 1684.450 2186.980 ;
        RECT 1408.590 2180.320 1408.910 2180.380 ;
        RECT 1683.670 2180.320 1683.990 2180.380 ;
        RECT 1408.590 2180.180 1683.990 2180.320 ;
        RECT 1408.590 2180.120 1408.910 2180.180 ;
        RECT 1683.670 2180.120 1683.990 2180.180 ;
        RECT 1408.590 2166.380 1408.910 2166.440 ;
        RECT 1676.770 2166.380 1677.090 2166.440 ;
        RECT 1408.590 2166.240 1677.090 2166.380 ;
        RECT 1408.590 2166.180 1408.910 2166.240 ;
        RECT 1676.770 2166.180 1677.090 2166.240 ;
        RECT 1408.590 2159.580 1408.910 2159.640 ;
        RECT 1669.870 2159.580 1670.190 2159.640 ;
        RECT 1408.590 2159.440 1670.190 2159.580 ;
        RECT 1408.590 2159.380 1408.910 2159.440 ;
        RECT 1669.870 2159.380 1670.190 2159.440 ;
        RECT 1408.590 2145.640 1408.910 2145.700 ;
        RECT 1662.970 2145.640 1663.290 2145.700 ;
        RECT 1408.590 2145.500 1663.290 2145.640 ;
        RECT 1408.590 2145.440 1408.910 2145.500 ;
        RECT 1662.970 2145.440 1663.290 2145.500 ;
        RECT 1408.590 2138.840 1408.910 2138.900 ;
        RECT 1656.070 2138.840 1656.390 2138.900 ;
        RECT 1408.590 2138.700 1656.390 2138.840 ;
        RECT 1408.590 2138.640 1408.910 2138.700 ;
        RECT 1656.070 2138.640 1656.390 2138.700 ;
        RECT 1408.590 2125.240 1408.910 2125.300 ;
        RECT 1649.630 2125.240 1649.950 2125.300 ;
        RECT 1408.590 2125.100 1649.950 2125.240 ;
        RECT 1408.590 2125.040 1408.910 2125.100 ;
        RECT 1649.630 2125.040 1649.950 2125.100 ;
        RECT 1408.590 2118.100 1408.910 2118.160 ;
        RECT 1649.170 2118.100 1649.490 2118.160 ;
        RECT 1408.590 2117.960 1649.490 2118.100 ;
        RECT 1408.590 2117.900 1408.910 2117.960 ;
        RECT 1649.170 2117.900 1649.490 2117.960 ;
        RECT 1408.590 2104.500 1408.910 2104.560 ;
        RECT 1642.270 2104.500 1642.590 2104.560 ;
        RECT 1408.590 2104.360 1642.590 2104.500 ;
        RECT 1408.590 2104.300 1408.910 2104.360 ;
        RECT 1642.270 2104.300 1642.590 2104.360 ;
        RECT 1408.590 2097.360 1408.910 2097.420 ;
        RECT 1635.370 2097.360 1635.690 2097.420 ;
        RECT 1408.590 2097.220 1635.690 2097.360 ;
        RECT 1408.590 2097.160 1408.910 2097.220 ;
        RECT 1635.370 2097.160 1635.690 2097.220 ;
        RECT 1408.590 2090.560 1408.910 2090.620 ;
        RECT 1628.470 2090.560 1628.790 2090.620 ;
        RECT 1408.590 2090.420 1628.790 2090.560 ;
        RECT 1408.590 2090.360 1408.910 2090.420 ;
        RECT 1628.470 2090.360 1628.790 2090.420 ;
        RECT 1408.590 2076.960 1408.910 2077.020 ;
        RECT 1621.570 2076.960 1621.890 2077.020 ;
        RECT 1408.590 2076.820 1621.890 2076.960 ;
        RECT 1408.590 2076.760 1408.910 2076.820 ;
        RECT 1621.570 2076.760 1621.890 2076.820 ;
        RECT 1408.590 2069.820 1408.910 2069.880 ;
        RECT 1614.670 2069.820 1614.990 2069.880 ;
        RECT 1408.590 2069.680 1614.990 2069.820 ;
        RECT 1408.590 2069.620 1408.910 2069.680 ;
        RECT 1614.670 2069.620 1614.990 2069.680 ;
        RECT 1426.530 2062.340 1426.850 2062.400 ;
        RECT 1580.170 2062.340 1580.490 2062.400 ;
        RECT 1426.530 2062.200 1580.490 2062.340 ;
        RECT 1426.530 2062.140 1426.850 2062.200 ;
        RECT 1580.170 2062.140 1580.490 2062.200 ;
        RECT 1408.130 2062.000 1408.450 2062.060 ;
        RECT 1624.790 2062.000 1625.110 2062.060 ;
        RECT 1408.130 2061.860 1625.110 2062.000 ;
        RECT 1408.130 2061.800 1408.450 2061.860 ;
        RECT 1624.790 2061.800 1625.110 2061.860 ;
        RECT 1407.670 2061.660 1407.990 2061.720 ;
        RECT 1631.690 2061.660 1632.010 2061.720 ;
        RECT 1407.670 2061.520 1632.010 2061.660 ;
        RECT 1407.670 2061.460 1407.990 2061.520 ;
        RECT 1631.690 2061.460 1632.010 2061.520 ;
        RECT 1409.985 2061.320 1410.275 2061.365 ;
        RECT 1638.590 2061.320 1638.910 2061.380 ;
        RECT 1409.985 2061.180 1638.910 2061.320 ;
        RECT 1409.985 2061.135 1410.275 2061.180 ;
        RECT 1638.590 2061.120 1638.910 2061.180 ;
        RECT 1415.490 2060.980 1415.810 2061.040 ;
        RECT 2192.890 2060.980 2193.210 2061.040 ;
        RECT 1415.490 2060.840 2193.210 2060.980 ;
        RECT 1415.490 2060.780 1415.810 2060.840 ;
        RECT 2192.890 2060.780 2193.210 2060.840 ;
        RECT 1415.030 2060.640 1415.350 2060.700 ;
        RECT 2192.430 2060.640 2192.750 2060.700 ;
        RECT 1415.030 2060.500 2192.750 2060.640 ;
        RECT 1415.030 2060.440 1415.350 2060.500 ;
        RECT 2192.430 2060.440 2192.750 2060.500 ;
        RECT 1415.950 2060.300 1416.270 2060.360 ;
        RECT 2193.350 2060.300 2193.670 2060.360 ;
        RECT 1415.950 2060.160 2193.670 2060.300 ;
        RECT 1415.950 2060.100 1416.270 2060.160 ;
        RECT 2193.350 2060.100 2193.670 2060.160 ;
        RECT 1416.410 2059.960 1416.730 2060.020 ;
        RECT 2228.770 2059.960 2229.090 2060.020 ;
        RECT 1416.410 2059.820 2229.090 2059.960 ;
        RECT 1416.410 2059.760 1416.730 2059.820 ;
        RECT 2228.770 2059.760 2229.090 2059.820 ;
        RECT 1426.990 2059.620 1427.310 2059.680 ;
        RECT 2266.490 2059.620 2266.810 2059.680 ;
        RECT 1426.990 2059.480 2266.810 2059.620 ;
        RECT 1426.990 2059.420 1427.310 2059.480 ;
        RECT 2266.490 2059.420 2266.810 2059.480 ;
        RECT 1408.590 2056.900 1408.910 2056.960 ;
        RECT 1409.970 2056.900 1410.290 2056.960 ;
        RECT 1408.590 2056.760 1410.290 2056.900 ;
        RECT 1408.590 2056.700 1408.910 2056.760 ;
        RECT 1409.970 2056.700 1410.290 2056.760 ;
        RECT 1409.970 2056.220 1410.290 2056.280 ;
        RECT 1607.770 2056.220 1608.090 2056.280 ;
        RECT 1409.970 2056.080 1608.090 2056.220 ;
        RECT 1409.970 2056.020 1410.290 2056.080 ;
        RECT 1607.770 2056.020 1608.090 2056.080 ;
        RECT 1426.070 2054.180 1426.390 2054.240 ;
        RECT 2190.590 2054.180 2190.910 2054.240 ;
        RECT 1426.070 2054.040 2190.910 2054.180 ;
        RECT 1426.070 2053.980 1426.390 2054.040 ;
        RECT 2190.590 2053.980 2190.910 2054.040 ;
        RECT 1425.610 2053.840 1425.930 2053.900 ;
        RECT 2191.050 2053.840 2191.370 2053.900 ;
        RECT 1425.610 2053.700 2191.370 2053.840 ;
        RECT 1425.610 2053.640 1425.930 2053.700 ;
        RECT 2191.050 2053.640 2191.370 2053.700 ;
        RECT 1425.150 2053.500 1425.470 2053.560 ;
        RECT 2191.510 2053.500 2191.830 2053.560 ;
        RECT 1425.150 2053.360 2191.830 2053.500 ;
        RECT 1425.150 2053.300 1425.470 2053.360 ;
        RECT 2191.510 2053.300 2191.830 2053.360 ;
        RECT 1416.870 2053.160 1417.190 2053.220 ;
        RECT 2193.810 2053.160 2194.130 2053.220 ;
        RECT 1416.870 2053.020 2194.130 2053.160 ;
        RECT 1416.870 2052.960 1417.190 2053.020 ;
        RECT 2193.810 2052.960 2194.130 2053.020 ;
        RECT 1409.970 2052.820 1410.290 2052.880 ;
        RECT 1409.775 2052.680 1410.290 2052.820 ;
        RECT 1409.970 2052.620 1410.290 2052.680 ;
        RECT 1414.570 2052.820 1414.890 2052.880 ;
        RECT 2191.970 2052.820 2192.290 2052.880 ;
        RECT 1414.570 2052.680 2192.290 2052.820 ;
        RECT 1414.570 2052.620 1414.890 2052.680 ;
        RECT 2191.970 2052.620 2192.290 2052.680 ;
        RECT 1407.670 2020.860 1407.990 2020.920 ;
        RECT 1409.970 2020.860 1410.290 2020.920 ;
        RECT 1407.670 2020.720 1410.290 2020.860 ;
        RECT 1407.670 2020.660 1407.990 2020.720 ;
        RECT 1409.970 2020.660 1410.290 2020.720 ;
        RECT 1407.670 1985.500 1407.990 1985.560 ;
        RECT 1417.330 1985.500 1417.650 1985.560 ;
        RECT 1407.670 1985.360 1417.650 1985.500 ;
        RECT 1407.670 1985.300 1407.990 1985.360 ;
        RECT 1417.330 1985.300 1417.650 1985.360 ;
        RECT 1409.510 1890.300 1409.830 1890.360 ;
        RECT 1426.990 1890.300 1427.310 1890.360 ;
        RECT 1409.510 1890.160 1427.310 1890.300 ;
        RECT 1409.510 1890.100 1409.830 1890.160 ;
        RECT 1426.990 1890.100 1427.310 1890.160 ;
        RECT 1414.110 1883.500 1414.430 1883.560 ;
        RECT 1473.450 1883.500 1473.770 1883.560 ;
        RECT 1414.110 1883.360 1473.770 1883.500 ;
        RECT 1414.110 1883.300 1414.430 1883.360 ;
        RECT 1473.450 1883.300 1473.770 1883.360 ;
        RECT 1414.110 1869.900 1414.430 1869.960 ;
        RECT 1459.190 1869.900 1459.510 1869.960 ;
        RECT 1414.110 1869.760 1459.510 1869.900 ;
        RECT 1414.110 1869.700 1414.430 1869.760 ;
        RECT 1459.190 1869.700 1459.510 1869.760 ;
        RECT 1414.110 1862.760 1414.430 1862.820 ;
        RECT 1452.290 1862.760 1452.610 1862.820 ;
        RECT 1414.110 1862.620 1452.610 1862.760 ;
        RECT 1414.110 1862.560 1414.430 1862.620 ;
        RECT 1452.290 1862.560 1452.610 1862.620 ;
        RECT 1411.810 1855.280 1412.130 1855.340 ;
        RECT 1438.490 1855.280 1438.810 1855.340 ;
        RECT 1411.810 1855.140 1438.810 1855.280 ;
        RECT 1411.810 1855.080 1412.130 1855.140 ;
        RECT 1438.490 1855.080 1438.810 1855.140 ;
        RECT 1411.350 1840.320 1411.670 1840.380 ;
        RECT 1431.590 1840.320 1431.910 1840.380 ;
        RECT 1411.350 1840.180 1431.910 1840.320 ;
        RECT 1411.350 1840.120 1411.670 1840.180 ;
        RECT 1431.590 1840.120 1431.910 1840.180 ;
        RECT 1408.590 1829.100 1408.910 1829.160 ;
        RECT 1424.690 1829.100 1425.010 1829.160 ;
        RECT 1408.590 1828.960 1425.010 1829.100 ;
        RECT 1408.590 1828.900 1408.910 1828.960 ;
        RECT 1424.690 1828.900 1425.010 1828.960 ;
        RECT 1414.110 1821.620 1414.430 1821.680 ;
        RECT 1472.990 1821.620 1473.310 1821.680 ;
        RECT 1414.110 1821.480 1473.310 1821.620 ;
        RECT 1414.110 1821.420 1414.430 1821.480 ;
        RECT 1472.990 1821.420 1473.310 1821.480 ;
        RECT 1409.510 1814.480 1409.830 1814.540 ;
        RECT 1426.530 1814.480 1426.850 1814.540 ;
        RECT 1409.510 1814.340 1426.850 1814.480 ;
        RECT 1409.510 1814.280 1409.830 1814.340 ;
        RECT 1426.530 1814.280 1426.850 1814.340 ;
        RECT 1409.510 1800.880 1409.830 1800.940 ;
        RECT 1426.070 1800.880 1426.390 1800.940 ;
        RECT 1409.510 1800.740 1426.390 1800.880 ;
        RECT 1409.510 1800.680 1409.830 1800.740 ;
        RECT 1426.070 1800.680 1426.390 1800.740 ;
        RECT 1408.590 1788.300 1408.910 1788.360 ;
        RECT 1425.610 1788.300 1425.930 1788.360 ;
        RECT 1408.590 1788.160 1425.930 1788.300 ;
        RECT 1408.590 1788.100 1408.910 1788.160 ;
        RECT 1425.610 1788.100 1425.930 1788.160 ;
        RECT 1410.430 1779.460 1410.750 1779.520 ;
        RECT 1425.150 1779.460 1425.470 1779.520 ;
        RECT 1410.430 1779.320 1425.470 1779.460 ;
        RECT 1410.430 1779.260 1410.750 1779.320 ;
        RECT 1425.150 1779.260 1425.470 1779.320 ;
        RECT 1407.670 1730.500 1407.990 1730.560 ;
        RECT 1416.410 1730.500 1416.730 1730.560 ;
        RECT 1407.670 1730.360 1416.730 1730.500 ;
        RECT 1407.670 1730.300 1407.990 1730.360 ;
        RECT 1416.410 1730.300 1416.730 1730.360 ;
        RECT 1414.110 1717.920 1414.430 1717.980 ;
        RECT 1514.390 1717.920 1514.710 1717.980 ;
        RECT 1414.110 1717.780 1514.710 1717.920 ;
        RECT 1414.110 1717.720 1414.430 1717.780 ;
        RECT 1514.390 1717.720 1514.710 1717.780 ;
        RECT 1407.670 1706.700 1407.990 1706.760 ;
        RECT 1416.870 1706.700 1417.190 1706.760 ;
        RECT 1407.670 1706.560 1417.190 1706.700 ;
        RECT 1407.670 1706.500 1407.990 1706.560 ;
        RECT 1416.870 1706.500 1417.190 1706.560 ;
        RECT 1408.590 1696.500 1408.910 1696.560 ;
        RECT 1421.010 1696.500 1421.330 1696.560 ;
        RECT 1408.590 1696.360 1421.330 1696.500 ;
        RECT 1408.590 1696.300 1408.910 1696.360 ;
        RECT 1421.010 1696.300 1421.330 1696.360 ;
        RECT 1407.670 1688.000 1407.990 1688.060 ;
        RECT 1420.550 1688.000 1420.870 1688.060 ;
        RECT 1407.670 1687.860 1420.870 1688.000 ;
        RECT 1407.670 1687.800 1407.990 1687.860 ;
        RECT 1420.550 1687.800 1420.870 1687.860 ;
        RECT 1408.130 1676.100 1408.450 1676.160 ;
        RECT 1420.090 1676.100 1420.410 1676.160 ;
        RECT 1408.130 1675.960 1420.410 1676.100 ;
        RECT 1408.130 1675.900 1408.450 1675.960 ;
        RECT 1420.090 1675.900 1420.410 1675.960 ;
        RECT 1407.670 1666.240 1407.990 1666.300 ;
        RECT 1419.630 1666.240 1419.950 1666.300 ;
        RECT 1407.670 1666.100 1419.950 1666.240 ;
        RECT 1407.670 1666.040 1407.990 1666.100 ;
        RECT 1419.630 1666.040 1419.950 1666.100 ;
        RECT 1407.670 1655.700 1407.990 1655.760 ;
        RECT 1419.170 1655.700 1419.490 1655.760 ;
        RECT 1407.670 1655.560 1419.490 1655.700 ;
        RECT 1407.670 1655.500 1407.990 1655.560 ;
        RECT 1419.170 1655.500 1419.490 1655.560 ;
        RECT 1407.670 1645.500 1407.990 1645.560 ;
        RECT 1418.710 1645.500 1419.030 1645.560 ;
        RECT 1407.670 1645.360 1419.030 1645.500 ;
        RECT 1407.670 1645.300 1407.990 1645.360 ;
        RECT 1418.710 1645.300 1419.030 1645.360 ;
        RECT 1407.670 1635.300 1407.990 1635.360 ;
        RECT 1418.250 1635.300 1418.570 1635.360 ;
        RECT 1407.670 1635.160 1418.570 1635.300 ;
        RECT 1407.670 1635.100 1407.990 1635.160 ;
        RECT 1418.250 1635.100 1418.570 1635.160 ;
        RECT 1407.670 1625.440 1407.990 1625.500 ;
        RECT 1417.790 1625.440 1418.110 1625.500 ;
        RECT 1407.670 1625.300 1418.110 1625.440 ;
        RECT 1407.670 1625.240 1407.990 1625.300 ;
        RECT 1417.790 1625.240 1418.110 1625.300 ;
      LAYER met1 ;
        RECT 1555.000 1605.000 1931.480 2051.235 ;
        RECT 2205.000 1605.000 2581.480 2051.235 ;
        RECT 1550.000 410.640 2646.500 1495.780 ;
      LAYER via ;
        RECT 1324.440 3266.760 1324.700 3267.020 ;
        RECT 1890.700 3266.760 1890.960 3267.020 ;
        RECT 1917.840 3266.760 1918.100 3267.020 ;
        RECT 2542.060 3266.760 2542.320 3267.020 ;
        RECT 1295.920 3264.380 1296.180 3264.640 ;
        RECT 1318.000 3264.380 1318.260 3264.640 ;
        RECT 1324.440 3264.380 1324.700 3264.640 ;
        RECT 1890.700 3264.380 1890.960 3264.640 ;
        RECT 1917.840 3264.380 1918.100 3264.640 ;
        RECT 2542.060 3264.040 2542.320 3264.300 ;
        RECT 2566.900 3264.040 2567.160 3264.300 ;
        RECT 646.400 3263.700 646.660 3263.960 ;
        RECT 668.480 3263.700 668.740 3263.960 ;
        RECT 697.000 3263.700 697.260 3263.960 ;
        RECT 2594.500 3263.700 2594.760 3263.960 ;
        RECT 688.260 3252.140 688.520 3252.400 ;
        RECT 1332.260 3252.480 1332.520 3252.740 ;
        RECT 1414.140 3252.140 1414.400 3252.400 ;
        RECT 2582.080 3252.140 2582.340 3252.400 ;
        RECT 697.000 2897.860 697.260 2898.120 ;
        RECT 938.500 2897.860 938.760 2898.120 ;
        RECT 1332.260 3251.120 1332.520 3251.380 ;
        RECT 1411.380 3250.780 1411.640 3251.040 ;
        RECT 1414.140 3250.780 1414.400 3251.040 ;
        RECT 1473.480 3229.360 1473.740 3229.620 ;
        RECT 1536.960 3229.360 1537.220 3229.620 ;
        RECT 1459.220 3222.220 1459.480 3222.480 ;
        RECT 1535.580 3222.220 1535.840 3222.480 ;
        RECT 1452.320 3215.420 1452.580 3215.680 ;
        RECT 1535.580 3215.420 1535.840 3215.680 ;
        RECT 1438.520 3208.620 1438.780 3208.880 ;
        RECT 1538.340 3208.620 1538.600 3208.880 ;
        RECT 1431.620 3201.480 1431.880 3201.740 ;
        RECT 1538.340 3201.480 1538.600 3201.740 ;
        RECT 1424.720 3194.680 1424.980 3194.940 ;
        RECT 1533.280 3194.680 1533.540 3194.940 ;
        RECT 1473.020 3187.880 1473.280 3188.140 ;
        RECT 1534.200 3187.880 1534.460 3188.140 ;
        RECT 1514.420 2898.200 1514.680 2898.460 ;
        RECT 1534.660 2898.200 1534.920 2898.460 ;
        RECT 1410.920 2894.460 1411.180 2894.720 ;
        RECT 1538.340 2894.460 1538.600 2894.720 ;
        RECT 1935.780 3251.120 1936.040 3251.380 ;
        RECT 1945.900 2901.260 1946.160 2901.520 ;
        RECT 2189.240 2901.260 2189.500 2901.520 ;
        RECT 330.840 2794.160 331.100 2794.420 ;
        RECT 1001.060 2794.160 1001.320 2794.420 ;
        RECT 1410.460 2794.160 1410.720 2794.420 ;
        RECT 337.280 2793.820 337.540 2794.080 ;
        RECT 1007.500 2793.820 1007.760 2794.080 ;
        RECT 1100.420 2793.820 1100.680 2794.080 ;
        RECT 1146.880 2793.820 1147.140 2794.080 ;
        RECT 397.540 2793.480 397.800 2793.740 ;
        RECT 444.460 2793.480 444.720 2793.740 ;
        RECT 492.760 2793.480 493.020 2793.740 ;
        RECT 524.500 2793.480 524.760 2793.740 ;
        RECT 627.540 2793.480 627.800 2793.740 ;
        RECT 1042.460 2793.480 1042.720 2793.740 ;
        RECT 1055.800 2793.480 1056.060 2793.740 ;
        RECT 1089.840 2793.480 1090.100 2793.740 ;
        RECT 1129.860 2793.480 1130.120 2793.740 ;
        RECT 1173.100 2793.480 1173.360 2793.740 ;
        RECT 392.480 2793.140 392.740 2793.400 ;
        RECT 439.400 2793.140 439.660 2793.400 ;
        RECT 485.400 2793.140 485.660 2793.400 ;
        RECT 386.960 2792.800 387.220 2793.060 ;
        RECT 433.420 2792.800 433.680 2793.060 ;
        RECT 379.600 2792.460 379.860 2792.720 ;
        RECT 426.980 2792.460 427.240 2792.720 ;
        RECT 474.360 2792.800 474.620 2793.060 ;
        RECT 510.240 2793.140 510.500 2793.400 ;
        RECT 700.220 2793.140 700.480 2793.400 ;
        RECT 1103.640 2793.140 1103.900 2793.400 ;
        RECT 1136.300 2793.140 1136.560 2793.400 ;
        RECT 1180.000 2793.140 1180.260 2793.400 ;
        RECT 1419.660 2794.160 1419.920 2794.420 ;
        RECT 1587.100 2794.160 1587.360 2794.420 ;
        RECT 1631.720 2794.160 1631.980 2794.420 ;
        RECT 1671.280 2794.160 1671.540 2794.420 ;
        RECT 1718.200 2794.160 1718.460 2794.420 ;
        RECT 1723.720 2794.160 1723.980 2794.420 ;
        RECT 1724.180 2794.160 1724.440 2794.420 ;
        RECT 1766.500 2794.160 1766.760 2794.420 ;
        RECT 2232.020 2794.160 2232.280 2794.420 ;
        RECT 2402.680 2794.160 2402.940 2794.420 ;
        RECT 1421.040 2793.820 1421.300 2794.080 ;
        RECT 1601.360 2793.820 1601.620 2794.080 ;
        RECT 1662.540 2793.820 1662.800 2794.080 ;
        RECT 1706.240 2793.820 1706.500 2794.080 ;
        RECT 1752.700 2793.820 1752.960 2794.080 ;
        RECT 2208.100 2793.820 2208.360 2794.080 ;
        RECT 2286.760 2793.820 2287.020 2794.080 ;
        RECT 2332.760 2793.820 2333.020 2794.080 ;
        RECT 2377.380 2793.820 2377.640 2794.080 ;
        RECT 2415.100 2793.820 2415.360 2794.080 ;
        RECT 1420.580 2793.480 1420.840 2793.740 ;
        RECT 1600.900 2793.480 1601.160 2793.740 ;
        RECT 1624.820 2793.480 1625.080 2793.740 ;
        RECT 1671.280 2793.480 1671.540 2793.740 ;
        RECT 1681.400 2793.480 1681.660 2793.740 ;
        RECT 1728.780 2793.480 1729.040 2793.740 ;
        RECT 1746.720 2793.480 1746.980 2793.740 ;
        RECT 2268.360 2793.480 2268.620 2793.740 ;
        RECT 2312.980 2793.480 2313.240 2793.740 ;
        RECT 2360.820 2793.480 2361.080 2793.740 ;
        RECT 2408.200 2793.480 2408.460 2793.740 ;
        RECT 1614.240 2793.140 1614.500 2793.400 ;
        RECT 1638.620 2793.140 1638.880 2793.400 ;
        RECT 403.980 2792.120 404.240 2792.380 ;
        RECT 433.420 2792.120 433.680 2792.380 ;
        RECT 478.500 2792.460 478.760 2792.720 ;
        RECT 513.920 2792.800 514.180 2793.060 ;
        RECT 524.040 2792.800 524.300 2793.060 ;
        RECT 720.920 2792.800 721.180 2793.060 ;
        RECT 1062.700 2792.800 1062.960 2793.060 ;
        RECT 1065.460 2792.800 1065.720 2793.060 ;
        RECT 1111.460 2792.800 1111.720 2793.060 ;
        RECT 1159.300 2792.800 1159.560 2793.060 ;
        RECT 1462.900 2792.800 1463.160 2793.060 ;
        RECT 1617.460 2792.800 1617.720 2793.060 ;
        RECT 1665.760 2792.800 1666.020 2793.060 ;
        RECT 1669.440 2792.800 1669.700 2793.060 ;
        RECT 1679.560 2793.140 1679.820 2793.400 ;
        RECT 1724.180 2793.140 1724.440 2793.400 ;
        RECT 1681.400 2792.800 1681.660 2793.060 ;
        RECT 1683.700 2792.800 1683.960 2793.060 ;
        RECT 1688.760 2792.800 1689.020 2793.060 ;
        RECT 1732.460 2793.140 1732.720 2793.400 ;
        RECT 1780.300 2793.140 1780.560 2793.400 ;
        RECT 2091.260 2793.140 2091.520 2793.400 ;
        RECT 2270.200 2793.140 2270.460 2793.400 ;
        RECT 2273.420 2793.140 2273.680 2793.400 ;
        RECT 1773.400 2792.800 1773.660 2793.060 ;
        RECT 2279.860 2792.800 2280.120 2793.060 ;
        RECT 2326.320 2793.140 2326.580 2793.400 ;
        RECT 2374.160 2793.140 2374.420 2793.400 ;
        RECT 2314.820 2792.800 2315.080 2793.060 ;
        RECT 2343.340 2792.800 2343.600 2793.060 ;
        RECT 2377.380 2792.800 2377.640 2793.060 ;
        RECT 2422.000 2792.800 2422.260 2793.060 ;
        RECT 520.820 2792.460 521.080 2792.720 ;
        RECT 542.440 2792.460 542.700 2792.720 ;
        RECT 741.620 2792.460 741.880 2792.720 ;
        RECT 1093.980 2792.460 1094.240 2792.720 ;
        RECT 1140.440 2792.460 1140.700 2792.720 ;
        RECT 1186.900 2792.460 1187.160 2792.720 ;
        RECT 1420.120 2792.460 1420.380 2792.720 ;
        RECT 1510.740 2792.460 1511.000 2792.720 ;
        RECT 1594.000 2792.460 1594.260 2792.720 ;
        RECT 2258.700 2792.460 2258.960 2792.720 ;
        RECT 2261.920 2792.460 2262.180 2792.720 ;
        RECT 449.060 2792.120 449.320 2792.380 ;
        RECT 496.900 2792.120 497.160 2792.380 ;
        RECT 500.580 2792.120 500.840 2792.380 ;
        RECT 502.880 2792.120 503.140 2792.380 ;
        RECT 700.680 2792.120 700.940 2792.380 ;
        RECT 1409.540 2792.120 1409.800 2792.380 ;
        RECT 1647.820 2792.120 1648.080 2792.380 ;
        RECT 1695.200 2792.120 1695.460 2792.380 ;
        RECT 368.560 2791.780 368.820 2792.040 ;
        RECT 414.560 2791.780 414.820 2792.040 ;
        RECT 488.160 2791.780 488.420 2792.040 ;
        RECT 693.320 2791.780 693.580 2792.040 ;
        RECT 1055.800 2791.780 1056.060 2792.040 ;
        RECT 1059.480 2791.780 1059.740 2792.040 ;
        RECT 1105.480 2791.780 1105.740 2792.040 ;
        RECT 1152.400 2791.780 1152.660 2792.040 ;
        RECT 407.200 2791.440 407.460 2791.700 ;
        RECT 409.960 2791.440 410.220 2791.700 ;
        RECT 455.500 2791.440 455.760 2791.700 ;
        RECT 461.480 2791.440 461.740 2791.700 ;
        RECT 687.340 2791.440 687.600 2791.700 ;
        RECT 1031.880 2791.440 1032.140 2791.700 ;
        RECT 1076.500 2791.440 1076.760 2791.700 ;
        RECT 1119.740 2791.440 1120.000 2791.700 ;
        RECT 1166.200 2791.440 1166.460 2791.700 ;
        RECT 1410.000 2791.780 1410.260 2792.040 ;
        RECT 1642.760 2791.780 1643.020 2792.040 ;
        RECT 1683.700 2791.780 1683.960 2792.040 ;
        RECT 1732.460 2792.120 1732.720 2792.380 ;
        RECT 1741.200 2792.120 1741.460 2792.380 ;
        RECT 1787.200 2792.120 1787.460 2792.380 ;
        RECT 1790.420 2792.120 1790.680 2792.380 ;
        RECT 2263.300 2792.120 2263.560 2792.380 ;
        RECT 2269.740 2792.460 2270.000 2792.720 ;
        RECT 2308.380 2792.460 2308.640 2792.720 ;
        RECT 2356.680 2792.460 2356.940 2792.720 ;
        RECT 2401.760 2792.460 2402.020 2792.720 ;
        RECT 2297.340 2792.120 2297.600 2792.380 ;
        RECT 2340.120 2792.120 2340.380 2792.380 ;
        RECT 2343.800 2792.120 2344.060 2792.380 ;
        RECT 2350.240 2792.120 2350.500 2792.380 ;
        RECT 2387.960 2792.120 2388.220 2792.380 ;
        RECT 1193.800 2791.440 1194.060 2791.700 ;
        RECT 1409.080 2791.440 1409.340 2791.700 ;
        RECT 1652.420 2791.440 1652.680 2791.700 ;
        RECT 371.320 2791.100 371.580 2791.360 ;
        RECT 686.880 2791.100 687.140 2791.360 ;
        RECT 1614.240 2791.100 1614.500 2791.360 ;
        RECT 1662.540 2791.100 1662.800 2791.360 ;
        RECT 1669.440 2791.440 1669.700 2791.700 ;
        RECT 1712.680 2791.440 1712.940 2791.700 ;
        RECT 1742.120 2791.780 1742.380 2792.040 ;
        RECT 1797.320 2791.780 1797.580 2792.040 ;
        RECT 2380.600 2791.780 2380.860 2792.040 ;
        RECT 2381.520 2791.780 2381.780 2792.040 ;
        RECT 2385.660 2791.780 2385.920 2792.040 ;
        RECT 2428.900 2791.780 2429.160 2792.040 ;
        RECT 1746.720 2791.440 1746.980 2791.700 ;
        RECT 1788.580 2791.440 1788.840 2791.700 ;
        RECT 1797.780 2791.440 1798.040 2791.700 ;
        RECT 2387.500 2791.440 2387.760 2791.700 ;
        RECT 1699.340 2791.100 1699.600 2791.360 ;
        RECT 1723.720 2791.100 1723.980 2791.360 ;
        RECT 1760.060 2791.100 1760.320 2791.360 ;
        RECT 1790.880 2791.100 1791.140 2791.360 ;
        RECT 2381.060 2791.100 2381.320 2791.360 ;
        RECT 2387.960 2791.100 2388.220 2791.360 ;
        RECT 2391.180 2791.100 2391.440 2791.360 ;
        RECT 2435.800 2791.100 2436.060 2791.360 ;
        RECT 362.580 2790.760 362.840 2791.020 ;
        RECT 407.200 2790.760 407.460 2791.020 ;
        RECT 419.160 2790.760 419.420 2791.020 ;
        RECT 748.520 2790.760 748.780 2791.020 ;
        RECT 1019.000 2790.760 1019.260 2791.020 ;
        RECT 1062.700 2790.760 1062.960 2791.020 ;
        RECT 1159.760 2790.760 1160.020 2791.020 ;
        RECT 1417.820 2790.760 1418.080 2791.020 ;
        RECT 2238.000 2790.760 2238.260 2791.020 ;
        RECT 384.200 2790.420 384.460 2790.680 ;
        RECT 727.820 2790.420 728.080 2790.680 ;
        RECT 1069.600 2790.420 1069.860 2790.680 ;
        RECT 1418.740 2790.420 1419.000 2790.680 ;
        RECT 2091.260 2790.420 2091.520 2790.680 ;
        RECT 2249.500 2790.420 2249.760 2790.680 ;
        RECT 406.280 2790.080 406.540 2790.340 ;
        RECT 762.780 2790.080 763.040 2790.340 ;
        RECT 1419.200 2790.080 1419.460 2790.340 ;
        RECT 2090.800 2790.080 2091.060 2790.340 ;
        RECT 2163.020 2790.080 2163.280 2790.340 ;
        RECT 2256.400 2790.080 2256.660 2790.340 ;
        RECT 396.620 2789.740 396.880 2790.000 ;
        RECT 762.320 2789.740 762.580 2790.000 ;
        RECT 1117.900 2789.740 1118.160 2790.000 ;
        RECT 1411.380 2789.740 1411.640 2790.000 ;
        RECT 2218.220 2789.740 2218.480 2790.000 ;
        RECT 2394.400 2790.760 2394.660 2791.020 ;
        RECT 2394.860 2790.760 2395.120 2791.020 ;
        RECT 2442.700 2790.760 2442.960 2791.020 ;
        RECT 375.000 2789.400 375.260 2789.660 ;
        RECT 421.000 2789.400 421.260 2789.660 ;
        RECT 449.060 2789.400 449.320 2789.660 ;
        RECT 468.840 2789.400 469.100 2789.660 ;
        RECT 686.420 2789.400 686.680 2789.660 ;
        RECT 1010.720 2789.400 1010.980 2789.660 ;
        RECT 1055.800 2789.400 1056.060 2789.660 ;
        RECT 1411.840 2789.400 1412.100 2789.660 ;
        RECT 2245.820 2789.400 2246.080 2789.660 ;
        RECT 2415.100 2790.420 2415.360 2790.680 ;
        RECT 538.300 2789.060 538.560 2789.320 ;
        RECT 1042.460 2789.060 1042.720 2789.320 ;
        RECT 1412.300 2789.060 1412.560 2789.320 ;
        RECT 446.760 2788.720 447.020 2788.980 ;
        RECT 485.400 2788.720 485.660 2788.980 ;
        RECT 531.400 2788.720 531.660 2788.980 ;
        RECT 606.840 2788.720 607.100 2788.980 ;
        RECT 1031.880 2788.720 1032.140 2788.980 ;
        RECT 1038.320 2788.720 1038.580 2788.980 ;
        RECT 1089.840 2788.720 1090.100 2788.980 ;
        RECT 1412.760 2788.720 1413.020 2788.980 ;
        RECT 455.500 2788.380 455.760 2788.640 ;
        RECT 500.120 2788.380 500.380 2788.640 ;
        RECT 500.580 2788.380 500.840 2788.640 ;
        RECT 541.520 2788.380 541.780 2788.640 ;
        RECT 586.140 2788.380 586.400 2788.640 ;
        RECT 1019.000 2788.380 1019.260 2788.640 ;
        RECT 1024.520 2788.380 1024.780 2788.640 ;
        RECT 1069.600 2788.380 1069.860 2788.640 ;
        RECT 1413.220 2788.380 1413.480 2788.640 ;
        RECT 462.400 2788.040 462.660 2788.300 ;
        RECT 504.260 2788.040 504.520 2788.300 ;
        RECT 421.000 2787.700 421.260 2787.960 ;
        RECT 467.920 2787.700 468.180 2787.960 ;
        RECT 537.380 2787.700 537.640 2787.960 ;
        RECT 648.700 2788.040 648.960 2788.300 ;
        RECT 1052.580 2788.040 1052.840 2788.300 ;
        RECT 1100.420 2788.040 1100.680 2788.300 ;
        RECT 1413.680 2788.040 1413.940 2788.300 ;
        RECT 2238.920 2789.060 2239.180 2789.320 ;
        RECT 2408.200 2790.080 2408.460 2790.340 ;
        RECT 2291.360 2789.740 2291.620 2790.000 ;
        RECT 2297.340 2789.740 2297.600 2790.000 ;
        RECT 2304.240 2789.740 2304.500 2790.000 ;
        RECT 2343.800 2789.740 2344.060 2790.000 ;
        RECT 2394.860 2789.740 2395.120 2790.000 ;
        RECT 2273.420 2789.400 2273.680 2789.660 ;
        RECT 2321.720 2789.400 2321.980 2789.660 ;
        RECT 2442.700 2789.400 2442.960 2789.660 ;
        RECT 2435.800 2789.060 2436.060 2789.320 ;
        RECT 2259.620 2788.720 2259.880 2788.980 ;
        RECT 2422.000 2788.720 2422.260 2788.980 ;
        RECT 2252.720 2788.380 2252.980 2788.640 ;
        RECT 2415.560 2788.380 2415.820 2788.640 ;
        RECT 2267.440 2788.040 2267.700 2788.300 ;
        RECT 2428.900 2788.040 2429.160 2788.300 ;
        RECT 707.120 2787.700 707.380 2787.960 ;
        RECT 1045.220 2787.700 1045.480 2787.960 ;
        RECT 1093.980 2787.700 1094.240 2787.960 ;
        RECT 1414.140 2787.700 1414.400 2787.960 ;
        RECT 2091.720 2787.700 2091.980 2787.960 ;
        RECT 2162.560 2787.700 2162.820 2787.960 ;
        RECT 2208.100 2787.700 2208.360 2787.960 ;
        RECT 2270.200 2787.700 2270.460 2787.960 ;
        RECT 2298.260 2787.700 2298.520 2787.960 ;
        RECT 2321.260 2787.700 2321.520 2787.960 ;
        RECT 2367.260 2787.700 2367.520 2787.960 ;
        RECT 2373.240 2787.700 2373.500 2787.960 ;
        RECT 2381.520 2787.700 2381.780 2787.960 ;
        RECT 2381.980 2787.700 2382.240 2787.960 ;
        RECT 2415.100 2787.700 2415.360 2787.960 ;
        RECT 658.820 2787.360 659.080 2787.620 ;
        RECT 1417.360 2787.360 1417.620 2787.620 ;
        RECT 482.640 2725.140 482.900 2725.400 ;
        RECT 948.160 2725.140 948.420 2725.400 ;
        RECT 470.680 2724.800 470.940 2725.060 ;
        RECT 942.180 2724.800 942.440 2725.060 ;
        RECT 510.240 2724.460 510.500 2724.720 ;
        RECT 989.560 2724.460 989.820 2724.720 ;
        RECT 460.560 2724.120 460.820 2724.380 ;
        RECT 942.640 2724.120 942.900 2724.380 ;
        RECT 449.980 2723.780 450.240 2724.040 ;
        RECT 943.100 2723.780 943.360 2724.040 ;
        RECT 530.940 2723.440 531.200 2723.700 ;
        RECT 1030.960 2723.440 1031.220 2723.700 ;
        RECT 439.860 2723.100 440.120 2723.360 ;
        RECT 943.560 2723.100 943.820 2723.360 ;
        RECT 551.640 2722.760 551.900 2723.020 ;
        RECT 1062.240 2722.760 1062.500 2723.020 ;
        RECT 429.280 2722.420 429.540 2722.680 ;
        RECT 944.020 2722.420 944.280 2722.680 ;
        RECT 419.160 2722.080 419.420 2722.340 ;
        RECT 944.480 2722.080 944.740 2722.340 ;
        RECT 408.580 2721.740 408.840 2722.000 ;
        RECT 979.900 2721.740 980.160 2722.000 ;
        RECT 433.880 2721.400 434.140 2721.660 ;
        RECT 865.360 2721.400 865.620 2721.660 ;
        RECT 441.240 2721.060 441.500 2721.320 ;
        RECT 875.480 2721.060 875.740 2721.320 ;
        RECT 434.340 2720.720 434.600 2720.980 ;
        RECT 854.780 2720.720 855.040 2720.980 ;
        RECT 427.440 2720.380 427.700 2720.640 ;
        RECT 844.200 2720.380 844.460 2720.640 ;
        RECT 413.640 2720.040 413.900 2720.300 ;
        RECT 823.500 2720.040 823.760 2720.300 ;
        RECT 365.340 2719.700 365.600 2719.960 ;
        RECT 740.700 2719.700 740.960 2719.960 ;
        RECT 289.440 2719.360 289.700 2719.620 ;
        RECT 564.060 2719.360 564.320 2719.620 ;
        RECT 288.980 2719.020 289.240 2719.280 ;
        RECT 553.940 2719.020 554.200 2719.280 ;
        RECT 1103.640 2718.680 1103.900 2718.940 ;
        RECT 358.440 2718.340 358.700 2718.600 ;
        RECT 377.300 2718.340 377.560 2718.600 ;
        RECT 379.140 2718.340 379.400 2718.600 ;
        RECT 727.820 2718.340 728.080 2718.600 ;
        RECT 762.780 2718.340 763.040 2718.600 ;
        RECT 813.380 2718.340 813.640 2718.600 ;
        RECT 1027.740 2718.340 1028.000 2718.600 ;
        RECT 1093.520 2718.340 1093.780 2718.600 ;
        RECT 1102.720 2718.340 1102.980 2718.600 ;
        RECT 1138.140 2718.340 1138.400 2718.600 ;
        RECT 1290.400 2718.340 1290.660 2718.600 ;
        RECT 392.940 2718.000 393.200 2718.260 ;
        RECT 782.100 2718.000 782.360 2718.260 ;
        RECT 1034.640 2718.000 1034.900 2718.260 ;
        RECT 1103.640 2718.000 1103.900 2718.260 ;
        RECT 1145.040 2718.000 1145.300 2718.260 ;
        RECT 1300.980 2718.000 1301.240 2718.260 ;
        RECT 305.080 2717.660 305.340 2717.920 ;
        RECT 310.140 2717.660 310.400 2717.920 ;
        RECT 325.780 2717.660 326.040 2717.920 ;
        RECT 330.840 2717.660 331.100 2717.920 ;
        RECT 351.540 2717.660 351.800 2717.920 ;
        RECT 356.600 2717.660 356.860 2717.920 ;
        RECT 399.840 2717.660 400.100 2717.920 ;
        RECT 762.320 2717.660 762.580 2717.920 ;
        RECT 792.680 2717.660 792.940 2717.920 ;
        RECT 1041.540 2717.660 1041.800 2717.920 ;
        RECT 1114.220 2717.660 1114.480 2717.920 ;
        RECT 1151.940 2717.660 1152.200 2717.920 ;
        RECT 1311.100 2717.660 1311.360 2717.920 ;
        RECT 287.140 2717.320 287.400 2717.580 ;
        RECT 512.540 2717.320 512.800 2717.580 ;
        RECT 636.740 2717.320 637.000 2717.580 ;
        RECT 1045.220 2717.320 1045.480 2717.580 ;
        RECT 1048.440 2717.320 1048.700 2717.580 ;
        RECT 1124.340 2717.320 1124.600 2717.580 ;
        RECT 1158.840 2717.320 1159.100 2717.580 ;
        RECT 1321.680 2717.320 1321.940 2717.580 ;
        RECT 287.600 2716.980 287.860 2717.240 ;
        RECT 522.660 2716.980 522.920 2717.240 ;
        RECT 616.040 2716.980 616.300 2717.240 ;
        RECT 1038.320 2716.980 1038.580 2717.240 ;
        RECT 1054.880 2716.980 1055.140 2717.240 ;
        RECT 1134.920 2716.980 1135.180 2717.240 ;
        RECT 1165.740 2716.980 1166.000 2717.240 ;
        RECT 1332.260 2716.980 1332.520 2717.240 ;
        RECT 288.060 2716.640 288.320 2716.900 ;
        RECT 533.240 2716.640 533.500 2716.900 ;
        RECT 595.340 2716.640 595.600 2716.900 ;
        RECT 1024.520 2716.640 1024.780 2716.900 ;
        RECT 1061.780 2716.640 1062.040 2716.900 ;
        RECT 1155.620 2716.640 1155.880 2716.900 ;
        RECT 1165.280 2716.640 1165.540 2716.900 ;
        RECT 1342.380 2716.640 1342.640 2716.900 ;
        RECT 455.040 2716.300 455.300 2716.560 ;
        RECT 896.180 2716.300 896.440 2716.560 ;
        RECT 1076.040 2716.300 1076.300 2716.560 ;
        RECT 1176.320 2716.300 1176.580 2716.560 ;
        RECT 1179.540 2716.300 1179.800 2716.560 ;
        RECT 1363.080 2716.300 1363.340 2716.560 ;
        RECT 288.520 2715.960 288.780 2716.220 ;
        RECT 543.360 2715.960 543.620 2716.220 ;
        RECT 574.640 2715.960 574.900 2716.220 ;
        RECT 1010.720 2715.960 1010.980 2716.220 ;
        RECT 1055.340 2715.960 1055.600 2716.220 ;
        RECT 1145.500 2715.960 1145.760 2716.220 ;
        RECT 1172.640 2715.960 1172.900 2716.220 ;
        RECT 1352.960 2715.960 1353.220 2716.220 ;
        RECT 468.380 2715.620 468.640 2715.880 ;
        RECT 916.880 2715.620 917.140 2715.880 ;
        RECT 1013.940 2715.620 1014.200 2715.880 ;
        RECT 1072.820 2715.620 1073.080 2715.880 ;
        RECT 1082.940 2715.620 1083.200 2715.880 ;
        RECT 1186.900 2715.620 1187.160 2715.880 ;
        RECT 1193.340 2715.620 1193.600 2715.880 ;
        RECT 1383.780 2715.620 1384.040 2715.880 ;
        RECT 286.220 2715.280 286.480 2715.540 ;
        RECT 398.460 2715.280 398.720 2715.540 ;
        RECT 475.280 2715.280 475.540 2715.540 ;
        RECT 937.580 2715.280 937.840 2715.540 ;
        RECT 1020.840 2715.280 1021.100 2715.540 ;
        RECT 1069.140 2715.280 1069.400 2715.540 ;
        RECT 1166.200 2715.280 1166.460 2715.540 ;
        RECT 1186.440 2715.280 1186.700 2715.540 ;
        RECT 1373.660 2715.280 1373.920 2715.540 ;
        RECT 337.740 2714.940 338.000 2715.200 ;
        RECT 491.840 2714.940 492.100 2715.200 ;
        RECT 496.440 2714.940 496.700 2715.200 ;
        RECT 968.860 2714.940 969.120 2715.200 ;
        RECT 1082.940 2714.940 1083.200 2715.200 ;
        RECT 1089.380 2714.940 1089.640 2715.200 ;
        RECT 1197.020 2714.940 1197.280 2715.200 ;
        RECT 1200.240 2714.940 1200.500 2715.200 ;
        RECT 1394.360 2714.940 1394.620 2715.200 ;
        RECT 286.680 2714.600 286.940 2714.860 ;
        RECT 501.960 2714.600 502.220 2714.860 ;
        RECT 542.900 2714.600 543.160 2714.860 ;
        RECT 720.000 2714.600 720.260 2714.860 ;
        RECT 720.920 2714.600 721.180 2714.860 ;
        RECT 1020.840 2714.600 1021.100 2714.860 ;
        RECT 1130.780 2714.600 1131.040 2714.860 ;
        RECT 1280.280 2714.600 1280.540 2714.860 ;
        RECT 527.720 2714.260 527.980 2714.520 ;
        RECT 699.300 2714.260 699.560 2714.520 ;
        RECT 700.680 2714.260 700.940 2714.520 ;
        RECT 979.440 2714.260 979.700 2714.520 ;
        RECT 1131.240 2714.260 1131.500 2714.520 ;
        RECT 1269.700 2714.260 1269.960 2714.520 ;
        RECT 520.820 2713.920 521.080 2714.180 ;
        RECT 688.720 2713.920 688.980 2714.180 ;
        RECT 693.320 2713.920 693.580 2714.180 ;
        RECT 958.740 2713.920 959.000 2714.180 ;
        RECT 1117.440 2713.920 1117.700 2714.180 ;
        RECT 1249.000 2713.920 1249.260 2714.180 ;
        RECT 513.920 2713.580 514.180 2713.840 ;
        RECT 678.600 2713.580 678.860 2713.840 ;
        RECT 686.420 2713.580 686.680 2713.840 ;
        RECT 927.460 2713.580 927.720 2713.840 ;
        RECT 1123.420 2713.580 1123.680 2713.840 ;
        RECT 1259.580 2713.580 1259.840 2713.840 ;
        RECT 351.080 2713.240 351.340 2713.500 ;
        RECT 367.180 2713.240 367.440 2713.500 ;
        RECT 500.120 2713.240 500.380 2713.500 ;
        RECT 657.440 2713.240 657.700 2713.500 ;
        RECT 658.820 2713.240 659.080 2713.500 ;
        RECT 886.060 2713.240 886.320 2713.500 ;
        RECT 1110.540 2713.240 1110.800 2713.500 ;
        RECT 1238.880 2713.240 1239.140 2713.500 ;
        RECT 507.020 2712.900 507.280 2713.160 ;
        RECT 668.020 2712.900 668.280 2713.160 ;
        RECT 687.340 2712.900 687.600 2713.160 ;
        RECT 906.760 2712.900 907.020 2713.160 ;
        RECT 1102.720 2712.900 1102.980 2713.160 ;
        RECT 1228.300 2712.900 1228.560 2713.160 ;
        RECT 541.520 2712.560 541.780 2712.820 ;
        RECT 730.120 2712.560 730.380 2712.820 ;
        RECT 534.620 2712.220 534.880 2712.480 ;
        RECT 709.420 2712.220 709.680 2712.480 ;
        RECT 761.400 2712.560 761.660 2712.820 ;
        RECT 771.980 2712.560 772.240 2712.820 ;
        RECT 748.520 2712.220 748.780 2712.480 ;
        RECT 834.080 2712.560 834.340 2712.820 ;
        RECT 1089.840 2712.560 1090.100 2712.820 ;
        RECT 1207.600 2712.560 1207.860 2712.820 ;
        RECT 1096.740 2712.220 1097.000 2712.480 ;
        RECT 1217.720 2712.220 1217.980 2712.480 ;
        RECT 686.880 2711.880 687.140 2712.140 ;
        RECT 750.820 2711.880 751.080 2712.140 ;
        RECT 802.800 2711.880 803.060 2712.140 ;
        RECT 1408.620 2697.600 1408.880 2697.860 ;
        RECT 2321.720 2697.600 2321.980 2697.860 ;
        RECT 1408.620 2690.800 1408.880 2691.060 ;
        RECT 2273.420 2690.800 2273.680 2691.060 ;
        RECT 1408.620 2676.860 1408.880 2677.120 ;
        RECT 2267.440 2676.860 2267.700 2677.120 ;
        RECT 1408.620 2670.060 1408.880 2670.320 ;
        RECT 2259.620 2670.060 2259.880 2670.320 ;
        RECT 1408.620 2656.120 1408.880 2656.380 ;
        RECT 2252.720 2656.120 2252.980 2656.380 ;
        RECT 1408.620 2649.320 1408.880 2649.580 ;
        RECT 2245.820 2649.320 2246.080 2649.580 ;
        RECT 1408.620 2635.380 1408.880 2635.640 ;
        RECT 2238.920 2635.380 2239.180 2635.640 ;
        RECT 1408.620 2628.580 1408.880 2628.840 ;
        RECT 2232.020 2628.580 2232.280 2628.840 ;
        RECT 1408.620 2614.640 1408.880 2614.900 ;
        RECT 2218.220 2614.640 2218.480 2614.900 ;
        RECT 1408.620 2607.840 1408.880 2608.100 ;
        RECT 1797.780 2607.840 1798.040 2608.100 ;
        RECT 1408.620 2594.240 1408.880 2594.500 ;
        RECT 1797.320 2594.240 1797.580 2594.500 ;
        RECT 1408.620 2587.100 1408.880 2587.360 ;
        RECT 1790.880 2587.100 1791.140 2587.360 ;
        RECT 1408.620 2573.500 1408.880 2573.760 ;
        RECT 1783.520 2573.500 1783.780 2573.760 ;
        RECT 1408.620 2566.360 1408.880 2566.620 ;
        RECT 2366.800 2566.360 2367.060 2566.620 ;
        RECT 1408.620 2552.760 1408.880 2553.020 ;
        RECT 2359.900 2552.760 2360.160 2553.020 ;
        RECT 1408.620 2545.960 1408.880 2546.220 ;
        RECT 2353.000 2545.960 2353.260 2546.220 ;
        RECT 1408.620 2532.020 1408.880 2532.280 ;
        RECT 2346.100 2532.020 2346.360 2532.280 ;
        RECT 1408.620 2525.220 1408.880 2525.480 ;
        RECT 2339.660 2525.220 2339.920 2525.480 ;
        RECT 1408.620 2511.280 1408.880 2511.540 ;
        RECT 2339.200 2511.280 2339.460 2511.540 ;
        RECT 1408.620 2504.480 1408.880 2504.740 ;
        RECT 2332.300 2504.480 2332.560 2504.740 ;
        RECT 1408.620 2497.340 1408.880 2497.600 ;
        RECT 2325.400 2497.340 2325.660 2497.600 ;
        RECT 1408.620 2483.740 1408.880 2484.000 ;
        RECT 2318.500 2483.740 2318.760 2484.000 ;
        RECT 1408.620 2476.940 1408.880 2477.200 ;
        RECT 2311.600 2476.940 2311.860 2477.200 ;
        RECT 1408.620 2463.000 1408.880 2463.260 ;
        RECT 2305.160 2463.000 2305.420 2463.260 ;
        RECT 1408.620 2456.200 1408.880 2456.460 ;
        RECT 2304.700 2456.200 2304.960 2456.460 ;
        RECT 1408.620 2442.260 1408.880 2442.520 ;
        RECT 2297.800 2442.260 2298.060 2442.520 ;
        RECT 1408.620 2435.460 1408.880 2435.720 ;
        RECT 2290.900 2435.460 2291.160 2435.720 ;
        RECT 1408.620 2421.520 1408.880 2421.780 ;
        RECT 2284.000 2421.520 2284.260 2421.780 ;
        RECT 1408.620 2414.720 1408.880 2414.980 ;
        RECT 2277.100 2414.720 2277.360 2414.980 ;
        RECT 1408.620 2400.780 1408.880 2401.040 ;
        RECT 2266.980 2400.780 2267.240 2401.040 ;
        RECT 1408.620 2393.980 1408.880 2394.240 ;
        RECT 1790.420 2393.980 1790.680 2394.240 ;
        RECT 1408.620 2380.040 1408.880 2380.300 ;
        RECT 2263.300 2380.040 2263.560 2380.300 ;
        RECT 1408.620 2373.240 1408.880 2373.500 ;
        RECT 1794.560 2373.240 1794.820 2373.500 ;
        RECT 1408.620 2359.640 1408.880 2359.900 ;
        RECT 1787.660 2359.640 1787.920 2359.900 ;
        RECT 1408.620 2352.500 1408.880 2352.760 ;
        RECT 1780.300 2352.500 1780.560 2352.760 ;
        RECT 1408.620 2338.900 1408.880 2339.160 ;
        RECT 1773.400 2338.900 1773.660 2339.160 ;
        RECT 1408.620 2331.760 1408.880 2332.020 ;
        RECT 1766.500 2331.760 1766.760 2332.020 ;
        RECT 1408.620 2318.160 1408.880 2318.420 ;
        RECT 1760.060 2318.160 1760.320 2318.420 ;
        RECT 1408.620 2311.360 1408.880 2311.620 ;
        RECT 1760.980 2311.360 1761.240 2311.620 ;
        RECT 1408.620 2297.420 1408.880 2297.680 ;
        RECT 1752.700 2297.420 1752.960 2297.680 ;
        RECT 1408.620 2290.620 1408.880 2290.880 ;
        RECT 1745.800 2290.620 1746.060 2290.880 ;
        RECT 1408.620 2276.680 1408.880 2276.940 ;
        RECT 1738.900 2276.680 1739.160 2276.940 ;
        RECT 1408.620 2269.880 1408.880 2270.140 ;
        RECT 1732.000 2269.880 1732.260 2270.140 ;
        RECT 1408.620 2262.740 1408.880 2263.000 ;
        RECT 1725.100 2262.740 1725.360 2263.000 ;
        RECT 1408.620 2249.140 1408.880 2249.400 ;
        RECT 1718.660 2249.140 1718.920 2249.400 ;
        RECT 1408.620 2242.340 1408.880 2242.600 ;
        RECT 1718.200 2242.340 1718.460 2242.600 ;
        RECT 1408.620 2228.400 1408.880 2228.660 ;
        RECT 1711.300 2228.400 1711.560 2228.660 ;
        RECT 1408.620 2221.600 1408.880 2221.860 ;
        RECT 1704.400 2221.600 1704.660 2221.860 ;
        RECT 1408.620 2207.660 1408.880 2207.920 ;
        RECT 1697.500 2207.660 1697.760 2207.920 ;
        RECT 1408.620 2200.860 1408.880 2201.120 ;
        RECT 1690.600 2200.860 1690.860 2201.120 ;
        RECT 1408.620 2186.920 1408.880 2187.180 ;
        RECT 1684.160 2186.920 1684.420 2187.180 ;
        RECT 1408.620 2180.120 1408.880 2180.380 ;
        RECT 1683.700 2180.120 1683.960 2180.380 ;
        RECT 1408.620 2166.180 1408.880 2166.440 ;
        RECT 1676.800 2166.180 1677.060 2166.440 ;
        RECT 1408.620 2159.380 1408.880 2159.640 ;
        RECT 1669.900 2159.380 1670.160 2159.640 ;
        RECT 1408.620 2145.440 1408.880 2145.700 ;
        RECT 1663.000 2145.440 1663.260 2145.700 ;
        RECT 1408.620 2138.640 1408.880 2138.900 ;
        RECT 1656.100 2138.640 1656.360 2138.900 ;
        RECT 1408.620 2125.040 1408.880 2125.300 ;
        RECT 1649.660 2125.040 1649.920 2125.300 ;
        RECT 1408.620 2117.900 1408.880 2118.160 ;
        RECT 1649.200 2117.900 1649.460 2118.160 ;
        RECT 1408.620 2104.300 1408.880 2104.560 ;
        RECT 1642.300 2104.300 1642.560 2104.560 ;
        RECT 1408.620 2097.160 1408.880 2097.420 ;
        RECT 1635.400 2097.160 1635.660 2097.420 ;
        RECT 1408.620 2090.360 1408.880 2090.620 ;
        RECT 1628.500 2090.360 1628.760 2090.620 ;
        RECT 1408.620 2076.760 1408.880 2077.020 ;
        RECT 1621.600 2076.760 1621.860 2077.020 ;
        RECT 1408.620 2069.620 1408.880 2069.880 ;
        RECT 1614.700 2069.620 1614.960 2069.880 ;
        RECT 1426.560 2062.140 1426.820 2062.400 ;
        RECT 1580.200 2062.140 1580.460 2062.400 ;
        RECT 1408.160 2061.800 1408.420 2062.060 ;
        RECT 1624.820 2061.800 1625.080 2062.060 ;
        RECT 1407.700 2061.460 1407.960 2061.720 ;
        RECT 1631.720 2061.460 1631.980 2061.720 ;
        RECT 1638.620 2061.120 1638.880 2061.380 ;
        RECT 1415.520 2060.780 1415.780 2061.040 ;
        RECT 2192.920 2060.780 2193.180 2061.040 ;
        RECT 1415.060 2060.440 1415.320 2060.700 ;
        RECT 2192.460 2060.440 2192.720 2060.700 ;
        RECT 1415.980 2060.100 1416.240 2060.360 ;
        RECT 2193.380 2060.100 2193.640 2060.360 ;
        RECT 1416.440 2059.760 1416.700 2060.020 ;
        RECT 2228.800 2059.760 2229.060 2060.020 ;
        RECT 1427.020 2059.420 1427.280 2059.680 ;
        RECT 2266.520 2059.420 2266.780 2059.680 ;
        RECT 1408.620 2056.700 1408.880 2056.960 ;
        RECT 1410.000 2056.700 1410.260 2056.960 ;
        RECT 1410.000 2056.020 1410.260 2056.280 ;
        RECT 1607.800 2056.020 1608.060 2056.280 ;
        RECT 1426.100 2053.980 1426.360 2054.240 ;
        RECT 2190.620 2053.980 2190.880 2054.240 ;
        RECT 1425.640 2053.640 1425.900 2053.900 ;
        RECT 2191.080 2053.640 2191.340 2053.900 ;
        RECT 1425.180 2053.300 1425.440 2053.560 ;
        RECT 2191.540 2053.300 2191.800 2053.560 ;
        RECT 1416.900 2052.960 1417.160 2053.220 ;
        RECT 2193.840 2052.960 2194.100 2053.220 ;
        RECT 1410.000 2052.620 1410.260 2052.880 ;
        RECT 1414.600 2052.620 1414.860 2052.880 ;
        RECT 2192.000 2052.620 2192.260 2052.880 ;
        RECT 1407.700 2020.660 1407.960 2020.920 ;
        RECT 1410.000 2020.660 1410.260 2020.920 ;
        RECT 1407.700 1985.300 1407.960 1985.560 ;
        RECT 1417.360 1985.300 1417.620 1985.560 ;
        RECT 1409.540 1890.100 1409.800 1890.360 ;
        RECT 1427.020 1890.100 1427.280 1890.360 ;
        RECT 1414.140 1883.300 1414.400 1883.560 ;
        RECT 1473.480 1883.300 1473.740 1883.560 ;
        RECT 1414.140 1869.700 1414.400 1869.960 ;
        RECT 1459.220 1869.700 1459.480 1869.960 ;
        RECT 1414.140 1862.560 1414.400 1862.820 ;
        RECT 1452.320 1862.560 1452.580 1862.820 ;
        RECT 1411.840 1855.080 1412.100 1855.340 ;
        RECT 1438.520 1855.080 1438.780 1855.340 ;
        RECT 1411.380 1840.120 1411.640 1840.380 ;
        RECT 1431.620 1840.120 1431.880 1840.380 ;
        RECT 1408.620 1828.900 1408.880 1829.160 ;
        RECT 1424.720 1828.900 1424.980 1829.160 ;
        RECT 1414.140 1821.420 1414.400 1821.680 ;
        RECT 1473.020 1821.420 1473.280 1821.680 ;
        RECT 1409.540 1814.280 1409.800 1814.540 ;
        RECT 1426.560 1814.280 1426.820 1814.540 ;
        RECT 1409.540 1800.680 1409.800 1800.940 ;
        RECT 1426.100 1800.680 1426.360 1800.940 ;
        RECT 1408.620 1788.100 1408.880 1788.360 ;
        RECT 1425.640 1788.100 1425.900 1788.360 ;
        RECT 1410.460 1779.260 1410.720 1779.520 ;
        RECT 1425.180 1779.260 1425.440 1779.520 ;
        RECT 1407.700 1730.300 1407.960 1730.560 ;
        RECT 1416.440 1730.300 1416.700 1730.560 ;
        RECT 1414.140 1717.720 1414.400 1717.980 ;
        RECT 1514.420 1717.720 1514.680 1717.980 ;
        RECT 1407.700 1706.500 1407.960 1706.760 ;
        RECT 1416.900 1706.500 1417.160 1706.760 ;
        RECT 1408.620 1696.300 1408.880 1696.560 ;
        RECT 1421.040 1696.300 1421.300 1696.560 ;
        RECT 1407.700 1687.800 1407.960 1688.060 ;
        RECT 1420.580 1687.800 1420.840 1688.060 ;
        RECT 1408.160 1675.900 1408.420 1676.160 ;
        RECT 1420.120 1675.900 1420.380 1676.160 ;
        RECT 1407.700 1666.040 1407.960 1666.300 ;
        RECT 1419.660 1666.040 1419.920 1666.300 ;
        RECT 1407.700 1655.500 1407.960 1655.760 ;
        RECT 1419.200 1655.500 1419.460 1655.760 ;
        RECT 1407.700 1645.300 1407.960 1645.560 ;
        RECT 1418.740 1645.300 1419.000 1645.560 ;
        RECT 1407.700 1635.100 1407.960 1635.360 ;
        RECT 1418.280 1635.100 1418.540 1635.360 ;
        RECT 1407.700 1625.240 1407.960 1625.500 ;
        RECT 1417.820 1625.240 1418.080 1625.500 ;
      LAYER met2 ;
        RECT 1324.440 3266.730 1324.700 3267.050 ;
        RECT 1890.700 3266.730 1890.960 3267.050 ;
        RECT 1917.840 3266.730 1918.100 3267.050 ;
        RECT 2542.060 3266.730 2542.320 3267.050 ;
        RECT 1324.500 3264.670 1324.640 3266.730 ;
        RECT 1890.760 3264.670 1890.900 3266.730 ;
        RECT 1917.900 3264.670 1918.040 3266.730 ;
        RECT 1295.920 3264.525 1296.180 3264.670 ;
        RECT 1318.000 3264.525 1318.260 3264.670 ;
        RECT 646.390 3264.155 646.670 3264.525 ;
        RECT 668.470 3264.155 668.750 3264.525 ;
        RECT 1295.910 3264.155 1296.190 3264.525 ;
        RECT 1317.990 3264.155 1318.270 3264.525 ;
        RECT 1324.440 3264.350 1324.700 3264.670 ;
        RECT 1890.700 3264.525 1890.960 3264.670 ;
        RECT 1917.840 3264.525 1918.100 3264.670 ;
        RECT 2542.120 3264.525 2542.260 3266.730 ;
        RECT 1890.690 3264.155 1890.970 3264.525 ;
        RECT 1917.830 3264.155 1918.110 3264.525 ;
        RECT 2542.050 3264.155 2542.330 3264.525 ;
        RECT 2566.890 3264.155 2567.170 3264.525 ;
        RECT 646.460 3263.990 646.600 3264.155 ;
        RECT 668.540 3263.990 668.680 3264.155 ;
        RECT 1917.900 3264.025 1918.040 3264.155 ;
        RECT 2542.060 3264.010 2542.320 3264.155 ;
        RECT 2566.900 3264.010 2567.160 3264.155 ;
        RECT 646.400 3263.670 646.660 3263.990 ;
        RECT 668.480 3263.670 668.740 3263.990 ;
        RECT 697.000 3263.670 697.260 3263.990 ;
        RECT 2542.120 3263.855 2542.260 3264.010 ;
        RECT 2594.500 3263.670 2594.760 3263.990 ;
        RECT 697.060 3252.850 697.200 3263.670 ;
        RECT 696.600 3252.710 697.200 3252.850 ;
        RECT 688.260 3252.110 688.520 3252.430 ;
        RECT 289.430 3230.155 289.710 3230.525 ;
        RECT 288.970 3224.715 289.250 3225.085 ;
        RECT 288.510 3215.875 288.790 3216.245 ;
        RECT 288.050 3209.755 288.330 3210.125 ;
        RECT 287.590 3201.595 287.870 3201.965 ;
        RECT 287.130 3196.155 287.410 3196.525 ;
        RECT 286.670 3187.995 286.950 3188.365 ;
        RECT 286.210 2898.315 286.490 2898.685 ;
        RECT 286.280 2715.570 286.420 2898.315 ;
        RECT 286.220 2715.250 286.480 2715.570 ;
        RECT 286.740 2714.890 286.880 3187.995 ;
        RECT 287.200 2717.610 287.340 3196.155 ;
        RECT 287.140 2717.290 287.400 2717.610 ;
        RECT 287.660 2717.270 287.800 3201.595 ;
        RECT 287.600 2716.950 287.860 2717.270 ;
        RECT 288.120 2716.930 288.260 3209.755 ;
        RECT 288.060 2716.610 288.320 2716.930 ;
        RECT 288.580 2716.250 288.720 3215.875 ;
        RECT 289.040 2719.310 289.180 3224.715 ;
        RECT 289.500 2719.650 289.640 3230.155 ;
      LAYER met2 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met2 ;
        RECT 688.320 3248.600 688.460 3252.110 ;
        RECT 696.600 3248.770 696.740 3252.710 ;
        RECT 1332.260 3252.450 1332.520 3252.770 ;
        RECT 1332.320 3251.410 1332.460 3252.450 ;
        RECT 1414.140 3252.110 1414.400 3252.430 ;
        RECT 2582.080 3252.110 2582.340 3252.430 ;
        RECT 696.600 3248.630 697.200 3248.770 ;
        RECT 688.250 3248.230 688.530 3248.600 ;
        RECT 697.060 2948.325 697.200 3248.630 ;
        RECT 941.710 3230.155 941.990 3230.525 ;
        RECT 696.990 2947.955 697.270 2948.325 ;
        RECT 696.990 2901.715 697.270 2902.085 ;
        RECT 697.060 2898.150 697.200 2901.715 ;
        RECT 697.000 2897.830 697.260 2898.150 ;
        RECT 938.500 2897.830 938.760 2898.150 ;
        RECT 938.560 2895.285 938.700 2897.830 ;
        RECT 938.490 2894.915 938.770 2895.285 ;
        RECT 330.840 2794.130 331.100 2794.450 ;
        RECT 337.730 2794.275 338.010 2794.645 ;
        RECT 344.630 2794.275 344.910 2794.645 ;
        RECT 351.070 2794.275 351.350 2794.645 ;
        RECT 358.430 2794.275 358.710 2794.645 ;
        RECT 362.570 2794.275 362.850 2794.645 ;
        RECT 365.330 2794.275 365.610 2794.645 ;
        RECT 368.550 2794.275 368.830 2794.645 ;
        RECT 371.310 2794.275 371.590 2794.645 ;
        RECT 374.990 2794.275 375.270 2794.645 ;
        RECT 379.130 2794.275 379.410 2794.645 ;
        RECT 384.190 2794.275 384.470 2794.645 ;
        RECT 386.950 2794.275 387.230 2794.645 ;
        RECT 392.930 2794.275 393.210 2794.645 ;
        RECT 396.610 2794.275 396.890 2794.645 ;
        RECT 399.830 2794.275 400.110 2794.645 ;
        RECT 403.970 2794.275 404.250 2794.645 ;
        RECT 406.270 2794.275 406.550 2794.645 ;
        RECT 409.950 2794.275 410.230 2794.645 ;
        RECT 413.630 2794.275 413.910 2794.645 ;
        RECT 419.150 2794.275 419.430 2794.645 ;
        RECT 420.990 2794.275 421.270 2794.645 ;
        RECT 427.430 2794.275 427.710 2794.645 ;
        RECT 433.870 2794.275 434.150 2794.645 ;
        RECT 439.390 2794.275 439.670 2794.645 ;
        RECT 441.230 2794.275 441.510 2794.645 ;
        RECT 444.450 2794.275 444.730 2794.645 ;
        RECT 446.750 2794.275 447.030 2794.645 ;
        RECT 449.050 2794.275 449.330 2794.645 ;
        RECT 455.030 2794.275 455.310 2794.645 ;
        RECT 461.470 2794.275 461.750 2794.645 ;
        RECT 462.390 2794.275 462.670 2794.645 ;
        RECT 468.370 2794.275 468.650 2794.645 ;
        RECT 474.350 2794.275 474.630 2794.645 ;
        RECT 475.270 2794.275 475.550 2794.645 ;
        RECT 478.490 2794.275 478.770 2794.645 ;
        RECT 482.630 2794.275 482.910 2794.645 ;
        RECT 485.390 2794.275 485.670 2794.645 ;
        RECT 488.150 2794.275 488.430 2794.645 ;
        RECT 492.750 2794.275 493.030 2794.645 ;
        RECT 496.430 2794.275 496.710 2794.645 ;
        RECT 502.870 2794.275 503.150 2794.645 ;
        RECT 510.230 2794.275 510.510 2794.645 ;
        RECT 524.030 2794.275 524.310 2794.645 ;
        RECT 537.370 2794.275 537.650 2794.645 ;
        RECT 542.430 2794.275 542.710 2794.645 ;
        RECT 310.130 2791.555 310.410 2791.925 ;
        RECT 289.440 2719.330 289.700 2719.650 ;
        RECT 288.980 2718.990 289.240 2719.310 ;
        RECT 310.200 2717.950 310.340 2791.555 ;
        RECT 317.030 2790.875 317.310 2791.245 ;
        RECT 305.080 2717.630 305.340 2717.950 ;
        RECT 310.140 2717.630 310.400 2717.950 ;
        RECT 288.520 2715.930 288.780 2716.250 ;
        RECT 286.680 2714.570 286.940 2714.890 ;
        RECT 305.140 2700.000 305.280 2717.630 ;
        RECT 317.100 2700.010 317.240 2790.875 ;
        RECT 330.900 2717.950 331.040 2794.130 ;
        RECT 337.280 2793.790 337.540 2794.110 ;
        RECT 325.780 2717.630 326.040 2717.950 ;
        RECT 330.840 2717.630 331.100 2717.950 ;
        RECT 315.330 2700.000 317.240 2700.010 ;
        RECT 325.840 2700.000 325.980 2717.630 ;
        RECT 337.340 2700.010 337.480 2793.790 ;
        RECT 337.800 2715.230 337.940 2794.275 ;
        RECT 337.740 2714.910 338.000 2715.230 ;
        RECT 344.700 2712.250 344.840 2794.275 ;
        RECT 351.140 2713.530 351.280 2794.275 ;
        RECT 351.530 2793.595 351.810 2793.965 ;
        RECT 351.600 2717.950 351.740 2793.595 ;
        RECT 358.500 2718.630 358.640 2794.275 ;
        RECT 362.640 2791.050 362.780 2794.275 ;
        RECT 362.580 2790.730 362.840 2791.050 ;
        RECT 365.400 2719.990 365.540 2794.275 ;
        RECT 368.620 2792.070 368.760 2794.275 ;
        RECT 368.560 2791.750 368.820 2792.070 ;
        RECT 371.380 2791.390 371.520 2794.275 ;
        RECT 371.320 2791.070 371.580 2791.390 ;
        RECT 375.060 2789.690 375.200 2794.275 ;
        RECT 375.000 2789.370 375.260 2789.690 ;
        RECT 365.340 2719.670 365.600 2719.990 ;
        RECT 379.200 2718.630 379.340 2794.275 ;
        RECT 379.590 2793.595 379.870 2793.965 ;
        RECT 379.660 2792.750 379.800 2793.595 ;
        RECT 379.600 2792.430 379.860 2792.750 ;
        RECT 384.260 2790.710 384.400 2794.275 ;
        RECT 387.020 2793.090 387.160 2794.275 ;
        RECT 392.470 2793.595 392.750 2793.965 ;
        RECT 392.540 2793.430 392.680 2793.595 ;
        RECT 392.480 2793.110 392.740 2793.430 ;
        RECT 386.960 2792.770 387.220 2793.090 ;
        RECT 384.200 2790.390 384.460 2790.710 ;
        RECT 358.440 2718.310 358.700 2718.630 ;
        RECT 377.300 2718.310 377.560 2718.630 ;
        RECT 379.140 2718.310 379.400 2718.630 ;
        RECT 351.540 2717.630 351.800 2717.950 ;
        RECT 356.600 2717.630 356.860 2717.950 ;
        RECT 351.080 2713.210 351.340 2713.530 ;
        RECT 344.700 2712.110 345.300 2712.250 ;
        RECT 336.030 2700.000 337.480 2700.010 ;
        RECT 305.080 2696.000 305.360 2700.000 ;
        RECT 315.200 2699.870 317.240 2700.000 ;
        RECT 315.200 2696.000 315.480 2699.870 ;
        RECT 325.780 2696.000 326.060 2700.000 ;
        RECT 335.900 2699.870 337.480 2700.000 ;
        RECT 345.160 2700.010 345.300 2712.110 ;
        RECT 345.160 2700.000 346.610 2700.010 ;
        RECT 356.660 2700.000 356.800 2717.630 ;
        RECT 367.180 2713.210 367.440 2713.530 ;
        RECT 367.240 2700.000 367.380 2713.210 ;
        RECT 377.360 2700.000 377.500 2718.310 ;
        RECT 393.000 2718.290 393.140 2794.275 ;
        RECT 396.680 2790.030 396.820 2794.275 ;
        RECT 397.530 2793.595 397.810 2793.965 ;
        RECT 397.540 2793.450 397.800 2793.595 ;
        RECT 396.620 2789.710 396.880 2790.030 ;
        RECT 392.940 2717.970 393.200 2718.290 ;
        RECT 399.900 2717.950 400.040 2794.275 ;
        RECT 404.040 2792.410 404.180 2794.275 ;
        RECT 403.980 2792.090 404.240 2792.410 ;
        RECT 406.340 2790.370 406.480 2794.275 ;
        RECT 410.020 2791.730 410.160 2794.275 ;
        RECT 407.200 2791.410 407.460 2791.730 ;
        RECT 409.960 2791.410 410.220 2791.730 ;
        RECT 407.260 2791.050 407.400 2791.410 ;
        RECT 407.200 2790.730 407.460 2791.050 ;
        RECT 406.280 2790.050 406.540 2790.370 ;
        RECT 408.580 2721.710 408.840 2722.030 ;
        RECT 399.840 2717.630 400.100 2717.950 ;
        RECT 398.460 2715.250 398.720 2715.570 ;
        RECT 387.870 2714.715 388.150 2715.085 ;
        RECT 387.940 2700.000 388.080 2714.715 ;
        RECT 398.520 2700.000 398.660 2715.250 ;
        RECT 408.640 2700.000 408.780 2721.710 ;
        RECT 413.700 2720.330 413.840 2794.275 ;
        RECT 414.550 2793.595 414.830 2793.965 ;
        RECT 414.620 2792.070 414.760 2793.595 ;
        RECT 414.560 2791.750 414.820 2792.070 ;
        RECT 419.220 2791.050 419.360 2794.275 ;
        RECT 419.160 2790.730 419.420 2791.050 ;
        RECT 421.060 2789.690 421.200 2794.275 ;
        RECT 426.970 2793.595 427.250 2793.965 ;
        RECT 427.040 2792.750 427.180 2793.595 ;
        RECT 426.980 2792.430 427.240 2792.750 ;
        RECT 421.000 2789.370 421.260 2789.690 ;
        RECT 421.060 2787.990 421.200 2789.370 ;
        RECT 421.000 2787.670 421.260 2787.990 ;
        RECT 419.160 2722.050 419.420 2722.370 ;
        RECT 413.640 2720.010 413.900 2720.330 ;
        RECT 419.220 2700.000 419.360 2722.050 ;
        RECT 427.500 2720.670 427.640 2794.275 ;
        RECT 433.410 2792.915 433.690 2793.285 ;
        RECT 433.420 2792.770 433.680 2792.915 ;
        RECT 433.480 2792.410 433.620 2792.770 ;
        RECT 433.420 2792.090 433.680 2792.410 ;
        RECT 429.280 2722.390 429.540 2722.710 ;
        RECT 427.440 2720.350 427.700 2720.670 ;
        RECT 429.340 2700.000 429.480 2722.390 ;
        RECT 433.940 2721.690 434.080 2794.275 ;
        RECT 434.330 2793.595 434.610 2793.965 ;
        RECT 433.880 2721.370 434.140 2721.690 ;
        RECT 434.400 2721.010 434.540 2793.595 ;
        RECT 439.460 2793.430 439.600 2794.275 ;
        RECT 439.400 2793.110 439.660 2793.430 ;
        RECT 439.860 2723.070 440.120 2723.390 ;
        RECT 434.340 2720.690 434.600 2721.010 ;
        RECT 439.920 2700.000 440.060 2723.070 ;
        RECT 441.300 2721.350 441.440 2794.275 ;
        RECT 444.520 2793.770 444.660 2794.275 ;
        RECT 444.460 2793.450 444.720 2793.770 ;
        RECT 446.820 2789.010 446.960 2794.275 ;
        RECT 449.120 2792.410 449.260 2794.275 ;
        RECT 449.060 2792.090 449.320 2792.410 ;
        RECT 449.120 2789.690 449.260 2792.090 ;
        RECT 449.060 2789.370 449.320 2789.690 ;
        RECT 446.760 2788.690 447.020 2789.010 ;
        RECT 449.980 2723.750 450.240 2724.070 ;
        RECT 441.240 2721.030 441.500 2721.350 ;
        RECT 450.040 2700.000 450.180 2723.750 ;
        RECT 455.100 2716.590 455.240 2794.275 ;
        RECT 455.490 2793.595 455.770 2793.965 ;
        RECT 455.560 2791.730 455.700 2793.595 ;
        RECT 461.540 2791.730 461.680 2794.275 ;
        RECT 455.500 2791.410 455.760 2791.730 ;
        RECT 461.480 2791.410 461.740 2791.730 ;
        RECT 455.560 2788.670 455.700 2791.410 ;
        RECT 455.500 2788.350 455.760 2788.670 ;
        RECT 462.460 2788.330 462.600 2794.275 ;
        RECT 467.910 2792.915 468.190 2793.285 ;
        RECT 462.400 2788.010 462.660 2788.330 ;
        RECT 467.980 2787.990 468.120 2792.915 ;
        RECT 467.920 2787.670 468.180 2787.990 ;
        RECT 460.560 2724.090 460.820 2724.410 ;
        RECT 455.040 2716.270 455.300 2716.590 ;
        RECT 460.620 2700.000 460.760 2724.090 ;
        RECT 468.440 2715.910 468.580 2794.275 ;
        RECT 468.830 2793.595 469.110 2793.965 ;
        RECT 468.900 2789.690 469.040 2793.595 ;
        RECT 474.420 2793.090 474.560 2794.275 ;
        RECT 474.360 2792.770 474.620 2793.090 ;
        RECT 468.840 2789.370 469.100 2789.690 ;
        RECT 470.680 2724.770 470.940 2725.090 ;
        RECT 468.380 2715.590 468.640 2715.910 ;
        RECT 470.740 2700.000 470.880 2724.770 ;
        RECT 475.340 2715.570 475.480 2794.275 ;
        RECT 478.560 2792.750 478.700 2794.275 ;
        RECT 478.500 2792.430 478.760 2792.750 ;
        RECT 482.700 2725.430 482.840 2794.275 ;
        RECT 485.460 2793.430 485.600 2794.275 ;
        RECT 485.400 2793.110 485.660 2793.430 ;
        RECT 485.460 2789.010 485.600 2793.110 ;
        RECT 488.220 2792.070 488.360 2794.275 ;
        RECT 492.820 2793.770 492.960 2794.275 ;
        RECT 492.760 2793.450 493.020 2793.770 ;
        RECT 488.160 2791.750 488.420 2792.070 ;
        RECT 485.400 2788.690 485.660 2789.010 ;
        RECT 482.640 2725.110 482.900 2725.430 ;
        RECT 481.250 2716.075 481.530 2716.445 ;
        RECT 475.280 2715.250 475.540 2715.570 ;
        RECT 481.320 2700.000 481.460 2716.075 ;
        RECT 496.500 2715.230 496.640 2794.275 ;
        RECT 496.890 2792.235 497.170 2792.605 ;
        RECT 502.940 2792.410 503.080 2794.275 ;
        RECT 510.300 2793.430 510.440 2794.275 ;
        RECT 510.240 2793.110 510.500 2793.430 ;
        RECT 524.100 2793.090 524.240 2794.275 ;
        RECT 524.490 2793.595 524.770 2793.965 ;
        RECT 524.500 2793.450 524.760 2793.595 ;
        RECT 513.920 2792.770 514.180 2793.090 ;
        RECT 524.040 2792.770 524.300 2793.090 ;
        RECT 496.900 2792.090 497.160 2792.235 ;
        RECT 500.580 2792.090 500.840 2792.410 ;
        RECT 502.880 2792.090 503.140 2792.410 ;
        RECT 500.110 2788.835 500.390 2789.205 ;
        RECT 500.180 2788.670 500.320 2788.835 ;
        RECT 500.640 2788.670 500.780 2792.090 ;
        RECT 500.120 2788.350 500.380 2788.670 ;
        RECT 500.580 2788.350 500.840 2788.670 ;
        RECT 491.840 2714.910 492.100 2715.230 ;
        RECT 496.440 2714.910 496.700 2715.230 ;
        RECT 491.900 2700.000 492.040 2714.910 ;
        RECT 500.180 2713.530 500.320 2788.350 ;
        RECT 504.250 2788.155 504.530 2788.525 ;
        RECT 507.010 2788.155 507.290 2788.525 ;
        RECT 504.260 2788.010 504.520 2788.155 ;
        RECT 501.960 2714.570 502.220 2714.890 ;
        RECT 500.120 2713.210 500.380 2713.530 ;
        RECT 502.020 2700.000 502.160 2714.570 ;
        RECT 507.080 2713.190 507.220 2788.155 ;
        RECT 513.980 2787.845 514.120 2792.770 ;
        RECT 520.820 2792.430 521.080 2792.750 ;
        RECT 520.880 2787.845 521.020 2792.430 ;
        RECT 531.400 2788.690 531.660 2789.010 ;
        RECT 531.460 2788.525 531.600 2788.690 ;
        RECT 531.390 2788.155 531.670 2788.525 ;
        RECT 534.610 2788.155 534.890 2788.525 ;
        RECT 510.230 2787.475 510.510 2787.845 ;
        RECT 513.910 2787.475 514.190 2787.845 ;
        RECT 517.130 2787.475 517.410 2787.845 ;
        RECT 520.810 2787.475 521.090 2787.845 ;
        RECT 527.710 2787.475 527.990 2787.845 ;
        RECT 530.930 2787.475 531.210 2787.845 ;
        RECT 510.300 2724.750 510.440 2787.475 ;
        RECT 510.240 2724.430 510.500 2724.750 ;
        RECT 512.540 2717.290 512.800 2717.610 ;
        RECT 507.020 2712.870 507.280 2713.190 ;
        RECT 512.600 2700.000 512.740 2717.290 ;
        RECT 513.980 2713.870 514.120 2787.475 ;
        RECT 517.200 2715.765 517.340 2787.475 ;
        RECT 517.130 2715.395 517.410 2715.765 ;
        RECT 520.880 2714.210 521.020 2787.475 ;
        RECT 522.660 2716.950 522.920 2717.270 ;
        RECT 520.820 2713.890 521.080 2714.210 ;
        RECT 513.920 2713.550 514.180 2713.870 ;
        RECT 522.720 2700.000 522.860 2716.950 ;
        RECT 527.780 2714.550 527.920 2787.475 ;
        RECT 531.000 2723.730 531.140 2787.475 ;
        RECT 530.940 2723.410 531.200 2723.730 ;
        RECT 533.240 2716.610 533.500 2716.930 ;
        RECT 527.720 2714.230 527.980 2714.550 ;
        RECT 533.300 2700.000 533.440 2716.610 ;
        RECT 534.680 2712.510 534.820 2788.155 ;
        RECT 537.440 2787.990 537.580 2794.275 ;
        RECT 542.500 2792.750 542.640 2794.275 ;
        RECT 627.540 2793.450 627.800 2793.770 ;
        RECT 541.510 2792.235 541.790 2792.605 ;
        RECT 542.440 2792.430 542.700 2792.750 ;
        RECT 538.300 2789.030 538.560 2789.350 ;
        RECT 537.380 2787.670 537.640 2787.990 ;
        RECT 538.360 2787.845 538.500 2789.030 ;
        RECT 541.580 2788.670 541.720 2792.235 ;
        RECT 606.840 2788.690 607.100 2789.010 ;
        RECT 541.520 2788.350 541.780 2788.670 ;
        RECT 586.140 2788.350 586.400 2788.670 ;
        RECT 538.290 2787.475 538.570 2787.845 ;
        RECT 541.580 2712.850 541.720 2788.350 ;
        RECT 542.430 2787.475 542.710 2787.845 ;
        RECT 551.630 2787.475 551.910 2787.845 ;
        RECT 542.500 2739.450 542.640 2787.475 ;
        RECT 542.500 2739.310 543.100 2739.450 ;
        RECT 542.960 2714.890 543.100 2739.310 ;
        RECT 551.700 2723.050 551.840 2787.475 ;
        RECT 551.640 2722.730 551.900 2723.050 ;
        RECT 564.060 2719.330 564.320 2719.650 ;
        RECT 553.940 2718.990 554.200 2719.310 ;
        RECT 543.360 2715.930 543.620 2716.250 ;
        RECT 542.900 2714.570 543.160 2714.890 ;
        RECT 541.520 2712.530 541.780 2712.850 ;
        RECT 534.620 2712.190 534.880 2712.510 ;
        RECT 543.420 2700.000 543.560 2715.930 ;
        RECT 554.000 2700.000 554.140 2718.990 ;
        RECT 564.120 2700.000 564.260 2719.330 ;
        RECT 574.640 2715.930 574.900 2716.250 ;
        RECT 574.700 2700.000 574.840 2715.930 ;
        RECT 586.200 2700.010 586.340 2788.350 ;
        RECT 595.340 2716.610 595.600 2716.930 ;
        RECT 585.350 2700.000 586.340 2700.010 ;
        RECT 595.400 2700.000 595.540 2716.610 ;
        RECT 606.900 2700.010 607.040 2788.690 ;
        RECT 616.040 2716.950 616.300 2717.270 ;
        RECT 606.050 2700.000 607.040 2700.010 ;
        RECT 616.100 2700.000 616.240 2716.950 ;
        RECT 627.600 2700.010 627.740 2793.450 ;
        RECT 700.220 2793.110 700.480 2793.430 ;
        RECT 693.320 2791.750 693.580 2792.070 ;
        RECT 687.340 2791.410 687.600 2791.730 ;
        RECT 686.880 2791.070 687.140 2791.390 ;
        RECT 686.420 2789.370 686.680 2789.690 ;
        RECT 648.700 2788.010 648.960 2788.330 ;
        RECT 648.760 2787.730 648.900 2788.010 ;
        RECT 648.300 2787.590 648.900 2787.730 ;
        RECT 636.740 2717.290 637.000 2717.610 ;
        RECT 626.750 2700.000 627.740 2700.010 ;
        RECT 636.800 2700.000 636.940 2717.290 ;
        RECT 648.300 2700.010 648.440 2787.590 ;
        RECT 658.820 2787.330 659.080 2787.650 ;
        RECT 658.880 2713.530 659.020 2787.330 ;
        RECT 686.480 2713.870 686.620 2789.370 ;
        RECT 678.600 2713.550 678.860 2713.870 ;
        RECT 686.420 2713.550 686.680 2713.870 ;
        RECT 657.440 2713.210 657.700 2713.530 ;
        RECT 658.820 2713.210 659.080 2713.530 ;
        RECT 647.450 2700.000 648.440 2700.010 ;
        RECT 657.500 2700.000 657.640 2713.210 ;
        RECT 668.020 2712.870 668.280 2713.190 ;
        RECT 668.080 2700.000 668.220 2712.870 ;
        RECT 678.660 2700.000 678.800 2713.550 ;
        RECT 686.940 2712.170 687.080 2791.070 ;
        RECT 687.400 2713.190 687.540 2791.410 ;
        RECT 693.380 2714.210 693.520 2791.750 ;
        RECT 700.280 2718.485 700.420 2793.110 ;
        RECT 720.920 2792.770 721.180 2793.090 ;
        RECT 700.680 2792.090 700.940 2792.410 ;
        RECT 700.210 2718.115 700.490 2718.485 ;
        RECT 700.740 2714.550 700.880 2792.090 ;
        RECT 707.120 2787.670 707.380 2787.990 ;
        RECT 707.180 2717.125 707.320 2787.670 ;
        RECT 707.110 2716.755 707.390 2717.125 ;
        RECT 720.980 2714.890 721.120 2792.770 ;
        RECT 741.620 2792.430 741.880 2792.750 ;
        RECT 727.820 2790.390 728.080 2790.710 ;
        RECT 727.880 2718.630 728.020 2790.390 ;
        RECT 740.700 2719.670 740.960 2719.990 ;
        RECT 727.820 2718.310 728.080 2718.630 ;
        RECT 720.000 2714.570 720.260 2714.890 ;
        RECT 720.920 2714.570 721.180 2714.890 ;
        RECT 699.300 2714.230 699.560 2714.550 ;
        RECT 700.680 2714.230 700.940 2714.550 ;
        RECT 688.720 2713.890 688.980 2714.210 ;
        RECT 693.320 2713.890 693.580 2714.210 ;
        RECT 687.340 2712.870 687.600 2713.190 ;
        RECT 686.880 2711.850 687.140 2712.170 ;
        RECT 688.780 2700.000 688.920 2713.890 ;
        RECT 699.360 2700.000 699.500 2714.230 ;
        RECT 709.420 2712.190 709.680 2712.510 ;
        RECT 709.480 2700.000 709.620 2712.190 ;
        RECT 720.060 2700.000 720.200 2714.570 ;
        RECT 730.120 2712.530 730.380 2712.850 ;
        RECT 730.180 2700.000 730.320 2712.530 ;
        RECT 740.760 2700.000 740.900 2719.670 ;
        RECT 741.680 2717.805 741.820 2792.430 ;
        RECT 748.520 2790.730 748.780 2791.050 ;
        RECT 741.610 2717.435 741.890 2717.805 ;
        RECT 748.580 2712.510 748.720 2790.730 ;
        RECT 762.780 2790.050 763.040 2790.370 ;
        RECT 762.320 2789.710 762.580 2790.030 ;
        RECT 762.380 2717.950 762.520 2789.710 ;
        RECT 762.840 2718.630 762.980 2790.050 ;
        RECT 865.360 2721.370 865.620 2721.690 ;
        RECT 854.780 2720.690 855.040 2721.010 ;
        RECT 844.200 2720.350 844.460 2720.670 ;
        RECT 823.500 2720.010 823.760 2720.330 ;
        RECT 762.780 2718.310 763.040 2718.630 ;
        RECT 813.380 2718.310 813.640 2718.630 ;
        RECT 782.100 2717.970 782.360 2718.290 ;
        RECT 762.320 2717.630 762.580 2717.950 ;
        RECT 761.400 2712.530 761.660 2712.850 ;
        RECT 771.980 2712.530 772.240 2712.850 ;
        RECT 748.520 2712.190 748.780 2712.510 ;
        RECT 750.820 2711.850 751.080 2712.170 ;
        RECT 750.880 2700.000 751.020 2711.850 ;
        RECT 761.460 2700.000 761.600 2712.530 ;
        RECT 772.040 2700.000 772.180 2712.530 ;
        RECT 782.160 2700.000 782.300 2717.970 ;
        RECT 792.680 2717.630 792.940 2717.950 ;
        RECT 792.740 2700.000 792.880 2717.630 ;
        RECT 802.800 2711.850 803.060 2712.170 ;
        RECT 802.860 2700.000 803.000 2711.850 ;
        RECT 813.440 2700.000 813.580 2718.310 ;
        RECT 823.560 2700.000 823.700 2720.010 ;
        RECT 834.080 2712.530 834.340 2712.850 ;
        RECT 834.140 2700.000 834.280 2712.530 ;
        RECT 844.260 2700.000 844.400 2720.350 ;
        RECT 854.840 2700.000 854.980 2720.690 ;
        RECT 865.420 2700.000 865.560 2721.370 ;
        RECT 875.480 2721.030 875.740 2721.350 ;
        RECT 875.540 2700.000 875.680 2721.030 ;
        RECT 896.180 2716.270 896.440 2716.590 ;
        RECT 941.780 2716.445 941.920 3230.155 ;
        RECT 942.170 3224.715 942.450 3225.085 ;
        RECT 942.240 2725.090 942.380 3224.715 ;
        RECT 942.630 3215.875 942.910 3216.245 ;
        RECT 942.180 2724.770 942.440 2725.090 ;
        RECT 942.700 2724.410 942.840 3215.875 ;
        RECT 943.090 3209.755 943.370 3210.125 ;
        RECT 942.640 2724.090 942.900 2724.410 ;
        RECT 943.160 2724.070 943.300 3209.755 ;
        RECT 943.550 3201.595 943.830 3201.965 ;
        RECT 943.100 2723.750 943.360 2724.070 ;
        RECT 943.620 2723.390 943.760 3201.595 ;
        RECT 944.010 3196.155 944.290 3196.525 ;
        RECT 943.560 2723.070 943.820 2723.390 ;
        RECT 944.080 2722.710 944.220 3196.155 ;
        RECT 944.470 3187.995 944.750 3188.365 ;
        RECT 944.020 2722.390 944.280 2722.710 ;
        RECT 944.540 2722.370 944.680 3187.995 ;
        RECT 944.930 2898.315 945.210 2898.685 ;
        RECT 944.480 2722.050 944.740 2722.370 ;
        RECT 886.060 2713.210 886.320 2713.530 ;
        RECT 886.120 2700.000 886.260 2713.210 ;
        RECT 896.240 2700.000 896.380 2716.270 ;
        RECT 941.710 2716.075 941.990 2716.445 ;
        RECT 916.880 2715.590 917.140 2715.910 ;
        RECT 906.760 2712.870 907.020 2713.190 ;
        RECT 906.820 2700.000 906.960 2712.870 ;
        RECT 916.940 2700.000 917.080 2715.590 ;
        RECT 937.580 2715.250 937.840 2715.570 ;
        RECT 927.460 2713.550 927.720 2713.870 ;
        RECT 927.520 2700.000 927.660 2713.550 ;
        RECT 937.640 2700.000 937.780 2715.250 ;
        RECT 945.000 2715.085 945.140 2898.315 ;
      LAYER met2 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met2 ;
        RECT 1332.260 3251.090 1332.520 3251.410 ;
        RECT 1332.320 3249.565 1332.460 3251.090 ;
        RECT 1414.200 3251.070 1414.340 3252.110 ;
        RECT 1411.380 3250.750 1411.640 3251.070 ;
        RECT 1414.140 3250.750 1414.400 3251.070 ;
        RECT 1332.250 3249.195 1332.530 3249.565 ;
        RECT 1411.440 3243.445 1411.580 3250.750 ;
        RECT 1411.370 3243.075 1411.650 3243.445 ;
        RECT 1536.950 3230.155 1537.230 3230.525 ;
        RECT 1537.020 3229.650 1537.160 3230.155 ;
        RECT 1473.480 3229.330 1473.740 3229.650 ;
        RECT 1536.960 3229.330 1537.220 3229.650 ;
        RECT 1459.220 3222.190 1459.480 3222.510 ;
        RECT 1452.320 3215.390 1452.580 3215.710 ;
        RECT 1438.520 3208.590 1438.780 3208.910 ;
        RECT 1431.620 3201.450 1431.880 3201.770 ;
        RECT 1424.720 3194.650 1424.980 3194.970 ;
        RECT 1410.910 2935.715 1411.190 2936.085 ;
        RECT 1410.980 2932.685 1411.120 2935.715 ;
        RECT 1410.910 2932.315 1411.190 2932.685 ;
        RECT 1410.980 2894.750 1411.120 2932.315 ;
        RECT 1410.920 2894.430 1411.180 2894.750 ;
        RECT 1146.870 2799.715 1147.150 2800.085 ;
        RECT 1129.850 2799.035 1130.130 2799.405 ;
        RECT 979.890 2794.275 980.170 2794.645 ;
        RECT 1001.050 2794.275 1001.330 2794.645 ;
        RECT 1007.490 2794.275 1007.770 2794.645 ;
        RECT 1013.930 2794.275 1014.210 2794.645 ;
        RECT 1018.990 2794.275 1019.270 2794.645 ;
        RECT 1020.830 2794.275 1021.110 2794.645 ;
        RECT 1027.730 2794.275 1028.010 2794.645 ;
        RECT 1031.870 2794.275 1032.150 2794.645 ;
        RECT 1042.450 2794.275 1042.730 2794.645 ;
        RECT 1059.470 2794.275 1059.750 2794.645 ;
        RECT 1065.450 2794.275 1065.730 2794.645 ;
        RECT 1069.590 2794.275 1069.870 2794.645 ;
        RECT 1076.490 2794.275 1076.770 2794.645 ;
        RECT 1093.970 2794.275 1094.250 2794.645 ;
        RECT 1100.410 2794.275 1100.690 2794.645 ;
        RECT 1105.470 2794.275 1105.750 2794.645 ;
        RECT 1111.450 2794.275 1111.730 2794.645 ;
        RECT 1117.890 2794.275 1118.170 2794.645 ;
        RECT 1119.730 2794.275 1120.010 2794.645 ;
        RECT 948.160 2725.110 948.420 2725.430 ;
        RECT 944.930 2714.715 945.210 2715.085 ;
        RECT 948.220 2700.000 948.360 2725.110 ;
        RECT 979.960 2722.030 980.100 2794.275 ;
        RECT 1001.060 2794.130 1001.320 2794.275 ;
        RECT 1007.560 2794.110 1007.700 2794.275 ;
        RECT 1007.500 2793.790 1007.760 2794.110 ;
        RECT 1010.710 2793.595 1010.990 2793.965 ;
        RECT 1010.780 2789.690 1010.920 2793.595 ;
        RECT 1010.720 2789.370 1010.980 2789.690 ;
        RECT 989.560 2724.430 989.820 2724.750 ;
        RECT 979.900 2721.710 980.160 2722.030 ;
        RECT 968.860 2714.910 969.120 2715.230 ;
        RECT 958.740 2713.890 959.000 2714.210 ;
        RECT 958.800 2700.000 958.940 2713.890 ;
        RECT 968.920 2700.000 969.060 2714.910 ;
        RECT 979.440 2714.230 979.700 2714.550 ;
        RECT 979.500 2700.000 979.640 2714.230 ;
        RECT 989.620 2700.000 989.760 2724.430 ;
        RECT 1000.130 2718.115 1000.410 2718.485 ;
        RECT 1000.200 2700.000 1000.340 2718.115 ;
        RECT 1010.780 2716.250 1010.920 2789.370 ;
        RECT 1010.720 2715.930 1010.980 2716.250 ;
        RECT 1014.000 2715.910 1014.140 2794.275 ;
        RECT 1019.060 2791.050 1019.200 2794.275 ;
        RECT 1019.000 2790.730 1019.260 2791.050 ;
        RECT 1019.060 2788.670 1019.200 2790.730 ;
        RECT 1019.000 2788.350 1019.260 2788.670 ;
        RECT 1010.250 2715.395 1010.530 2715.765 ;
        RECT 1013.940 2715.590 1014.200 2715.910 ;
        RECT 1020.900 2715.570 1021.040 2794.275 ;
        RECT 1024.510 2792.915 1024.790 2793.285 ;
        RECT 1024.580 2788.670 1024.720 2792.915 ;
        RECT 1024.520 2788.350 1024.780 2788.670 ;
        RECT 1024.580 2716.930 1024.720 2788.350 ;
        RECT 1027.800 2718.630 1027.940 2794.275 ;
        RECT 1031.940 2791.730 1032.080 2794.275 ;
        RECT 1042.520 2793.770 1042.660 2794.275 ;
        RECT 1042.460 2793.450 1042.720 2793.770 ;
        RECT 1055.800 2793.450 1056.060 2793.770 ;
        RECT 1031.880 2791.410 1032.140 2791.730 ;
        RECT 1031.940 2789.010 1032.080 2791.410 ;
        RECT 1042.520 2789.350 1042.660 2793.450 ;
        RECT 1055.860 2793.285 1056.000 2793.450 ;
        RECT 1052.570 2792.915 1052.850 2793.285 ;
        RECT 1055.790 2792.915 1056.070 2793.285 ;
        RECT 1042.460 2789.030 1042.720 2789.350 ;
        RECT 1031.880 2788.690 1032.140 2789.010 ;
        RECT 1038.320 2788.690 1038.580 2789.010 ;
        RECT 1038.380 2788.525 1038.520 2788.690 ;
        RECT 1038.310 2788.155 1038.590 2788.525 ;
        RECT 1045.210 2788.155 1045.490 2788.525 ;
        RECT 1052.640 2788.330 1052.780 2792.915 ;
        RECT 1059.540 2792.070 1059.680 2794.275 ;
        RECT 1065.520 2793.090 1065.660 2794.275 ;
        RECT 1062.700 2792.770 1062.960 2793.090 ;
        RECT 1065.460 2792.770 1065.720 2793.090 ;
        RECT 1055.800 2791.750 1056.060 2792.070 ;
        RECT 1059.480 2791.750 1059.740 2792.070 ;
        RECT 1055.860 2789.690 1056.000 2791.750 ;
        RECT 1062.760 2791.050 1062.900 2792.770 ;
        RECT 1062.700 2790.730 1062.960 2791.050 ;
        RECT 1069.660 2790.710 1069.800 2794.275 ;
        RECT 1076.560 2791.730 1076.700 2794.275 ;
        RECT 1089.830 2793.595 1090.110 2793.965 ;
        RECT 1089.840 2793.450 1090.100 2793.595 ;
        RECT 1076.500 2791.410 1076.760 2791.730 ;
        RECT 1069.600 2790.390 1069.860 2790.710 ;
        RECT 1055.800 2789.370 1056.060 2789.690 ;
        RECT 1069.660 2788.670 1069.800 2790.390 ;
        RECT 1089.900 2789.010 1090.040 2793.450 ;
        RECT 1094.040 2792.750 1094.180 2794.275 ;
        RECT 1100.480 2794.110 1100.620 2794.275 ;
        RECT 1100.420 2793.790 1100.680 2794.110 ;
        RECT 1093.980 2792.430 1094.240 2792.750 ;
        RECT 1089.840 2788.690 1090.100 2789.010 ;
        RECT 1034.630 2787.475 1034.910 2787.845 ;
        RECT 1030.960 2723.410 1031.220 2723.730 ;
        RECT 1027.740 2718.310 1028.000 2718.630 ;
        RECT 1024.520 2716.610 1024.780 2716.930 ;
        RECT 1010.320 2700.000 1010.460 2715.395 ;
        RECT 1020.840 2715.250 1021.100 2715.570 ;
        RECT 1020.840 2714.570 1021.100 2714.890 ;
        RECT 1020.900 2700.000 1021.040 2714.570 ;
        RECT 1031.020 2700.000 1031.160 2723.410 ;
        RECT 1034.700 2718.290 1034.840 2787.475 ;
        RECT 1034.640 2717.970 1034.900 2718.290 ;
        RECT 1038.380 2717.270 1038.520 2788.155 ;
        RECT 1045.280 2787.990 1045.420 2788.155 ;
        RECT 1052.580 2788.010 1052.840 2788.330 ;
        RECT 1054.870 2788.155 1055.150 2788.525 ;
        RECT 1069.600 2788.350 1069.860 2788.670 ;
        RECT 1089.370 2788.155 1089.650 2788.525 ;
        RECT 1041.530 2787.475 1041.810 2787.845 ;
        RECT 1045.220 2787.670 1045.480 2787.990 ;
        RECT 1041.600 2717.950 1041.740 2787.475 ;
        RECT 1041.540 2717.630 1041.800 2717.950 ;
        RECT 1045.280 2717.610 1045.420 2787.670 ;
        RECT 1048.430 2787.475 1048.710 2787.845 ;
        RECT 1048.500 2717.610 1048.640 2787.475 ;
        RECT 1045.220 2717.290 1045.480 2717.610 ;
        RECT 1048.440 2717.290 1048.700 2717.610 ;
        RECT 1052.110 2717.435 1052.390 2717.805 ;
        RECT 1038.320 2716.950 1038.580 2717.270 ;
        RECT 1041.530 2716.755 1041.810 2717.125 ;
        RECT 1041.600 2700.000 1041.740 2716.755 ;
        RECT 1052.180 2700.000 1052.320 2717.435 ;
        RECT 1054.940 2717.270 1055.080 2788.155 ;
        RECT 1055.330 2787.475 1055.610 2787.845 ;
        RECT 1062.230 2787.475 1062.510 2787.845 ;
        RECT 1069.130 2787.475 1069.410 2787.845 ;
        RECT 1076.030 2787.475 1076.310 2787.845 ;
        RECT 1082.930 2787.475 1083.210 2787.845 ;
        RECT 1054.880 2716.950 1055.140 2717.270 ;
        RECT 1055.400 2716.250 1055.540 2787.475 ;
        RECT 1062.300 2727.890 1062.440 2787.475 ;
        RECT 1061.840 2727.750 1062.440 2727.890 ;
        RECT 1061.840 2716.930 1061.980 2727.750 ;
        RECT 1062.240 2722.730 1062.500 2723.050 ;
        RECT 1061.780 2716.610 1062.040 2716.930 ;
        RECT 1055.340 2715.930 1055.600 2716.250 ;
        RECT 1062.300 2700.000 1062.440 2722.730 ;
        RECT 1069.200 2715.570 1069.340 2787.475 ;
        RECT 1076.100 2716.590 1076.240 2787.475 ;
        RECT 1076.040 2716.270 1076.300 2716.590 ;
        RECT 1083.000 2715.910 1083.140 2787.475 ;
        RECT 1072.820 2715.590 1073.080 2715.910 ;
        RECT 1082.940 2715.590 1083.200 2715.910 ;
        RECT 1069.140 2715.250 1069.400 2715.570 ;
        RECT 1072.880 2700.000 1073.020 2715.590 ;
        RECT 1089.440 2715.230 1089.580 2788.155 ;
        RECT 1094.040 2787.990 1094.180 2792.430 ;
        RECT 1100.480 2788.330 1100.620 2793.790 ;
        RECT 1103.640 2793.285 1103.900 2793.430 ;
        RECT 1103.630 2792.915 1103.910 2793.285 ;
        RECT 1105.540 2792.070 1105.680 2794.275 ;
        RECT 1111.520 2793.090 1111.660 2794.275 ;
        RECT 1111.460 2792.770 1111.720 2793.090 ;
        RECT 1105.480 2791.750 1105.740 2792.070 ;
        RECT 1117.960 2790.030 1118.100 2794.275 ;
        RECT 1119.800 2791.730 1119.940 2794.275 ;
        RECT 1129.920 2793.770 1130.060 2799.035 ;
        RECT 1136.290 2796.315 1136.570 2796.685 ;
        RECT 1129.860 2793.450 1130.120 2793.770 ;
        RECT 1136.360 2793.430 1136.500 2796.315 ;
        RECT 1140.430 2794.275 1140.710 2794.645 ;
        RECT 1136.300 2793.110 1136.560 2793.430 ;
        RECT 1140.500 2792.750 1140.640 2794.275 ;
        RECT 1146.940 2794.110 1147.080 2799.715 ;
        RECT 1179.530 2794.275 1179.810 2794.645 ;
        RECT 1186.430 2794.275 1186.710 2794.645 ;
        RECT 1200.230 2794.275 1200.510 2794.645 ;
        RECT 1146.880 2793.790 1147.140 2794.110 ;
        RECT 1159.750 2793.595 1160.030 2793.965 ;
        RECT 1166.190 2793.595 1166.470 2793.965 ;
        RECT 1173.090 2793.595 1173.370 2793.965 ;
        RECT 1159.290 2792.915 1159.570 2793.285 ;
        RECT 1159.300 2792.770 1159.560 2792.915 ;
        RECT 1140.440 2792.430 1140.700 2792.750 ;
        RECT 1152.390 2792.235 1152.670 2792.605 ;
        RECT 1152.460 2792.070 1152.600 2792.235 ;
        RECT 1152.400 2791.750 1152.660 2792.070 ;
        RECT 1119.740 2791.410 1120.000 2791.730 ;
        RECT 1159.820 2791.050 1159.960 2793.595 ;
        RECT 1166.260 2791.730 1166.400 2793.595 ;
        RECT 1173.100 2793.450 1173.360 2793.595 ;
        RECT 1166.200 2791.410 1166.460 2791.730 ;
        RECT 1159.760 2790.730 1160.020 2791.050 ;
        RECT 1117.900 2789.710 1118.160 2790.030 ;
        RECT 1100.420 2788.010 1100.680 2788.330 ;
        RECT 1131.230 2788.155 1131.510 2788.525 ;
        RECT 1165.730 2788.155 1166.010 2788.525 ;
        RECT 1089.830 2787.475 1090.110 2787.845 ;
        RECT 1093.980 2787.670 1094.240 2787.990 ;
        RECT 1096.730 2787.475 1097.010 2787.845 ;
        RECT 1103.630 2787.475 1103.910 2787.845 ;
        RECT 1110.530 2787.475 1110.810 2787.845 ;
        RECT 1117.430 2787.475 1117.710 2787.845 ;
        RECT 1124.330 2787.475 1124.610 2787.845 ;
        RECT 1130.770 2787.475 1131.050 2787.845 ;
        RECT 1082.940 2714.910 1083.200 2715.230 ;
        RECT 1089.380 2714.910 1089.640 2715.230 ;
        RECT 1083.000 2700.000 1083.140 2714.910 ;
        RECT 1089.900 2712.850 1090.040 2787.475 ;
        RECT 1093.520 2718.310 1093.780 2718.630 ;
        RECT 1089.840 2712.530 1090.100 2712.850 ;
        RECT 1093.580 2700.000 1093.720 2718.310 ;
        RECT 1096.800 2712.510 1096.940 2787.475 ;
        RECT 1103.700 2718.970 1103.840 2787.475 ;
        RECT 1103.640 2718.650 1103.900 2718.970 ;
        RECT 1102.720 2718.310 1102.980 2718.630 ;
        RECT 1102.780 2713.190 1102.920 2718.310 ;
        RECT 1103.640 2717.970 1103.900 2718.290 ;
        RECT 1102.720 2712.870 1102.980 2713.190 ;
        RECT 1096.740 2712.190 1097.000 2712.510 ;
        RECT 1103.700 2700.000 1103.840 2717.970 ;
        RECT 1110.600 2713.530 1110.740 2787.475 ;
        RECT 1114.220 2717.630 1114.480 2717.950 ;
        RECT 1110.540 2713.210 1110.800 2713.530 ;
        RECT 1114.280 2700.000 1114.420 2717.630 ;
        RECT 1117.500 2714.210 1117.640 2787.475 ;
        RECT 1124.400 2726.530 1124.540 2787.475 ;
        RECT 1123.480 2726.390 1124.540 2726.530 ;
        RECT 1117.440 2713.890 1117.700 2714.210 ;
        RECT 1123.480 2713.870 1123.620 2726.390 ;
        RECT 1124.340 2717.290 1124.600 2717.610 ;
        RECT 1123.420 2713.550 1123.680 2713.870 ;
        RECT 1124.400 2700.000 1124.540 2717.290 ;
        RECT 1130.840 2714.890 1130.980 2787.475 ;
        RECT 1130.780 2714.570 1131.040 2714.890 ;
        RECT 1131.300 2714.550 1131.440 2788.155 ;
        RECT 1138.130 2787.475 1138.410 2787.845 ;
        RECT 1145.030 2787.475 1145.310 2787.845 ;
        RECT 1151.930 2787.475 1152.210 2787.845 ;
        RECT 1158.830 2787.475 1159.110 2787.845 ;
        RECT 1165.270 2787.475 1165.550 2787.845 ;
        RECT 1138.200 2718.630 1138.340 2787.475 ;
        RECT 1138.140 2718.310 1138.400 2718.630 ;
        RECT 1145.100 2718.290 1145.240 2787.475 ;
        RECT 1145.040 2717.970 1145.300 2718.290 ;
        RECT 1152.000 2717.950 1152.140 2787.475 ;
        RECT 1151.940 2717.630 1152.200 2717.950 ;
        RECT 1158.900 2717.610 1159.040 2787.475 ;
        RECT 1158.840 2717.290 1159.100 2717.610 ;
        RECT 1134.920 2716.950 1135.180 2717.270 ;
        RECT 1131.240 2714.230 1131.500 2714.550 ;
        RECT 1134.980 2700.000 1135.120 2716.950 ;
        RECT 1165.340 2716.930 1165.480 2787.475 ;
        RECT 1165.800 2717.270 1165.940 2788.155 ;
        RECT 1172.630 2787.475 1172.910 2787.845 ;
        RECT 1165.740 2716.950 1166.000 2717.270 ;
        RECT 1155.620 2716.610 1155.880 2716.930 ;
        RECT 1165.280 2716.610 1165.540 2716.930 ;
        RECT 1145.500 2715.930 1145.760 2716.250 ;
        RECT 1145.560 2700.000 1145.700 2715.930 ;
        RECT 1155.680 2700.000 1155.820 2716.610 ;
        RECT 1172.700 2716.250 1172.840 2787.475 ;
        RECT 1179.600 2716.590 1179.740 2794.275 ;
        RECT 1179.990 2793.595 1180.270 2793.965 ;
        RECT 1180.060 2793.430 1180.200 2793.595 ;
        RECT 1180.000 2793.110 1180.260 2793.430 ;
        RECT 1176.320 2716.270 1176.580 2716.590 ;
        RECT 1179.540 2716.270 1179.800 2716.590 ;
        RECT 1172.640 2715.930 1172.900 2716.250 ;
        RECT 1166.200 2715.250 1166.460 2715.570 ;
        RECT 1166.260 2700.000 1166.400 2715.250 ;
        RECT 1176.380 2700.000 1176.520 2716.270 ;
        RECT 1186.500 2715.570 1186.640 2794.275 ;
        RECT 1186.890 2792.915 1187.170 2793.285 ;
        RECT 1186.960 2792.750 1187.100 2792.915 ;
        RECT 1186.900 2792.430 1187.160 2792.750 ;
        RECT 1193.790 2791.555 1194.070 2791.925 ;
        RECT 1193.800 2791.410 1194.060 2791.555 ;
        RECT 1193.330 2790.195 1193.610 2790.565 ;
        RECT 1193.400 2715.910 1193.540 2790.195 ;
        RECT 1186.900 2715.590 1187.160 2715.910 ;
        RECT 1193.340 2715.590 1193.600 2715.910 ;
        RECT 1186.440 2715.250 1186.700 2715.570 ;
        RECT 1186.960 2700.000 1187.100 2715.590 ;
        RECT 1200.300 2715.230 1200.440 2794.275 ;
        RECT 1410.460 2794.130 1410.720 2794.450 ;
        RECT 1409.540 2792.090 1409.800 2792.410 ;
        RECT 1409.080 2791.410 1409.340 2791.730 ;
        RECT 1290.400 2718.310 1290.660 2718.630 ;
        RECT 1197.020 2714.910 1197.280 2715.230 ;
        RECT 1200.240 2714.910 1200.500 2715.230 ;
        RECT 1197.080 2700.000 1197.220 2714.910 ;
        RECT 1280.280 2714.570 1280.540 2714.890 ;
        RECT 1269.700 2714.230 1269.960 2714.550 ;
        RECT 1249.000 2713.890 1249.260 2714.210 ;
        RECT 1238.880 2713.210 1239.140 2713.530 ;
        RECT 1228.300 2712.870 1228.560 2713.190 ;
        RECT 1207.600 2712.530 1207.860 2712.850 ;
        RECT 1207.660 2700.000 1207.800 2712.530 ;
        RECT 1217.720 2712.190 1217.980 2712.510 ;
        RECT 1217.780 2700.000 1217.920 2712.190 ;
        RECT 1228.360 2700.000 1228.500 2712.870 ;
        RECT 1238.940 2700.000 1239.080 2713.210 ;
        RECT 1249.060 2700.000 1249.200 2713.890 ;
        RECT 1259.580 2713.550 1259.840 2713.870 ;
        RECT 1259.640 2700.000 1259.780 2713.550 ;
        RECT 1269.760 2700.000 1269.900 2714.230 ;
        RECT 1280.340 2700.000 1280.480 2714.570 ;
        RECT 1290.460 2700.000 1290.600 2718.310 ;
        RECT 1300.980 2717.970 1301.240 2718.290 ;
        RECT 1301.040 2700.000 1301.180 2717.970 ;
        RECT 1311.100 2717.630 1311.360 2717.950 ;
        RECT 1311.160 2700.000 1311.300 2717.630 ;
        RECT 1321.680 2717.290 1321.940 2717.610 ;
        RECT 1321.740 2700.000 1321.880 2717.290 ;
        RECT 1332.260 2716.950 1332.520 2717.270 ;
        RECT 1332.320 2700.000 1332.460 2716.950 ;
        RECT 1342.380 2716.610 1342.640 2716.930 ;
        RECT 1342.440 2700.000 1342.580 2716.610 ;
        RECT 1363.080 2716.270 1363.340 2716.590 ;
        RECT 1352.960 2715.930 1353.220 2716.250 ;
        RECT 1353.020 2700.000 1353.160 2715.930 ;
        RECT 1363.140 2700.000 1363.280 2716.270 ;
        RECT 1383.780 2715.590 1384.040 2715.910 ;
        RECT 1373.660 2715.250 1373.920 2715.570 ;
        RECT 1373.720 2700.000 1373.860 2715.250 ;
        RECT 1383.840 2700.000 1383.980 2715.590 ;
        RECT 1394.360 2714.910 1394.620 2715.230 ;
        RECT 1394.420 2700.000 1394.560 2714.910 ;
        RECT 345.160 2699.870 346.760 2700.000 ;
        RECT 335.900 2696.000 336.180 2699.870 ;
        RECT 346.480 2696.000 346.760 2699.870 ;
        RECT 356.600 2696.000 356.880 2700.000 ;
        RECT 367.180 2696.000 367.460 2700.000 ;
        RECT 377.300 2696.000 377.580 2700.000 ;
        RECT 387.880 2696.000 388.160 2700.000 ;
        RECT 398.460 2696.000 398.740 2700.000 ;
        RECT 408.580 2696.000 408.860 2700.000 ;
        RECT 419.160 2696.000 419.440 2700.000 ;
        RECT 429.280 2696.000 429.560 2700.000 ;
        RECT 439.860 2696.000 440.140 2700.000 ;
        RECT 449.980 2696.000 450.260 2700.000 ;
        RECT 460.560 2696.000 460.840 2700.000 ;
        RECT 470.680 2696.000 470.960 2700.000 ;
        RECT 481.260 2696.000 481.540 2700.000 ;
        RECT 491.840 2696.000 492.120 2700.000 ;
        RECT 501.960 2696.000 502.240 2700.000 ;
        RECT 512.540 2696.000 512.820 2700.000 ;
        RECT 522.660 2696.000 522.940 2700.000 ;
        RECT 533.240 2696.000 533.520 2700.000 ;
        RECT 543.360 2696.000 543.640 2700.000 ;
        RECT 553.940 2696.000 554.220 2700.000 ;
        RECT 564.060 2696.000 564.340 2700.000 ;
        RECT 574.640 2696.000 574.920 2700.000 ;
        RECT 585.220 2699.870 586.340 2700.000 ;
        RECT 585.220 2696.000 585.500 2699.870 ;
        RECT 595.340 2696.000 595.620 2700.000 ;
        RECT 605.920 2699.870 607.040 2700.000 ;
        RECT 605.920 2696.000 606.200 2699.870 ;
        RECT 616.040 2696.000 616.320 2700.000 ;
        RECT 626.620 2699.870 627.740 2700.000 ;
        RECT 626.620 2696.000 626.900 2699.870 ;
        RECT 636.740 2696.000 637.020 2700.000 ;
        RECT 647.320 2699.870 648.440 2700.000 ;
        RECT 647.320 2696.000 647.600 2699.870 ;
        RECT 657.440 2696.000 657.720 2700.000 ;
        RECT 668.020 2696.000 668.300 2700.000 ;
        RECT 678.600 2696.000 678.880 2700.000 ;
        RECT 688.720 2696.000 689.000 2700.000 ;
        RECT 699.300 2696.000 699.580 2700.000 ;
        RECT 709.420 2696.000 709.700 2700.000 ;
        RECT 720.000 2696.000 720.280 2700.000 ;
        RECT 730.120 2696.000 730.400 2700.000 ;
        RECT 740.700 2696.000 740.980 2700.000 ;
        RECT 750.820 2696.000 751.100 2700.000 ;
        RECT 761.400 2696.000 761.680 2700.000 ;
        RECT 771.980 2696.000 772.260 2700.000 ;
        RECT 782.100 2696.000 782.380 2700.000 ;
        RECT 792.680 2696.000 792.960 2700.000 ;
        RECT 802.800 2696.000 803.080 2700.000 ;
        RECT 813.380 2696.000 813.660 2700.000 ;
        RECT 823.500 2696.000 823.780 2700.000 ;
        RECT 834.080 2696.000 834.360 2700.000 ;
        RECT 844.200 2696.000 844.480 2700.000 ;
        RECT 854.780 2696.000 855.060 2700.000 ;
        RECT 865.360 2696.000 865.640 2700.000 ;
        RECT 875.480 2696.000 875.760 2700.000 ;
        RECT 886.060 2696.000 886.340 2700.000 ;
        RECT 896.180 2696.000 896.460 2700.000 ;
        RECT 906.760 2696.000 907.040 2700.000 ;
        RECT 916.880 2696.000 917.160 2700.000 ;
        RECT 927.460 2696.000 927.740 2700.000 ;
        RECT 937.580 2696.000 937.860 2700.000 ;
        RECT 948.160 2696.000 948.440 2700.000 ;
        RECT 958.740 2696.000 959.020 2700.000 ;
        RECT 968.860 2696.000 969.140 2700.000 ;
        RECT 979.440 2696.000 979.720 2700.000 ;
        RECT 989.560 2696.000 989.840 2700.000 ;
        RECT 1000.140 2696.000 1000.420 2700.000 ;
        RECT 1010.260 2696.000 1010.540 2700.000 ;
        RECT 1020.840 2696.000 1021.120 2700.000 ;
        RECT 1030.960 2696.000 1031.240 2700.000 ;
        RECT 1041.540 2696.000 1041.820 2700.000 ;
        RECT 1052.120 2696.000 1052.400 2700.000 ;
        RECT 1062.240 2696.000 1062.520 2700.000 ;
        RECT 1072.820 2696.000 1073.100 2700.000 ;
        RECT 1082.940 2696.000 1083.220 2700.000 ;
        RECT 1093.520 2696.000 1093.800 2700.000 ;
        RECT 1103.640 2696.000 1103.920 2700.000 ;
        RECT 1114.220 2696.000 1114.500 2700.000 ;
        RECT 1124.340 2696.000 1124.620 2700.000 ;
        RECT 1134.920 2696.000 1135.200 2700.000 ;
        RECT 1145.500 2696.000 1145.780 2700.000 ;
        RECT 1155.620 2696.000 1155.900 2700.000 ;
        RECT 1166.200 2696.000 1166.480 2700.000 ;
        RECT 1176.320 2696.000 1176.600 2700.000 ;
        RECT 1186.900 2696.000 1187.180 2700.000 ;
        RECT 1197.020 2696.000 1197.300 2700.000 ;
        RECT 1207.600 2696.000 1207.880 2700.000 ;
        RECT 1217.720 2696.000 1218.000 2700.000 ;
        RECT 1228.300 2696.000 1228.580 2700.000 ;
        RECT 1238.880 2696.000 1239.160 2700.000 ;
        RECT 1249.000 2696.000 1249.280 2700.000 ;
        RECT 1259.580 2696.000 1259.860 2700.000 ;
        RECT 1269.700 2696.000 1269.980 2700.000 ;
        RECT 1280.280 2696.000 1280.560 2700.000 ;
        RECT 1290.400 2696.000 1290.680 2700.000 ;
        RECT 1300.980 2696.000 1301.260 2700.000 ;
        RECT 1311.100 2696.000 1311.380 2700.000 ;
        RECT 1321.680 2696.000 1321.960 2700.000 ;
        RECT 1332.260 2696.000 1332.540 2700.000 ;
        RECT 1342.380 2696.000 1342.660 2700.000 ;
        RECT 1352.960 2696.000 1353.240 2700.000 ;
        RECT 1363.080 2696.000 1363.360 2700.000 ;
        RECT 1373.660 2696.000 1373.940 2700.000 ;
        RECT 1383.780 2696.000 1384.060 2700.000 ;
        RECT 1394.360 2696.000 1394.640 2700.000 ;
        RECT 1408.620 2697.570 1408.880 2697.890 ;
      LAYER met2 ;
        RECT 300.030 2695.720 304.800 2696.000 ;
        RECT 305.640 2695.720 314.920 2696.000 ;
        RECT 315.760 2695.720 325.500 2696.000 ;
        RECT 326.340 2695.720 335.620 2696.000 ;
        RECT 336.460 2695.720 346.200 2696.000 ;
        RECT 347.040 2695.720 356.320 2696.000 ;
        RECT 357.160 2695.720 366.900 2696.000 ;
        RECT 367.740 2695.720 377.020 2696.000 ;
        RECT 377.860 2695.720 387.600 2696.000 ;
        RECT 388.440 2695.720 398.180 2696.000 ;
        RECT 399.020 2695.720 408.300 2696.000 ;
        RECT 409.140 2695.720 418.880 2696.000 ;
        RECT 419.720 2695.720 429.000 2696.000 ;
        RECT 429.840 2695.720 439.580 2696.000 ;
        RECT 440.420 2695.720 449.700 2696.000 ;
        RECT 450.540 2695.720 460.280 2696.000 ;
        RECT 461.120 2695.720 470.400 2696.000 ;
        RECT 471.240 2695.720 480.980 2696.000 ;
        RECT 481.820 2695.720 491.560 2696.000 ;
        RECT 492.400 2695.720 501.680 2696.000 ;
        RECT 502.520 2695.720 512.260 2696.000 ;
        RECT 513.100 2695.720 522.380 2696.000 ;
        RECT 523.220 2695.720 532.960 2696.000 ;
        RECT 533.800 2695.720 543.080 2696.000 ;
        RECT 543.920 2695.720 553.660 2696.000 ;
        RECT 554.500 2695.720 563.780 2696.000 ;
        RECT 564.620 2695.720 574.360 2696.000 ;
        RECT 575.200 2695.720 584.940 2696.000 ;
        RECT 585.780 2695.720 595.060 2696.000 ;
        RECT 595.900 2695.720 605.640 2696.000 ;
        RECT 606.480 2695.720 615.760 2696.000 ;
        RECT 616.600 2695.720 626.340 2696.000 ;
        RECT 627.180 2695.720 636.460 2696.000 ;
        RECT 637.300 2695.720 647.040 2696.000 ;
        RECT 647.880 2695.720 657.160 2696.000 ;
        RECT 658.000 2695.720 667.740 2696.000 ;
        RECT 668.580 2695.720 678.320 2696.000 ;
        RECT 679.160 2695.720 688.440 2696.000 ;
        RECT 689.280 2695.720 699.020 2696.000 ;
        RECT 699.860 2695.720 709.140 2696.000 ;
        RECT 709.980 2695.720 719.720 2696.000 ;
        RECT 720.560 2695.720 729.840 2696.000 ;
        RECT 730.680 2695.720 740.420 2696.000 ;
        RECT 741.260 2695.720 750.540 2696.000 ;
        RECT 751.380 2695.720 761.120 2696.000 ;
        RECT 761.960 2695.720 771.700 2696.000 ;
        RECT 772.540 2695.720 781.820 2696.000 ;
        RECT 782.660 2695.720 792.400 2696.000 ;
        RECT 793.240 2695.720 802.520 2696.000 ;
        RECT 803.360 2695.720 813.100 2696.000 ;
        RECT 813.940 2695.720 823.220 2696.000 ;
        RECT 824.060 2695.720 833.800 2696.000 ;
        RECT 834.640 2695.720 843.920 2696.000 ;
        RECT 844.760 2695.720 854.500 2696.000 ;
        RECT 855.340 2695.720 865.080 2696.000 ;
        RECT 865.920 2695.720 875.200 2696.000 ;
        RECT 876.040 2695.720 885.780 2696.000 ;
        RECT 886.620 2695.720 895.900 2696.000 ;
        RECT 896.740 2695.720 906.480 2696.000 ;
        RECT 907.320 2695.720 916.600 2696.000 ;
        RECT 917.440 2695.720 927.180 2696.000 ;
        RECT 928.020 2695.720 937.300 2696.000 ;
        RECT 938.140 2695.720 947.880 2696.000 ;
        RECT 948.720 2695.720 958.460 2696.000 ;
        RECT 959.300 2695.720 968.580 2696.000 ;
        RECT 969.420 2695.720 979.160 2696.000 ;
        RECT 980.000 2695.720 989.280 2696.000 ;
        RECT 990.120 2695.720 999.860 2696.000 ;
        RECT 1000.700 2695.720 1009.980 2696.000 ;
        RECT 1010.820 2695.720 1020.560 2696.000 ;
        RECT 1021.400 2695.720 1030.680 2696.000 ;
        RECT 1031.520 2695.720 1041.260 2696.000 ;
        RECT 1042.100 2695.720 1051.840 2696.000 ;
        RECT 1052.680 2695.720 1061.960 2696.000 ;
        RECT 1062.800 2695.720 1072.540 2696.000 ;
        RECT 1073.380 2695.720 1082.660 2696.000 ;
        RECT 1083.500 2695.720 1093.240 2696.000 ;
        RECT 1094.080 2695.720 1103.360 2696.000 ;
        RECT 1104.200 2695.720 1113.940 2696.000 ;
        RECT 1114.780 2695.720 1124.060 2696.000 ;
        RECT 1124.900 2695.720 1134.640 2696.000 ;
        RECT 1135.480 2695.720 1145.220 2696.000 ;
        RECT 1146.060 2695.720 1155.340 2696.000 ;
        RECT 1156.180 2695.720 1165.920 2696.000 ;
        RECT 1166.760 2695.720 1176.040 2696.000 ;
        RECT 1176.880 2695.720 1186.620 2696.000 ;
        RECT 1187.460 2695.720 1196.740 2696.000 ;
        RECT 1197.580 2695.720 1207.320 2696.000 ;
        RECT 1208.160 2695.720 1217.440 2696.000 ;
        RECT 1218.280 2695.720 1228.020 2696.000 ;
        RECT 1228.860 2695.720 1238.600 2696.000 ;
        RECT 1239.440 2695.720 1248.720 2696.000 ;
        RECT 1249.560 2695.720 1259.300 2696.000 ;
        RECT 1260.140 2695.720 1269.420 2696.000 ;
        RECT 1270.260 2695.720 1280.000 2696.000 ;
        RECT 1280.840 2695.720 1290.120 2696.000 ;
        RECT 1290.960 2695.720 1300.700 2696.000 ;
        RECT 1301.540 2695.720 1310.820 2696.000 ;
        RECT 1311.660 2695.720 1321.400 2696.000 ;
        RECT 1322.240 2695.720 1331.980 2696.000 ;
        RECT 1332.820 2695.720 1342.100 2696.000 ;
        RECT 1342.940 2695.720 1352.680 2696.000 ;
        RECT 1353.520 2695.720 1362.800 2696.000 ;
        RECT 1363.640 2695.720 1373.380 2696.000 ;
        RECT 1374.220 2695.720 1383.500 2696.000 ;
        RECT 1384.340 2695.720 1394.080 2696.000 ;
        RECT 1394.920 2695.720 1396.470 2696.000 ;
        RECT 300.030 1604.280 1396.470 2695.720 ;
      LAYER met2 ;
        RECT 1408.680 2695.365 1408.820 2697.570 ;
        RECT 1408.610 2694.995 1408.890 2695.365 ;
        RECT 1408.620 2690.770 1408.880 2691.090 ;
        RECT 1408.680 2685.165 1408.820 2690.770 ;
        RECT 1408.610 2684.795 1408.890 2685.165 ;
        RECT 1408.620 2676.830 1408.880 2677.150 ;
        RECT 1408.680 2674.965 1408.820 2676.830 ;
        RECT 1408.610 2674.595 1408.890 2674.965 ;
        RECT 1408.620 2670.030 1408.880 2670.350 ;
        RECT 1408.680 2664.765 1408.820 2670.030 ;
        RECT 1408.610 2664.395 1408.890 2664.765 ;
        RECT 1408.620 2656.090 1408.880 2656.410 ;
        RECT 1408.680 2654.565 1408.820 2656.090 ;
        RECT 1408.610 2654.195 1408.890 2654.565 ;
        RECT 1408.620 2649.290 1408.880 2649.610 ;
        RECT 1408.680 2644.365 1408.820 2649.290 ;
        RECT 1408.610 2643.995 1408.890 2644.365 ;
        RECT 1408.620 2635.350 1408.880 2635.670 ;
        RECT 1408.680 2634.165 1408.820 2635.350 ;
        RECT 1408.610 2633.795 1408.890 2634.165 ;
        RECT 1408.620 2628.550 1408.880 2628.870 ;
        RECT 1408.680 2623.965 1408.820 2628.550 ;
        RECT 1408.610 2623.595 1408.890 2623.965 ;
        RECT 1408.620 2614.610 1408.880 2614.930 ;
        RECT 1408.680 2613.765 1408.820 2614.610 ;
        RECT 1408.610 2613.395 1408.890 2613.765 ;
        RECT 1408.620 2607.810 1408.880 2608.130 ;
        RECT 1408.680 2603.565 1408.820 2607.810 ;
        RECT 1408.610 2603.195 1408.890 2603.565 ;
        RECT 1408.620 2594.210 1408.880 2594.530 ;
        RECT 1408.680 2593.365 1408.820 2594.210 ;
        RECT 1408.610 2592.995 1408.890 2593.365 ;
        RECT 1408.620 2587.070 1408.880 2587.390 ;
        RECT 1408.680 2583.165 1408.820 2587.070 ;
        RECT 1408.610 2582.795 1408.890 2583.165 ;
        RECT 1408.620 2573.470 1408.880 2573.790 ;
        RECT 1408.680 2572.965 1408.820 2573.470 ;
        RECT 1408.610 2572.595 1408.890 2572.965 ;
        RECT 1408.620 2566.330 1408.880 2566.650 ;
        RECT 1408.680 2562.765 1408.820 2566.330 ;
        RECT 1408.610 2562.395 1408.890 2562.765 ;
        RECT 1408.620 2552.730 1408.880 2553.050 ;
        RECT 1408.680 2552.565 1408.820 2552.730 ;
        RECT 1408.610 2552.195 1408.890 2552.565 ;
        RECT 1408.620 2545.930 1408.880 2546.250 ;
        RECT 1408.680 2542.365 1408.820 2545.930 ;
        RECT 1408.610 2541.995 1408.890 2542.365 ;
        RECT 1408.620 2532.165 1408.880 2532.310 ;
        RECT 1408.610 2531.795 1408.890 2532.165 ;
        RECT 1408.620 2525.190 1408.880 2525.510 ;
        RECT 1408.680 2521.965 1408.820 2525.190 ;
        RECT 1408.610 2521.595 1408.890 2521.965 ;
        RECT 1408.610 2511.395 1408.890 2511.765 ;
        RECT 1408.620 2511.250 1408.880 2511.395 ;
        RECT 1408.620 2504.450 1408.880 2504.770 ;
        RECT 1408.680 2501.565 1408.820 2504.450 ;
        RECT 1408.610 2501.195 1408.890 2501.565 ;
        RECT 1408.620 2497.310 1408.880 2497.630 ;
        RECT 1408.680 2491.365 1408.820 2497.310 ;
        RECT 1408.610 2490.995 1408.890 2491.365 ;
        RECT 1408.620 2483.710 1408.880 2484.030 ;
        RECT 1408.680 2481.165 1408.820 2483.710 ;
        RECT 1408.610 2480.795 1408.890 2481.165 ;
        RECT 1408.620 2476.910 1408.880 2477.230 ;
        RECT 1408.680 2470.965 1408.820 2476.910 ;
        RECT 1408.610 2470.595 1408.890 2470.965 ;
        RECT 1408.620 2462.970 1408.880 2463.290 ;
        RECT 1408.680 2460.765 1408.820 2462.970 ;
        RECT 1408.610 2460.395 1408.890 2460.765 ;
        RECT 1408.620 2456.170 1408.880 2456.490 ;
        RECT 1408.680 2450.565 1408.820 2456.170 ;
        RECT 1408.610 2450.195 1408.890 2450.565 ;
        RECT 1408.620 2442.230 1408.880 2442.550 ;
        RECT 1408.680 2440.365 1408.820 2442.230 ;
        RECT 1408.610 2439.995 1408.890 2440.365 ;
        RECT 1408.620 2435.430 1408.880 2435.750 ;
        RECT 1408.680 2430.165 1408.820 2435.430 ;
        RECT 1408.610 2429.795 1408.890 2430.165 ;
        RECT 1408.620 2421.490 1408.880 2421.810 ;
        RECT 1408.680 2419.965 1408.820 2421.490 ;
        RECT 1408.610 2419.595 1408.890 2419.965 ;
        RECT 1408.620 2414.690 1408.880 2415.010 ;
        RECT 1408.680 2409.765 1408.820 2414.690 ;
        RECT 1408.610 2409.395 1408.890 2409.765 ;
        RECT 1408.620 2400.750 1408.880 2401.070 ;
        RECT 1408.680 2399.565 1408.820 2400.750 ;
        RECT 1408.610 2399.195 1408.890 2399.565 ;
        RECT 1408.620 2393.950 1408.880 2394.270 ;
        RECT 1408.680 2389.365 1408.820 2393.950 ;
        RECT 1408.610 2388.995 1408.890 2389.365 ;
        RECT 1408.620 2380.010 1408.880 2380.330 ;
        RECT 1408.680 2379.165 1408.820 2380.010 ;
        RECT 1408.610 2378.795 1408.890 2379.165 ;
        RECT 1408.620 2373.210 1408.880 2373.530 ;
        RECT 1408.680 2368.965 1408.820 2373.210 ;
        RECT 1408.610 2368.595 1408.890 2368.965 ;
        RECT 1408.620 2359.610 1408.880 2359.930 ;
        RECT 1408.680 2358.765 1408.820 2359.610 ;
        RECT 1408.610 2358.395 1408.890 2358.765 ;
        RECT 1408.620 2352.470 1408.880 2352.790 ;
        RECT 1408.680 2348.565 1408.820 2352.470 ;
        RECT 1408.610 2348.195 1408.890 2348.565 ;
        RECT 1408.620 2338.870 1408.880 2339.190 ;
        RECT 1408.680 2338.365 1408.820 2338.870 ;
        RECT 1408.610 2337.995 1408.890 2338.365 ;
        RECT 1408.620 2331.730 1408.880 2332.050 ;
        RECT 1408.680 2328.165 1408.820 2331.730 ;
        RECT 1408.610 2327.795 1408.890 2328.165 ;
        RECT 1408.620 2318.130 1408.880 2318.450 ;
        RECT 1408.680 2317.965 1408.820 2318.130 ;
        RECT 1408.610 2317.595 1408.890 2317.965 ;
        RECT 1408.620 2311.330 1408.880 2311.650 ;
        RECT 1408.680 2307.765 1408.820 2311.330 ;
        RECT 1408.610 2307.395 1408.890 2307.765 ;
        RECT 1408.620 2297.565 1408.880 2297.710 ;
        RECT 1408.610 2297.195 1408.890 2297.565 ;
        RECT 1408.620 2290.590 1408.880 2290.910 ;
        RECT 1408.680 2287.365 1408.820 2290.590 ;
        RECT 1408.610 2286.995 1408.890 2287.365 ;
        RECT 1408.610 2276.795 1408.890 2277.165 ;
        RECT 1408.620 2276.650 1408.880 2276.795 ;
        RECT 1408.620 2269.850 1408.880 2270.170 ;
        RECT 1408.680 2266.965 1408.820 2269.850 ;
        RECT 1408.610 2266.595 1408.890 2266.965 ;
        RECT 1408.620 2262.710 1408.880 2263.030 ;
        RECT 1408.680 2256.765 1408.820 2262.710 ;
        RECT 1408.610 2256.395 1408.890 2256.765 ;
        RECT 1408.620 2249.110 1408.880 2249.430 ;
        RECT 1408.680 2246.565 1408.820 2249.110 ;
        RECT 1408.610 2246.195 1408.890 2246.565 ;
        RECT 1408.620 2242.310 1408.880 2242.630 ;
        RECT 1408.680 2236.365 1408.820 2242.310 ;
        RECT 1408.610 2235.995 1408.890 2236.365 ;
        RECT 1408.620 2228.370 1408.880 2228.690 ;
        RECT 1408.680 2226.165 1408.820 2228.370 ;
        RECT 1408.610 2225.795 1408.890 2226.165 ;
        RECT 1408.620 2221.570 1408.880 2221.890 ;
        RECT 1408.680 2215.965 1408.820 2221.570 ;
        RECT 1408.610 2215.595 1408.890 2215.965 ;
        RECT 1408.620 2207.630 1408.880 2207.950 ;
        RECT 1408.680 2205.765 1408.820 2207.630 ;
        RECT 1408.610 2205.395 1408.890 2205.765 ;
        RECT 1408.620 2200.830 1408.880 2201.150 ;
        RECT 1408.680 2195.565 1408.820 2200.830 ;
        RECT 1408.610 2195.195 1408.890 2195.565 ;
        RECT 1408.620 2186.890 1408.880 2187.210 ;
        RECT 1408.680 2185.365 1408.820 2186.890 ;
        RECT 1408.610 2184.995 1408.890 2185.365 ;
        RECT 1408.620 2180.090 1408.880 2180.410 ;
        RECT 1408.680 2175.165 1408.820 2180.090 ;
        RECT 1408.610 2174.795 1408.890 2175.165 ;
        RECT 1408.620 2166.150 1408.880 2166.470 ;
        RECT 1408.680 2164.965 1408.820 2166.150 ;
        RECT 1408.610 2164.595 1408.890 2164.965 ;
        RECT 1408.620 2159.350 1408.880 2159.670 ;
        RECT 1408.680 2155.445 1408.820 2159.350 ;
        RECT 1408.610 2155.075 1408.890 2155.445 ;
        RECT 1408.620 2145.410 1408.880 2145.730 ;
        RECT 1408.680 2145.245 1408.820 2145.410 ;
        RECT 1408.610 2144.875 1408.890 2145.245 ;
        RECT 1408.620 2138.610 1408.880 2138.930 ;
        RECT 1408.680 2135.045 1408.820 2138.610 ;
        RECT 1408.610 2134.675 1408.890 2135.045 ;
        RECT 1408.620 2125.010 1408.880 2125.330 ;
        RECT 1408.680 2124.845 1408.820 2125.010 ;
        RECT 1408.610 2124.475 1408.890 2124.845 ;
        RECT 1408.620 2117.870 1408.880 2118.190 ;
        RECT 1408.680 2114.645 1408.820 2117.870 ;
        RECT 1408.610 2114.275 1408.890 2114.645 ;
        RECT 1408.620 2104.445 1408.880 2104.590 ;
        RECT 1408.610 2104.075 1408.890 2104.445 ;
        RECT 1408.620 2097.130 1408.880 2097.450 ;
        RECT 1408.680 2094.245 1408.820 2097.130 ;
        RECT 1408.610 2093.875 1408.890 2094.245 ;
        RECT 1408.620 2090.330 1408.880 2090.650 ;
        RECT 1408.680 2084.045 1408.820 2090.330 ;
        RECT 1408.610 2083.675 1408.890 2084.045 ;
        RECT 1408.620 2076.730 1408.880 2077.050 ;
        RECT 1408.680 2073.845 1408.820 2076.730 ;
        RECT 1408.610 2073.475 1408.890 2073.845 ;
        RECT 1408.620 2069.590 1408.880 2069.910 ;
        RECT 1408.680 2063.645 1408.820 2069.590 ;
        RECT 1408.610 2063.275 1408.890 2063.645 ;
        RECT 1408.160 2061.770 1408.420 2062.090 ;
        RECT 1407.700 2061.430 1407.960 2061.750 ;
        RECT 1407.760 2021.370 1407.900 2061.430 ;
        RECT 1408.220 2022.050 1408.360 2061.770 ;
        RECT 1408.620 2056.670 1408.880 2056.990 ;
        RECT 1408.680 2022.845 1408.820 2056.670 ;
        RECT 1409.140 2043.245 1409.280 2791.410 ;
        RECT 1409.070 2042.875 1409.350 2043.245 ;
        RECT 1409.600 2033.045 1409.740 2792.090 ;
        RECT 1410.000 2791.750 1410.260 2792.070 ;
        RECT 1410.060 2056.990 1410.200 2791.750 ;
        RECT 1410.000 2056.670 1410.260 2056.990 ;
        RECT 1410.000 2055.990 1410.260 2056.310 ;
        RECT 1410.060 2053.445 1410.200 2055.990 ;
        RECT 1409.990 2053.075 1410.270 2053.445 ;
        RECT 1410.000 2052.590 1410.260 2052.910 ;
        RECT 1409.530 2032.675 1409.810 2033.045 ;
        RECT 1408.610 2022.475 1408.890 2022.845 ;
        RECT 1408.220 2021.910 1408.820 2022.050 ;
        RECT 1407.760 2021.230 1408.360 2021.370 ;
        RECT 1407.700 2020.630 1407.960 2020.950 ;
        RECT 1407.760 2012.645 1407.900 2020.630 ;
        RECT 1407.690 2012.275 1407.970 2012.645 ;
        RECT 1408.220 2002.445 1408.360 2021.230 ;
        RECT 1408.150 2002.075 1408.430 2002.445 ;
        RECT 1408.680 1992.245 1408.820 2021.910 ;
        RECT 1410.060 2020.950 1410.200 2052.590 ;
        RECT 1410.000 2020.630 1410.260 2020.950 ;
        RECT 1408.610 1991.875 1408.890 1992.245 ;
        RECT 1407.700 1985.270 1407.960 1985.590 ;
        RECT 1407.760 1982.045 1407.900 1985.270 ;
        RECT 1407.690 1981.675 1407.970 1982.045 ;
        RECT 1410.520 1971.845 1410.660 2794.130 ;
        RECT 1410.450 1971.475 1410.730 1971.845 ;
        RECT 1409.540 1890.245 1409.800 1890.390 ;
        RECT 1409.530 1889.875 1409.810 1890.245 ;
        RECT 1408.620 1829.045 1408.880 1829.190 ;
        RECT 1408.610 1828.675 1408.890 1829.045 ;
        RECT 1409.540 1814.250 1409.800 1814.570 ;
        RECT 1409.600 1808.645 1409.740 1814.250 ;
        RECT 1409.530 1808.275 1409.810 1808.645 ;
        RECT 1409.540 1800.650 1409.800 1800.970 ;
        RECT 1409.600 1798.445 1409.740 1800.650 ;
        RECT 1409.530 1798.075 1409.810 1798.445 ;
        RECT 1408.620 1788.245 1408.880 1788.390 ;
        RECT 1408.610 1787.875 1408.890 1788.245 ;
        RECT 1410.460 1779.230 1410.720 1779.550 ;
        RECT 1410.520 1778.045 1410.660 1779.230 ;
        RECT 1410.450 1777.675 1410.730 1778.045 ;
        RECT 1407.700 1730.270 1407.960 1730.590 ;
        RECT 1407.760 1727.045 1407.900 1730.270 ;
        RECT 1407.690 1726.675 1407.970 1727.045 ;
        RECT 1407.700 1706.645 1407.960 1706.790 ;
        RECT 1407.690 1706.275 1407.970 1706.645 ;
        RECT 1408.620 1696.445 1408.880 1696.590 ;
        RECT 1408.610 1696.075 1408.890 1696.445 ;
        RECT 1407.700 1687.770 1407.960 1688.090 ;
        RECT 1407.760 1686.245 1407.900 1687.770 ;
        RECT 1407.690 1685.875 1407.970 1686.245 ;
        RECT 1408.160 1676.045 1408.420 1676.190 ;
        RECT 1408.150 1675.675 1408.430 1676.045 ;
        RECT 1407.700 1666.010 1407.960 1666.330 ;
        RECT 1407.760 1665.845 1407.900 1666.010 ;
        RECT 1407.690 1665.475 1407.970 1665.845 ;
        RECT 1407.700 1655.645 1407.960 1655.790 ;
        RECT 1407.690 1655.275 1407.970 1655.645 ;
        RECT 1407.700 1645.445 1407.960 1645.590 ;
        RECT 1407.690 1645.075 1407.970 1645.445 ;
        RECT 1407.700 1635.245 1407.960 1635.390 ;
        RECT 1407.690 1634.875 1407.970 1635.245 ;
        RECT 1407.700 1625.210 1407.960 1625.530 ;
        RECT 1407.760 1625.045 1407.900 1625.210 ;
        RECT 1407.690 1624.675 1407.970 1625.045 ;
        RECT 1410.980 1605.325 1411.120 2894.430 ;
        RECT 1419.660 2794.130 1419.920 2794.450 ;
        RECT 1417.820 2790.730 1418.080 2791.050 ;
        RECT 1418.270 2790.875 1418.550 2791.245 ;
        RECT 1411.380 2789.710 1411.640 2790.030 ;
        RECT 1411.440 1900.445 1411.580 2789.710 ;
        RECT 1411.840 2789.370 1412.100 2789.690 ;
        RECT 1411.900 1910.645 1412.040 2789.370 ;
        RECT 1412.300 2789.030 1412.560 2789.350 ;
        RECT 1412.360 1920.845 1412.500 2789.030 ;
        RECT 1412.760 2788.690 1413.020 2789.010 ;
        RECT 1412.820 1931.045 1412.960 2788.690 ;
        RECT 1413.220 2788.350 1413.480 2788.670 ;
        RECT 1413.280 1941.245 1413.420 2788.350 ;
        RECT 1413.680 2788.010 1413.940 2788.330 ;
        RECT 1413.740 1951.445 1413.880 2788.010 ;
        RECT 1414.140 2787.670 1414.400 2787.990 ;
        RECT 1414.200 1961.645 1414.340 2787.670 ;
        RECT 1417.360 2787.330 1417.620 2787.650 ;
        RECT 1415.520 2060.750 1415.780 2061.070 ;
        RECT 1415.060 2060.410 1415.320 2060.730 ;
        RECT 1414.600 2052.590 1414.860 2052.910 ;
        RECT 1414.130 1961.275 1414.410 1961.645 ;
        RECT 1413.670 1951.075 1413.950 1951.445 ;
        RECT 1413.210 1940.875 1413.490 1941.245 ;
        RECT 1412.750 1930.675 1413.030 1931.045 ;
        RECT 1412.290 1920.475 1412.570 1920.845 ;
        RECT 1411.830 1910.275 1412.110 1910.645 ;
        RECT 1411.370 1900.075 1411.650 1900.445 ;
        RECT 1414.140 1883.270 1414.400 1883.590 ;
        RECT 1414.200 1880.045 1414.340 1883.270 ;
        RECT 1414.130 1879.675 1414.410 1880.045 ;
        RECT 1414.140 1869.845 1414.400 1869.990 ;
        RECT 1414.130 1869.475 1414.410 1869.845 ;
        RECT 1414.140 1862.530 1414.400 1862.850 ;
        RECT 1414.200 1859.645 1414.340 1862.530 ;
        RECT 1414.130 1859.275 1414.410 1859.645 ;
        RECT 1411.840 1855.050 1412.100 1855.370 ;
        RECT 1411.900 1849.445 1412.040 1855.050 ;
        RECT 1411.830 1849.075 1412.110 1849.445 ;
        RECT 1411.380 1840.090 1411.640 1840.410 ;
        RECT 1411.440 1839.245 1411.580 1840.090 ;
        RECT 1411.370 1838.875 1411.650 1839.245 ;
        RECT 1414.140 1821.390 1414.400 1821.710 ;
        RECT 1414.200 1818.845 1414.340 1821.390 ;
        RECT 1414.130 1818.475 1414.410 1818.845 ;
        RECT 1414.130 1767.730 1414.410 1767.845 ;
        RECT 1414.660 1767.730 1414.800 2052.590 ;
        RECT 1414.130 1767.590 1414.800 1767.730 ;
        RECT 1414.130 1767.475 1414.410 1767.590 ;
        RECT 1414.130 1757.530 1414.410 1757.645 ;
        RECT 1415.120 1757.530 1415.260 2060.410 ;
        RECT 1414.130 1757.390 1415.260 1757.530 ;
        RECT 1414.130 1757.275 1414.410 1757.390 ;
        RECT 1414.130 1747.330 1414.410 1747.445 ;
        RECT 1415.580 1747.330 1415.720 2060.750 ;
        RECT 1415.980 2060.070 1416.240 2060.390 ;
        RECT 1414.130 1747.190 1415.720 1747.330 ;
        RECT 1414.130 1747.075 1414.410 1747.190 ;
        RECT 1414.130 1738.490 1414.410 1738.605 ;
        RECT 1416.040 1738.490 1416.180 2060.070 ;
        RECT 1416.440 2059.730 1416.700 2060.050 ;
        RECT 1414.130 1738.350 1416.180 1738.490 ;
        RECT 1414.130 1738.235 1414.410 1738.350 ;
        RECT 1416.500 1730.590 1416.640 2059.730 ;
        RECT 1416.900 2052.930 1417.160 2053.250 ;
        RECT 1416.440 1730.270 1416.700 1730.590 ;
        RECT 1414.140 1717.690 1414.400 1718.010 ;
        RECT 1414.200 1716.845 1414.340 1717.690 ;
        RECT 1414.130 1716.475 1414.410 1716.845 ;
        RECT 1416.960 1706.790 1417.100 2052.930 ;
        RECT 1417.420 1985.590 1417.560 2787.330 ;
        RECT 1417.360 1985.270 1417.620 1985.590 ;
        RECT 1416.900 1706.470 1417.160 1706.790 ;
        RECT 1417.880 1625.530 1418.020 2790.730 ;
        RECT 1418.340 1635.390 1418.480 2790.875 ;
        RECT 1418.740 2790.390 1419.000 2790.710 ;
        RECT 1418.800 1645.590 1418.940 2790.390 ;
        RECT 1419.200 2790.050 1419.460 2790.370 ;
        RECT 1419.260 1655.790 1419.400 2790.050 ;
        RECT 1419.720 1666.330 1419.860 2794.130 ;
        RECT 1421.040 2793.790 1421.300 2794.110 ;
        RECT 1420.580 2793.450 1420.840 2793.770 ;
        RECT 1420.120 2792.430 1420.380 2792.750 ;
        RECT 1420.180 1676.190 1420.320 2792.430 ;
        RECT 1420.640 1688.090 1420.780 2793.450 ;
        RECT 1421.100 1696.590 1421.240 2793.790 ;
        RECT 1424.780 1829.190 1424.920 3194.650 ;
        RECT 1426.560 2062.110 1426.820 2062.430 ;
        RECT 1426.100 2053.950 1426.360 2054.270 ;
        RECT 1425.640 2053.610 1425.900 2053.930 ;
        RECT 1425.180 2053.270 1425.440 2053.590 ;
        RECT 1424.720 1828.870 1424.980 1829.190 ;
        RECT 1425.240 1779.550 1425.380 2053.270 ;
        RECT 1425.700 1788.390 1425.840 2053.610 ;
        RECT 1426.160 1800.970 1426.300 2053.950 ;
        RECT 1426.620 1814.570 1426.760 2062.110 ;
        RECT 1427.020 2059.390 1427.280 2059.710 ;
        RECT 1427.080 1890.390 1427.220 2059.390 ;
        RECT 1427.020 1890.070 1427.280 1890.390 ;
        RECT 1431.680 1840.410 1431.820 3201.450 ;
        RECT 1438.580 1855.370 1438.720 3208.590 ;
        RECT 1452.380 1862.850 1452.520 3215.390 ;
        RECT 1459.280 1869.990 1459.420 3222.190 ;
        RECT 1473.020 3187.850 1473.280 3188.170 ;
        RECT 1462.890 2792.915 1463.170 2793.285 ;
        RECT 1462.900 2792.770 1463.160 2792.915 ;
        RECT 1459.220 1869.670 1459.480 1869.990 ;
        RECT 1452.320 1862.530 1452.580 1862.850 ;
        RECT 1438.520 1855.050 1438.780 1855.370 ;
        RECT 1431.620 1840.090 1431.880 1840.410 ;
        RECT 1473.080 1821.710 1473.220 3187.850 ;
        RECT 1473.540 1883.590 1473.680 3229.330 ;
        RECT 1535.570 3224.715 1535.850 3225.085 ;
        RECT 1535.640 3222.510 1535.780 3224.715 ;
        RECT 1535.580 3222.190 1535.840 3222.510 ;
        RECT 1535.570 3217.235 1535.850 3217.605 ;
        RECT 1535.640 3215.710 1535.780 3217.235 ;
        RECT 1535.580 3215.390 1535.840 3215.710 ;
        RECT 1538.330 3210.435 1538.610 3210.805 ;
        RECT 1538.400 3208.910 1538.540 3210.435 ;
        RECT 1538.340 3208.590 1538.600 3208.910 ;
        RECT 1538.330 3202.275 1538.610 3202.645 ;
        RECT 1538.400 3201.770 1538.540 3202.275 ;
        RECT 1538.340 3201.450 1538.600 3201.770 ;
        RECT 1533.270 3196.835 1533.550 3197.205 ;
        RECT 1533.340 3194.970 1533.480 3196.835 ;
        RECT 1533.280 3194.650 1533.540 3194.970 ;
        RECT 1534.190 3189.355 1534.470 3189.725 ;
        RECT 1534.260 3188.170 1534.400 3189.355 ;
        RECT 1534.200 3187.850 1534.460 3188.170 ;
        RECT 1534.650 2899.675 1534.930 2900.045 ;
        RECT 1534.720 2898.490 1534.860 2899.675 ;
        RECT 1514.420 2898.170 1514.680 2898.490 ;
        RECT 1534.660 2898.170 1534.920 2898.490 ;
        RECT 1510.730 2792.915 1511.010 2793.285 ;
        RECT 1510.800 2792.750 1510.940 2792.915 ;
        RECT 1510.740 2792.430 1511.000 2792.750 ;
        RECT 1473.480 1883.270 1473.740 1883.590 ;
        RECT 1473.020 1821.390 1473.280 1821.710 ;
        RECT 1426.560 1814.250 1426.820 1814.570 ;
        RECT 1426.100 1800.650 1426.360 1800.970 ;
        RECT 1425.640 1788.070 1425.900 1788.390 ;
        RECT 1425.180 1779.230 1425.440 1779.550 ;
        RECT 1514.480 1718.010 1514.620 2898.170 ;
        RECT 1538.340 2894.605 1538.600 2894.750 ;
        RECT 1538.330 2894.235 1538.610 2894.605 ;
      LAYER met2 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met2 ;
        RECT 1935.780 3251.090 1936.040 3251.410 ;
        RECT 1935.840 3249.565 1935.980 3251.090 ;
        RECT 1935.770 3249.195 1936.050 3249.565 ;
        RECT 2190.610 3230.155 2190.890 3230.525 ;
        RECT 1945.890 2904.435 1946.170 2904.805 ;
        RECT 1945.960 2901.550 1946.100 2904.435 ;
        RECT 1945.900 2901.230 1946.160 2901.550 ;
        RECT 2189.240 2901.230 2189.500 2901.550 ;
        RECT 2189.300 2895.965 2189.440 2901.230 ;
        RECT 2189.230 2895.595 2189.510 2895.965 ;
        RECT 1742.110 2796.315 1742.390 2796.685 ;
        RECT 1788.570 2796.315 1788.850 2796.685 ;
        RECT 1580.190 2794.275 1580.470 2794.645 ;
        RECT 1587.090 2794.275 1587.370 2794.645 ;
        RECT 1601.350 2794.275 1601.630 2794.645 ;
        RECT 1614.230 2794.275 1614.510 2794.645 ;
        RECT 1617.450 2794.275 1617.730 2794.645 ;
        RECT 1580.260 2062.430 1580.400 2794.275 ;
        RECT 1587.100 2794.130 1587.360 2794.275 ;
        RECT 1601.420 2794.110 1601.560 2794.275 ;
        RECT 1600.890 2793.595 1601.170 2793.965 ;
        RECT 1601.360 2793.790 1601.620 2794.110 ;
        RECT 1600.900 2793.450 1601.160 2793.595 ;
        RECT 1614.300 2793.430 1614.440 2794.275 ;
        RECT 1593.990 2792.915 1594.270 2793.285 ;
        RECT 1614.240 2793.110 1614.500 2793.430 ;
        RECT 1594.060 2792.750 1594.200 2792.915 ;
        RECT 1594.000 2792.430 1594.260 2792.750 ;
        RECT 1614.300 2791.390 1614.440 2793.110 ;
        RECT 1617.520 2793.090 1617.660 2794.275 ;
        RECT 1631.720 2794.130 1631.980 2794.450 ;
        RECT 1642.750 2794.275 1643.030 2794.645 ;
        RECT 1647.810 2794.275 1648.090 2794.645 ;
        RECT 1652.410 2794.275 1652.690 2794.645 ;
        RECT 1662.530 2794.275 1662.810 2794.645 ;
        RECT 1665.750 2794.275 1666.030 2794.645 ;
        RECT 1671.270 2794.275 1671.550 2794.645 ;
        RECT 1679.550 2794.275 1679.830 2794.645 ;
        RECT 1681.390 2794.275 1681.670 2794.645 ;
        RECT 1688.750 2794.275 1689.030 2794.645 ;
        RECT 1695.190 2794.275 1695.470 2794.645 ;
        RECT 1699.330 2794.275 1699.610 2794.645 ;
        RECT 1706.230 2794.275 1706.510 2794.645 ;
        RECT 1712.670 2794.275 1712.950 2794.645 ;
        RECT 1718.190 2794.275 1718.470 2794.645 ;
        RECT 1624.820 2793.450 1625.080 2793.770 ;
        RECT 1617.460 2792.770 1617.720 2793.090 ;
        RECT 1614.240 2791.070 1614.500 2791.390 ;
        RECT 1624.880 2788.525 1625.020 2793.450 ;
        RECT 1631.780 2788.525 1631.920 2794.130 ;
        RECT 1638.620 2793.110 1638.880 2793.430 ;
        RECT 1638.680 2788.525 1638.820 2793.110 ;
        RECT 1642.820 2792.070 1642.960 2794.275 ;
        RECT 1647.880 2792.410 1648.020 2794.275 ;
        RECT 1647.820 2792.090 1648.080 2792.410 ;
        RECT 1642.760 2791.750 1643.020 2792.070 ;
        RECT 1652.480 2791.730 1652.620 2794.275 ;
        RECT 1662.600 2794.110 1662.740 2794.275 ;
        RECT 1662.540 2793.790 1662.800 2794.110 ;
        RECT 1652.420 2791.410 1652.680 2791.730 ;
        RECT 1662.600 2791.390 1662.740 2793.790 ;
        RECT 1665.820 2793.090 1665.960 2794.275 ;
        RECT 1671.280 2794.130 1671.540 2794.275 ;
        RECT 1671.340 2793.770 1671.480 2794.130 ;
        RECT 1671.280 2793.450 1671.540 2793.770 ;
        RECT 1679.620 2793.430 1679.760 2794.275 ;
        RECT 1681.460 2793.770 1681.600 2794.275 ;
        RECT 1681.400 2793.450 1681.660 2793.770 ;
        RECT 1679.560 2793.110 1679.820 2793.430 ;
        RECT 1681.460 2793.090 1681.600 2793.450 ;
        RECT 1688.820 2793.090 1688.960 2794.275 ;
        RECT 1665.760 2792.770 1666.020 2793.090 ;
        RECT 1669.440 2792.770 1669.700 2793.090 ;
        RECT 1681.400 2792.770 1681.660 2793.090 ;
        RECT 1683.700 2792.770 1683.960 2793.090 ;
        RECT 1688.760 2792.770 1689.020 2793.090 ;
        RECT 1669.500 2791.730 1669.640 2792.770 ;
        RECT 1683.760 2792.070 1683.900 2792.770 ;
        RECT 1695.260 2792.410 1695.400 2794.275 ;
        RECT 1695.200 2792.090 1695.460 2792.410 ;
        RECT 1683.700 2791.750 1683.960 2792.070 ;
        RECT 1669.440 2791.410 1669.700 2791.730 ;
        RECT 1699.400 2791.390 1699.540 2794.275 ;
        RECT 1706.300 2794.110 1706.440 2794.275 ;
        RECT 1706.240 2793.790 1706.500 2794.110 ;
        RECT 1712.740 2791.730 1712.880 2794.275 ;
        RECT 1718.200 2794.130 1718.460 2794.275 ;
        RECT 1723.720 2794.130 1723.980 2794.450 ;
        RECT 1724.170 2794.275 1724.450 2794.645 ;
        RECT 1728.770 2794.275 1729.050 2794.645 ;
        RECT 1732.450 2794.275 1732.730 2794.645 ;
        RECT 1741.190 2794.275 1741.470 2794.645 ;
        RECT 1724.180 2794.130 1724.440 2794.275 ;
        RECT 1712.680 2791.410 1712.940 2791.730 ;
        RECT 1723.780 2791.390 1723.920 2794.130 ;
        RECT 1724.240 2793.430 1724.380 2794.130 ;
        RECT 1728.840 2793.770 1728.980 2794.275 ;
        RECT 1728.780 2793.450 1729.040 2793.770 ;
        RECT 1732.520 2793.430 1732.660 2794.275 ;
        RECT 1724.180 2793.110 1724.440 2793.430 ;
        RECT 1732.460 2793.110 1732.720 2793.430 ;
        RECT 1732.520 2792.410 1732.660 2793.110 ;
        RECT 1741.260 2792.410 1741.400 2794.275 ;
        RECT 1732.460 2792.090 1732.720 2792.410 ;
        RECT 1741.200 2792.090 1741.460 2792.410 ;
        RECT 1742.180 2792.070 1742.320 2796.315 ;
        RECT 1746.710 2794.275 1746.990 2794.645 ;
        RECT 1752.690 2794.275 1752.970 2794.645 ;
        RECT 1760.050 2794.275 1760.330 2794.645 ;
        RECT 1766.490 2794.275 1766.770 2794.645 ;
        RECT 1746.780 2793.770 1746.920 2794.275 ;
        RECT 1752.760 2794.110 1752.900 2794.275 ;
        RECT 1752.700 2793.790 1752.960 2794.110 ;
        RECT 1746.720 2793.450 1746.980 2793.770 ;
        RECT 1742.120 2791.750 1742.380 2792.070 ;
        RECT 1746.780 2791.730 1746.920 2793.450 ;
        RECT 1746.720 2791.410 1746.980 2791.730 ;
        RECT 1760.120 2791.390 1760.260 2794.275 ;
        RECT 1766.500 2794.130 1766.760 2794.275 ;
        RECT 1773.390 2793.595 1773.670 2793.965 ;
        RECT 1780.290 2793.595 1780.570 2793.965 ;
        RECT 1773.460 2793.090 1773.600 2793.595 ;
        RECT 1780.360 2793.430 1780.500 2793.595 ;
        RECT 1780.300 2793.110 1780.560 2793.430 ;
        RECT 1773.400 2792.770 1773.660 2793.090 ;
        RECT 1787.190 2792.235 1787.470 2792.605 ;
        RECT 1787.200 2792.090 1787.460 2792.235 ;
        RECT 1783.510 2791.555 1783.790 2791.925 ;
        RECT 1788.640 2791.730 1788.780 2796.315 ;
        RECT 2091.260 2793.110 2091.520 2793.430 ;
        RECT 1790.420 2792.090 1790.680 2792.410 ;
        RECT 1662.540 2791.070 1662.800 2791.390 ;
        RECT 1699.340 2791.070 1699.600 2791.390 ;
        RECT 1723.720 2791.070 1723.980 2791.390 ;
        RECT 1760.060 2791.070 1760.320 2791.390 ;
        RECT 1624.810 2788.155 1625.090 2788.525 ;
        RECT 1631.710 2788.155 1631.990 2788.525 ;
        RECT 1638.610 2788.155 1638.890 2788.525 ;
        RECT 1649.650 2788.155 1649.930 2788.525 ;
        RECT 1684.150 2788.155 1684.430 2788.525 ;
        RECT 1718.650 2788.155 1718.930 2788.525 ;
        RECT 1760.050 2788.155 1760.330 2788.525 ;
        RECT 1607.790 2787.475 1608.070 2787.845 ;
        RECT 1614.690 2787.475 1614.970 2787.845 ;
        RECT 1621.590 2787.475 1621.870 2787.845 ;
        RECT 1580.200 2062.110 1580.460 2062.430 ;
        RECT 1607.860 2056.310 1608.000 2787.475 ;
        RECT 1614.760 2069.910 1614.900 2787.475 ;
        RECT 1621.660 2077.050 1621.800 2787.475 ;
        RECT 1621.600 2076.730 1621.860 2077.050 ;
        RECT 1614.700 2069.590 1614.960 2069.910 ;
        RECT 1624.880 2062.090 1625.020 2788.155 ;
        RECT 1628.490 2787.475 1628.770 2787.845 ;
        RECT 1628.560 2090.650 1628.700 2787.475 ;
        RECT 1628.500 2090.330 1628.760 2090.650 ;
        RECT 1624.820 2061.770 1625.080 2062.090 ;
        RECT 1631.780 2061.750 1631.920 2788.155 ;
        RECT 1635.390 2787.475 1635.670 2787.845 ;
        RECT 1635.460 2097.450 1635.600 2787.475 ;
        RECT 1635.400 2097.130 1635.660 2097.450 ;
        RECT 1631.720 2061.430 1631.980 2061.750 ;
        RECT 1638.680 2061.410 1638.820 2788.155 ;
        RECT 1642.290 2787.475 1642.570 2787.845 ;
        RECT 1649.190 2787.475 1649.470 2787.845 ;
        RECT 1642.360 2104.590 1642.500 2787.475 ;
        RECT 1649.260 2118.190 1649.400 2787.475 ;
        RECT 1649.720 2125.330 1649.860 2788.155 ;
        RECT 1656.090 2787.475 1656.370 2787.845 ;
        RECT 1662.990 2787.475 1663.270 2787.845 ;
        RECT 1669.890 2787.475 1670.170 2787.845 ;
        RECT 1676.790 2787.475 1677.070 2787.845 ;
        RECT 1683.690 2787.475 1683.970 2787.845 ;
        RECT 1656.160 2138.930 1656.300 2787.475 ;
        RECT 1663.060 2145.730 1663.200 2787.475 ;
        RECT 1669.960 2159.670 1670.100 2787.475 ;
        RECT 1676.860 2166.470 1677.000 2787.475 ;
        RECT 1683.760 2180.410 1683.900 2787.475 ;
        RECT 1684.220 2187.210 1684.360 2788.155 ;
        RECT 1690.590 2787.475 1690.870 2787.845 ;
        RECT 1697.490 2787.475 1697.770 2787.845 ;
        RECT 1704.390 2787.475 1704.670 2787.845 ;
        RECT 1711.290 2787.475 1711.570 2787.845 ;
        RECT 1718.190 2787.475 1718.470 2787.845 ;
        RECT 1690.660 2201.150 1690.800 2787.475 ;
        RECT 1697.560 2207.950 1697.700 2787.475 ;
        RECT 1704.460 2221.890 1704.600 2787.475 ;
        RECT 1711.360 2228.690 1711.500 2787.475 ;
        RECT 1718.260 2242.630 1718.400 2787.475 ;
        RECT 1718.720 2249.430 1718.860 2788.155 ;
        RECT 1725.090 2787.475 1725.370 2787.845 ;
        RECT 1731.990 2787.475 1732.270 2787.845 ;
        RECT 1738.890 2787.475 1739.170 2787.845 ;
        RECT 1745.790 2787.475 1746.070 2787.845 ;
        RECT 1752.690 2787.475 1752.970 2787.845 ;
        RECT 1725.160 2263.030 1725.300 2787.475 ;
        RECT 1732.060 2270.170 1732.200 2787.475 ;
        RECT 1738.960 2276.970 1739.100 2787.475 ;
        RECT 1745.860 2290.910 1746.000 2787.475 ;
        RECT 1752.760 2297.710 1752.900 2787.475 ;
        RECT 1760.120 2318.450 1760.260 2788.155 ;
        RECT 1766.490 2787.475 1766.770 2787.845 ;
        RECT 1773.390 2787.475 1773.670 2787.845 ;
        RECT 1780.290 2787.475 1780.570 2787.845 ;
        RECT 1760.970 2777.275 1761.250 2777.645 ;
        RECT 1760.060 2318.130 1760.320 2318.450 ;
        RECT 1761.040 2311.650 1761.180 2777.275 ;
        RECT 1766.560 2332.050 1766.700 2787.475 ;
        RECT 1773.460 2339.190 1773.600 2787.475 ;
        RECT 1780.360 2352.790 1780.500 2787.475 ;
        RECT 1783.580 2573.790 1783.720 2791.555 ;
        RECT 1788.580 2791.410 1788.840 2791.730 ;
        RECT 1787.650 2787.475 1787.930 2787.845 ;
        RECT 1783.520 2573.470 1783.780 2573.790 ;
        RECT 1787.720 2359.930 1787.860 2787.475 ;
        RECT 1790.480 2394.270 1790.620 2792.090 ;
        RECT 1797.320 2791.750 1797.580 2792.070 ;
        RECT 1790.880 2791.070 1791.140 2791.390 ;
        RECT 1790.940 2587.390 1791.080 2791.070 ;
        RECT 1794.550 2777.275 1794.830 2777.645 ;
        RECT 1790.880 2587.070 1791.140 2587.390 ;
        RECT 1790.420 2393.950 1790.680 2394.270 ;
        RECT 1794.620 2373.530 1794.760 2777.275 ;
        RECT 1797.380 2594.530 1797.520 2791.750 ;
        RECT 1797.780 2791.410 1798.040 2791.730 ;
        RECT 1797.840 2608.130 1797.980 2791.410 ;
        RECT 2091.320 2790.710 2091.460 2793.110 ;
        RECT 2091.260 2790.390 2091.520 2790.710 ;
        RECT 2090.800 2790.050 2091.060 2790.370 ;
        RECT 2163.020 2790.050 2163.280 2790.370 ;
        RECT 2090.860 2789.770 2091.000 2790.050 ;
        RECT 2090.860 2789.630 2091.920 2789.770 ;
        RECT 2091.780 2787.990 2091.920 2789.630 ;
        RECT 2163.080 2788.410 2163.220 2790.050 ;
        RECT 2162.620 2788.270 2163.220 2788.410 ;
        RECT 2162.620 2787.990 2162.760 2788.270 ;
        RECT 2091.720 2787.670 2091.980 2787.990 ;
        RECT 2162.560 2787.670 2162.820 2787.990 ;
        RECT 1797.780 2607.810 1798.040 2608.130 ;
        RECT 1797.320 2594.210 1797.580 2594.530 ;
        RECT 1794.560 2373.210 1794.820 2373.530 ;
        RECT 1787.660 2359.610 1787.920 2359.930 ;
        RECT 1780.300 2352.470 1780.560 2352.790 ;
        RECT 1773.400 2338.870 1773.660 2339.190 ;
        RECT 1766.500 2331.730 1766.760 2332.050 ;
        RECT 1760.980 2311.330 1761.240 2311.650 ;
        RECT 1752.700 2297.390 1752.960 2297.710 ;
        RECT 1745.800 2290.590 1746.060 2290.910 ;
        RECT 1738.900 2276.650 1739.160 2276.970 ;
        RECT 1732.000 2269.850 1732.260 2270.170 ;
        RECT 1725.100 2262.710 1725.360 2263.030 ;
        RECT 1718.660 2249.110 1718.920 2249.430 ;
        RECT 1718.200 2242.310 1718.460 2242.630 ;
        RECT 1711.300 2228.370 1711.560 2228.690 ;
        RECT 1704.400 2221.570 1704.660 2221.890 ;
        RECT 1697.500 2207.630 1697.760 2207.950 ;
        RECT 1690.600 2200.830 1690.860 2201.150 ;
        RECT 1684.160 2186.890 1684.420 2187.210 ;
        RECT 1683.700 2180.090 1683.960 2180.410 ;
        RECT 1676.800 2166.150 1677.060 2166.470 ;
        RECT 1669.900 2159.350 1670.160 2159.670 ;
        RECT 1663.000 2145.410 1663.260 2145.730 ;
        RECT 1656.100 2138.610 1656.360 2138.930 ;
        RECT 1649.660 2125.010 1649.920 2125.330 ;
        RECT 1649.200 2117.870 1649.460 2118.190 ;
        RECT 1642.300 2104.270 1642.560 2104.590 ;
        RECT 1638.620 2061.090 1638.880 2061.410 ;
        RECT 1607.800 2055.990 1608.060 2056.310 ;
        RECT 2190.680 2054.270 2190.820 3230.155 ;
        RECT 2191.070 3224.715 2191.350 3225.085 ;
        RECT 2190.620 2053.950 2190.880 2054.270 ;
        RECT 2191.140 2053.930 2191.280 3224.715 ;
        RECT 2191.530 3215.875 2191.810 3216.245 ;
        RECT 2191.080 2053.610 2191.340 2053.930 ;
        RECT 2191.600 2053.590 2191.740 3215.875 ;
        RECT 2191.990 3209.755 2192.270 3210.125 ;
        RECT 2191.540 2053.270 2191.800 2053.590 ;
        RECT 2192.060 2052.910 2192.200 3209.755 ;
        RECT 2192.450 3201.595 2192.730 3201.965 ;
        RECT 2192.520 2060.730 2192.660 3201.595 ;
        RECT 2192.910 3196.155 2193.190 3196.525 ;
        RECT 2192.980 2061.070 2193.120 3196.155 ;
        RECT 2193.370 3187.995 2193.650 3188.365 ;
        RECT 2192.920 2060.750 2193.180 2061.070 ;
        RECT 2192.460 2060.410 2192.720 2060.730 ;
        RECT 2193.440 2060.390 2193.580 3187.995 ;
        RECT 2193.830 2898.315 2194.110 2898.685 ;
        RECT 2193.380 2060.070 2193.640 2060.390 ;
        RECT 2193.900 2053.250 2194.040 2898.315 ;
      LAYER met2 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met2 ;
        RECT 2582.140 3249.565 2582.280 3252.110 ;
        RECT 2582.070 3249.195 2582.350 3249.565 ;
        RECT 2594.560 2946.965 2594.700 3263.670 ;
        RECT 2594.490 2946.595 2594.770 2946.965 ;
        RECT 2594.560 2938.805 2594.700 2946.595 ;
        RECT 2594.490 2938.435 2594.770 2938.805 ;
        RECT 2228.790 2794.275 2229.070 2794.645 ;
        RECT 2208.100 2793.790 2208.360 2794.110 ;
        RECT 2208.160 2787.990 2208.300 2793.790 ;
        RECT 2218.220 2789.710 2218.480 2790.030 ;
        RECT 2208.100 2787.670 2208.360 2787.990 ;
        RECT 2218.280 2614.930 2218.420 2789.710 ;
        RECT 2218.220 2614.610 2218.480 2614.930 ;
        RECT 2228.860 2060.050 2229.000 2794.275 ;
        RECT 2232.020 2794.130 2232.280 2794.450 ;
        RECT 2237.990 2794.275 2238.270 2794.645 ;
        RECT 2268.350 2794.275 2268.630 2794.645 ;
        RECT 2273.410 2794.275 2273.690 2794.645 ;
        RECT 2279.850 2794.275 2280.130 2794.645 ;
        RECT 2286.750 2794.275 2287.030 2794.645 ;
        RECT 2291.350 2794.275 2291.630 2794.645 ;
        RECT 2304.230 2794.275 2304.510 2794.645 ;
        RECT 2308.370 2794.275 2308.650 2794.645 ;
        RECT 2312.970 2794.275 2313.250 2794.645 ;
        RECT 2321.250 2794.275 2321.530 2794.645 ;
        RECT 2326.310 2794.275 2326.590 2794.645 ;
        RECT 2332.290 2794.275 2332.570 2794.645 ;
        RECT 2339.190 2794.275 2339.470 2794.645 ;
        RECT 2343.330 2794.275 2343.610 2794.645 ;
        RECT 2346.090 2794.275 2346.370 2794.645 ;
        RECT 2352.990 2794.275 2353.270 2794.645 ;
        RECT 2359.890 2794.275 2360.170 2794.645 ;
        RECT 2366.790 2794.275 2367.070 2794.645 ;
        RECT 2374.150 2794.275 2374.430 2794.645 ;
        RECT 2377.370 2794.275 2377.650 2794.645 ;
        RECT 2385.650 2794.275 2385.930 2794.645 ;
        RECT 2391.170 2794.275 2391.450 2794.645 ;
        RECT 2394.850 2794.275 2395.130 2794.645 ;
        RECT 2402.670 2794.275 2402.950 2794.645 ;
        RECT 2415.090 2794.275 2415.370 2794.645 ;
        RECT 2232.080 2628.870 2232.220 2794.130 ;
        RECT 2238.060 2791.050 2238.200 2794.275 ;
        RECT 2263.290 2793.595 2263.570 2793.965 ;
        RECT 2268.420 2793.770 2268.560 2794.275 ;
        RECT 2249.490 2792.235 2249.770 2792.605 ;
        RECT 2258.700 2792.490 2258.960 2792.750 ;
        RECT 2261.920 2792.490 2262.180 2792.750 ;
        RECT 2258.700 2792.430 2262.180 2792.490 ;
        RECT 2258.760 2792.350 2262.120 2792.430 ;
        RECT 2263.360 2792.410 2263.500 2793.595 ;
        RECT 2268.360 2793.450 2268.620 2793.770 ;
        RECT 2273.480 2793.430 2273.620 2794.275 ;
        RECT 2266.510 2792.915 2266.790 2793.285 ;
        RECT 2269.730 2792.915 2270.010 2793.285 ;
        RECT 2270.200 2793.110 2270.460 2793.430 ;
        RECT 2273.420 2793.110 2273.680 2793.430 ;
        RECT 2238.000 2790.730 2238.260 2791.050 ;
        RECT 2249.560 2790.710 2249.700 2792.235 ;
        RECT 2263.300 2792.090 2263.560 2792.410 ;
        RECT 2249.500 2790.390 2249.760 2790.710 ;
        RECT 2256.390 2790.195 2256.670 2790.565 ;
        RECT 2256.400 2790.050 2256.660 2790.195 ;
        RECT 2245.820 2789.370 2246.080 2789.690 ;
        RECT 2238.920 2789.030 2239.180 2789.350 ;
        RECT 2238.980 2635.670 2239.120 2789.030 ;
        RECT 2245.880 2649.610 2246.020 2789.370 ;
        RECT 2259.620 2788.690 2259.880 2789.010 ;
        RECT 2252.720 2788.350 2252.980 2788.670 ;
        RECT 2252.780 2656.410 2252.920 2788.350 ;
        RECT 2259.680 2670.350 2259.820 2788.690 ;
        RECT 2263.290 2787.475 2263.570 2787.845 ;
        RECT 2259.620 2670.030 2259.880 2670.350 ;
        RECT 2252.720 2656.090 2252.980 2656.410 ;
        RECT 2245.820 2649.290 2246.080 2649.610 ;
        RECT 2238.920 2635.350 2239.180 2635.670 ;
        RECT 2232.020 2628.550 2232.280 2628.870 ;
        RECT 2263.360 2380.330 2263.500 2787.475 ;
        RECT 2263.300 2380.010 2263.560 2380.330 ;
        RECT 2228.800 2059.730 2229.060 2060.050 ;
        RECT 2266.580 2059.710 2266.720 2792.915 ;
        RECT 2269.800 2792.750 2269.940 2792.915 ;
        RECT 2269.740 2792.430 2270.000 2792.750 ;
        RECT 2267.440 2788.010 2267.700 2788.330 ;
        RECT 2266.970 2787.475 2267.250 2787.845 ;
        RECT 2267.040 2401.070 2267.180 2787.475 ;
        RECT 2267.500 2677.150 2267.640 2788.010 ;
        RECT 2270.260 2787.990 2270.400 2793.110 ;
        RECT 2279.920 2793.090 2280.060 2794.275 ;
        RECT 2286.820 2794.110 2286.960 2794.275 ;
        RECT 2286.760 2793.790 2287.020 2794.110 ;
        RECT 2279.860 2792.770 2280.120 2793.090 ;
        RECT 2291.420 2790.030 2291.560 2794.275 ;
        RECT 2298.250 2792.915 2298.530 2793.285 ;
        RECT 2297.340 2792.090 2297.600 2792.410 ;
        RECT 2297.400 2790.030 2297.540 2792.090 ;
        RECT 2291.360 2789.710 2291.620 2790.030 ;
        RECT 2297.340 2789.710 2297.600 2790.030 ;
        RECT 2273.420 2789.370 2273.680 2789.690 ;
        RECT 2270.200 2787.670 2270.460 2787.990 ;
        RECT 2273.480 2691.090 2273.620 2789.370 ;
        RECT 2298.320 2787.990 2298.460 2792.915 ;
        RECT 2304.300 2790.030 2304.440 2794.275 ;
        RECT 2308.440 2792.750 2308.580 2794.275 ;
        RECT 2313.040 2793.770 2313.180 2794.275 ;
        RECT 2312.980 2793.450 2313.240 2793.770 ;
        RECT 2314.810 2792.915 2315.090 2793.285 ;
        RECT 2314.820 2792.770 2315.080 2792.915 ;
        RECT 2308.380 2792.430 2308.640 2792.750 ;
        RECT 2304.240 2789.710 2304.500 2790.030 ;
        RECT 2305.150 2788.155 2305.430 2788.525 ;
        RECT 2277.090 2787.475 2277.370 2787.845 ;
        RECT 2283.990 2787.475 2284.270 2787.845 ;
        RECT 2290.890 2787.475 2291.170 2787.845 ;
        RECT 2297.790 2787.475 2298.070 2787.845 ;
        RECT 2298.260 2787.670 2298.520 2787.990 ;
        RECT 2304.690 2787.475 2304.970 2787.845 ;
        RECT 2273.420 2690.770 2273.680 2691.090 ;
        RECT 2267.440 2676.830 2267.700 2677.150 ;
        RECT 2277.160 2415.010 2277.300 2787.475 ;
        RECT 2284.060 2421.810 2284.200 2787.475 ;
        RECT 2290.960 2435.750 2291.100 2787.475 ;
        RECT 2297.860 2442.550 2298.000 2787.475 ;
        RECT 2304.760 2456.490 2304.900 2787.475 ;
        RECT 2305.220 2463.290 2305.360 2788.155 ;
        RECT 2321.320 2787.990 2321.460 2794.275 ;
        RECT 2326.380 2793.430 2326.520 2794.275 ;
        RECT 2326.320 2793.110 2326.580 2793.430 ;
        RECT 2321.720 2789.370 2321.980 2789.690 ;
        RECT 2311.590 2787.475 2311.870 2787.845 ;
        RECT 2318.490 2787.475 2318.770 2787.845 ;
        RECT 2321.260 2787.670 2321.520 2787.990 ;
        RECT 2311.660 2477.230 2311.800 2787.475 ;
        RECT 2318.560 2484.030 2318.700 2787.475 ;
        RECT 2321.780 2697.890 2321.920 2789.370 ;
        RECT 2325.390 2787.475 2325.670 2787.845 ;
        RECT 2321.720 2697.570 2321.980 2697.890 ;
        RECT 2325.460 2497.630 2325.600 2787.475 ;
        RECT 2332.360 2504.770 2332.500 2794.275 ;
        RECT 2332.760 2793.965 2333.020 2794.110 ;
        RECT 2332.750 2793.595 2333.030 2793.965 ;
        RECT 2339.260 2511.570 2339.400 2794.275 ;
        RECT 2339.650 2793.595 2339.930 2793.965 ;
        RECT 2339.720 2525.510 2339.860 2793.595 ;
        RECT 2340.110 2792.915 2340.390 2793.285 ;
        RECT 2343.400 2793.090 2343.540 2794.275 ;
        RECT 2340.180 2792.410 2340.320 2792.915 ;
        RECT 2343.340 2792.770 2343.600 2793.090 ;
        RECT 2340.120 2792.090 2340.380 2792.410 ;
        RECT 2343.800 2792.090 2344.060 2792.410 ;
        RECT 2343.860 2790.030 2344.000 2792.090 ;
        RECT 2343.800 2789.710 2344.060 2790.030 ;
        RECT 2346.160 2532.310 2346.300 2794.275 ;
        RECT 2350.230 2793.595 2350.510 2793.965 ;
        RECT 2350.300 2792.410 2350.440 2793.595 ;
        RECT 2350.240 2792.090 2350.500 2792.410 ;
        RECT 2353.060 2546.250 2353.200 2794.275 ;
        RECT 2356.670 2793.595 2356.950 2793.965 ;
        RECT 2356.740 2792.750 2356.880 2793.595 ;
        RECT 2356.680 2792.430 2356.940 2792.750 ;
        RECT 2359.960 2553.050 2360.100 2794.275 ;
        RECT 2360.810 2793.595 2361.090 2793.965 ;
        RECT 2360.820 2793.450 2361.080 2793.595 ;
        RECT 2366.860 2566.650 2367.000 2794.275 ;
        RECT 2374.220 2793.430 2374.360 2794.275 ;
        RECT 2377.440 2794.110 2377.580 2794.275 ;
        RECT 2377.380 2793.790 2377.640 2794.110 ;
        RECT 2367.250 2792.915 2367.530 2793.285 ;
        RECT 2374.160 2793.110 2374.420 2793.430 ;
        RECT 2377.440 2793.090 2377.580 2793.790 ;
        RECT 2367.320 2787.990 2367.460 2792.915 ;
        RECT 2377.380 2792.770 2377.640 2793.090 ;
        RECT 2380.590 2792.235 2380.870 2792.605 ;
        RECT 2380.660 2792.070 2380.800 2792.235 ;
        RECT 2385.720 2792.070 2385.860 2794.275 ;
        RECT 2387.960 2792.090 2388.220 2792.410 ;
        RECT 2380.600 2791.750 2380.860 2792.070 ;
        RECT 2381.050 2791.555 2381.330 2791.925 ;
        RECT 2381.520 2791.750 2381.780 2792.070 ;
        RECT 2385.660 2791.750 2385.920 2792.070 ;
        RECT 2381.120 2791.390 2381.260 2791.555 ;
        RECT 2381.060 2791.070 2381.320 2791.390 ;
        RECT 2381.580 2787.990 2381.720 2791.750 ;
        RECT 2387.490 2791.555 2387.770 2791.925 ;
        RECT 2387.500 2791.410 2387.760 2791.555 ;
        RECT 2388.020 2791.390 2388.160 2792.090 ;
        RECT 2391.240 2791.390 2391.380 2794.275 ;
        RECT 2387.960 2791.070 2388.220 2791.390 ;
        RECT 2391.180 2791.070 2391.440 2791.390 ;
        RECT 2394.390 2790.875 2394.670 2791.245 ;
        RECT 2394.920 2791.050 2395.060 2794.275 ;
        RECT 2402.680 2794.130 2402.940 2794.275 ;
        RECT 2415.160 2794.110 2415.300 2794.275 ;
        RECT 2401.750 2793.595 2402.030 2793.965 ;
        RECT 2408.190 2793.595 2408.470 2793.965 ;
        RECT 2415.100 2793.790 2415.360 2794.110 ;
        RECT 2401.820 2792.750 2401.960 2793.595 ;
        RECT 2408.200 2793.450 2408.460 2793.595 ;
        RECT 2421.990 2792.915 2422.270 2793.285 ;
        RECT 2442.690 2792.915 2442.970 2793.285 ;
        RECT 2422.000 2792.770 2422.260 2792.915 ;
        RECT 2401.760 2792.430 2402.020 2792.750 ;
        RECT 2408.190 2792.235 2408.470 2792.605 ;
        RECT 2428.890 2792.235 2429.170 2792.605 ;
        RECT 2435.790 2792.235 2436.070 2792.605 ;
        RECT 2394.400 2790.730 2394.660 2790.875 ;
        RECT 2394.860 2790.730 2395.120 2791.050 ;
        RECT 2394.920 2790.030 2395.060 2790.730 ;
        RECT 2408.260 2790.370 2408.400 2792.235 ;
        RECT 2428.960 2792.070 2429.100 2792.235 ;
        RECT 2428.900 2791.750 2429.160 2792.070 ;
        RECT 2435.860 2791.390 2436.000 2792.235 ;
        RECT 2415.090 2790.875 2415.370 2791.245 ;
        RECT 2421.990 2790.875 2422.270 2791.245 ;
        RECT 2428.890 2790.875 2429.170 2791.245 ;
        RECT 2435.800 2791.070 2436.060 2791.390 ;
        RECT 2442.760 2791.050 2442.900 2792.915 ;
        RECT 2415.160 2790.710 2415.300 2790.875 ;
        RECT 2415.100 2790.390 2415.360 2790.710 ;
        RECT 2408.200 2790.050 2408.460 2790.370 ;
        RECT 2415.550 2790.195 2415.830 2790.565 ;
        RECT 2394.860 2789.710 2395.120 2790.030 ;
        RECT 2415.620 2788.670 2415.760 2790.195 ;
        RECT 2422.060 2789.010 2422.200 2790.875 ;
        RECT 2422.000 2788.690 2422.260 2789.010 ;
        RECT 2415.090 2788.155 2415.370 2788.525 ;
        RECT 2415.560 2788.350 2415.820 2788.670 ;
        RECT 2428.960 2788.330 2429.100 2790.875 ;
        RECT 2442.700 2790.730 2442.960 2791.050 ;
        RECT 2442.690 2790.195 2442.970 2790.565 ;
        RECT 2435.790 2789.515 2436.070 2789.885 ;
        RECT 2442.760 2789.690 2442.900 2790.195 ;
        RECT 2435.860 2789.350 2436.000 2789.515 ;
        RECT 2442.700 2789.370 2442.960 2789.690 ;
        RECT 2435.800 2789.030 2436.060 2789.350 ;
        RECT 2415.160 2787.990 2415.300 2788.155 ;
        RECT 2428.900 2788.010 2429.160 2788.330 ;
        RECT 2367.260 2787.670 2367.520 2787.990 ;
        RECT 2373.240 2787.845 2373.500 2787.990 ;
        RECT 2373.230 2787.475 2373.510 2787.845 ;
        RECT 2381.520 2787.670 2381.780 2787.990 ;
        RECT 2381.980 2787.845 2382.240 2787.990 ;
        RECT 2381.970 2787.475 2382.250 2787.845 ;
        RECT 2415.100 2787.670 2415.360 2787.990 ;
        RECT 2366.800 2566.330 2367.060 2566.650 ;
        RECT 2359.900 2552.730 2360.160 2553.050 ;
        RECT 2353.000 2545.930 2353.260 2546.250 ;
        RECT 2346.100 2531.990 2346.360 2532.310 ;
        RECT 2339.660 2525.190 2339.920 2525.510 ;
        RECT 2339.200 2511.250 2339.460 2511.570 ;
        RECT 2332.300 2504.450 2332.560 2504.770 ;
        RECT 2325.400 2497.310 2325.660 2497.630 ;
        RECT 2318.500 2483.710 2318.760 2484.030 ;
        RECT 2311.600 2476.910 2311.860 2477.230 ;
        RECT 2305.160 2462.970 2305.420 2463.290 ;
        RECT 2304.700 2456.170 2304.960 2456.490 ;
        RECT 2297.800 2442.230 2298.060 2442.550 ;
        RECT 2290.900 2435.430 2291.160 2435.750 ;
        RECT 2284.000 2421.490 2284.260 2421.810 ;
        RECT 2277.100 2414.690 2277.360 2415.010 ;
        RECT 2266.980 2400.750 2267.240 2401.070 ;
        RECT 2266.520 2059.390 2266.780 2059.710 ;
        RECT 2193.840 2052.930 2194.100 2053.250 ;
        RECT 2192.000 2052.590 2192.260 2052.910 ;
        RECT 1514.420 1717.690 1514.680 1718.010 ;
        RECT 1421.040 1696.270 1421.300 1696.590 ;
        RECT 1420.580 1687.770 1420.840 1688.090 ;
        RECT 1420.120 1675.870 1420.380 1676.190 ;
        RECT 1419.660 1666.010 1419.920 1666.330 ;
        RECT 1419.200 1655.470 1419.460 1655.790 ;
        RECT 1418.740 1645.270 1419.000 1645.590 ;
        RECT 1418.280 1635.070 1418.540 1635.390 ;
        RECT 1417.820 1625.210 1418.080 1625.530 ;
        RECT 1410.910 1604.955 1411.190 1605.325 ;
      LAYER met2 ;
        RECT 1555.000 1605.000 1931.480 2051.235 ;
        RECT 2205.000 1605.000 2581.480 2051.235 ;
        RECT 300.030 1604.000 300.660 1604.280 ;
        RECT 301.500 1604.000 302.500 1604.280 ;
        RECT 303.340 1604.000 304.800 1604.280 ;
        RECT 305.640 1604.000 307.100 1604.280 ;
        RECT 307.940 1604.000 309.400 1604.280 ;
        RECT 310.240 1604.000 311.700 1604.280 ;
        RECT 312.540 1604.000 314.000 1604.280 ;
        RECT 314.840 1604.000 316.300 1604.280 ;
        RECT 317.140 1604.000 318.600 1604.280 ;
        RECT 319.440 1604.000 320.440 1604.280 ;
        RECT 321.280 1604.000 322.740 1604.280 ;
        RECT 323.580 1604.000 325.040 1604.280 ;
        RECT 325.880 1604.000 327.340 1604.280 ;
        RECT 328.180 1604.000 329.640 1604.280 ;
        RECT 330.480 1604.000 331.940 1604.280 ;
        RECT 332.780 1604.000 334.240 1604.280 ;
        RECT 335.080 1604.000 336.540 1604.280 ;
        RECT 337.380 1604.000 338.380 1604.280 ;
        RECT 339.220 1604.000 340.680 1604.280 ;
        RECT 341.520 1604.000 342.980 1604.280 ;
        RECT 343.820 1604.000 345.280 1604.280 ;
        RECT 346.120 1604.000 347.580 1604.280 ;
        RECT 348.420 1604.000 349.880 1604.280 ;
        RECT 350.720 1604.000 352.180 1604.280 ;
        RECT 353.020 1604.000 354.480 1604.280 ;
        RECT 355.320 1604.000 356.320 1604.280 ;
        RECT 357.160 1604.000 358.620 1604.280 ;
        RECT 359.460 1604.000 360.920 1604.280 ;
        RECT 361.760 1604.000 363.220 1604.280 ;
        RECT 364.060 1604.000 365.520 1604.280 ;
        RECT 366.360 1604.000 367.820 1604.280 ;
        RECT 368.660 1604.000 370.120 1604.280 ;
        RECT 370.960 1604.000 372.420 1604.280 ;
        RECT 373.260 1604.000 374.720 1604.280 ;
        RECT 375.560 1604.000 376.560 1604.280 ;
        RECT 377.400 1604.000 378.860 1604.280 ;
        RECT 379.700 1604.000 381.160 1604.280 ;
        RECT 382.000 1604.000 383.460 1604.280 ;
        RECT 384.300 1604.000 385.760 1604.280 ;
        RECT 386.600 1604.000 388.060 1604.280 ;
        RECT 388.900 1604.000 390.360 1604.280 ;
        RECT 391.200 1604.000 392.660 1604.280 ;
        RECT 393.500 1604.000 394.500 1604.280 ;
        RECT 395.340 1604.000 396.800 1604.280 ;
        RECT 397.640 1604.000 399.100 1604.280 ;
        RECT 399.940 1604.000 401.400 1604.280 ;
        RECT 402.240 1604.000 403.700 1604.280 ;
        RECT 404.540 1604.000 406.000 1604.280 ;
        RECT 406.840 1604.000 408.300 1604.280 ;
        RECT 409.140 1604.000 410.600 1604.280 ;
        RECT 411.440 1604.000 412.440 1604.280 ;
        RECT 413.280 1604.000 414.740 1604.280 ;
        RECT 415.580 1604.000 417.040 1604.280 ;
        RECT 417.880 1604.000 419.340 1604.280 ;
        RECT 420.180 1604.000 421.640 1604.280 ;
        RECT 422.480 1604.000 423.940 1604.280 ;
        RECT 424.780 1604.000 426.240 1604.280 ;
        RECT 427.080 1604.000 428.540 1604.280 ;
        RECT 429.380 1604.000 430.840 1604.280 ;
        RECT 431.680 1604.000 432.680 1604.280 ;
        RECT 433.520 1604.000 434.980 1604.280 ;
        RECT 435.820 1604.000 437.280 1604.280 ;
        RECT 438.120 1604.000 439.580 1604.280 ;
        RECT 440.420 1604.000 441.880 1604.280 ;
        RECT 442.720 1604.000 444.180 1604.280 ;
        RECT 445.020 1604.000 446.480 1604.280 ;
        RECT 447.320 1604.000 448.780 1604.280 ;
        RECT 449.620 1604.000 450.620 1604.280 ;
        RECT 451.460 1604.000 452.920 1604.280 ;
        RECT 453.760 1604.000 455.220 1604.280 ;
        RECT 456.060 1604.000 457.520 1604.280 ;
        RECT 458.360 1604.000 459.820 1604.280 ;
        RECT 460.660 1604.000 462.120 1604.280 ;
        RECT 462.960 1604.000 464.420 1604.280 ;
        RECT 465.260 1604.000 466.720 1604.280 ;
        RECT 467.560 1604.000 468.560 1604.280 ;
        RECT 469.400 1604.000 470.860 1604.280 ;
        RECT 471.700 1604.000 473.160 1604.280 ;
        RECT 474.000 1604.000 475.460 1604.280 ;
        RECT 476.300 1604.000 477.760 1604.280 ;
        RECT 478.600 1604.000 480.060 1604.280 ;
        RECT 480.900 1604.000 482.360 1604.280 ;
        RECT 483.200 1604.000 484.660 1604.280 ;
        RECT 485.500 1604.000 486.960 1604.280 ;
        RECT 487.800 1604.000 488.800 1604.280 ;
        RECT 489.640 1604.000 491.100 1604.280 ;
        RECT 491.940 1604.000 493.400 1604.280 ;
        RECT 494.240 1604.000 495.700 1604.280 ;
        RECT 496.540 1604.000 498.000 1604.280 ;
        RECT 498.840 1604.000 500.300 1604.280 ;
        RECT 501.140 1604.000 502.600 1604.280 ;
        RECT 503.440 1604.000 504.900 1604.280 ;
        RECT 505.740 1604.000 506.740 1604.280 ;
        RECT 507.580 1604.000 509.040 1604.280 ;
        RECT 509.880 1604.000 511.340 1604.280 ;
        RECT 512.180 1604.000 513.640 1604.280 ;
        RECT 514.480 1604.000 515.940 1604.280 ;
        RECT 516.780 1604.000 518.240 1604.280 ;
        RECT 519.080 1604.000 520.540 1604.280 ;
        RECT 521.380 1604.000 522.840 1604.280 ;
        RECT 523.680 1604.000 524.680 1604.280 ;
        RECT 525.520 1604.000 526.980 1604.280 ;
        RECT 527.820 1604.000 529.280 1604.280 ;
        RECT 530.120 1604.000 531.580 1604.280 ;
        RECT 532.420 1604.000 533.880 1604.280 ;
        RECT 534.720 1604.000 536.180 1604.280 ;
        RECT 537.020 1604.000 538.480 1604.280 ;
        RECT 539.320 1604.000 540.780 1604.280 ;
        RECT 541.620 1604.000 542.620 1604.280 ;
        RECT 543.460 1604.000 544.920 1604.280 ;
        RECT 545.760 1604.000 547.220 1604.280 ;
        RECT 548.060 1604.000 549.520 1604.280 ;
        RECT 550.360 1604.000 551.820 1604.280 ;
        RECT 552.660 1604.000 554.120 1604.280 ;
        RECT 554.960 1604.000 556.420 1604.280 ;
        RECT 557.260 1604.000 558.720 1604.280 ;
        RECT 559.560 1604.000 561.020 1604.280 ;
        RECT 561.860 1604.000 562.860 1604.280 ;
        RECT 563.700 1604.000 565.160 1604.280 ;
        RECT 566.000 1604.000 567.460 1604.280 ;
        RECT 568.300 1604.000 569.760 1604.280 ;
        RECT 570.600 1604.000 572.060 1604.280 ;
        RECT 572.900 1604.000 574.360 1604.280 ;
        RECT 575.200 1604.000 576.660 1604.280 ;
        RECT 577.500 1604.000 578.960 1604.280 ;
        RECT 579.800 1604.000 580.800 1604.280 ;
        RECT 581.640 1604.000 583.100 1604.280 ;
        RECT 583.940 1604.000 585.400 1604.280 ;
        RECT 586.240 1604.000 587.700 1604.280 ;
        RECT 588.540 1604.000 590.000 1604.280 ;
        RECT 590.840 1604.000 592.300 1604.280 ;
        RECT 593.140 1604.000 594.600 1604.280 ;
        RECT 595.440 1604.000 596.900 1604.280 ;
        RECT 597.740 1604.000 598.740 1604.280 ;
        RECT 599.580 1604.000 601.040 1604.280 ;
        RECT 601.880 1604.000 603.340 1604.280 ;
        RECT 604.180 1604.000 605.640 1604.280 ;
        RECT 606.480 1604.000 607.940 1604.280 ;
        RECT 608.780 1604.000 610.240 1604.280 ;
        RECT 611.080 1604.000 612.540 1604.280 ;
        RECT 613.380 1604.000 614.840 1604.280 ;
        RECT 615.680 1604.000 617.140 1604.280 ;
        RECT 617.980 1604.000 618.980 1604.280 ;
        RECT 619.820 1604.000 621.280 1604.280 ;
        RECT 622.120 1604.000 623.580 1604.280 ;
        RECT 624.420 1604.000 625.880 1604.280 ;
        RECT 626.720 1604.000 628.180 1604.280 ;
        RECT 629.020 1604.000 630.480 1604.280 ;
        RECT 631.320 1604.000 632.780 1604.280 ;
        RECT 633.620 1604.000 635.080 1604.280 ;
        RECT 635.920 1604.000 636.920 1604.280 ;
        RECT 637.760 1604.000 639.220 1604.280 ;
        RECT 640.060 1604.000 641.520 1604.280 ;
        RECT 642.360 1604.000 643.820 1604.280 ;
        RECT 644.660 1604.000 646.120 1604.280 ;
        RECT 646.960 1604.000 648.420 1604.280 ;
        RECT 649.260 1604.000 650.720 1604.280 ;
        RECT 651.560 1604.000 653.020 1604.280 ;
        RECT 653.860 1604.000 654.860 1604.280 ;
        RECT 655.700 1604.000 657.160 1604.280 ;
        RECT 658.000 1604.000 659.460 1604.280 ;
        RECT 660.300 1604.000 661.760 1604.280 ;
        RECT 662.600 1604.000 664.060 1604.280 ;
        RECT 664.900 1604.000 666.360 1604.280 ;
        RECT 667.200 1604.000 668.660 1604.280 ;
        RECT 669.500 1604.000 670.960 1604.280 ;
        RECT 671.800 1604.000 673.260 1604.280 ;
        RECT 674.100 1604.000 675.100 1604.280 ;
        RECT 675.940 1604.000 677.400 1604.280 ;
        RECT 678.240 1604.000 679.700 1604.280 ;
        RECT 680.540 1604.000 682.000 1604.280 ;
        RECT 682.840 1604.000 684.300 1604.280 ;
        RECT 685.140 1604.000 686.600 1604.280 ;
        RECT 687.440 1604.000 688.900 1604.280 ;
        RECT 689.740 1604.000 691.200 1604.280 ;
        RECT 692.040 1604.000 693.040 1604.280 ;
        RECT 693.880 1604.000 695.340 1604.280 ;
        RECT 696.180 1604.000 697.640 1604.280 ;
        RECT 698.480 1604.000 699.940 1604.280 ;
        RECT 700.780 1604.000 702.240 1604.280 ;
        RECT 703.080 1604.000 704.540 1604.280 ;
        RECT 705.380 1604.000 706.840 1604.280 ;
        RECT 707.680 1604.000 709.140 1604.280 ;
        RECT 709.980 1604.000 710.980 1604.280 ;
        RECT 711.820 1604.000 713.280 1604.280 ;
        RECT 714.120 1604.000 715.580 1604.280 ;
        RECT 716.420 1604.000 717.880 1604.280 ;
        RECT 718.720 1604.000 720.180 1604.280 ;
        RECT 721.020 1604.000 722.480 1604.280 ;
        RECT 723.320 1604.000 724.780 1604.280 ;
        RECT 725.620 1604.000 727.080 1604.280 ;
        RECT 727.920 1604.000 729.380 1604.280 ;
        RECT 730.220 1604.000 731.220 1604.280 ;
        RECT 732.060 1604.000 733.520 1604.280 ;
        RECT 734.360 1604.000 735.820 1604.280 ;
        RECT 736.660 1604.000 738.120 1604.280 ;
        RECT 738.960 1604.000 740.420 1604.280 ;
        RECT 741.260 1604.000 742.720 1604.280 ;
        RECT 743.560 1604.000 745.020 1604.280 ;
        RECT 745.860 1604.000 747.320 1604.280 ;
        RECT 748.160 1604.000 749.160 1604.280 ;
        RECT 750.000 1604.000 751.460 1604.280 ;
        RECT 752.300 1604.000 753.760 1604.280 ;
        RECT 754.600 1604.000 756.060 1604.280 ;
        RECT 756.900 1604.000 758.360 1604.280 ;
        RECT 759.200 1604.000 760.660 1604.280 ;
        RECT 761.500 1604.000 762.960 1604.280 ;
        RECT 763.800 1604.000 765.260 1604.280 ;
        RECT 766.100 1604.000 767.100 1604.280 ;
        RECT 767.940 1604.000 769.400 1604.280 ;
        RECT 770.240 1604.000 771.700 1604.280 ;
        RECT 772.540 1604.000 774.000 1604.280 ;
        RECT 774.840 1604.000 776.300 1604.280 ;
        RECT 777.140 1604.000 778.600 1604.280 ;
        RECT 779.440 1604.000 780.900 1604.280 ;
        RECT 781.740 1604.000 783.200 1604.280 ;
        RECT 784.040 1604.000 785.040 1604.280 ;
        RECT 785.880 1604.000 787.340 1604.280 ;
        RECT 788.180 1604.000 789.640 1604.280 ;
        RECT 790.480 1604.000 791.940 1604.280 ;
        RECT 792.780 1604.000 794.240 1604.280 ;
        RECT 795.080 1604.000 796.540 1604.280 ;
        RECT 797.380 1604.000 798.840 1604.280 ;
        RECT 799.680 1604.000 801.140 1604.280 ;
        RECT 801.980 1604.000 803.440 1604.280 ;
        RECT 804.280 1604.000 805.280 1604.280 ;
        RECT 806.120 1604.000 807.580 1604.280 ;
        RECT 808.420 1604.000 809.880 1604.280 ;
        RECT 810.720 1604.000 812.180 1604.280 ;
        RECT 813.020 1604.000 814.480 1604.280 ;
        RECT 815.320 1604.000 816.780 1604.280 ;
        RECT 817.620 1604.000 819.080 1604.280 ;
        RECT 819.920 1604.000 821.380 1604.280 ;
        RECT 822.220 1604.000 823.220 1604.280 ;
        RECT 824.060 1604.000 825.520 1604.280 ;
        RECT 826.360 1604.000 827.820 1604.280 ;
        RECT 828.660 1604.000 830.120 1604.280 ;
        RECT 830.960 1604.000 832.420 1604.280 ;
        RECT 833.260 1604.000 834.720 1604.280 ;
        RECT 835.560 1604.000 837.020 1604.280 ;
        RECT 837.860 1604.000 839.320 1604.280 ;
        RECT 840.160 1604.000 841.160 1604.280 ;
        RECT 842.000 1604.000 843.460 1604.280 ;
        RECT 844.300 1604.000 845.760 1604.280 ;
        RECT 846.600 1604.000 848.060 1604.280 ;
        RECT 848.900 1604.000 850.360 1604.280 ;
        RECT 851.200 1604.000 852.660 1604.280 ;
        RECT 853.500 1604.000 854.960 1604.280 ;
        RECT 855.800 1604.000 857.260 1604.280 ;
        RECT 858.100 1604.000 859.560 1604.280 ;
        RECT 860.400 1604.000 861.400 1604.280 ;
        RECT 862.240 1604.000 863.700 1604.280 ;
        RECT 864.540 1604.000 866.000 1604.280 ;
        RECT 866.840 1604.000 868.300 1604.280 ;
        RECT 869.140 1604.000 870.600 1604.280 ;
        RECT 871.440 1604.000 872.900 1604.280 ;
        RECT 873.740 1604.000 875.200 1604.280 ;
        RECT 876.040 1604.000 877.500 1604.280 ;
        RECT 878.340 1604.000 879.340 1604.280 ;
        RECT 880.180 1604.000 881.640 1604.280 ;
        RECT 882.480 1604.000 883.940 1604.280 ;
        RECT 884.780 1604.000 886.240 1604.280 ;
        RECT 887.080 1604.000 888.540 1604.280 ;
        RECT 889.380 1604.000 890.840 1604.280 ;
        RECT 891.680 1604.000 893.140 1604.280 ;
        RECT 893.980 1604.000 895.440 1604.280 ;
        RECT 896.280 1604.000 897.280 1604.280 ;
        RECT 898.120 1604.000 899.580 1604.280 ;
        RECT 900.420 1604.000 901.880 1604.280 ;
        RECT 902.720 1604.000 904.180 1604.280 ;
        RECT 905.020 1604.000 906.480 1604.280 ;
        RECT 907.320 1604.000 908.780 1604.280 ;
        RECT 909.620 1604.000 911.080 1604.280 ;
        RECT 911.920 1604.000 913.380 1604.280 ;
        RECT 914.220 1604.000 915.680 1604.280 ;
        RECT 916.520 1604.000 917.520 1604.280 ;
        RECT 918.360 1604.000 919.820 1604.280 ;
        RECT 920.660 1604.000 922.120 1604.280 ;
        RECT 922.960 1604.000 924.420 1604.280 ;
        RECT 925.260 1604.000 926.720 1604.280 ;
        RECT 927.560 1604.000 929.020 1604.280 ;
        RECT 929.860 1604.000 931.320 1604.280 ;
        RECT 932.160 1604.000 933.620 1604.280 ;
        RECT 934.460 1604.000 935.460 1604.280 ;
        RECT 936.300 1604.000 937.760 1604.280 ;
        RECT 938.600 1604.000 940.060 1604.280 ;
        RECT 940.900 1604.000 942.360 1604.280 ;
        RECT 943.200 1604.000 944.660 1604.280 ;
        RECT 945.500 1604.000 946.960 1604.280 ;
        RECT 947.800 1604.000 949.260 1604.280 ;
        RECT 950.100 1604.000 951.560 1604.280 ;
        RECT 952.400 1604.000 953.400 1604.280 ;
        RECT 954.240 1604.000 955.700 1604.280 ;
        RECT 956.540 1604.000 958.000 1604.280 ;
        RECT 958.840 1604.000 960.300 1604.280 ;
        RECT 961.140 1604.000 962.600 1604.280 ;
        RECT 963.440 1604.000 964.900 1604.280 ;
        RECT 965.740 1604.000 967.200 1604.280 ;
        RECT 968.040 1604.000 969.500 1604.280 ;
        RECT 970.340 1604.000 971.340 1604.280 ;
        RECT 972.180 1604.000 973.640 1604.280 ;
        RECT 974.480 1604.000 975.940 1604.280 ;
        RECT 976.780 1604.000 978.240 1604.280 ;
        RECT 979.080 1604.000 980.540 1604.280 ;
        RECT 981.380 1604.000 982.840 1604.280 ;
        RECT 983.680 1604.000 985.140 1604.280 ;
        RECT 985.980 1604.000 987.440 1604.280 ;
        RECT 988.280 1604.000 989.740 1604.280 ;
        RECT 990.580 1604.000 991.580 1604.280 ;
        RECT 992.420 1604.000 993.880 1604.280 ;
        RECT 994.720 1604.000 996.180 1604.280 ;
        RECT 997.020 1604.000 998.480 1604.280 ;
        RECT 999.320 1604.000 1000.780 1604.280 ;
        RECT 1001.620 1604.000 1003.080 1604.280 ;
        RECT 1003.920 1604.000 1005.380 1604.280 ;
        RECT 1006.220 1604.000 1007.680 1604.280 ;
        RECT 1008.520 1604.000 1009.520 1604.280 ;
        RECT 1010.360 1604.000 1011.820 1604.280 ;
        RECT 1012.660 1604.000 1014.120 1604.280 ;
        RECT 1014.960 1604.000 1016.420 1604.280 ;
        RECT 1017.260 1604.000 1018.720 1604.280 ;
        RECT 1019.560 1604.000 1021.020 1604.280 ;
        RECT 1021.860 1604.000 1023.320 1604.280 ;
        RECT 1024.160 1604.000 1025.620 1604.280 ;
        RECT 1026.460 1604.000 1027.460 1604.280 ;
        RECT 1028.300 1604.000 1029.760 1604.280 ;
        RECT 1030.600 1604.000 1032.060 1604.280 ;
        RECT 1032.900 1604.000 1034.360 1604.280 ;
        RECT 1035.200 1604.000 1036.660 1604.280 ;
        RECT 1037.500 1604.000 1038.960 1604.280 ;
        RECT 1039.800 1604.000 1041.260 1604.280 ;
        RECT 1042.100 1604.000 1043.560 1604.280 ;
        RECT 1044.400 1604.000 1045.860 1604.280 ;
        RECT 1046.700 1604.000 1047.700 1604.280 ;
        RECT 1048.540 1604.000 1050.000 1604.280 ;
        RECT 1050.840 1604.000 1052.300 1604.280 ;
        RECT 1053.140 1604.000 1054.600 1604.280 ;
        RECT 1055.440 1604.000 1056.900 1604.280 ;
        RECT 1057.740 1604.000 1059.200 1604.280 ;
        RECT 1060.040 1604.000 1061.500 1604.280 ;
        RECT 1062.340 1604.000 1063.800 1604.280 ;
        RECT 1064.640 1604.000 1065.640 1604.280 ;
        RECT 1066.480 1604.000 1067.940 1604.280 ;
        RECT 1068.780 1604.000 1070.240 1604.280 ;
        RECT 1071.080 1604.000 1072.540 1604.280 ;
        RECT 1073.380 1604.000 1074.840 1604.280 ;
        RECT 1075.680 1604.000 1077.140 1604.280 ;
        RECT 1077.980 1604.000 1079.440 1604.280 ;
        RECT 1080.280 1604.000 1081.740 1604.280 ;
        RECT 1082.580 1604.000 1083.580 1604.280 ;
        RECT 1084.420 1604.000 1085.880 1604.280 ;
        RECT 1086.720 1604.000 1088.180 1604.280 ;
        RECT 1089.020 1604.000 1090.480 1604.280 ;
        RECT 1091.320 1604.000 1092.780 1604.280 ;
        RECT 1093.620 1604.000 1095.080 1604.280 ;
        RECT 1095.920 1604.000 1097.380 1604.280 ;
        RECT 1098.220 1604.000 1099.680 1604.280 ;
        RECT 1100.520 1604.000 1101.980 1604.280 ;
        RECT 1102.820 1604.000 1103.820 1604.280 ;
        RECT 1104.660 1604.000 1106.120 1604.280 ;
        RECT 1106.960 1604.000 1108.420 1604.280 ;
        RECT 1109.260 1604.000 1110.720 1604.280 ;
        RECT 1111.560 1604.000 1113.020 1604.280 ;
        RECT 1113.860 1604.000 1115.320 1604.280 ;
        RECT 1116.160 1604.000 1117.620 1604.280 ;
        RECT 1118.460 1604.000 1119.920 1604.280 ;
        RECT 1120.760 1604.000 1121.760 1604.280 ;
        RECT 1122.600 1604.000 1124.060 1604.280 ;
        RECT 1124.900 1604.000 1126.360 1604.280 ;
        RECT 1127.200 1604.000 1128.660 1604.280 ;
        RECT 1129.500 1604.000 1130.960 1604.280 ;
        RECT 1131.800 1604.000 1133.260 1604.280 ;
        RECT 1134.100 1604.000 1135.560 1604.280 ;
        RECT 1136.400 1604.000 1137.860 1604.280 ;
        RECT 1138.700 1604.000 1139.700 1604.280 ;
        RECT 1140.540 1604.000 1142.000 1604.280 ;
        RECT 1142.840 1604.000 1144.300 1604.280 ;
        RECT 1145.140 1604.000 1146.600 1604.280 ;
        RECT 1147.440 1604.000 1148.900 1604.280 ;
        RECT 1149.740 1604.000 1151.200 1604.280 ;
        RECT 1152.040 1604.000 1153.500 1604.280 ;
        RECT 1154.340 1604.000 1155.800 1604.280 ;
        RECT 1156.640 1604.000 1158.100 1604.280 ;
        RECT 1158.940 1604.000 1159.940 1604.280 ;
        RECT 1160.780 1604.000 1162.240 1604.280 ;
        RECT 1163.080 1604.000 1164.540 1604.280 ;
        RECT 1165.380 1604.000 1166.840 1604.280 ;
        RECT 1167.680 1604.000 1169.140 1604.280 ;
        RECT 1169.980 1604.000 1171.440 1604.280 ;
        RECT 1172.280 1604.000 1173.740 1604.280 ;
        RECT 1174.580 1604.000 1176.040 1604.280 ;
        RECT 1176.880 1604.000 1177.880 1604.280 ;
        RECT 1178.720 1604.000 1180.180 1604.280 ;
        RECT 1181.020 1604.000 1182.480 1604.280 ;
        RECT 1183.320 1604.000 1184.780 1604.280 ;
        RECT 1185.620 1604.000 1187.080 1604.280 ;
        RECT 1187.920 1604.000 1189.380 1604.280 ;
        RECT 1190.220 1604.000 1191.680 1604.280 ;
        RECT 1192.520 1604.000 1193.980 1604.280 ;
        RECT 1194.820 1604.000 1195.820 1604.280 ;
        RECT 1196.660 1604.000 1198.120 1604.280 ;
        RECT 1198.960 1604.000 1200.420 1604.280 ;
        RECT 1201.260 1604.000 1202.720 1604.280 ;
        RECT 1203.560 1604.000 1205.020 1604.280 ;
        RECT 1205.860 1604.000 1207.320 1604.280 ;
        RECT 1208.160 1604.000 1209.620 1604.280 ;
        RECT 1210.460 1604.000 1211.920 1604.280 ;
        RECT 1212.760 1604.000 1213.760 1604.280 ;
        RECT 1214.600 1604.000 1216.060 1604.280 ;
        RECT 1216.900 1604.000 1218.360 1604.280 ;
        RECT 1219.200 1604.000 1220.660 1604.280 ;
        RECT 1221.500 1604.000 1222.960 1604.280 ;
        RECT 1223.800 1604.000 1225.260 1604.280 ;
        RECT 1226.100 1604.000 1227.560 1604.280 ;
        RECT 1228.400 1604.000 1229.860 1604.280 ;
        RECT 1230.700 1604.000 1232.160 1604.280 ;
        RECT 1233.000 1604.000 1234.000 1604.280 ;
        RECT 1234.840 1604.000 1236.300 1604.280 ;
        RECT 1237.140 1604.000 1238.600 1604.280 ;
        RECT 1239.440 1604.000 1240.900 1604.280 ;
        RECT 1241.740 1604.000 1243.200 1604.280 ;
        RECT 1244.040 1604.000 1245.500 1604.280 ;
        RECT 1246.340 1604.000 1247.800 1604.280 ;
        RECT 1248.640 1604.000 1250.100 1604.280 ;
        RECT 1250.940 1604.000 1251.940 1604.280 ;
        RECT 1252.780 1604.000 1254.240 1604.280 ;
        RECT 1255.080 1604.000 1256.540 1604.280 ;
        RECT 1257.380 1604.000 1258.840 1604.280 ;
        RECT 1259.680 1604.000 1261.140 1604.280 ;
        RECT 1261.980 1604.000 1263.440 1604.280 ;
        RECT 1264.280 1604.000 1265.740 1604.280 ;
        RECT 1266.580 1604.000 1268.040 1604.280 ;
        RECT 1268.880 1604.000 1269.880 1604.280 ;
        RECT 1270.720 1604.000 1272.180 1604.280 ;
        RECT 1273.020 1604.000 1274.480 1604.280 ;
        RECT 1275.320 1604.000 1276.780 1604.280 ;
        RECT 1277.620 1604.000 1279.080 1604.280 ;
        RECT 1279.920 1604.000 1281.380 1604.280 ;
        RECT 1282.220 1604.000 1283.680 1604.280 ;
        RECT 1284.520 1604.000 1285.980 1604.280 ;
        RECT 1286.820 1604.000 1288.280 1604.280 ;
        RECT 1289.120 1604.000 1290.120 1604.280 ;
        RECT 1290.960 1604.000 1292.420 1604.280 ;
        RECT 1293.260 1604.000 1294.720 1604.280 ;
        RECT 1295.560 1604.000 1297.020 1604.280 ;
        RECT 1297.860 1604.000 1299.320 1604.280 ;
        RECT 1300.160 1604.000 1301.620 1604.280 ;
        RECT 1302.460 1604.000 1303.920 1604.280 ;
        RECT 1304.760 1604.000 1306.220 1604.280 ;
        RECT 1307.060 1604.000 1308.060 1604.280 ;
        RECT 1308.900 1604.000 1310.360 1604.280 ;
        RECT 1311.200 1604.000 1312.660 1604.280 ;
        RECT 1313.500 1604.000 1314.960 1604.280 ;
        RECT 1315.800 1604.000 1317.260 1604.280 ;
        RECT 1318.100 1604.000 1319.560 1604.280 ;
        RECT 1320.400 1604.000 1321.860 1604.280 ;
        RECT 1322.700 1604.000 1324.160 1604.280 ;
        RECT 1325.000 1604.000 1326.000 1604.280 ;
        RECT 1326.840 1604.000 1328.300 1604.280 ;
        RECT 1329.140 1604.000 1330.600 1604.280 ;
        RECT 1331.440 1604.000 1332.900 1604.280 ;
        RECT 1333.740 1604.000 1335.200 1604.280 ;
        RECT 1336.040 1604.000 1337.500 1604.280 ;
        RECT 1338.340 1604.000 1339.800 1604.280 ;
        RECT 1340.640 1604.000 1342.100 1604.280 ;
        RECT 1342.940 1604.000 1344.400 1604.280 ;
        RECT 1345.240 1604.000 1346.240 1604.280 ;
        RECT 1347.080 1604.000 1348.540 1604.280 ;
        RECT 1349.380 1604.000 1350.840 1604.280 ;
        RECT 1351.680 1604.000 1353.140 1604.280 ;
        RECT 1353.980 1604.000 1355.440 1604.280 ;
        RECT 1356.280 1604.000 1357.740 1604.280 ;
        RECT 1358.580 1604.000 1360.040 1604.280 ;
        RECT 1360.880 1604.000 1362.340 1604.280 ;
        RECT 1363.180 1604.000 1364.180 1604.280 ;
        RECT 1365.020 1604.000 1366.480 1604.280 ;
        RECT 1367.320 1604.000 1368.780 1604.280 ;
        RECT 1369.620 1604.000 1371.080 1604.280 ;
        RECT 1371.920 1604.000 1373.380 1604.280 ;
        RECT 1374.220 1604.000 1375.680 1604.280 ;
        RECT 1376.520 1604.000 1377.980 1604.280 ;
        RECT 1378.820 1604.000 1380.280 1604.280 ;
        RECT 1381.120 1604.000 1382.120 1604.280 ;
        RECT 1382.960 1604.000 1384.420 1604.280 ;
        RECT 1385.260 1604.000 1386.720 1604.280 ;
        RECT 1387.560 1604.000 1389.020 1604.280 ;
        RECT 1389.860 1604.000 1391.320 1604.280 ;
        RECT 1392.160 1604.000 1393.620 1604.280 ;
        RECT 1394.460 1604.000 1395.920 1604.280 ;
      LAYER met2 ;
        RECT 1555.080 1496.000 1555.360 1500.000 ;
        RECT 1565.200 1496.000 1565.480 1500.000 ;
        RECT 1575.780 1496.000 1576.060 1500.000 ;
        RECT 1585.900 1496.000 1586.180 1500.000 ;
        RECT 1596.480 1496.000 1596.760 1500.000 ;
        RECT 1606.600 1496.000 1606.880 1500.000 ;
        RECT 1617.180 1496.000 1617.460 1500.000 ;
        RECT 1627.300 1496.000 1627.580 1500.000 ;
        RECT 1637.880 1496.000 1638.160 1500.000 ;
        RECT 1648.460 1496.000 1648.740 1500.000 ;
        RECT 1658.580 1496.000 1658.860 1500.000 ;
        RECT 1669.160 1496.000 1669.440 1500.000 ;
        RECT 1679.280 1496.000 1679.560 1500.000 ;
        RECT 1689.860 1496.000 1690.140 1500.000 ;
        RECT 1699.980 1496.000 1700.260 1500.000 ;
        RECT 1710.560 1496.000 1710.840 1500.000 ;
        RECT 1720.680 1496.000 1720.960 1500.000 ;
        RECT 1731.260 1496.000 1731.540 1500.000 ;
        RECT 1741.840 1496.000 1742.120 1500.000 ;
        RECT 1751.960 1496.000 1752.240 1500.000 ;
        RECT 1762.540 1496.000 1762.820 1500.000 ;
        RECT 1772.660 1496.000 1772.940 1500.000 ;
        RECT 1783.240 1496.000 1783.520 1500.000 ;
        RECT 1793.360 1496.000 1793.640 1500.000 ;
        RECT 1803.940 1496.000 1804.220 1500.000 ;
        RECT 1814.060 1496.000 1814.340 1500.000 ;
        RECT 1824.640 1496.000 1824.920 1500.000 ;
        RECT 1835.220 1496.000 1835.500 1500.000 ;
        RECT 1845.340 1496.000 1845.620 1500.000 ;
        RECT 1855.920 1496.000 1856.200 1500.000 ;
        RECT 1866.040 1496.000 1866.320 1500.000 ;
        RECT 1876.620 1496.000 1876.900 1500.000 ;
        RECT 1886.740 1496.000 1887.020 1500.000 ;
        RECT 1897.320 1496.000 1897.600 1500.000 ;
        RECT 1907.440 1496.000 1907.720 1500.000 ;
        RECT 1918.020 1496.000 1918.300 1500.000 ;
        RECT 1928.600 1496.000 1928.880 1500.000 ;
        RECT 1938.720 1496.000 1939.000 1500.000 ;
        RECT 1949.300 1496.000 1949.580 1500.000 ;
        RECT 1959.420 1496.000 1959.700 1500.000 ;
        RECT 1970.000 1496.000 1970.280 1500.000 ;
        RECT 1980.120 1496.000 1980.400 1500.000 ;
        RECT 1990.700 1496.000 1990.980 1500.000 ;
        RECT 2000.820 1496.000 2001.100 1500.000 ;
        RECT 2011.400 1496.000 2011.680 1500.000 ;
        RECT 2021.980 1496.000 2022.260 1500.000 ;
        RECT 2032.100 1496.000 2032.380 1500.000 ;
        RECT 2042.680 1496.000 2042.960 1500.000 ;
        RECT 2052.800 1496.000 2053.080 1500.000 ;
        RECT 2063.380 1496.000 2063.660 1500.000 ;
        RECT 2073.500 1496.000 2073.780 1500.000 ;
        RECT 2084.080 1496.000 2084.360 1500.000 ;
        RECT 2094.200 1496.000 2094.480 1500.000 ;
        RECT 2104.780 1496.000 2105.060 1500.000 ;
        RECT 2115.360 1496.000 2115.640 1500.000 ;
        RECT 2125.480 1496.000 2125.760 1500.000 ;
        RECT 2136.060 1496.000 2136.340 1500.000 ;
        RECT 2146.180 1496.000 2146.460 1500.000 ;
        RECT 2156.760 1496.000 2157.040 1500.000 ;
        RECT 2166.880 1496.000 2167.160 1500.000 ;
        RECT 2177.460 1496.000 2177.740 1500.000 ;
        RECT 2187.580 1496.000 2187.860 1500.000 ;
        RECT 2198.160 1496.000 2198.440 1500.000 ;
        RECT 2208.740 1496.000 2209.020 1500.000 ;
        RECT 2218.860 1496.000 2219.140 1500.000 ;
        RECT 2229.440 1496.000 2229.720 1500.000 ;
        RECT 2239.560 1496.000 2239.840 1500.000 ;
        RECT 2250.140 1496.000 2250.420 1500.000 ;
        RECT 2260.260 1496.000 2260.540 1500.000 ;
        RECT 2270.840 1496.000 2271.120 1500.000 ;
        RECT 2280.960 1496.000 2281.240 1500.000 ;
        RECT 2291.540 1496.000 2291.820 1500.000 ;
        RECT 2302.120 1496.000 2302.400 1500.000 ;
        RECT 2312.240 1496.000 2312.520 1500.000 ;
        RECT 2322.820 1496.000 2323.100 1500.000 ;
        RECT 2332.940 1496.000 2333.220 1500.000 ;
        RECT 2343.520 1496.000 2343.800 1500.000 ;
        RECT 2353.640 1496.000 2353.920 1500.000 ;
        RECT 2364.220 1496.000 2364.500 1500.000 ;
        RECT 2374.340 1496.000 2374.620 1500.000 ;
        RECT 2384.920 1496.000 2385.200 1500.000 ;
        RECT 2395.500 1496.000 2395.780 1500.000 ;
        RECT 2405.620 1496.000 2405.900 1500.000 ;
        RECT 2416.200 1496.000 2416.480 1500.000 ;
        RECT 2426.320 1496.000 2426.600 1500.000 ;
        RECT 2436.900 1496.000 2437.180 1500.000 ;
        RECT 2447.020 1496.000 2447.300 1500.000 ;
        RECT 2457.600 1496.000 2457.880 1500.000 ;
        RECT 2467.720 1496.000 2468.000 1500.000 ;
        RECT 2478.300 1496.000 2478.580 1500.000 ;
        RECT 2488.880 1496.000 2489.160 1500.000 ;
        RECT 2499.000 1496.000 2499.280 1500.000 ;
        RECT 2509.580 1496.000 2509.860 1500.000 ;
        RECT 2519.700 1496.000 2519.980 1500.000 ;
        RECT 2530.280 1496.000 2530.560 1500.000 ;
        RECT 2540.400 1496.000 2540.680 1500.000 ;
        RECT 2550.980 1496.000 2551.260 1500.000 ;
        RECT 2561.100 1496.000 2561.380 1500.000 ;
        RECT 2571.680 1496.000 2571.960 1500.000 ;
        RECT 2582.260 1496.000 2582.540 1500.000 ;
        RECT 2592.380 1496.000 2592.660 1500.000 ;
        RECT 2602.960 1496.000 2603.240 1500.000 ;
        RECT 2613.080 1496.000 2613.360 1500.000 ;
        RECT 2623.660 1496.000 2623.940 1500.000 ;
        RECT 2633.780 1496.000 2634.060 1500.000 ;
        RECT 2644.360 1496.000 2644.640 1500.000 ;
      LAYER met2 ;
        RECT 1550.030 1495.720 1554.800 1496.000 ;
        RECT 1555.640 1495.720 1564.920 1496.000 ;
        RECT 1565.760 1495.720 1575.500 1496.000 ;
        RECT 1576.340 1495.720 1585.620 1496.000 ;
        RECT 1586.460 1495.720 1596.200 1496.000 ;
        RECT 1597.040 1495.720 1606.320 1496.000 ;
        RECT 1607.160 1495.720 1616.900 1496.000 ;
        RECT 1617.740 1495.720 1627.020 1496.000 ;
        RECT 1627.860 1495.720 1637.600 1496.000 ;
        RECT 1638.440 1495.720 1648.180 1496.000 ;
        RECT 1649.020 1495.720 1658.300 1496.000 ;
        RECT 1659.140 1495.720 1668.880 1496.000 ;
        RECT 1669.720 1495.720 1679.000 1496.000 ;
        RECT 1679.840 1495.720 1689.580 1496.000 ;
        RECT 1690.420 1495.720 1699.700 1496.000 ;
        RECT 1700.540 1495.720 1710.280 1496.000 ;
        RECT 1711.120 1495.720 1720.400 1496.000 ;
        RECT 1721.240 1495.720 1730.980 1496.000 ;
        RECT 1731.820 1495.720 1741.560 1496.000 ;
        RECT 1742.400 1495.720 1751.680 1496.000 ;
        RECT 1752.520 1495.720 1762.260 1496.000 ;
        RECT 1763.100 1495.720 1772.380 1496.000 ;
        RECT 1773.220 1495.720 1782.960 1496.000 ;
        RECT 1783.800 1495.720 1793.080 1496.000 ;
        RECT 1793.920 1495.720 1803.660 1496.000 ;
        RECT 1804.500 1495.720 1813.780 1496.000 ;
        RECT 1814.620 1495.720 1824.360 1496.000 ;
        RECT 1825.200 1495.720 1834.940 1496.000 ;
        RECT 1835.780 1495.720 1845.060 1496.000 ;
        RECT 1845.900 1495.720 1855.640 1496.000 ;
        RECT 1856.480 1495.720 1865.760 1496.000 ;
        RECT 1866.600 1495.720 1876.340 1496.000 ;
        RECT 1877.180 1495.720 1886.460 1496.000 ;
        RECT 1887.300 1495.720 1897.040 1496.000 ;
        RECT 1897.880 1495.720 1907.160 1496.000 ;
        RECT 1908.000 1495.720 1917.740 1496.000 ;
        RECT 1918.580 1495.720 1928.320 1496.000 ;
        RECT 1929.160 1495.720 1938.440 1496.000 ;
        RECT 1939.280 1495.720 1949.020 1496.000 ;
        RECT 1949.860 1495.720 1959.140 1496.000 ;
        RECT 1959.980 1495.720 1969.720 1496.000 ;
        RECT 1970.560 1495.720 1979.840 1496.000 ;
        RECT 1980.680 1495.720 1990.420 1496.000 ;
        RECT 1991.260 1495.720 2000.540 1496.000 ;
        RECT 2001.380 1495.720 2011.120 1496.000 ;
        RECT 2011.960 1495.720 2021.700 1496.000 ;
        RECT 2022.540 1495.720 2031.820 1496.000 ;
        RECT 2032.660 1495.720 2042.400 1496.000 ;
        RECT 2043.240 1495.720 2052.520 1496.000 ;
        RECT 2053.360 1495.720 2063.100 1496.000 ;
        RECT 2063.940 1495.720 2073.220 1496.000 ;
        RECT 2074.060 1495.720 2083.800 1496.000 ;
        RECT 2084.640 1495.720 2093.920 1496.000 ;
        RECT 2094.760 1495.720 2104.500 1496.000 ;
        RECT 2105.340 1495.720 2115.080 1496.000 ;
        RECT 2115.920 1495.720 2125.200 1496.000 ;
        RECT 2126.040 1495.720 2135.780 1496.000 ;
        RECT 2136.620 1495.720 2145.900 1496.000 ;
        RECT 2146.740 1495.720 2156.480 1496.000 ;
        RECT 2157.320 1495.720 2166.600 1496.000 ;
        RECT 2167.440 1495.720 2177.180 1496.000 ;
        RECT 2178.020 1495.720 2187.300 1496.000 ;
        RECT 2188.140 1495.720 2197.880 1496.000 ;
        RECT 2198.720 1495.720 2208.460 1496.000 ;
        RECT 2209.300 1495.720 2218.580 1496.000 ;
        RECT 2219.420 1495.720 2229.160 1496.000 ;
        RECT 2230.000 1495.720 2239.280 1496.000 ;
        RECT 2240.120 1495.720 2249.860 1496.000 ;
        RECT 2250.700 1495.720 2259.980 1496.000 ;
        RECT 2260.820 1495.720 2270.560 1496.000 ;
        RECT 2271.400 1495.720 2280.680 1496.000 ;
        RECT 2281.520 1495.720 2291.260 1496.000 ;
        RECT 2292.100 1495.720 2301.840 1496.000 ;
        RECT 2302.680 1495.720 2311.960 1496.000 ;
        RECT 2312.800 1495.720 2322.540 1496.000 ;
        RECT 2323.380 1495.720 2332.660 1496.000 ;
        RECT 2333.500 1495.720 2343.240 1496.000 ;
        RECT 2344.080 1495.720 2353.360 1496.000 ;
        RECT 2354.200 1495.720 2363.940 1496.000 ;
        RECT 2364.780 1495.720 2374.060 1496.000 ;
        RECT 2374.900 1495.720 2384.640 1496.000 ;
        RECT 2385.480 1495.720 2395.220 1496.000 ;
        RECT 2396.060 1495.720 2405.340 1496.000 ;
        RECT 2406.180 1495.720 2415.920 1496.000 ;
        RECT 2416.760 1495.720 2426.040 1496.000 ;
        RECT 2426.880 1495.720 2436.620 1496.000 ;
        RECT 2437.460 1495.720 2446.740 1496.000 ;
        RECT 2447.580 1495.720 2457.320 1496.000 ;
        RECT 2458.160 1495.720 2467.440 1496.000 ;
        RECT 2468.280 1495.720 2478.020 1496.000 ;
        RECT 2478.860 1495.720 2488.600 1496.000 ;
        RECT 2489.440 1495.720 2498.720 1496.000 ;
        RECT 2499.560 1495.720 2509.300 1496.000 ;
        RECT 2510.140 1495.720 2519.420 1496.000 ;
        RECT 2520.260 1495.720 2530.000 1496.000 ;
        RECT 2530.840 1495.720 2540.120 1496.000 ;
        RECT 2540.960 1495.720 2550.700 1496.000 ;
        RECT 2551.540 1495.720 2560.820 1496.000 ;
        RECT 2561.660 1495.720 2571.400 1496.000 ;
        RECT 2572.240 1495.720 2581.980 1496.000 ;
        RECT 2582.820 1495.720 2592.100 1496.000 ;
        RECT 2592.940 1495.720 2602.680 1496.000 ;
        RECT 2603.520 1495.720 2612.800 1496.000 ;
        RECT 2613.640 1495.720 2623.380 1496.000 ;
        RECT 2624.220 1495.720 2633.500 1496.000 ;
        RECT 2634.340 1495.720 2644.080 1496.000 ;
        RECT 2644.920 1495.720 2646.470 1496.000 ;
        RECT 1550.030 404.280 2646.470 1495.720 ;
        RECT 1550.030 404.000 1550.660 404.280 ;
        RECT 1551.500 404.000 1552.500 404.280 ;
        RECT 1553.340 404.000 1554.800 404.280 ;
        RECT 1555.640 404.000 1557.100 404.280 ;
        RECT 1557.940 404.000 1559.400 404.280 ;
        RECT 1560.240 404.000 1561.700 404.280 ;
        RECT 1562.540 404.000 1564.000 404.280 ;
        RECT 1564.840 404.000 1566.300 404.280 ;
        RECT 1567.140 404.000 1568.600 404.280 ;
        RECT 1569.440 404.000 1570.440 404.280 ;
        RECT 1571.280 404.000 1572.740 404.280 ;
        RECT 1573.580 404.000 1575.040 404.280 ;
        RECT 1575.880 404.000 1577.340 404.280 ;
        RECT 1578.180 404.000 1579.640 404.280 ;
        RECT 1580.480 404.000 1581.940 404.280 ;
        RECT 1582.780 404.000 1584.240 404.280 ;
        RECT 1585.080 404.000 1586.540 404.280 ;
        RECT 1587.380 404.000 1588.380 404.280 ;
        RECT 1589.220 404.000 1590.680 404.280 ;
        RECT 1591.520 404.000 1592.980 404.280 ;
        RECT 1593.820 404.000 1595.280 404.280 ;
        RECT 1596.120 404.000 1597.580 404.280 ;
        RECT 1598.420 404.000 1599.880 404.280 ;
        RECT 1600.720 404.000 1602.180 404.280 ;
        RECT 1603.020 404.000 1604.480 404.280 ;
        RECT 1605.320 404.000 1606.320 404.280 ;
        RECT 1607.160 404.000 1608.620 404.280 ;
        RECT 1609.460 404.000 1610.920 404.280 ;
        RECT 1611.760 404.000 1613.220 404.280 ;
        RECT 1614.060 404.000 1615.520 404.280 ;
        RECT 1616.360 404.000 1617.820 404.280 ;
        RECT 1618.660 404.000 1620.120 404.280 ;
        RECT 1620.960 404.000 1622.420 404.280 ;
        RECT 1623.260 404.000 1624.720 404.280 ;
        RECT 1625.560 404.000 1626.560 404.280 ;
        RECT 1627.400 404.000 1628.860 404.280 ;
        RECT 1629.700 404.000 1631.160 404.280 ;
        RECT 1632.000 404.000 1633.460 404.280 ;
        RECT 1634.300 404.000 1635.760 404.280 ;
        RECT 1636.600 404.000 1638.060 404.280 ;
        RECT 1638.900 404.000 1640.360 404.280 ;
        RECT 1641.200 404.000 1642.660 404.280 ;
        RECT 1643.500 404.000 1644.500 404.280 ;
        RECT 1645.340 404.000 1646.800 404.280 ;
        RECT 1647.640 404.000 1649.100 404.280 ;
        RECT 1649.940 404.000 1651.400 404.280 ;
        RECT 1652.240 404.000 1653.700 404.280 ;
        RECT 1654.540 404.000 1656.000 404.280 ;
        RECT 1656.840 404.000 1658.300 404.280 ;
        RECT 1659.140 404.000 1660.600 404.280 ;
        RECT 1661.440 404.000 1662.440 404.280 ;
        RECT 1663.280 404.000 1664.740 404.280 ;
        RECT 1665.580 404.000 1667.040 404.280 ;
        RECT 1667.880 404.000 1669.340 404.280 ;
        RECT 1670.180 404.000 1671.640 404.280 ;
        RECT 1672.480 404.000 1673.940 404.280 ;
        RECT 1674.780 404.000 1676.240 404.280 ;
        RECT 1677.080 404.000 1678.540 404.280 ;
        RECT 1679.380 404.000 1680.840 404.280 ;
        RECT 1681.680 404.000 1682.680 404.280 ;
        RECT 1683.520 404.000 1684.980 404.280 ;
        RECT 1685.820 404.000 1687.280 404.280 ;
        RECT 1688.120 404.000 1689.580 404.280 ;
        RECT 1690.420 404.000 1691.880 404.280 ;
        RECT 1692.720 404.000 1694.180 404.280 ;
        RECT 1695.020 404.000 1696.480 404.280 ;
        RECT 1697.320 404.000 1698.780 404.280 ;
        RECT 1699.620 404.000 1700.620 404.280 ;
        RECT 1701.460 404.000 1702.920 404.280 ;
        RECT 1703.760 404.000 1705.220 404.280 ;
        RECT 1706.060 404.000 1707.520 404.280 ;
        RECT 1708.360 404.000 1709.820 404.280 ;
        RECT 1710.660 404.000 1712.120 404.280 ;
        RECT 1712.960 404.000 1714.420 404.280 ;
        RECT 1715.260 404.000 1716.720 404.280 ;
        RECT 1717.560 404.000 1718.560 404.280 ;
        RECT 1719.400 404.000 1720.860 404.280 ;
        RECT 1721.700 404.000 1723.160 404.280 ;
        RECT 1724.000 404.000 1725.460 404.280 ;
        RECT 1726.300 404.000 1727.760 404.280 ;
        RECT 1728.600 404.000 1730.060 404.280 ;
        RECT 1730.900 404.000 1732.360 404.280 ;
        RECT 1733.200 404.000 1734.660 404.280 ;
        RECT 1735.500 404.000 1736.960 404.280 ;
        RECT 1737.800 404.000 1738.800 404.280 ;
        RECT 1739.640 404.000 1741.100 404.280 ;
        RECT 1741.940 404.000 1743.400 404.280 ;
        RECT 1744.240 404.000 1745.700 404.280 ;
        RECT 1746.540 404.000 1748.000 404.280 ;
        RECT 1748.840 404.000 1750.300 404.280 ;
        RECT 1751.140 404.000 1752.600 404.280 ;
        RECT 1753.440 404.000 1754.900 404.280 ;
        RECT 1755.740 404.000 1756.740 404.280 ;
        RECT 1757.580 404.000 1759.040 404.280 ;
        RECT 1759.880 404.000 1761.340 404.280 ;
        RECT 1762.180 404.000 1763.640 404.280 ;
        RECT 1764.480 404.000 1765.940 404.280 ;
        RECT 1766.780 404.000 1768.240 404.280 ;
        RECT 1769.080 404.000 1770.540 404.280 ;
        RECT 1771.380 404.000 1772.840 404.280 ;
        RECT 1773.680 404.000 1774.680 404.280 ;
        RECT 1775.520 404.000 1776.980 404.280 ;
        RECT 1777.820 404.000 1779.280 404.280 ;
        RECT 1780.120 404.000 1781.580 404.280 ;
        RECT 1782.420 404.000 1783.880 404.280 ;
        RECT 1784.720 404.000 1786.180 404.280 ;
        RECT 1787.020 404.000 1788.480 404.280 ;
        RECT 1789.320 404.000 1790.780 404.280 ;
        RECT 1791.620 404.000 1792.620 404.280 ;
        RECT 1793.460 404.000 1794.920 404.280 ;
        RECT 1795.760 404.000 1797.220 404.280 ;
        RECT 1798.060 404.000 1799.520 404.280 ;
        RECT 1800.360 404.000 1801.820 404.280 ;
        RECT 1802.660 404.000 1804.120 404.280 ;
        RECT 1804.960 404.000 1806.420 404.280 ;
        RECT 1807.260 404.000 1808.720 404.280 ;
        RECT 1809.560 404.000 1811.020 404.280 ;
        RECT 1811.860 404.000 1812.860 404.280 ;
        RECT 1813.700 404.000 1815.160 404.280 ;
        RECT 1816.000 404.000 1817.460 404.280 ;
        RECT 1818.300 404.000 1819.760 404.280 ;
        RECT 1820.600 404.000 1822.060 404.280 ;
        RECT 1822.900 404.000 1824.360 404.280 ;
        RECT 1825.200 404.000 1826.660 404.280 ;
        RECT 1827.500 404.000 1828.960 404.280 ;
        RECT 1829.800 404.000 1830.800 404.280 ;
        RECT 1831.640 404.000 1833.100 404.280 ;
        RECT 1833.940 404.000 1835.400 404.280 ;
        RECT 1836.240 404.000 1837.700 404.280 ;
        RECT 1838.540 404.000 1840.000 404.280 ;
        RECT 1840.840 404.000 1842.300 404.280 ;
        RECT 1843.140 404.000 1844.600 404.280 ;
        RECT 1845.440 404.000 1846.900 404.280 ;
        RECT 1847.740 404.000 1848.740 404.280 ;
        RECT 1849.580 404.000 1851.040 404.280 ;
        RECT 1851.880 404.000 1853.340 404.280 ;
        RECT 1854.180 404.000 1855.640 404.280 ;
        RECT 1856.480 404.000 1857.940 404.280 ;
        RECT 1858.780 404.000 1860.240 404.280 ;
        RECT 1861.080 404.000 1862.540 404.280 ;
        RECT 1863.380 404.000 1864.840 404.280 ;
        RECT 1865.680 404.000 1867.140 404.280 ;
        RECT 1867.980 404.000 1868.980 404.280 ;
        RECT 1869.820 404.000 1871.280 404.280 ;
        RECT 1872.120 404.000 1873.580 404.280 ;
        RECT 1874.420 404.000 1875.880 404.280 ;
        RECT 1876.720 404.000 1878.180 404.280 ;
        RECT 1879.020 404.000 1880.480 404.280 ;
        RECT 1881.320 404.000 1882.780 404.280 ;
        RECT 1883.620 404.000 1885.080 404.280 ;
        RECT 1885.920 404.000 1886.920 404.280 ;
        RECT 1887.760 404.000 1889.220 404.280 ;
        RECT 1890.060 404.000 1891.520 404.280 ;
        RECT 1892.360 404.000 1893.820 404.280 ;
        RECT 1894.660 404.000 1896.120 404.280 ;
        RECT 1896.960 404.000 1898.420 404.280 ;
        RECT 1899.260 404.000 1900.720 404.280 ;
        RECT 1901.560 404.000 1903.020 404.280 ;
        RECT 1903.860 404.000 1904.860 404.280 ;
        RECT 1905.700 404.000 1907.160 404.280 ;
        RECT 1908.000 404.000 1909.460 404.280 ;
        RECT 1910.300 404.000 1911.760 404.280 ;
        RECT 1912.600 404.000 1914.060 404.280 ;
        RECT 1914.900 404.000 1916.360 404.280 ;
        RECT 1917.200 404.000 1918.660 404.280 ;
        RECT 1919.500 404.000 1920.960 404.280 ;
        RECT 1921.800 404.000 1923.260 404.280 ;
        RECT 1924.100 404.000 1925.100 404.280 ;
        RECT 1925.940 404.000 1927.400 404.280 ;
        RECT 1928.240 404.000 1929.700 404.280 ;
        RECT 1930.540 404.000 1932.000 404.280 ;
        RECT 1932.840 404.000 1934.300 404.280 ;
        RECT 1935.140 404.000 1936.600 404.280 ;
        RECT 1937.440 404.000 1938.900 404.280 ;
        RECT 1939.740 404.000 1941.200 404.280 ;
        RECT 1942.040 404.000 1943.040 404.280 ;
        RECT 1943.880 404.000 1945.340 404.280 ;
        RECT 1946.180 404.000 1947.640 404.280 ;
        RECT 1948.480 404.000 1949.940 404.280 ;
        RECT 1950.780 404.000 1952.240 404.280 ;
        RECT 1953.080 404.000 1954.540 404.280 ;
        RECT 1955.380 404.000 1956.840 404.280 ;
        RECT 1957.680 404.000 1959.140 404.280 ;
        RECT 1959.980 404.000 1960.980 404.280 ;
        RECT 1961.820 404.000 1963.280 404.280 ;
        RECT 1964.120 404.000 1965.580 404.280 ;
        RECT 1966.420 404.000 1967.880 404.280 ;
        RECT 1968.720 404.000 1970.180 404.280 ;
        RECT 1971.020 404.000 1972.480 404.280 ;
        RECT 1973.320 404.000 1974.780 404.280 ;
        RECT 1975.620 404.000 1977.080 404.280 ;
        RECT 1977.920 404.000 1979.380 404.280 ;
        RECT 1980.220 404.000 1981.220 404.280 ;
        RECT 1982.060 404.000 1983.520 404.280 ;
        RECT 1984.360 404.000 1985.820 404.280 ;
        RECT 1986.660 404.000 1988.120 404.280 ;
        RECT 1988.960 404.000 1990.420 404.280 ;
        RECT 1991.260 404.000 1992.720 404.280 ;
        RECT 1993.560 404.000 1995.020 404.280 ;
        RECT 1995.860 404.000 1997.320 404.280 ;
        RECT 1998.160 404.000 1999.160 404.280 ;
        RECT 2000.000 404.000 2001.460 404.280 ;
        RECT 2002.300 404.000 2003.760 404.280 ;
        RECT 2004.600 404.000 2006.060 404.280 ;
        RECT 2006.900 404.000 2008.360 404.280 ;
        RECT 2009.200 404.000 2010.660 404.280 ;
        RECT 2011.500 404.000 2012.960 404.280 ;
        RECT 2013.800 404.000 2015.260 404.280 ;
        RECT 2016.100 404.000 2017.100 404.280 ;
        RECT 2017.940 404.000 2019.400 404.280 ;
        RECT 2020.240 404.000 2021.700 404.280 ;
        RECT 2022.540 404.000 2024.000 404.280 ;
        RECT 2024.840 404.000 2026.300 404.280 ;
        RECT 2027.140 404.000 2028.600 404.280 ;
        RECT 2029.440 404.000 2030.900 404.280 ;
        RECT 2031.740 404.000 2033.200 404.280 ;
        RECT 2034.040 404.000 2035.040 404.280 ;
        RECT 2035.880 404.000 2037.340 404.280 ;
        RECT 2038.180 404.000 2039.640 404.280 ;
        RECT 2040.480 404.000 2041.940 404.280 ;
        RECT 2042.780 404.000 2044.240 404.280 ;
        RECT 2045.080 404.000 2046.540 404.280 ;
        RECT 2047.380 404.000 2048.840 404.280 ;
        RECT 2049.680 404.000 2051.140 404.280 ;
        RECT 2051.980 404.000 2053.440 404.280 ;
        RECT 2054.280 404.000 2055.280 404.280 ;
        RECT 2056.120 404.000 2057.580 404.280 ;
        RECT 2058.420 404.000 2059.880 404.280 ;
        RECT 2060.720 404.000 2062.180 404.280 ;
        RECT 2063.020 404.000 2064.480 404.280 ;
        RECT 2065.320 404.000 2066.780 404.280 ;
        RECT 2067.620 404.000 2069.080 404.280 ;
        RECT 2069.920 404.000 2071.380 404.280 ;
        RECT 2072.220 404.000 2073.220 404.280 ;
        RECT 2074.060 404.000 2075.520 404.280 ;
        RECT 2076.360 404.000 2077.820 404.280 ;
        RECT 2078.660 404.000 2080.120 404.280 ;
        RECT 2080.960 404.000 2082.420 404.280 ;
        RECT 2083.260 404.000 2084.720 404.280 ;
        RECT 2085.560 404.000 2087.020 404.280 ;
        RECT 2087.860 404.000 2089.320 404.280 ;
        RECT 2090.160 404.000 2091.160 404.280 ;
        RECT 2092.000 404.000 2093.460 404.280 ;
        RECT 2094.300 404.000 2095.760 404.280 ;
        RECT 2096.600 404.000 2098.060 404.280 ;
        RECT 2098.900 404.000 2100.360 404.280 ;
        RECT 2101.200 404.000 2102.660 404.280 ;
        RECT 2103.500 404.000 2104.960 404.280 ;
        RECT 2105.800 404.000 2107.260 404.280 ;
        RECT 2108.100 404.000 2109.560 404.280 ;
        RECT 2110.400 404.000 2111.400 404.280 ;
        RECT 2112.240 404.000 2113.700 404.280 ;
        RECT 2114.540 404.000 2116.000 404.280 ;
        RECT 2116.840 404.000 2118.300 404.280 ;
        RECT 2119.140 404.000 2120.600 404.280 ;
        RECT 2121.440 404.000 2122.900 404.280 ;
        RECT 2123.740 404.000 2125.200 404.280 ;
        RECT 2126.040 404.000 2127.500 404.280 ;
        RECT 2128.340 404.000 2129.340 404.280 ;
        RECT 2130.180 404.000 2131.640 404.280 ;
        RECT 2132.480 404.000 2133.940 404.280 ;
        RECT 2134.780 404.000 2136.240 404.280 ;
        RECT 2137.080 404.000 2138.540 404.280 ;
        RECT 2139.380 404.000 2140.840 404.280 ;
        RECT 2141.680 404.000 2143.140 404.280 ;
        RECT 2143.980 404.000 2145.440 404.280 ;
        RECT 2146.280 404.000 2147.280 404.280 ;
        RECT 2148.120 404.000 2149.580 404.280 ;
        RECT 2150.420 404.000 2151.880 404.280 ;
        RECT 2152.720 404.000 2154.180 404.280 ;
        RECT 2155.020 404.000 2156.480 404.280 ;
        RECT 2157.320 404.000 2158.780 404.280 ;
        RECT 2159.620 404.000 2161.080 404.280 ;
        RECT 2161.920 404.000 2163.380 404.280 ;
        RECT 2164.220 404.000 2165.680 404.280 ;
        RECT 2166.520 404.000 2167.520 404.280 ;
        RECT 2168.360 404.000 2169.820 404.280 ;
        RECT 2170.660 404.000 2172.120 404.280 ;
        RECT 2172.960 404.000 2174.420 404.280 ;
        RECT 2175.260 404.000 2176.720 404.280 ;
        RECT 2177.560 404.000 2179.020 404.280 ;
        RECT 2179.860 404.000 2181.320 404.280 ;
        RECT 2182.160 404.000 2183.620 404.280 ;
        RECT 2184.460 404.000 2185.460 404.280 ;
        RECT 2186.300 404.000 2187.760 404.280 ;
        RECT 2188.600 404.000 2190.060 404.280 ;
        RECT 2190.900 404.000 2192.360 404.280 ;
        RECT 2193.200 404.000 2194.660 404.280 ;
        RECT 2195.500 404.000 2196.960 404.280 ;
        RECT 2197.800 404.000 2199.260 404.280 ;
        RECT 2200.100 404.000 2201.560 404.280 ;
        RECT 2202.400 404.000 2203.400 404.280 ;
        RECT 2204.240 404.000 2205.700 404.280 ;
        RECT 2206.540 404.000 2208.000 404.280 ;
        RECT 2208.840 404.000 2210.300 404.280 ;
        RECT 2211.140 404.000 2212.600 404.280 ;
        RECT 2213.440 404.000 2214.900 404.280 ;
        RECT 2215.740 404.000 2217.200 404.280 ;
        RECT 2218.040 404.000 2219.500 404.280 ;
        RECT 2220.340 404.000 2221.340 404.280 ;
        RECT 2222.180 404.000 2223.640 404.280 ;
        RECT 2224.480 404.000 2225.940 404.280 ;
        RECT 2226.780 404.000 2228.240 404.280 ;
        RECT 2229.080 404.000 2230.540 404.280 ;
        RECT 2231.380 404.000 2232.840 404.280 ;
        RECT 2233.680 404.000 2235.140 404.280 ;
        RECT 2235.980 404.000 2237.440 404.280 ;
        RECT 2238.280 404.000 2239.740 404.280 ;
        RECT 2240.580 404.000 2241.580 404.280 ;
        RECT 2242.420 404.000 2243.880 404.280 ;
        RECT 2244.720 404.000 2246.180 404.280 ;
        RECT 2247.020 404.000 2248.480 404.280 ;
        RECT 2249.320 404.000 2250.780 404.280 ;
        RECT 2251.620 404.000 2253.080 404.280 ;
        RECT 2253.920 404.000 2255.380 404.280 ;
        RECT 2256.220 404.000 2257.680 404.280 ;
        RECT 2258.520 404.000 2259.520 404.280 ;
        RECT 2260.360 404.000 2261.820 404.280 ;
        RECT 2262.660 404.000 2264.120 404.280 ;
        RECT 2264.960 404.000 2266.420 404.280 ;
        RECT 2267.260 404.000 2268.720 404.280 ;
        RECT 2269.560 404.000 2271.020 404.280 ;
        RECT 2271.860 404.000 2273.320 404.280 ;
        RECT 2274.160 404.000 2275.620 404.280 ;
        RECT 2276.460 404.000 2277.460 404.280 ;
        RECT 2278.300 404.000 2279.760 404.280 ;
        RECT 2280.600 404.000 2282.060 404.280 ;
        RECT 2282.900 404.000 2284.360 404.280 ;
        RECT 2285.200 404.000 2286.660 404.280 ;
        RECT 2287.500 404.000 2288.960 404.280 ;
        RECT 2289.800 404.000 2291.260 404.280 ;
        RECT 2292.100 404.000 2293.560 404.280 ;
        RECT 2294.400 404.000 2295.860 404.280 ;
        RECT 2296.700 404.000 2297.700 404.280 ;
        RECT 2298.540 404.000 2300.000 404.280 ;
        RECT 2300.840 404.000 2302.300 404.280 ;
        RECT 2303.140 404.000 2304.600 404.280 ;
        RECT 2305.440 404.000 2306.900 404.280 ;
        RECT 2307.740 404.000 2309.200 404.280 ;
        RECT 2310.040 404.000 2311.500 404.280 ;
        RECT 2312.340 404.000 2313.800 404.280 ;
        RECT 2314.640 404.000 2315.640 404.280 ;
        RECT 2316.480 404.000 2317.940 404.280 ;
        RECT 2318.780 404.000 2320.240 404.280 ;
        RECT 2321.080 404.000 2322.540 404.280 ;
        RECT 2323.380 404.000 2324.840 404.280 ;
        RECT 2325.680 404.000 2327.140 404.280 ;
        RECT 2327.980 404.000 2329.440 404.280 ;
        RECT 2330.280 404.000 2331.740 404.280 ;
        RECT 2332.580 404.000 2333.580 404.280 ;
        RECT 2334.420 404.000 2335.880 404.280 ;
        RECT 2336.720 404.000 2338.180 404.280 ;
        RECT 2339.020 404.000 2340.480 404.280 ;
        RECT 2341.320 404.000 2342.780 404.280 ;
        RECT 2343.620 404.000 2345.080 404.280 ;
        RECT 2345.920 404.000 2347.380 404.280 ;
        RECT 2348.220 404.000 2349.680 404.280 ;
        RECT 2350.520 404.000 2351.980 404.280 ;
        RECT 2352.820 404.000 2353.820 404.280 ;
        RECT 2354.660 404.000 2356.120 404.280 ;
        RECT 2356.960 404.000 2358.420 404.280 ;
        RECT 2359.260 404.000 2360.720 404.280 ;
        RECT 2361.560 404.000 2363.020 404.280 ;
        RECT 2363.860 404.000 2365.320 404.280 ;
        RECT 2366.160 404.000 2367.620 404.280 ;
        RECT 2368.460 404.000 2369.920 404.280 ;
        RECT 2370.760 404.000 2371.760 404.280 ;
        RECT 2372.600 404.000 2374.060 404.280 ;
        RECT 2374.900 404.000 2376.360 404.280 ;
        RECT 2377.200 404.000 2378.660 404.280 ;
        RECT 2379.500 404.000 2380.960 404.280 ;
        RECT 2381.800 404.000 2383.260 404.280 ;
        RECT 2384.100 404.000 2385.560 404.280 ;
        RECT 2386.400 404.000 2387.860 404.280 ;
        RECT 2388.700 404.000 2389.700 404.280 ;
        RECT 2390.540 404.000 2392.000 404.280 ;
        RECT 2392.840 404.000 2394.300 404.280 ;
        RECT 2395.140 404.000 2396.600 404.280 ;
        RECT 2397.440 404.000 2398.900 404.280 ;
        RECT 2399.740 404.000 2401.200 404.280 ;
        RECT 2402.040 404.000 2403.500 404.280 ;
        RECT 2404.340 404.000 2405.800 404.280 ;
        RECT 2406.640 404.000 2408.100 404.280 ;
        RECT 2408.940 404.000 2409.940 404.280 ;
        RECT 2410.780 404.000 2412.240 404.280 ;
        RECT 2413.080 404.000 2414.540 404.280 ;
        RECT 2415.380 404.000 2416.840 404.280 ;
        RECT 2417.680 404.000 2419.140 404.280 ;
        RECT 2419.980 404.000 2421.440 404.280 ;
        RECT 2422.280 404.000 2423.740 404.280 ;
        RECT 2424.580 404.000 2426.040 404.280 ;
        RECT 2426.880 404.000 2427.880 404.280 ;
        RECT 2428.720 404.000 2430.180 404.280 ;
        RECT 2431.020 404.000 2432.480 404.280 ;
        RECT 2433.320 404.000 2434.780 404.280 ;
        RECT 2435.620 404.000 2437.080 404.280 ;
        RECT 2437.920 404.000 2439.380 404.280 ;
        RECT 2440.220 404.000 2441.680 404.280 ;
        RECT 2442.520 404.000 2443.980 404.280 ;
        RECT 2444.820 404.000 2445.820 404.280 ;
        RECT 2446.660 404.000 2448.120 404.280 ;
        RECT 2448.960 404.000 2450.420 404.280 ;
        RECT 2451.260 404.000 2452.720 404.280 ;
        RECT 2453.560 404.000 2455.020 404.280 ;
        RECT 2455.860 404.000 2457.320 404.280 ;
        RECT 2458.160 404.000 2459.620 404.280 ;
        RECT 2460.460 404.000 2461.920 404.280 ;
        RECT 2462.760 404.000 2463.760 404.280 ;
        RECT 2464.600 404.000 2466.060 404.280 ;
        RECT 2466.900 404.000 2468.360 404.280 ;
        RECT 2469.200 404.000 2470.660 404.280 ;
        RECT 2471.500 404.000 2472.960 404.280 ;
        RECT 2473.800 404.000 2475.260 404.280 ;
        RECT 2476.100 404.000 2477.560 404.280 ;
        RECT 2478.400 404.000 2479.860 404.280 ;
        RECT 2480.700 404.000 2482.160 404.280 ;
        RECT 2483.000 404.000 2484.000 404.280 ;
        RECT 2484.840 404.000 2486.300 404.280 ;
        RECT 2487.140 404.000 2488.600 404.280 ;
        RECT 2489.440 404.000 2490.900 404.280 ;
        RECT 2491.740 404.000 2493.200 404.280 ;
        RECT 2494.040 404.000 2495.500 404.280 ;
        RECT 2496.340 404.000 2497.800 404.280 ;
        RECT 2498.640 404.000 2500.100 404.280 ;
        RECT 2500.940 404.000 2501.940 404.280 ;
        RECT 2502.780 404.000 2504.240 404.280 ;
        RECT 2505.080 404.000 2506.540 404.280 ;
        RECT 2507.380 404.000 2508.840 404.280 ;
        RECT 2509.680 404.000 2511.140 404.280 ;
        RECT 2511.980 404.000 2513.440 404.280 ;
        RECT 2514.280 404.000 2515.740 404.280 ;
        RECT 2516.580 404.000 2518.040 404.280 ;
        RECT 2518.880 404.000 2519.880 404.280 ;
        RECT 2520.720 404.000 2522.180 404.280 ;
        RECT 2523.020 404.000 2524.480 404.280 ;
        RECT 2525.320 404.000 2526.780 404.280 ;
        RECT 2527.620 404.000 2529.080 404.280 ;
        RECT 2529.920 404.000 2531.380 404.280 ;
        RECT 2532.220 404.000 2533.680 404.280 ;
        RECT 2534.520 404.000 2535.980 404.280 ;
        RECT 2536.820 404.000 2538.280 404.280 ;
        RECT 2539.120 404.000 2540.120 404.280 ;
        RECT 2540.960 404.000 2542.420 404.280 ;
        RECT 2543.260 404.000 2544.720 404.280 ;
        RECT 2545.560 404.000 2547.020 404.280 ;
        RECT 2547.860 404.000 2549.320 404.280 ;
        RECT 2550.160 404.000 2551.620 404.280 ;
        RECT 2552.460 404.000 2553.920 404.280 ;
        RECT 2554.760 404.000 2556.220 404.280 ;
        RECT 2557.060 404.000 2558.060 404.280 ;
        RECT 2558.900 404.000 2560.360 404.280 ;
        RECT 2561.200 404.000 2562.660 404.280 ;
        RECT 2563.500 404.000 2564.960 404.280 ;
        RECT 2565.800 404.000 2567.260 404.280 ;
        RECT 2568.100 404.000 2569.560 404.280 ;
        RECT 2570.400 404.000 2571.860 404.280 ;
        RECT 2572.700 404.000 2574.160 404.280 ;
        RECT 2575.000 404.000 2576.000 404.280 ;
        RECT 2576.840 404.000 2578.300 404.280 ;
        RECT 2579.140 404.000 2580.600 404.280 ;
        RECT 2581.440 404.000 2582.900 404.280 ;
        RECT 2583.740 404.000 2585.200 404.280 ;
        RECT 2586.040 404.000 2587.500 404.280 ;
        RECT 2588.340 404.000 2589.800 404.280 ;
        RECT 2590.640 404.000 2592.100 404.280 ;
        RECT 2592.940 404.000 2594.400 404.280 ;
        RECT 2595.240 404.000 2596.240 404.280 ;
        RECT 2597.080 404.000 2598.540 404.280 ;
        RECT 2599.380 404.000 2600.840 404.280 ;
        RECT 2601.680 404.000 2603.140 404.280 ;
        RECT 2603.980 404.000 2605.440 404.280 ;
        RECT 2606.280 404.000 2607.740 404.280 ;
        RECT 2608.580 404.000 2610.040 404.280 ;
        RECT 2610.880 404.000 2612.340 404.280 ;
        RECT 2613.180 404.000 2614.180 404.280 ;
        RECT 2615.020 404.000 2616.480 404.280 ;
        RECT 2617.320 404.000 2618.780 404.280 ;
        RECT 2619.620 404.000 2621.080 404.280 ;
        RECT 2621.920 404.000 2623.380 404.280 ;
        RECT 2624.220 404.000 2625.680 404.280 ;
        RECT 2626.520 404.000 2627.980 404.280 ;
        RECT 2628.820 404.000 2630.280 404.280 ;
        RECT 2631.120 404.000 2632.120 404.280 ;
        RECT 2632.960 404.000 2634.420 404.280 ;
        RECT 2635.260 404.000 2636.720 404.280 ;
        RECT 2637.560 404.000 2639.020 404.280 ;
        RECT 2639.860 404.000 2641.320 404.280 ;
        RECT 2642.160 404.000 2643.620 404.280 ;
        RECT 2644.460 404.000 2645.920 404.280 ;
      LAYER met2 ;
        RECT 1550.940 400.000 1551.220 404.000 ;
        RECT 1552.780 400.000 1553.060 404.000 ;
        RECT 1555.080 400.000 1555.360 404.000 ;
        RECT 1557.380 400.000 1557.660 404.000 ;
        RECT 1559.680 400.000 1559.960 404.000 ;
        RECT 1561.980 400.000 1562.260 404.000 ;
        RECT 1564.280 400.000 1564.560 404.000 ;
        RECT 1566.580 400.000 1566.860 404.000 ;
        RECT 1568.880 400.000 1569.160 404.000 ;
        RECT 1570.720 400.000 1571.000 404.000 ;
        RECT 1573.020 400.000 1573.300 404.000 ;
        RECT 1575.320 400.000 1575.600 404.000 ;
        RECT 1577.620 400.000 1577.900 404.000 ;
        RECT 1579.920 400.000 1580.200 404.000 ;
        RECT 1582.220 400.000 1582.500 404.000 ;
        RECT 1584.520 400.000 1584.800 404.000 ;
        RECT 1586.820 400.000 1587.100 404.000 ;
        RECT 1588.660 400.000 1588.940 404.000 ;
        RECT 1590.960 400.000 1591.240 404.000 ;
        RECT 1593.260 400.000 1593.540 404.000 ;
        RECT 1595.560 400.000 1595.840 404.000 ;
        RECT 1597.860 400.000 1598.140 404.000 ;
        RECT 1600.160 400.000 1600.440 404.000 ;
        RECT 1602.460 400.000 1602.740 404.000 ;
        RECT 1604.760 400.000 1605.040 404.000 ;
        RECT 1606.600 400.000 1606.880 404.000 ;
        RECT 1608.900 400.000 1609.180 404.000 ;
        RECT 1611.200 400.000 1611.480 404.000 ;
        RECT 1613.500 400.000 1613.780 404.000 ;
        RECT 1615.800 400.000 1616.080 404.000 ;
        RECT 1618.100 400.000 1618.380 404.000 ;
        RECT 1620.400 400.000 1620.680 404.000 ;
        RECT 1622.700 400.000 1622.980 404.000 ;
        RECT 1625.000 400.000 1625.280 404.000 ;
        RECT 1626.840 400.000 1627.120 404.000 ;
        RECT 1629.140 400.000 1629.420 404.000 ;
        RECT 1631.440 400.000 1631.720 404.000 ;
        RECT 1633.740 400.000 1634.020 404.000 ;
        RECT 1636.040 400.000 1636.320 404.000 ;
        RECT 1638.340 400.000 1638.620 404.000 ;
        RECT 1640.640 400.000 1640.920 404.000 ;
        RECT 1642.940 400.000 1643.220 404.000 ;
        RECT 1644.780 400.000 1645.060 404.000 ;
        RECT 1647.080 400.000 1647.360 404.000 ;
        RECT 1649.380 400.000 1649.660 404.000 ;
        RECT 1651.680 400.000 1651.960 404.000 ;
        RECT 1653.980 400.000 1654.260 404.000 ;
        RECT 1656.280 400.000 1656.560 404.000 ;
        RECT 1658.580 400.000 1658.860 404.000 ;
        RECT 1660.880 400.000 1661.160 404.000 ;
        RECT 1662.720 400.000 1663.000 404.000 ;
        RECT 1665.020 400.000 1665.300 404.000 ;
        RECT 1667.320 400.000 1667.600 404.000 ;
        RECT 1669.620 400.000 1669.900 404.000 ;
        RECT 1671.920 400.000 1672.200 404.000 ;
        RECT 1674.220 400.000 1674.500 404.000 ;
        RECT 1676.520 400.000 1676.800 404.000 ;
        RECT 1678.820 400.000 1679.100 404.000 ;
        RECT 1681.120 400.000 1681.400 404.000 ;
        RECT 1682.960 400.000 1683.240 404.000 ;
        RECT 1685.260 400.000 1685.540 404.000 ;
        RECT 1687.560 400.000 1687.840 404.000 ;
        RECT 1689.860 400.000 1690.140 404.000 ;
        RECT 1692.160 400.000 1692.440 404.000 ;
        RECT 1694.460 400.000 1694.740 404.000 ;
        RECT 1696.760 400.000 1697.040 404.000 ;
        RECT 1699.060 400.000 1699.340 404.000 ;
        RECT 1700.900 400.000 1701.180 404.000 ;
        RECT 1703.200 400.000 1703.480 404.000 ;
        RECT 1705.500 400.000 1705.780 404.000 ;
        RECT 1707.800 400.000 1708.080 404.000 ;
        RECT 1710.100 400.000 1710.380 404.000 ;
        RECT 1712.400 400.000 1712.680 404.000 ;
        RECT 1714.700 400.000 1714.980 404.000 ;
        RECT 1717.000 400.000 1717.280 404.000 ;
        RECT 1718.840 400.000 1719.120 404.000 ;
        RECT 1721.140 400.000 1721.420 404.000 ;
        RECT 1723.440 400.000 1723.720 404.000 ;
        RECT 1725.740 400.000 1726.020 404.000 ;
        RECT 1728.040 400.000 1728.320 404.000 ;
        RECT 1730.340 400.000 1730.620 404.000 ;
        RECT 1732.640 400.000 1732.920 404.000 ;
        RECT 1734.940 400.000 1735.220 404.000 ;
        RECT 1737.240 400.000 1737.520 404.000 ;
        RECT 1739.080 400.000 1739.360 404.000 ;
        RECT 1741.380 400.000 1741.660 404.000 ;
        RECT 1743.680 400.000 1743.960 404.000 ;
        RECT 1745.980 400.000 1746.260 404.000 ;
        RECT 1748.280 400.000 1748.560 404.000 ;
        RECT 1750.580 400.000 1750.860 404.000 ;
        RECT 1752.880 400.000 1753.160 404.000 ;
        RECT 1755.180 400.000 1755.460 404.000 ;
        RECT 1757.020 400.000 1757.300 404.000 ;
        RECT 1759.320 400.000 1759.600 404.000 ;
        RECT 1761.620 400.000 1761.900 404.000 ;
        RECT 1763.920 400.000 1764.200 404.000 ;
        RECT 1766.220 400.000 1766.500 404.000 ;
        RECT 1768.520 400.000 1768.800 404.000 ;
        RECT 1770.820 400.000 1771.100 404.000 ;
        RECT 1773.120 400.000 1773.400 404.000 ;
        RECT 1774.960 400.000 1775.240 404.000 ;
        RECT 1777.260 400.000 1777.540 404.000 ;
        RECT 1779.560 400.000 1779.840 404.000 ;
        RECT 1781.860 400.000 1782.140 404.000 ;
        RECT 1784.160 400.000 1784.440 404.000 ;
        RECT 1786.460 400.000 1786.740 404.000 ;
        RECT 1788.760 400.000 1789.040 404.000 ;
        RECT 1791.060 400.000 1791.340 404.000 ;
        RECT 1792.900 400.000 1793.180 404.000 ;
        RECT 1795.200 400.000 1795.480 404.000 ;
        RECT 1797.500 400.000 1797.780 404.000 ;
        RECT 1799.800 400.000 1800.080 404.000 ;
        RECT 1802.100 400.000 1802.380 404.000 ;
        RECT 1804.400 400.000 1804.680 404.000 ;
        RECT 1806.700 400.000 1806.980 404.000 ;
        RECT 1809.000 400.000 1809.280 404.000 ;
        RECT 1811.300 400.000 1811.580 404.000 ;
        RECT 1813.140 400.000 1813.420 404.000 ;
        RECT 1815.440 400.000 1815.720 404.000 ;
        RECT 1817.740 400.000 1818.020 404.000 ;
        RECT 1820.040 400.000 1820.320 404.000 ;
        RECT 1822.340 400.000 1822.620 404.000 ;
        RECT 1824.640 400.000 1824.920 404.000 ;
        RECT 1826.940 400.000 1827.220 404.000 ;
        RECT 1829.240 400.000 1829.520 404.000 ;
        RECT 1831.080 400.000 1831.360 404.000 ;
        RECT 1833.380 400.000 1833.660 404.000 ;
        RECT 1835.680 400.000 1835.960 404.000 ;
        RECT 1837.980 400.000 1838.260 404.000 ;
        RECT 1840.280 400.000 1840.560 404.000 ;
        RECT 1842.580 400.000 1842.860 404.000 ;
        RECT 1844.880 400.000 1845.160 404.000 ;
        RECT 1847.180 400.000 1847.460 404.000 ;
        RECT 1849.020 400.000 1849.300 404.000 ;
        RECT 1851.320 400.000 1851.600 404.000 ;
        RECT 1853.620 400.000 1853.900 404.000 ;
        RECT 1855.920 400.000 1856.200 404.000 ;
        RECT 1858.220 400.000 1858.500 404.000 ;
        RECT 1860.520 400.000 1860.800 404.000 ;
        RECT 1862.820 400.000 1863.100 404.000 ;
        RECT 1865.120 400.000 1865.400 404.000 ;
        RECT 1867.420 400.000 1867.700 404.000 ;
        RECT 1869.260 400.000 1869.540 404.000 ;
        RECT 1871.560 400.000 1871.840 404.000 ;
        RECT 1873.860 400.000 1874.140 404.000 ;
        RECT 1876.160 400.000 1876.440 404.000 ;
        RECT 1878.460 400.000 1878.740 404.000 ;
        RECT 1880.760 400.000 1881.040 404.000 ;
        RECT 1883.060 400.000 1883.340 404.000 ;
        RECT 1885.360 400.000 1885.640 404.000 ;
        RECT 1887.200 400.000 1887.480 404.000 ;
        RECT 1889.500 400.000 1889.780 404.000 ;
        RECT 1891.800 400.000 1892.080 404.000 ;
        RECT 1894.100 400.000 1894.380 404.000 ;
        RECT 1896.400 400.000 1896.680 404.000 ;
        RECT 1898.700 400.000 1898.980 404.000 ;
        RECT 1901.000 400.000 1901.280 404.000 ;
        RECT 1903.300 400.000 1903.580 404.000 ;
        RECT 1905.140 400.000 1905.420 404.000 ;
        RECT 1907.440 400.000 1907.720 404.000 ;
        RECT 1909.740 400.000 1910.020 404.000 ;
        RECT 1912.040 400.000 1912.320 404.000 ;
        RECT 1914.340 400.000 1914.620 404.000 ;
        RECT 1916.640 400.000 1916.920 404.000 ;
        RECT 1918.940 400.000 1919.220 404.000 ;
        RECT 1921.240 400.000 1921.520 404.000 ;
        RECT 1923.540 400.000 1923.820 404.000 ;
        RECT 1925.380 400.000 1925.660 404.000 ;
        RECT 1927.680 400.000 1927.960 404.000 ;
        RECT 1929.980 400.000 1930.260 404.000 ;
        RECT 1932.280 400.000 1932.560 404.000 ;
        RECT 1934.580 400.000 1934.860 404.000 ;
        RECT 1936.880 400.000 1937.160 404.000 ;
        RECT 1939.180 400.000 1939.460 404.000 ;
        RECT 1941.480 400.000 1941.760 404.000 ;
        RECT 1943.320 400.000 1943.600 404.000 ;
        RECT 1945.620 400.000 1945.900 404.000 ;
        RECT 1947.920 400.000 1948.200 404.000 ;
        RECT 1950.220 400.000 1950.500 404.000 ;
        RECT 1952.520 400.000 1952.800 404.000 ;
        RECT 1954.820 400.000 1955.100 404.000 ;
        RECT 1957.120 400.000 1957.400 404.000 ;
        RECT 1959.420 400.000 1959.700 404.000 ;
        RECT 1961.260 400.000 1961.540 404.000 ;
        RECT 1963.560 400.000 1963.840 404.000 ;
        RECT 1965.860 400.000 1966.140 404.000 ;
        RECT 1968.160 400.000 1968.440 404.000 ;
        RECT 1970.460 400.000 1970.740 404.000 ;
        RECT 1972.760 400.000 1973.040 404.000 ;
        RECT 1975.060 400.000 1975.340 404.000 ;
        RECT 1977.360 400.000 1977.640 404.000 ;
        RECT 1979.660 400.000 1979.940 404.000 ;
        RECT 1981.500 400.000 1981.780 404.000 ;
        RECT 1983.800 400.000 1984.080 404.000 ;
        RECT 1986.100 400.000 1986.380 404.000 ;
        RECT 1988.400 400.000 1988.680 404.000 ;
        RECT 1990.700 400.000 1990.980 404.000 ;
        RECT 1993.000 400.000 1993.280 404.000 ;
        RECT 1995.300 400.000 1995.580 404.000 ;
        RECT 1997.600 400.000 1997.880 404.000 ;
        RECT 1999.440 400.000 1999.720 404.000 ;
        RECT 2001.740 400.000 2002.020 404.000 ;
        RECT 2004.040 400.000 2004.320 404.000 ;
        RECT 2006.340 400.000 2006.620 404.000 ;
        RECT 2008.640 400.000 2008.920 404.000 ;
        RECT 2010.940 400.000 2011.220 404.000 ;
        RECT 2013.240 400.000 2013.520 404.000 ;
        RECT 2015.540 400.000 2015.820 404.000 ;
        RECT 2017.380 400.000 2017.660 404.000 ;
        RECT 2019.680 400.000 2019.960 404.000 ;
        RECT 2021.980 400.000 2022.260 404.000 ;
        RECT 2024.280 400.000 2024.560 404.000 ;
        RECT 2026.580 400.000 2026.860 404.000 ;
        RECT 2028.880 400.000 2029.160 404.000 ;
        RECT 2031.180 400.000 2031.460 404.000 ;
        RECT 2033.480 400.000 2033.760 404.000 ;
        RECT 2035.320 400.000 2035.600 404.000 ;
        RECT 2037.620 400.000 2037.900 404.000 ;
        RECT 2039.920 400.000 2040.200 404.000 ;
        RECT 2042.220 400.000 2042.500 404.000 ;
        RECT 2044.520 400.000 2044.800 404.000 ;
        RECT 2046.820 400.000 2047.100 404.000 ;
        RECT 2049.120 400.000 2049.400 404.000 ;
        RECT 2051.420 400.000 2051.700 404.000 ;
        RECT 2053.720 400.000 2054.000 404.000 ;
        RECT 2055.560 400.000 2055.840 404.000 ;
        RECT 2057.860 400.000 2058.140 404.000 ;
        RECT 2060.160 400.000 2060.440 404.000 ;
        RECT 2062.460 400.000 2062.740 404.000 ;
        RECT 2064.760 400.000 2065.040 404.000 ;
        RECT 2067.060 400.000 2067.340 404.000 ;
        RECT 2069.360 400.000 2069.640 404.000 ;
        RECT 2071.660 400.000 2071.940 404.000 ;
        RECT 2073.500 400.000 2073.780 404.000 ;
        RECT 2075.800 400.000 2076.080 404.000 ;
        RECT 2078.100 400.000 2078.380 404.000 ;
        RECT 2080.400 400.000 2080.680 404.000 ;
        RECT 2082.700 400.000 2082.980 404.000 ;
        RECT 2085.000 400.000 2085.280 404.000 ;
        RECT 2087.300 400.000 2087.580 404.000 ;
        RECT 2089.600 400.000 2089.880 404.000 ;
        RECT 2091.440 400.000 2091.720 404.000 ;
        RECT 2093.740 400.000 2094.020 404.000 ;
        RECT 2096.040 400.000 2096.320 404.000 ;
        RECT 2098.340 400.000 2098.620 404.000 ;
        RECT 2100.640 400.000 2100.920 404.000 ;
        RECT 2102.940 400.000 2103.220 404.000 ;
        RECT 2105.240 400.000 2105.520 404.000 ;
        RECT 2107.540 400.000 2107.820 404.000 ;
        RECT 2109.840 400.000 2110.120 404.000 ;
        RECT 2111.680 400.000 2111.960 404.000 ;
        RECT 2113.980 400.000 2114.260 404.000 ;
        RECT 2116.280 400.000 2116.560 404.000 ;
        RECT 2118.580 400.000 2118.860 404.000 ;
        RECT 2120.880 400.000 2121.160 404.000 ;
        RECT 2123.180 400.000 2123.460 404.000 ;
        RECT 2125.480 400.000 2125.760 404.000 ;
        RECT 2127.780 400.000 2128.060 404.000 ;
        RECT 2129.620 400.000 2129.900 404.000 ;
        RECT 2131.920 400.000 2132.200 404.000 ;
        RECT 2134.220 400.000 2134.500 404.000 ;
        RECT 2136.520 400.000 2136.800 404.000 ;
        RECT 2138.820 400.000 2139.100 404.000 ;
        RECT 2141.120 400.000 2141.400 404.000 ;
        RECT 2143.420 400.000 2143.700 404.000 ;
        RECT 2145.720 400.000 2146.000 404.000 ;
        RECT 2147.560 400.000 2147.840 404.000 ;
        RECT 2149.860 400.000 2150.140 404.000 ;
        RECT 2152.160 400.000 2152.440 404.000 ;
        RECT 2154.460 400.000 2154.740 404.000 ;
        RECT 2156.760 400.000 2157.040 404.000 ;
        RECT 2159.060 400.000 2159.340 404.000 ;
        RECT 2161.360 400.000 2161.640 404.000 ;
        RECT 2163.660 400.000 2163.940 404.000 ;
        RECT 2165.960 400.000 2166.240 404.000 ;
        RECT 2167.800 400.000 2168.080 404.000 ;
        RECT 2170.100 400.000 2170.380 404.000 ;
        RECT 2172.400 400.000 2172.680 404.000 ;
        RECT 2174.700 400.000 2174.980 404.000 ;
        RECT 2177.000 400.000 2177.280 404.000 ;
        RECT 2179.300 400.000 2179.580 404.000 ;
        RECT 2181.600 400.000 2181.880 404.000 ;
        RECT 2183.900 400.000 2184.180 404.000 ;
        RECT 2185.740 400.000 2186.020 404.000 ;
        RECT 2188.040 400.000 2188.320 404.000 ;
        RECT 2190.340 400.000 2190.620 404.000 ;
        RECT 2192.640 400.000 2192.920 404.000 ;
        RECT 2194.940 400.000 2195.220 404.000 ;
        RECT 2197.240 400.000 2197.520 404.000 ;
        RECT 2199.540 400.000 2199.820 404.000 ;
        RECT 2201.840 400.000 2202.120 404.000 ;
        RECT 2203.680 400.000 2203.960 404.000 ;
        RECT 2205.980 400.000 2206.260 404.000 ;
        RECT 2208.280 400.000 2208.560 404.000 ;
        RECT 2210.580 400.000 2210.860 404.000 ;
        RECT 2212.880 400.000 2213.160 404.000 ;
        RECT 2215.180 400.000 2215.460 404.000 ;
        RECT 2217.480 400.000 2217.760 404.000 ;
        RECT 2219.780 400.000 2220.060 404.000 ;
        RECT 2221.620 400.000 2221.900 404.000 ;
        RECT 2223.920 400.000 2224.200 404.000 ;
        RECT 2226.220 400.000 2226.500 404.000 ;
        RECT 2228.520 400.000 2228.800 404.000 ;
        RECT 2230.820 400.000 2231.100 404.000 ;
        RECT 2233.120 400.000 2233.400 404.000 ;
        RECT 2235.420 400.000 2235.700 404.000 ;
        RECT 2237.720 400.000 2238.000 404.000 ;
        RECT 2240.020 400.000 2240.300 404.000 ;
        RECT 2241.860 400.000 2242.140 404.000 ;
        RECT 2244.160 400.000 2244.440 404.000 ;
        RECT 2246.460 400.000 2246.740 404.000 ;
        RECT 2248.760 400.000 2249.040 404.000 ;
        RECT 2251.060 400.000 2251.340 404.000 ;
        RECT 2253.360 400.000 2253.640 404.000 ;
        RECT 2255.660 400.000 2255.940 404.000 ;
        RECT 2257.960 400.000 2258.240 404.000 ;
        RECT 2259.800 400.000 2260.080 404.000 ;
        RECT 2262.100 400.000 2262.380 404.000 ;
        RECT 2264.400 400.000 2264.680 404.000 ;
        RECT 2266.700 400.000 2266.980 404.000 ;
        RECT 2269.000 400.000 2269.280 404.000 ;
        RECT 2271.300 400.000 2271.580 404.000 ;
        RECT 2273.600 400.000 2273.880 404.000 ;
        RECT 2275.900 400.000 2276.180 404.000 ;
        RECT 2277.740 400.000 2278.020 404.000 ;
        RECT 2280.040 400.000 2280.320 404.000 ;
        RECT 2282.340 400.000 2282.620 404.000 ;
        RECT 2284.640 400.000 2284.920 404.000 ;
        RECT 2286.940 400.000 2287.220 404.000 ;
        RECT 2289.240 400.000 2289.520 404.000 ;
        RECT 2291.540 400.000 2291.820 404.000 ;
        RECT 2293.840 400.000 2294.120 404.000 ;
        RECT 2296.140 400.000 2296.420 404.000 ;
        RECT 2297.980 400.000 2298.260 404.000 ;
        RECT 2300.280 400.000 2300.560 404.000 ;
        RECT 2302.580 400.000 2302.860 404.000 ;
        RECT 2304.880 400.000 2305.160 404.000 ;
        RECT 2307.180 400.000 2307.460 404.000 ;
        RECT 2309.480 400.000 2309.760 404.000 ;
        RECT 2311.780 400.000 2312.060 404.000 ;
        RECT 2314.080 400.000 2314.360 404.000 ;
        RECT 2315.920 400.000 2316.200 404.000 ;
        RECT 2318.220 400.000 2318.500 404.000 ;
        RECT 2320.520 400.000 2320.800 404.000 ;
        RECT 2322.820 400.000 2323.100 404.000 ;
        RECT 2325.120 400.000 2325.400 404.000 ;
        RECT 2327.420 400.000 2327.700 404.000 ;
        RECT 2329.720 400.000 2330.000 404.000 ;
        RECT 2332.020 400.000 2332.300 404.000 ;
        RECT 2333.860 400.000 2334.140 404.000 ;
        RECT 2336.160 400.000 2336.440 404.000 ;
        RECT 2338.460 400.000 2338.740 404.000 ;
        RECT 2340.760 400.000 2341.040 404.000 ;
        RECT 2343.060 400.000 2343.340 404.000 ;
        RECT 2345.360 400.000 2345.640 404.000 ;
        RECT 2347.660 400.000 2347.940 404.000 ;
        RECT 2349.960 400.000 2350.240 404.000 ;
        RECT 2352.260 400.000 2352.540 404.000 ;
        RECT 2354.100 400.000 2354.380 404.000 ;
        RECT 2356.400 400.000 2356.680 404.000 ;
        RECT 2358.700 400.000 2358.980 404.000 ;
        RECT 2361.000 400.000 2361.280 404.000 ;
        RECT 2363.300 400.000 2363.580 404.000 ;
        RECT 2365.600 400.000 2365.880 404.000 ;
        RECT 2367.900 400.000 2368.180 404.000 ;
        RECT 2370.200 400.000 2370.480 404.000 ;
        RECT 2372.040 400.000 2372.320 404.000 ;
        RECT 2374.340 400.000 2374.620 404.000 ;
        RECT 2376.640 400.000 2376.920 404.000 ;
        RECT 2378.940 400.000 2379.220 404.000 ;
        RECT 2381.240 400.000 2381.520 404.000 ;
        RECT 2383.540 400.000 2383.820 404.000 ;
        RECT 2385.840 400.000 2386.120 404.000 ;
        RECT 2388.140 400.000 2388.420 404.000 ;
        RECT 2389.980 400.000 2390.260 404.000 ;
        RECT 2392.280 400.000 2392.560 404.000 ;
        RECT 2394.580 400.000 2394.860 404.000 ;
        RECT 2396.880 400.000 2397.160 404.000 ;
        RECT 2399.180 400.000 2399.460 404.000 ;
        RECT 2401.480 400.000 2401.760 404.000 ;
        RECT 2403.780 400.000 2404.060 404.000 ;
        RECT 2406.080 400.000 2406.360 404.000 ;
        RECT 2408.380 400.000 2408.660 404.000 ;
        RECT 2410.220 400.000 2410.500 404.000 ;
        RECT 2412.520 400.000 2412.800 404.000 ;
        RECT 2414.820 400.000 2415.100 404.000 ;
        RECT 2417.120 400.000 2417.400 404.000 ;
        RECT 2419.420 400.000 2419.700 404.000 ;
        RECT 2421.720 400.000 2422.000 404.000 ;
        RECT 2424.020 400.000 2424.300 404.000 ;
        RECT 2426.320 400.000 2426.600 404.000 ;
        RECT 2428.160 400.000 2428.440 404.000 ;
        RECT 2430.460 400.000 2430.740 404.000 ;
        RECT 2432.760 400.000 2433.040 404.000 ;
        RECT 2435.060 400.000 2435.340 404.000 ;
        RECT 2437.360 400.000 2437.640 404.000 ;
        RECT 2439.660 400.000 2439.940 404.000 ;
        RECT 2441.960 400.000 2442.240 404.000 ;
        RECT 2444.260 400.000 2444.540 404.000 ;
        RECT 2446.100 400.000 2446.380 404.000 ;
        RECT 2448.400 400.000 2448.680 404.000 ;
        RECT 2450.700 400.000 2450.980 404.000 ;
        RECT 2453.000 400.000 2453.280 404.000 ;
        RECT 2455.300 400.000 2455.580 404.000 ;
        RECT 2457.600 400.000 2457.880 404.000 ;
        RECT 2459.900 400.000 2460.180 404.000 ;
        RECT 2462.200 400.000 2462.480 404.000 ;
        RECT 2464.040 400.000 2464.320 404.000 ;
        RECT 2466.340 400.000 2466.620 404.000 ;
        RECT 2468.640 400.000 2468.920 404.000 ;
        RECT 2470.940 400.000 2471.220 404.000 ;
        RECT 2473.240 400.000 2473.520 404.000 ;
        RECT 2475.540 400.000 2475.820 404.000 ;
        RECT 2477.840 400.000 2478.120 404.000 ;
        RECT 2480.140 400.000 2480.420 404.000 ;
        RECT 2482.440 400.000 2482.720 404.000 ;
        RECT 2484.280 400.000 2484.560 404.000 ;
        RECT 2486.580 400.000 2486.860 404.000 ;
        RECT 2488.880 400.000 2489.160 404.000 ;
        RECT 2491.180 400.000 2491.460 404.000 ;
        RECT 2493.480 400.000 2493.760 404.000 ;
        RECT 2495.780 400.000 2496.060 404.000 ;
        RECT 2498.080 400.000 2498.360 404.000 ;
        RECT 2500.380 400.000 2500.660 404.000 ;
        RECT 2502.220 400.000 2502.500 404.000 ;
        RECT 2504.520 400.000 2504.800 404.000 ;
        RECT 2506.820 400.000 2507.100 404.000 ;
        RECT 2509.120 400.000 2509.400 404.000 ;
        RECT 2511.420 400.000 2511.700 404.000 ;
        RECT 2513.720 400.000 2514.000 404.000 ;
        RECT 2516.020 400.000 2516.300 404.000 ;
        RECT 2518.320 400.000 2518.600 404.000 ;
        RECT 2520.160 400.000 2520.440 404.000 ;
        RECT 2522.460 400.000 2522.740 404.000 ;
        RECT 2524.760 400.000 2525.040 404.000 ;
        RECT 2527.060 400.000 2527.340 404.000 ;
        RECT 2529.360 400.000 2529.640 404.000 ;
        RECT 2531.660 400.000 2531.940 404.000 ;
        RECT 2533.960 400.000 2534.240 404.000 ;
        RECT 2536.260 400.000 2536.540 404.000 ;
        RECT 2538.560 400.000 2538.840 404.000 ;
        RECT 2540.400 400.000 2540.680 404.000 ;
        RECT 2542.700 400.000 2542.980 404.000 ;
        RECT 2545.000 400.000 2545.280 404.000 ;
        RECT 2547.300 400.000 2547.580 404.000 ;
        RECT 2549.600 400.000 2549.880 404.000 ;
        RECT 2551.900 400.000 2552.180 404.000 ;
        RECT 2554.200 400.000 2554.480 404.000 ;
        RECT 2556.500 400.000 2556.780 404.000 ;
        RECT 2558.340 400.000 2558.620 404.000 ;
        RECT 2560.640 400.000 2560.920 404.000 ;
        RECT 2562.940 400.000 2563.220 404.000 ;
        RECT 2565.240 400.000 2565.520 404.000 ;
        RECT 2567.540 400.000 2567.820 404.000 ;
        RECT 2569.840 400.000 2570.120 404.000 ;
        RECT 2572.140 400.000 2572.420 404.000 ;
        RECT 2574.440 400.000 2574.720 404.000 ;
        RECT 2576.280 400.000 2576.560 404.000 ;
        RECT 2578.580 400.000 2578.860 404.000 ;
        RECT 2580.880 400.000 2581.160 404.000 ;
        RECT 2583.180 400.000 2583.460 404.000 ;
        RECT 2585.480 400.000 2585.760 404.000 ;
        RECT 2587.780 400.000 2588.060 404.000 ;
        RECT 2590.080 400.000 2590.360 404.000 ;
        RECT 2592.380 400.000 2592.660 404.000 ;
        RECT 2594.680 400.000 2594.960 404.000 ;
        RECT 2596.520 400.000 2596.800 404.000 ;
        RECT 2598.820 400.000 2599.100 404.000 ;
        RECT 2601.120 400.000 2601.400 404.000 ;
        RECT 2603.420 400.000 2603.700 404.000 ;
        RECT 2605.720 400.000 2606.000 404.000 ;
        RECT 2608.020 400.000 2608.300 404.000 ;
        RECT 2610.320 400.000 2610.600 404.000 ;
        RECT 2612.620 400.000 2612.900 404.000 ;
        RECT 2614.460 400.000 2614.740 404.000 ;
        RECT 2616.760 400.000 2617.040 404.000 ;
        RECT 2619.060 400.000 2619.340 404.000 ;
        RECT 2621.360 400.000 2621.640 404.000 ;
        RECT 2623.660 400.000 2623.940 404.000 ;
        RECT 2625.960 400.000 2626.240 404.000 ;
        RECT 2628.260 400.000 2628.540 404.000 ;
        RECT 2630.560 400.000 2630.840 404.000 ;
        RECT 2632.400 400.000 2632.680 404.000 ;
        RECT 2634.700 400.000 2634.980 404.000 ;
        RECT 2637.000 400.000 2637.280 404.000 ;
        RECT 2639.300 400.000 2639.580 404.000 ;
        RECT 2641.600 400.000 2641.880 404.000 ;
        RECT 2643.900 400.000 2644.180 404.000 ;
        RECT 2646.200 400.000 2646.480 404.000 ;
        RECT 2648.500 400.000 2648.780 404.000 ;
      LAYER via2 ;
        RECT 646.390 3264.200 646.670 3264.480 ;
        RECT 668.470 3264.200 668.750 3264.480 ;
        RECT 1295.910 3264.200 1296.190 3264.480 ;
        RECT 1317.990 3264.200 1318.270 3264.480 ;
        RECT 1890.690 3264.200 1890.970 3264.480 ;
        RECT 1917.830 3264.200 1918.110 3264.480 ;
        RECT 2542.050 3264.200 2542.330 3264.480 ;
        RECT 2566.890 3264.200 2567.170 3264.480 ;
        RECT 289.430 3230.200 289.710 3230.480 ;
        RECT 288.970 3224.760 289.250 3225.040 ;
        RECT 288.510 3215.920 288.790 3216.200 ;
        RECT 288.050 3209.800 288.330 3210.080 ;
        RECT 287.590 3201.640 287.870 3201.920 ;
        RECT 287.130 3196.200 287.410 3196.480 ;
        RECT 286.670 3188.040 286.950 3188.320 ;
        RECT 286.210 2898.360 286.490 2898.640 ;
        RECT 688.250 3248.275 688.530 3248.555 ;
        RECT 941.710 3230.200 941.990 3230.480 ;
        RECT 696.990 2948.000 697.270 2948.280 ;
        RECT 696.990 2901.760 697.270 2902.040 ;
        RECT 938.490 2894.960 938.770 2895.240 ;
        RECT 337.730 2794.320 338.010 2794.600 ;
        RECT 344.630 2794.320 344.910 2794.600 ;
        RECT 351.070 2794.320 351.350 2794.600 ;
        RECT 358.430 2794.320 358.710 2794.600 ;
        RECT 362.570 2794.320 362.850 2794.600 ;
        RECT 365.330 2794.320 365.610 2794.600 ;
        RECT 368.550 2794.320 368.830 2794.600 ;
        RECT 371.310 2794.320 371.590 2794.600 ;
        RECT 374.990 2794.320 375.270 2794.600 ;
        RECT 379.130 2794.320 379.410 2794.600 ;
        RECT 384.190 2794.320 384.470 2794.600 ;
        RECT 386.950 2794.320 387.230 2794.600 ;
        RECT 392.930 2794.320 393.210 2794.600 ;
        RECT 396.610 2794.320 396.890 2794.600 ;
        RECT 399.830 2794.320 400.110 2794.600 ;
        RECT 403.970 2794.320 404.250 2794.600 ;
        RECT 406.270 2794.320 406.550 2794.600 ;
        RECT 409.950 2794.320 410.230 2794.600 ;
        RECT 413.630 2794.320 413.910 2794.600 ;
        RECT 419.150 2794.320 419.430 2794.600 ;
        RECT 420.990 2794.320 421.270 2794.600 ;
        RECT 427.430 2794.320 427.710 2794.600 ;
        RECT 433.870 2794.320 434.150 2794.600 ;
        RECT 439.390 2794.320 439.670 2794.600 ;
        RECT 441.230 2794.320 441.510 2794.600 ;
        RECT 444.450 2794.320 444.730 2794.600 ;
        RECT 446.750 2794.320 447.030 2794.600 ;
        RECT 449.050 2794.320 449.330 2794.600 ;
        RECT 455.030 2794.320 455.310 2794.600 ;
        RECT 461.470 2794.320 461.750 2794.600 ;
        RECT 462.390 2794.320 462.670 2794.600 ;
        RECT 468.370 2794.320 468.650 2794.600 ;
        RECT 474.350 2794.320 474.630 2794.600 ;
        RECT 475.270 2794.320 475.550 2794.600 ;
        RECT 478.490 2794.320 478.770 2794.600 ;
        RECT 482.630 2794.320 482.910 2794.600 ;
        RECT 485.390 2794.320 485.670 2794.600 ;
        RECT 488.150 2794.320 488.430 2794.600 ;
        RECT 492.750 2794.320 493.030 2794.600 ;
        RECT 496.430 2794.320 496.710 2794.600 ;
        RECT 502.870 2794.320 503.150 2794.600 ;
        RECT 510.230 2794.320 510.510 2794.600 ;
        RECT 524.030 2794.320 524.310 2794.600 ;
        RECT 537.370 2794.320 537.650 2794.600 ;
        RECT 542.430 2794.320 542.710 2794.600 ;
        RECT 310.130 2791.600 310.410 2791.880 ;
        RECT 317.030 2790.920 317.310 2791.200 ;
        RECT 351.530 2793.640 351.810 2793.920 ;
        RECT 379.590 2793.640 379.870 2793.920 ;
        RECT 392.470 2793.640 392.750 2793.920 ;
        RECT 397.530 2793.640 397.810 2793.920 ;
        RECT 387.870 2714.760 388.150 2715.040 ;
        RECT 414.550 2793.640 414.830 2793.920 ;
        RECT 426.970 2793.640 427.250 2793.920 ;
        RECT 433.410 2792.960 433.690 2793.240 ;
        RECT 434.330 2793.640 434.610 2793.920 ;
        RECT 455.490 2793.640 455.770 2793.920 ;
        RECT 467.910 2792.960 468.190 2793.240 ;
        RECT 468.830 2793.640 469.110 2793.920 ;
        RECT 481.250 2716.120 481.530 2716.400 ;
        RECT 496.890 2792.280 497.170 2792.560 ;
        RECT 524.490 2793.640 524.770 2793.920 ;
        RECT 500.110 2788.880 500.390 2789.160 ;
        RECT 504.250 2788.200 504.530 2788.480 ;
        RECT 507.010 2788.200 507.290 2788.480 ;
        RECT 531.390 2788.200 531.670 2788.480 ;
        RECT 534.610 2788.200 534.890 2788.480 ;
        RECT 510.230 2787.520 510.510 2787.800 ;
        RECT 513.910 2787.520 514.190 2787.800 ;
        RECT 517.130 2787.520 517.410 2787.800 ;
        RECT 520.810 2787.520 521.090 2787.800 ;
        RECT 527.710 2787.520 527.990 2787.800 ;
        RECT 530.930 2787.520 531.210 2787.800 ;
        RECT 517.130 2715.440 517.410 2715.720 ;
        RECT 541.510 2792.280 541.790 2792.560 ;
        RECT 538.290 2787.520 538.570 2787.800 ;
        RECT 542.430 2787.520 542.710 2787.800 ;
        RECT 551.630 2787.520 551.910 2787.800 ;
        RECT 700.210 2718.160 700.490 2718.440 ;
        RECT 707.110 2716.800 707.390 2717.080 ;
        RECT 741.610 2717.480 741.890 2717.760 ;
        RECT 942.170 3224.760 942.450 3225.040 ;
        RECT 942.630 3215.920 942.910 3216.200 ;
        RECT 943.090 3209.800 943.370 3210.080 ;
        RECT 943.550 3201.640 943.830 3201.920 ;
        RECT 944.010 3196.200 944.290 3196.480 ;
        RECT 944.470 3188.040 944.750 3188.320 ;
        RECT 944.930 2898.360 945.210 2898.640 ;
        RECT 941.710 2716.120 941.990 2716.400 ;
        RECT 1332.250 3249.240 1332.530 3249.520 ;
        RECT 1411.370 3243.120 1411.650 3243.400 ;
        RECT 1536.950 3230.200 1537.230 3230.480 ;
        RECT 1410.910 2935.760 1411.190 2936.040 ;
        RECT 1410.910 2932.360 1411.190 2932.640 ;
        RECT 1146.870 2799.760 1147.150 2800.040 ;
        RECT 1129.850 2799.080 1130.130 2799.360 ;
        RECT 979.890 2794.320 980.170 2794.600 ;
        RECT 1001.050 2794.320 1001.330 2794.600 ;
        RECT 1007.490 2794.320 1007.770 2794.600 ;
        RECT 1013.930 2794.320 1014.210 2794.600 ;
        RECT 1018.990 2794.320 1019.270 2794.600 ;
        RECT 1020.830 2794.320 1021.110 2794.600 ;
        RECT 1027.730 2794.320 1028.010 2794.600 ;
        RECT 1031.870 2794.320 1032.150 2794.600 ;
        RECT 1042.450 2794.320 1042.730 2794.600 ;
        RECT 1059.470 2794.320 1059.750 2794.600 ;
        RECT 1065.450 2794.320 1065.730 2794.600 ;
        RECT 1069.590 2794.320 1069.870 2794.600 ;
        RECT 1076.490 2794.320 1076.770 2794.600 ;
        RECT 1093.970 2794.320 1094.250 2794.600 ;
        RECT 1100.410 2794.320 1100.690 2794.600 ;
        RECT 1105.470 2794.320 1105.750 2794.600 ;
        RECT 1111.450 2794.320 1111.730 2794.600 ;
        RECT 1117.890 2794.320 1118.170 2794.600 ;
        RECT 1119.730 2794.320 1120.010 2794.600 ;
        RECT 944.930 2714.760 945.210 2715.040 ;
        RECT 1010.710 2793.640 1010.990 2793.920 ;
        RECT 1000.130 2718.160 1000.410 2718.440 ;
        RECT 1010.250 2715.440 1010.530 2715.720 ;
        RECT 1024.510 2792.960 1024.790 2793.240 ;
        RECT 1052.570 2792.960 1052.850 2793.240 ;
        RECT 1055.790 2792.960 1056.070 2793.240 ;
        RECT 1038.310 2788.200 1038.590 2788.480 ;
        RECT 1045.210 2788.200 1045.490 2788.480 ;
        RECT 1089.830 2793.640 1090.110 2793.920 ;
        RECT 1034.630 2787.520 1034.910 2787.800 ;
        RECT 1054.870 2788.200 1055.150 2788.480 ;
        RECT 1089.370 2788.200 1089.650 2788.480 ;
        RECT 1041.530 2787.520 1041.810 2787.800 ;
        RECT 1048.430 2787.520 1048.710 2787.800 ;
        RECT 1052.110 2717.480 1052.390 2717.760 ;
        RECT 1041.530 2716.800 1041.810 2717.080 ;
        RECT 1055.330 2787.520 1055.610 2787.800 ;
        RECT 1062.230 2787.520 1062.510 2787.800 ;
        RECT 1069.130 2787.520 1069.410 2787.800 ;
        RECT 1076.030 2787.520 1076.310 2787.800 ;
        RECT 1082.930 2787.520 1083.210 2787.800 ;
        RECT 1103.630 2792.960 1103.910 2793.240 ;
        RECT 1136.290 2796.360 1136.570 2796.640 ;
        RECT 1140.430 2794.320 1140.710 2794.600 ;
        RECT 1179.530 2794.320 1179.810 2794.600 ;
        RECT 1186.430 2794.320 1186.710 2794.600 ;
        RECT 1200.230 2794.320 1200.510 2794.600 ;
        RECT 1159.750 2793.640 1160.030 2793.920 ;
        RECT 1166.190 2793.640 1166.470 2793.920 ;
        RECT 1173.090 2793.640 1173.370 2793.920 ;
        RECT 1159.290 2792.960 1159.570 2793.240 ;
        RECT 1152.390 2792.280 1152.670 2792.560 ;
        RECT 1131.230 2788.200 1131.510 2788.480 ;
        RECT 1165.730 2788.200 1166.010 2788.480 ;
        RECT 1089.830 2787.520 1090.110 2787.800 ;
        RECT 1096.730 2787.520 1097.010 2787.800 ;
        RECT 1103.630 2787.520 1103.910 2787.800 ;
        RECT 1110.530 2787.520 1110.810 2787.800 ;
        RECT 1117.430 2787.520 1117.710 2787.800 ;
        RECT 1124.330 2787.520 1124.610 2787.800 ;
        RECT 1130.770 2787.520 1131.050 2787.800 ;
        RECT 1138.130 2787.520 1138.410 2787.800 ;
        RECT 1145.030 2787.520 1145.310 2787.800 ;
        RECT 1151.930 2787.520 1152.210 2787.800 ;
        RECT 1158.830 2787.520 1159.110 2787.800 ;
        RECT 1165.270 2787.520 1165.550 2787.800 ;
        RECT 1172.630 2787.520 1172.910 2787.800 ;
        RECT 1179.990 2793.640 1180.270 2793.920 ;
        RECT 1186.890 2792.960 1187.170 2793.240 ;
        RECT 1193.790 2791.600 1194.070 2791.880 ;
        RECT 1193.330 2790.240 1193.610 2790.520 ;
        RECT 1408.610 2695.040 1408.890 2695.320 ;
        RECT 1408.610 2684.840 1408.890 2685.120 ;
        RECT 1408.610 2674.640 1408.890 2674.920 ;
        RECT 1408.610 2664.440 1408.890 2664.720 ;
        RECT 1408.610 2654.240 1408.890 2654.520 ;
        RECT 1408.610 2644.040 1408.890 2644.320 ;
        RECT 1408.610 2633.840 1408.890 2634.120 ;
        RECT 1408.610 2623.640 1408.890 2623.920 ;
        RECT 1408.610 2613.440 1408.890 2613.720 ;
        RECT 1408.610 2603.240 1408.890 2603.520 ;
        RECT 1408.610 2593.040 1408.890 2593.320 ;
        RECT 1408.610 2582.840 1408.890 2583.120 ;
        RECT 1408.610 2572.640 1408.890 2572.920 ;
        RECT 1408.610 2562.440 1408.890 2562.720 ;
        RECT 1408.610 2552.240 1408.890 2552.520 ;
        RECT 1408.610 2542.040 1408.890 2542.320 ;
        RECT 1408.610 2531.840 1408.890 2532.120 ;
        RECT 1408.610 2521.640 1408.890 2521.920 ;
        RECT 1408.610 2511.440 1408.890 2511.720 ;
        RECT 1408.610 2501.240 1408.890 2501.520 ;
        RECT 1408.610 2491.040 1408.890 2491.320 ;
        RECT 1408.610 2480.840 1408.890 2481.120 ;
        RECT 1408.610 2470.640 1408.890 2470.920 ;
        RECT 1408.610 2460.440 1408.890 2460.720 ;
        RECT 1408.610 2450.240 1408.890 2450.520 ;
        RECT 1408.610 2440.040 1408.890 2440.320 ;
        RECT 1408.610 2429.840 1408.890 2430.120 ;
        RECT 1408.610 2419.640 1408.890 2419.920 ;
        RECT 1408.610 2409.440 1408.890 2409.720 ;
        RECT 1408.610 2399.240 1408.890 2399.520 ;
        RECT 1408.610 2389.040 1408.890 2389.320 ;
        RECT 1408.610 2378.840 1408.890 2379.120 ;
        RECT 1408.610 2368.640 1408.890 2368.920 ;
        RECT 1408.610 2358.440 1408.890 2358.720 ;
        RECT 1408.610 2348.240 1408.890 2348.520 ;
        RECT 1408.610 2338.040 1408.890 2338.320 ;
        RECT 1408.610 2327.840 1408.890 2328.120 ;
        RECT 1408.610 2317.640 1408.890 2317.920 ;
        RECT 1408.610 2307.440 1408.890 2307.720 ;
        RECT 1408.610 2297.240 1408.890 2297.520 ;
        RECT 1408.610 2287.040 1408.890 2287.320 ;
        RECT 1408.610 2276.840 1408.890 2277.120 ;
        RECT 1408.610 2266.640 1408.890 2266.920 ;
        RECT 1408.610 2256.440 1408.890 2256.720 ;
        RECT 1408.610 2246.240 1408.890 2246.520 ;
        RECT 1408.610 2236.040 1408.890 2236.320 ;
        RECT 1408.610 2225.840 1408.890 2226.120 ;
        RECT 1408.610 2215.640 1408.890 2215.920 ;
        RECT 1408.610 2205.440 1408.890 2205.720 ;
        RECT 1408.610 2195.240 1408.890 2195.520 ;
        RECT 1408.610 2185.040 1408.890 2185.320 ;
        RECT 1408.610 2174.840 1408.890 2175.120 ;
        RECT 1408.610 2164.640 1408.890 2164.920 ;
        RECT 1408.610 2155.120 1408.890 2155.400 ;
        RECT 1408.610 2144.920 1408.890 2145.200 ;
        RECT 1408.610 2134.720 1408.890 2135.000 ;
        RECT 1408.610 2124.520 1408.890 2124.800 ;
        RECT 1408.610 2114.320 1408.890 2114.600 ;
        RECT 1408.610 2104.120 1408.890 2104.400 ;
        RECT 1408.610 2093.920 1408.890 2094.200 ;
        RECT 1408.610 2083.720 1408.890 2084.000 ;
        RECT 1408.610 2073.520 1408.890 2073.800 ;
        RECT 1408.610 2063.320 1408.890 2063.600 ;
        RECT 1409.070 2042.920 1409.350 2043.200 ;
        RECT 1409.990 2053.120 1410.270 2053.400 ;
        RECT 1409.530 2032.720 1409.810 2033.000 ;
        RECT 1408.610 2022.520 1408.890 2022.800 ;
        RECT 1407.690 2012.320 1407.970 2012.600 ;
        RECT 1408.150 2002.120 1408.430 2002.400 ;
        RECT 1408.610 1991.920 1408.890 1992.200 ;
        RECT 1407.690 1981.720 1407.970 1982.000 ;
        RECT 1410.450 1971.520 1410.730 1971.800 ;
        RECT 1409.530 1889.920 1409.810 1890.200 ;
        RECT 1408.610 1828.720 1408.890 1829.000 ;
        RECT 1409.530 1808.320 1409.810 1808.600 ;
        RECT 1409.530 1798.120 1409.810 1798.400 ;
        RECT 1408.610 1787.920 1408.890 1788.200 ;
        RECT 1410.450 1777.720 1410.730 1778.000 ;
        RECT 1407.690 1726.720 1407.970 1727.000 ;
        RECT 1407.690 1706.320 1407.970 1706.600 ;
        RECT 1408.610 1696.120 1408.890 1696.400 ;
        RECT 1407.690 1685.920 1407.970 1686.200 ;
        RECT 1408.150 1675.720 1408.430 1676.000 ;
        RECT 1407.690 1665.520 1407.970 1665.800 ;
        RECT 1407.690 1655.320 1407.970 1655.600 ;
        RECT 1407.690 1645.120 1407.970 1645.400 ;
        RECT 1407.690 1634.920 1407.970 1635.200 ;
        RECT 1407.690 1624.720 1407.970 1625.000 ;
        RECT 1418.270 2790.920 1418.550 2791.200 ;
        RECT 1414.130 1961.320 1414.410 1961.600 ;
        RECT 1413.670 1951.120 1413.950 1951.400 ;
        RECT 1413.210 1940.920 1413.490 1941.200 ;
        RECT 1412.750 1930.720 1413.030 1931.000 ;
        RECT 1412.290 1920.520 1412.570 1920.800 ;
        RECT 1411.830 1910.320 1412.110 1910.600 ;
        RECT 1411.370 1900.120 1411.650 1900.400 ;
        RECT 1414.130 1879.720 1414.410 1880.000 ;
        RECT 1414.130 1869.520 1414.410 1869.800 ;
        RECT 1414.130 1859.320 1414.410 1859.600 ;
        RECT 1411.830 1849.120 1412.110 1849.400 ;
        RECT 1411.370 1838.920 1411.650 1839.200 ;
        RECT 1414.130 1818.520 1414.410 1818.800 ;
        RECT 1414.130 1767.520 1414.410 1767.800 ;
        RECT 1414.130 1757.320 1414.410 1757.600 ;
        RECT 1414.130 1747.120 1414.410 1747.400 ;
        RECT 1414.130 1738.280 1414.410 1738.560 ;
        RECT 1414.130 1716.520 1414.410 1716.800 ;
        RECT 1462.890 2792.960 1463.170 2793.240 ;
        RECT 1535.570 3224.760 1535.850 3225.040 ;
        RECT 1535.570 3217.280 1535.850 3217.560 ;
        RECT 1538.330 3210.480 1538.610 3210.760 ;
        RECT 1538.330 3202.320 1538.610 3202.600 ;
        RECT 1533.270 3196.880 1533.550 3197.160 ;
        RECT 1534.190 3189.400 1534.470 3189.680 ;
        RECT 1534.650 2899.720 1534.930 2900.000 ;
        RECT 1510.730 2792.960 1511.010 2793.240 ;
        RECT 1538.330 2894.280 1538.610 2894.560 ;
        RECT 1935.770 3249.240 1936.050 3249.520 ;
        RECT 2190.610 3230.200 2190.890 3230.480 ;
        RECT 1945.890 2904.480 1946.170 2904.760 ;
        RECT 2189.230 2895.640 2189.510 2895.920 ;
        RECT 1742.110 2796.360 1742.390 2796.640 ;
        RECT 1788.570 2796.360 1788.850 2796.640 ;
        RECT 1580.190 2794.320 1580.470 2794.600 ;
        RECT 1587.090 2794.320 1587.370 2794.600 ;
        RECT 1601.350 2794.320 1601.630 2794.600 ;
        RECT 1614.230 2794.320 1614.510 2794.600 ;
        RECT 1617.450 2794.320 1617.730 2794.600 ;
        RECT 1600.890 2793.640 1601.170 2793.920 ;
        RECT 1593.990 2792.960 1594.270 2793.240 ;
        RECT 1642.750 2794.320 1643.030 2794.600 ;
        RECT 1647.810 2794.320 1648.090 2794.600 ;
        RECT 1652.410 2794.320 1652.690 2794.600 ;
        RECT 1662.530 2794.320 1662.810 2794.600 ;
        RECT 1665.750 2794.320 1666.030 2794.600 ;
        RECT 1671.270 2794.320 1671.550 2794.600 ;
        RECT 1679.550 2794.320 1679.830 2794.600 ;
        RECT 1681.390 2794.320 1681.670 2794.600 ;
        RECT 1688.750 2794.320 1689.030 2794.600 ;
        RECT 1695.190 2794.320 1695.470 2794.600 ;
        RECT 1699.330 2794.320 1699.610 2794.600 ;
        RECT 1706.230 2794.320 1706.510 2794.600 ;
        RECT 1712.670 2794.320 1712.950 2794.600 ;
        RECT 1718.190 2794.320 1718.470 2794.600 ;
        RECT 1724.170 2794.320 1724.450 2794.600 ;
        RECT 1728.770 2794.320 1729.050 2794.600 ;
        RECT 1732.450 2794.320 1732.730 2794.600 ;
        RECT 1741.190 2794.320 1741.470 2794.600 ;
        RECT 1746.710 2794.320 1746.990 2794.600 ;
        RECT 1752.690 2794.320 1752.970 2794.600 ;
        RECT 1760.050 2794.320 1760.330 2794.600 ;
        RECT 1766.490 2794.320 1766.770 2794.600 ;
        RECT 1773.390 2793.640 1773.670 2793.920 ;
        RECT 1780.290 2793.640 1780.570 2793.920 ;
        RECT 1787.190 2792.280 1787.470 2792.560 ;
        RECT 1783.510 2791.600 1783.790 2791.880 ;
        RECT 1624.810 2788.200 1625.090 2788.480 ;
        RECT 1631.710 2788.200 1631.990 2788.480 ;
        RECT 1638.610 2788.200 1638.890 2788.480 ;
        RECT 1649.650 2788.200 1649.930 2788.480 ;
        RECT 1684.150 2788.200 1684.430 2788.480 ;
        RECT 1718.650 2788.200 1718.930 2788.480 ;
        RECT 1760.050 2788.200 1760.330 2788.480 ;
        RECT 1607.790 2787.520 1608.070 2787.800 ;
        RECT 1614.690 2787.520 1614.970 2787.800 ;
        RECT 1621.590 2787.520 1621.870 2787.800 ;
        RECT 1628.490 2787.520 1628.770 2787.800 ;
        RECT 1635.390 2787.520 1635.670 2787.800 ;
        RECT 1642.290 2787.520 1642.570 2787.800 ;
        RECT 1649.190 2787.520 1649.470 2787.800 ;
        RECT 1656.090 2787.520 1656.370 2787.800 ;
        RECT 1662.990 2787.520 1663.270 2787.800 ;
        RECT 1669.890 2787.520 1670.170 2787.800 ;
        RECT 1676.790 2787.520 1677.070 2787.800 ;
        RECT 1683.690 2787.520 1683.970 2787.800 ;
        RECT 1690.590 2787.520 1690.870 2787.800 ;
        RECT 1697.490 2787.520 1697.770 2787.800 ;
        RECT 1704.390 2787.520 1704.670 2787.800 ;
        RECT 1711.290 2787.520 1711.570 2787.800 ;
        RECT 1718.190 2787.520 1718.470 2787.800 ;
        RECT 1725.090 2787.520 1725.370 2787.800 ;
        RECT 1731.990 2787.520 1732.270 2787.800 ;
        RECT 1738.890 2787.520 1739.170 2787.800 ;
        RECT 1745.790 2787.520 1746.070 2787.800 ;
        RECT 1752.690 2787.520 1752.970 2787.800 ;
        RECT 1766.490 2787.520 1766.770 2787.800 ;
        RECT 1773.390 2787.520 1773.670 2787.800 ;
        RECT 1780.290 2787.520 1780.570 2787.800 ;
        RECT 1760.970 2777.320 1761.250 2777.600 ;
        RECT 1787.650 2787.520 1787.930 2787.800 ;
        RECT 1794.550 2777.320 1794.830 2777.600 ;
        RECT 2191.070 3224.760 2191.350 3225.040 ;
        RECT 2191.530 3215.920 2191.810 3216.200 ;
        RECT 2191.990 3209.800 2192.270 3210.080 ;
        RECT 2192.450 3201.640 2192.730 3201.920 ;
        RECT 2192.910 3196.200 2193.190 3196.480 ;
        RECT 2193.370 3188.040 2193.650 3188.320 ;
        RECT 2193.830 2898.360 2194.110 2898.640 ;
        RECT 2582.070 3249.240 2582.350 3249.520 ;
        RECT 2594.490 2946.640 2594.770 2946.920 ;
        RECT 2594.490 2938.480 2594.770 2938.760 ;
        RECT 2228.790 2794.320 2229.070 2794.600 ;
        RECT 2237.990 2794.320 2238.270 2794.600 ;
        RECT 2268.350 2794.320 2268.630 2794.600 ;
        RECT 2273.410 2794.320 2273.690 2794.600 ;
        RECT 2279.850 2794.320 2280.130 2794.600 ;
        RECT 2286.750 2794.320 2287.030 2794.600 ;
        RECT 2291.350 2794.320 2291.630 2794.600 ;
        RECT 2304.230 2794.320 2304.510 2794.600 ;
        RECT 2308.370 2794.320 2308.650 2794.600 ;
        RECT 2312.970 2794.320 2313.250 2794.600 ;
        RECT 2321.250 2794.320 2321.530 2794.600 ;
        RECT 2326.310 2794.320 2326.590 2794.600 ;
        RECT 2332.290 2794.320 2332.570 2794.600 ;
        RECT 2339.190 2794.320 2339.470 2794.600 ;
        RECT 2343.330 2794.320 2343.610 2794.600 ;
        RECT 2346.090 2794.320 2346.370 2794.600 ;
        RECT 2352.990 2794.320 2353.270 2794.600 ;
        RECT 2359.890 2794.320 2360.170 2794.600 ;
        RECT 2366.790 2794.320 2367.070 2794.600 ;
        RECT 2374.150 2794.320 2374.430 2794.600 ;
        RECT 2377.370 2794.320 2377.650 2794.600 ;
        RECT 2385.650 2794.320 2385.930 2794.600 ;
        RECT 2391.170 2794.320 2391.450 2794.600 ;
        RECT 2394.850 2794.320 2395.130 2794.600 ;
        RECT 2402.670 2794.320 2402.950 2794.600 ;
        RECT 2415.090 2794.320 2415.370 2794.600 ;
        RECT 2263.290 2793.640 2263.570 2793.920 ;
        RECT 2249.490 2792.280 2249.770 2792.560 ;
        RECT 2266.510 2792.960 2266.790 2793.240 ;
        RECT 2269.730 2792.960 2270.010 2793.240 ;
        RECT 2256.390 2790.240 2256.670 2790.520 ;
        RECT 2263.290 2787.520 2263.570 2787.800 ;
        RECT 2266.970 2787.520 2267.250 2787.800 ;
        RECT 2298.250 2792.960 2298.530 2793.240 ;
        RECT 2314.810 2792.960 2315.090 2793.240 ;
        RECT 2305.150 2788.200 2305.430 2788.480 ;
        RECT 2277.090 2787.520 2277.370 2787.800 ;
        RECT 2283.990 2787.520 2284.270 2787.800 ;
        RECT 2290.890 2787.520 2291.170 2787.800 ;
        RECT 2297.790 2787.520 2298.070 2787.800 ;
        RECT 2304.690 2787.520 2304.970 2787.800 ;
        RECT 2311.590 2787.520 2311.870 2787.800 ;
        RECT 2318.490 2787.520 2318.770 2787.800 ;
        RECT 2325.390 2787.520 2325.670 2787.800 ;
        RECT 2332.750 2793.640 2333.030 2793.920 ;
        RECT 2339.650 2793.640 2339.930 2793.920 ;
        RECT 2340.110 2792.960 2340.390 2793.240 ;
        RECT 2350.230 2793.640 2350.510 2793.920 ;
        RECT 2356.670 2793.640 2356.950 2793.920 ;
        RECT 2360.810 2793.640 2361.090 2793.920 ;
        RECT 2367.250 2792.960 2367.530 2793.240 ;
        RECT 2380.590 2792.280 2380.870 2792.560 ;
        RECT 2381.050 2791.600 2381.330 2791.880 ;
        RECT 2387.490 2791.600 2387.770 2791.880 ;
        RECT 2394.390 2790.920 2394.670 2791.200 ;
        RECT 2401.750 2793.640 2402.030 2793.920 ;
        RECT 2408.190 2793.640 2408.470 2793.920 ;
        RECT 2421.990 2792.960 2422.270 2793.240 ;
        RECT 2442.690 2792.960 2442.970 2793.240 ;
        RECT 2408.190 2792.280 2408.470 2792.560 ;
        RECT 2428.890 2792.280 2429.170 2792.560 ;
        RECT 2435.790 2792.280 2436.070 2792.560 ;
        RECT 2415.090 2790.920 2415.370 2791.200 ;
        RECT 2421.990 2790.920 2422.270 2791.200 ;
        RECT 2428.890 2790.920 2429.170 2791.200 ;
        RECT 2415.550 2790.240 2415.830 2790.520 ;
        RECT 2415.090 2788.200 2415.370 2788.480 ;
        RECT 2442.690 2790.240 2442.970 2790.520 ;
        RECT 2435.790 2789.560 2436.070 2789.840 ;
        RECT 2373.230 2787.520 2373.510 2787.800 ;
        RECT 2381.970 2787.520 2382.250 2787.800 ;
        RECT 1410.910 1605.000 1411.190 1605.280 ;
      LAYER met3 ;
        RECT 646.365 3264.500 646.695 3264.505 ;
        RECT 668.445 3264.500 668.775 3264.505 ;
        RECT 1295.885 3264.500 1296.215 3264.505 ;
        RECT 1317.965 3264.500 1318.295 3264.505 ;
        RECT 646.110 3264.490 646.695 3264.500 ;
        RECT 668.190 3264.490 668.775 3264.500 ;
        RECT 1295.630 3264.490 1296.215 3264.500 ;
        RECT 645.910 3264.190 646.695 3264.490 ;
        RECT 667.990 3264.190 668.775 3264.490 ;
        RECT 1295.430 3264.190 1296.215 3264.490 ;
        RECT 646.110 3264.180 646.695 3264.190 ;
        RECT 668.190 3264.180 668.775 3264.190 ;
        RECT 1295.630 3264.180 1296.215 3264.190 ;
        RECT 1317.710 3264.490 1318.295 3264.500 ;
        RECT 1890.665 3264.500 1890.995 3264.505 ;
        RECT 1917.805 3264.500 1918.135 3264.505 ;
        RECT 1890.665 3264.490 1891.250 3264.500 ;
        RECT 1917.550 3264.490 1918.135 3264.500 ;
        RECT 1317.710 3264.190 1318.520 3264.490 ;
        RECT 1890.665 3264.190 1891.450 3264.490 ;
        RECT 1917.350 3264.190 1918.135 3264.490 ;
        RECT 1317.710 3264.180 1318.295 3264.190 ;
        RECT 646.365 3264.175 646.695 3264.180 ;
        RECT 668.445 3264.175 668.775 3264.180 ;
        RECT 1295.885 3264.175 1296.215 3264.180 ;
        RECT 1317.965 3264.175 1318.295 3264.180 ;
        RECT 1890.665 3264.180 1891.250 3264.190 ;
        RECT 1917.550 3264.180 1918.135 3264.190 ;
        RECT 1890.665 3264.175 1890.995 3264.180 ;
        RECT 1917.805 3264.175 1918.135 3264.180 ;
        RECT 2542.025 3264.500 2542.355 3264.505 ;
        RECT 2566.865 3264.500 2567.195 3264.505 ;
        RECT 2542.025 3264.490 2542.610 3264.500 ;
        RECT 2566.865 3264.490 2567.450 3264.500 ;
        RECT 2542.025 3264.190 2542.810 3264.490 ;
        RECT 2566.865 3264.190 2567.650 3264.490 ;
        RECT 2542.025 3264.180 2542.610 3264.190 ;
        RECT 2566.865 3264.180 2567.450 3264.190 ;
        RECT 2542.025 3264.175 2542.355 3264.180 ;
        RECT 2566.865 3264.175 2567.195 3264.180 ;
        RECT 659.280 3251.235 661.020 3252.140 ;
        RECT 1309.280 3251.235 1311.020 3252.140 ;
        RECT 1909.280 3251.235 1911.020 3252.140 ;
        RECT 2559.280 3251.235 2561.020 3252.140 ;
        RECT 300.000 3232.785 304.600 3233.085 ;
        RECT 289.405 3230.490 289.735 3230.505 ;
        RECT 300.230 3230.490 300.530 3232.785 ;
        RECT 289.405 3230.190 300.530 3230.490 ;
        RECT 289.405 3230.175 289.735 3230.190 ;
        RECT 300.000 3227.145 304.600 3227.445 ;
        RECT 288.945 3225.050 289.275 3225.065 ;
        RECT 300.230 3225.050 300.530 3227.145 ;
        RECT 288.945 3224.750 300.530 3225.050 ;
        RECT 288.945 3224.735 289.275 3224.750 ;
        RECT 300.000 3218.645 304.600 3218.945 ;
        RECT 288.485 3216.210 288.815 3216.225 ;
        RECT 300.230 3216.210 300.530 3218.645 ;
        RECT 288.485 3215.910 300.530 3216.210 ;
        RECT 288.485 3215.895 288.815 3215.910 ;
        RECT 300.000 3213.005 304.600 3213.305 ;
        RECT 288.025 3210.090 288.355 3210.105 ;
        RECT 300.230 3210.090 300.530 3213.005 ;
        RECT 288.025 3209.790 300.530 3210.090 ;
        RECT 288.025 3209.775 288.355 3209.790 ;
        RECT 300.000 3204.505 304.600 3204.805 ;
        RECT 287.565 3201.930 287.895 3201.945 ;
        RECT 300.230 3201.930 300.530 3204.505 ;
        RECT 287.565 3201.630 300.530 3201.930 ;
        RECT 287.565 3201.615 287.895 3201.630 ;
        RECT 300.000 3198.865 304.600 3199.165 ;
        RECT 287.105 3196.490 287.435 3196.505 ;
        RECT 300.230 3196.490 300.530 3198.865 ;
        RECT 287.105 3196.190 300.530 3196.490 ;
        RECT 287.105 3196.175 287.435 3196.190 ;
        RECT 300.000 3190.365 304.600 3190.665 ;
        RECT 286.645 3188.330 286.975 3188.345 ;
        RECT 300.230 3188.330 300.530 3190.365 ;
        RECT 286.645 3188.030 300.530 3188.330 ;
        RECT 286.645 3188.015 286.975 3188.030 ;
        RECT 300.000 2901.125 304.600 2901.425 ;
        RECT 286.185 2898.650 286.515 2898.665 ;
        RECT 300.230 2898.650 300.530 2901.125 ;
        RECT 286.185 2898.350 300.530 2898.650 ;
        RECT 286.185 2898.335 286.515 2898.350 ;
        RECT 302.950 2894.940 303.330 2895.260 ;
        RECT 302.990 2892.925 303.290 2894.940 ;
        RECT 300.000 2892.625 304.600 2892.925 ;
      LAYER met3 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met3 ;
        RECT 688.225 3248.565 688.555 3248.580 ;
        RECT 681.880 3248.265 688.555 3248.565 ;
        RECT 688.225 3248.250 688.555 3248.265 ;
        RECT 950.000 3232.785 954.600 3233.085 ;
        RECT 941.685 3230.490 942.015 3230.505 ;
        RECT 950.670 3230.490 950.970 3232.785 ;
        RECT 941.685 3230.190 950.970 3230.490 ;
        RECT 941.685 3230.175 942.015 3230.190 ;
        RECT 950.000 3227.145 954.600 3227.445 ;
        RECT 942.145 3225.050 942.475 3225.065 ;
        RECT 950.670 3225.050 950.970 3227.145 ;
        RECT 942.145 3224.750 950.970 3225.050 ;
        RECT 942.145 3224.735 942.475 3224.750 ;
        RECT 950.000 3218.645 954.600 3218.945 ;
        RECT 942.605 3216.210 942.935 3216.225 ;
        RECT 950.670 3216.210 950.970 3218.645 ;
        RECT 942.605 3215.910 950.970 3216.210 ;
        RECT 942.605 3215.895 942.935 3215.910 ;
        RECT 950.000 3213.005 954.600 3213.305 ;
        RECT 943.065 3210.090 943.395 3210.105 ;
        RECT 950.670 3210.090 950.970 3213.005 ;
        RECT 943.065 3209.790 950.970 3210.090 ;
        RECT 943.065 3209.775 943.395 3209.790 ;
        RECT 950.000 3204.505 954.600 3204.805 ;
        RECT 943.525 3201.930 943.855 3201.945 ;
        RECT 950.670 3201.930 950.970 3204.505 ;
        RECT 943.525 3201.630 950.970 3201.930 ;
        RECT 943.525 3201.615 943.855 3201.630 ;
        RECT 950.000 3198.865 954.600 3199.165 ;
        RECT 943.985 3196.490 944.315 3196.505 ;
        RECT 950.670 3196.490 950.970 3198.865 ;
        RECT 943.985 3196.190 950.970 3196.490 ;
        RECT 943.985 3196.175 944.315 3196.190 ;
        RECT 950.000 3190.365 954.600 3190.665 ;
        RECT 944.445 3188.330 944.775 3188.345 ;
        RECT 950.670 3188.330 950.970 3190.365 ;
        RECT 944.445 3188.030 950.970 3188.330 ;
        RECT 944.445 3188.015 944.775 3188.030 ;
        RECT 696.965 2948.290 697.295 2948.305 ;
        RECT 684.790 2947.990 697.295 2948.290 ;
        RECT 684.790 2947.210 685.090 2947.990 ;
        RECT 696.965 2947.975 697.295 2947.990 ;
        RECT 681.880 2946.910 686.480 2947.210 ;
        RECT 684.790 2938.710 685.090 2946.910 ;
        RECT 681.880 2938.410 686.480 2938.710 ;
        RECT 684.790 2933.070 685.090 2938.410 ;
        RECT 681.880 2932.770 686.480 2933.070 ;
        RECT 685.710 2924.570 686.010 2932.770 ;
        RECT 681.880 2924.270 686.480 2924.570 ;
        RECT 685.710 2918.930 686.010 2924.270 ;
        RECT 681.880 2918.630 686.480 2918.930 ;
        RECT 685.710 2910.430 686.010 2918.630 ;
        RECT 681.880 2910.130 686.480 2910.430 ;
        RECT 685.710 2904.790 686.010 2910.130 ;
        RECT 681.880 2904.490 686.480 2904.790 ;
        RECT 685.710 2902.050 686.010 2904.490 ;
        RECT 687.510 2902.050 687.890 2902.060 ;
        RECT 696.965 2902.050 697.295 2902.065 ;
        RECT 685.710 2901.750 697.295 2902.050 ;
        RECT 687.510 2901.740 687.890 2901.750 ;
        RECT 696.965 2901.735 697.295 2901.750 ;
        RECT 950.000 2901.125 954.600 2901.425 ;
        RECT 944.905 2898.650 945.235 2898.665 ;
        RECT 950.670 2898.650 950.970 2901.125 ;
        RECT 944.905 2898.350 950.970 2898.650 ;
        RECT 944.905 2898.335 945.235 2898.350 ;
        RECT 938.465 2895.250 938.795 2895.265 ;
        RECT 950.630 2895.250 951.010 2895.260 ;
        RECT 938.465 2894.950 951.010 2895.250 ;
        RECT 938.465 2894.935 938.795 2894.950 ;
        RECT 950.630 2894.940 951.010 2894.950 ;
        RECT 950.670 2892.925 950.970 2894.940 ;
        RECT 950.000 2892.625 954.600 2892.925 ;
      LAYER met3 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met3 ;
        RECT 1332.225 3249.530 1332.555 3249.545 ;
        RECT 1332.225 3249.215 1332.770 3249.530 ;
        RECT 1332.470 3248.565 1332.770 3249.215 ;
        RECT 1331.880 3248.265 1336.480 3248.565 ;
        RECT 1411.345 3243.420 1411.675 3243.425 ;
        RECT 1411.345 3243.410 1411.930 3243.420 ;
        RECT 1411.345 3243.110 1412.130 3243.410 ;
        RECT 1411.345 3243.100 1411.930 3243.110 ;
        RECT 1411.345 3243.095 1411.675 3243.100 ;
        RECT 1550.000 3232.785 1554.600 3233.085 ;
        RECT 1536.925 3230.490 1537.255 3230.505 ;
        RECT 1550.510 3230.490 1550.810 3232.785 ;
        RECT 1536.925 3230.190 1550.810 3230.490 ;
        RECT 1536.925 3230.175 1537.255 3230.190 ;
        RECT 1550.000 3227.145 1554.600 3227.445 ;
        RECT 1535.545 3225.050 1535.875 3225.065 ;
        RECT 1550.510 3225.050 1550.810 3227.145 ;
        RECT 1535.545 3224.750 1550.810 3225.050 ;
        RECT 1535.545 3224.735 1535.875 3224.750 ;
        RECT 1550.000 3218.645 1554.600 3218.945 ;
        RECT 1535.545 3217.570 1535.875 3217.585 ;
        RECT 1550.510 3217.570 1550.810 3218.645 ;
        RECT 1535.545 3217.270 1550.810 3217.570 ;
        RECT 1535.545 3217.255 1535.875 3217.270 ;
        RECT 1550.000 3213.005 1554.600 3213.305 ;
        RECT 1538.305 3210.770 1538.635 3210.785 ;
        RECT 1550.510 3210.770 1550.810 3213.005 ;
        RECT 1538.305 3210.470 1550.810 3210.770 ;
        RECT 1538.305 3210.455 1538.635 3210.470 ;
        RECT 1550.000 3204.505 1554.600 3204.805 ;
        RECT 1538.305 3202.610 1538.635 3202.625 ;
        RECT 1550.510 3202.610 1550.810 3204.505 ;
        RECT 1538.305 3202.310 1550.810 3202.610 ;
        RECT 1538.305 3202.295 1538.635 3202.310 ;
        RECT 1550.000 3198.865 1554.600 3199.165 ;
        RECT 1533.245 3197.170 1533.575 3197.185 ;
        RECT 1550.510 3197.170 1550.810 3198.865 ;
        RECT 1533.245 3196.870 1550.810 3197.170 ;
        RECT 1533.245 3196.855 1533.575 3196.870 ;
        RECT 1550.000 3190.365 1554.600 3190.665 ;
        RECT 1534.165 3189.690 1534.495 3189.705 ;
        RECT 1550.510 3189.690 1550.810 3190.365 ;
        RECT 1534.165 3189.390 1550.810 3189.690 ;
        RECT 1534.165 3189.375 1534.495 3189.390 ;
        RECT 1331.880 2946.910 1336.480 2947.210 ;
        RECT 1335.230 2938.710 1335.530 2946.910 ;
        RECT 1331.880 2938.410 1336.480 2938.710 ;
        RECT 1335.230 2933.330 1335.530 2938.410 ;
        RECT 1410.885 2936.050 1411.215 2936.065 ;
        RECT 1413.390 2936.050 1413.770 2936.060 ;
        RECT 1410.885 2935.750 1413.770 2936.050 ;
        RECT 1410.885 2935.735 1411.215 2935.750 ;
        RECT 1413.390 2935.740 1413.770 2935.750 ;
        RECT 1335.230 2933.070 1336.450 2933.330 ;
        RECT 1331.880 2932.770 1338.290 2933.070 ;
        RECT 1335.230 2924.570 1335.530 2932.770 ;
        RECT 1337.990 2932.650 1338.290 2932.770 ;
        RECT 1410.885 2932.650 1411.215 2932.665 ;
        RECT 1337.990 2932.350 1411.215 2932.650 ;
        RECT 1410.885 2932.335 1411.215 2932.350 ;
        RECT 1331.880 2924.270 1336.480 2924.570 ;
        RECT 1335.230 2918.930 1335.530 2924.270 ;
        RECT 1331.880 2918.630 1336.480 2918.930 ;
        RECT 1336.150 2910.430 1336.450 2918.630 ;
        RECT 1331.880 2910.130 1336.480 2910.430 ;
        RECT 1336.150 2904.790 1336.450 2910.130 ;
        RECT 1331.880 2904.770 1336.480 2904.790 ;
        RECT 1345.310 2904.770 1345.690 2904.780 ;
        RECT 1331.880 2904.490 1345.690 2904.770 ;
        RECT 1336.150 2904.470 1345.690 2904.490 ;
        RECT 1345.310 2904.460 1345.690 2904.470 ;
        RECT 1550.000 2901.125 1554.600 2901.425 ;
        RECT 1534.625 2900.010 1534.955 2900.025 ;
        RECT 1550.510 2900.010 1550.810 2901.125 ;
        RECT 1534.625 2899.710 1550.810 2900.010 ;
        RECT 1534.625 2899.695 1534.955 2899.710 ;
        RECT 1538.305 2894.570 1538.635 2894.585 ;
        RECT 1538.305 2894.270 1550.810 2894.570 ;
        RECT 1538.305 2894.255 1538.635 2894.270 ;
        RECT 1550.510 2892.925 1550.810 2894.270 ;
        RECT 1550.000 2892.625 1554.600 2892.925 ;
      LAYER met3 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met3 ;
        RECT 1935.745 3249.530 1936.075 3249.545 ;
        RECT 1935.745 3249.215 1936.290 3249.530 ;
        RECT 1935.990 3248.565 1936.290 3249.215 ;
        RECT 1931.880 3248.265 1936.480 3248.565 ;
        RECT 2200.000 3232.785 2204.600 3233.085 ;
        RECT 2190.585 3230.490 2190.915 3230.505 ;
        RECT 2200.030 3230.490 2200.330 3232.785 ;
        RECT 2190.585 3230.190 2200.330 3230.490 ;
        RECT 2190.585 3230.175 2190.915 3230.190 ;
        RECT 2200.000 3227.145 2204.600 3227.445 ;
        RECT 2191.045 3225.050 2191.375 3225.065 ;
        RECT 2200.030 3225.050 2200.330 3227.145 ;
        RECT 2191.045 3224.750 2200.330 3225.050 ;
        RECT 2191.045 3224.735 2191.375 3224.750 ;
        RECT 2200.000 3218.645 2204.600 3218.945 ;
        RECT 2191.505 3216.210 2191.835 3216.225 ;
        RECT 2200.030 3216.210 2200.330 3218.645 ;
        RECT 2191.505 3215.910 2200.330 3216.210 ;
        RECT 2191.505 3215.895 2191.835 3215.910 ;
        RECT 2200.000 3213.005 2204.600 3213.305 ;
        RECT 2191.965 3210.090 2192.295 3210.105 ;
        RECT 2200.030 3210.090 2200.330 3213.005 ;
        RECT 2191.965 3209.790 2200.330 3210.090 ;
        RECT 2191.965 3209.775 2192.295 3209.790 ;
        RECT 2200.000 3204.505 2204.600 3204.805 ;
        RECT 2192.425 3201.930 2192.755 3201.945 ;
        RECT 2200.030 3201.930 2200.330 3204.505 ;
        RECT 2192.425 3201.630 2200.330 3201.930 ;
        RECT 2192.425 3201.615 2192.755 3201.630 ;
        RECT 2200.000 3198.865 2204.600 3199.165 ;
        RECT 2192.885 3196.490 2193.215 3196.505 ;
        RECT 2200.030 3196.490 2200.330 3198.865 ;
        RECT 2192.885 3196.190 2200.330 3196.490 ;
        RECT 2192.885 3196.175 2193.215 3196.190 ;
        RECT 2200.000 3190.365 2204.600 3190.665 ;
        RECT 2193.345 3188.330 2193.675 3188.345 ;
        RECT 2200.030 3188.330 2200.330 3190.365 ;
        RECT 2193.345 3188.030 2200.330 3188.330 ;
        RECT 2193.345 3188.015 2193.675 3188.030 ;
        RECT 1931.880 2946.910 1936.480 2947.210 ;
        RECT 1935.990 2938.710 1936.290 2946.910 ;
        RECT 1931.880 2938.410 1936.480 2938.710 ;
        RECT 1935.990 2936.050 1936.290 2938.410 ;
        RECT 1937.790 2936.050 1938.170 2936.060 ;
        RECT 1935.990 2935.750 1938.170 2936.050 ;
        RECT 1935.990 2933.070 1936.290 2935.750 ;
        RECT 1937.790 2935.740 1938.170 2935.750 ;
        RECT 1931.880 2932.770 1936.480 2933.070 ;
        RECT 1935.990 2924.570 1936.290 2932.770 ;
        RECT 1931.880 2924.270 1936.480 2924.570 ;
        RECT 1935.990 2918.930 1936.290 2924.270 ;
        RECT 1931.880 2918.630 1936.480 2918.930 ;
        RECT 1935.990 2910.430 1936.290 2918.630 ;
        RECT 1931.880 2910.130 1936.480 2910.430 ;
        RECT 1935.990 2904.790 1936.290 2910.130 ;
        RECT 1931.880 2904.770 1936.480 2904.790 ;
        RECT 1945.865 2904.770 1946.195 2904.785 ;
        RECT 1931.880 2904.490 1946.195 2904.770 ;
        RECT 1935.990 2904.470 1946.195 2904.490 ;
        RECT 1945.865 2904.455 1946.195 2904.470 ;
        RECT 2200.000 2901.125 2204.600 2901.425 ;
        RECT 2193.805 2898.650 2194.135 2898.665 ;
        RECT 2200.030 2898.650 2200.330 2901.125 ;
        RECT 2193.805 2898.350 2200.330 2898.650 ;
        RECT 2193.805 2898.335 2194.135 2898.350 ;
        RECT 2189.205 2895.930 2189.535 2895.945 ;
        RECT 2199.990 2895.930 2200.370 2895.940 ;
        RECT 2189.205 2895.630 2200.370 2895.930 ;
        RECT 2189.205 2895.615 2189.535 2895.630 ;
        RECT 2199.990 2895.620 2200.370 2895.630 ;
        RECT 2200.030 2892.925 2200.330 2895.620 ;
        RECT 2200.000 2892.625 2204.600 2892.925 ;
      LAYER met3 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met3 ;
        RECT 2582.045 3249.530 2582.375 3249.545 ;
        RECT 2582.045 3249.230 2583.050 3249.530 ;
        RECT 2582.045 3249.215 2582.375 3249.230 ;
        RECT 2582.750 3248.565 2583.050 3249.230 ;
        RECT 2581.880 3248.265 2586.480 3248.565 ;
        RECT 2581.880 2946.930 2586.480 2947.210 ;
        RECT 2594.465 2946.930 2594.795 2946.945 ;
        RECT 2581.880 2946.910 2594.795 2946.930 ;
        RECT 2585.510 2946.630 2594.795 2946.910 ;
        RECT 2594.465 2946.615 2594.795 2946.630 ;
        RECT 2594.465 2938.770 2594.795 2938.785 ;
        RECT 2585.510 2938.710 2594.795 2938.770 ;
        RECT 2581.880 2938.470 2594.795 2938.710 ;
        RECT 2581.880 2938.410 2586.480 2938.470 ;
        RECT 2594.465 2938.455 2594.795 2938.470 ;
        RECT 2585.510 2933.070 2585.810 2938.410 ;
        RECT 2581.880 2932.770 2586.480 2933.070 ;
        RECT 2585.510 2924.570 2585.810 2932.770 ;
        RECT 2581.880 2924.270 2586.480 2924.570 ;
        RECT 2585.510 2918.930 2585.810 2924.270 ;
        RECT 2581.880 2918.630 2586.480 2918.930 ;
        RECT 2585.510 2910.430 2585.810 2918.630 ;
        RECT 2581.880 2910.130 2586.480 2910.430 ;
        RECT 2585.510 2904.790 2585.810 2910.130 ;
        RECT 2581.880 2904.770 2586.480 2904.790 ;
        RECT 2594.670 2904.770 2595.050 2904.780 ;
        RECT 2581.880 2904.490 2595.050 2904.770 ;
        RECT 2585.510 2904.470 2595.050 2904.490 ;
        RECT 2594.670 2904.460 2595.050 2904.470 ;
        RECT 1146.845 2800.060 1147.175 2800.065 ;
        RECT 1146.590 2800.050 1147.175 2800.060 ;
        RECT 1146.390 2799.750 1147.175 2800.050 ;
        RECT 1146.590 2799.740 1147.175 2799.750 ;
        RECT 1146.845 2799.735 1147.175 2799.740 ;
        RECT 1129.110 2799.370 1129.490 2799.380 ;
        RECT 1129.825 2799.370 1130.155 2799.385 ;
        RECT 1129.110 2799.070 1130.155 2799.370 ;
        RECT 1129.110 2799.060 1129.490 2799.070 ;
        RECT 1129.825 2799.055 1130.155 2799.070 ;
        RECT 1135.550 2796.650 1135.930 2796.660 ;
        RECT 1136.265 2796.650 1136.595 2796.665 ;
        RECT 1135.550 2796.350 1136.595 2796.650 ;
        RECT 1135.550 2796.340 1135.930 2796.350 ;
        RECT 1136.265 2796.335 1136.595 2796.350 ;
        RECT 1742.085 2796.650 1742.415 2796.665 ;
        RECT 1759.310 2796.650 1759.690 2796.660 ;
        RECT 1742.085 2796.350 1759.690 2796.650 ;
        RECT 1742.085 2796.335 1742.415 2796.350 ;
        RECT 1759.310 2796.340 1759.690 2796.350 ;
        RECT 1788.545 2796.650 1788.875 2796.665 ;
        RECT 1794.270 2796.650 1794.650 2796.660 ;
        RECT 1788.545 2796.350 1794.650 2796.650 ;
        RECT 1788.545 2796.335 1788.875 2796.350 ;
        RECT 1794.270 2796.340 1794.650 2796.350 ;
        RECT 336.990 2794.610 337.370 2794.620 ;
        RECT 337.705 2794.610 338.035 2794.625 ;
        RECT 336.990 2794.310 338.035 2794.610 ;
        RECT 336.990 2794.300 337.370 2794.310 ;
        RECT 337.705 2794.295 338.035 2794.310 ;
        RECT 342.510 2794.610 342.890 2794.620 ;
        RECT 344.605 2794.610 344.935 2794.625 ;
        RECT 351.045 2794.620 351.375 2794.625 ;
        RECT 358.405 2794.620 358.735 2794.625 ;
        RECT 342.510 2794.310 344.935 2794.610 ;
        RECT 342.510 2794.300 342.890 2794.310 ;
        RECT 344.605 2794.295 344.935 2794.310 ;
        RECT 350.790 2794.610 351.375 2794.620 ;
        RECT 358.150 2794.610 358.735 2794.620 ;
        RECT 361.830 2794.610 362.210 2794.620 ;
        RECT 362.545 2794.610 362.875 2794.625 ;
        RECT 350.790 2794.310 351.600 2794.610 ;
        RECT 358.150 2794.310 358.960 2794.610 ;
        RECT 361.830 2794.310 362.875 2794.610 ;
        RECT 350.790 2794.300 351.375 2794.310 ;
        RECT 358.150 2794.300 358.735 2794.310 ;
        RECT 361.830 2794.300 362.210 2794.310 ;
        RECT 351.045 2794.295 351.375 2794.300 ;
        RECT 358.405 2794.295 358.735 2794.300 ;
        RECT 362.545 2794.295 362.875 2794.310 ;
        RECT 364.590 2794.610 364.970 2794.620 ;
        RECT 365.305 2794.610 365.635 2794.625 ;
        RECT 368.525 2794.620 368.855 2794.625 ;
        RECT 371.285 2794.620 371.615 2794.625 ;
        RECT 374.965 2794.620 375.295 2794.625 ;
        RECT 368.270 2794.610 368.855 2794.620 ;
        RECT 371.030 2794.610 371.615 2794.620 ;
        RECT 374.710 2794.610 375.295 2794.620 ;
        RECT 364.590 2794.310 365.635 2794.610 ;
        RECT 368.070 2794.310 368.855 2794.610 ;
        RECT 370.830 2794.310 371.615 2794.610 ;
        RECT 374.510 2794.310 375.295 2794.610 ;
        RECT 364.590 2794.300 364.970 2794.310 ;
        RECT 365.305 2794.295 365.635 2794.310 ;
        RECT 368.270 2794.300 368.855 2794.310 ;
        RECT 371.030 2794.300 371.615 2794.310 ;
        RECT 374.710 2794.300 375.295 2794.310 ;
        RECT 378.390 2794.610 378.770 2794.620 ;
        RECT 379.105 2794.610 379.435 2794.625 ;
        RECT 384.165 2794.620 384.495 2794.625 ;
        RECT 386.925 2794.620 387.255 2794.625 ;
        RECT 383.910 2794.610 384.495 2794.620 ;
        RECT 386.670 2794.610 387.255 2794.620 ;
        RECT 378.390 2794.310 379.435 2794.610 ;
        RECT 383.710 2794.310 384.495 2794.610 ;
        RECT 386.470 2794.310 387.255 2794.610 ;
        RECT 378.390 2794.300 378.770 2794.310 ;
        RECT 368.525 2794.295 368.855 2794.300 ;
        RECT 371.285 2794.295 371.615 2794.300 ;
        RECT 374.965 2794.295 375.295 2794.300 ;
        RECT 379.105 2794.295 379.435 2794.310 ;
        RECT 383.910 2794.300 384.495 2794.310 ;
        RECT 386.670 2794.300 387.255 2794.310 ;
        RECT 390.350 2794.610 390.730 2794.620 ;
        RECT 392.905 2794.610 393.235 2794.625 ;
        RECT 390.350 2794.310 393.235 2794.610 ;
        RECT 390.350 2794.300 390.730 2794.310 ;
        RECT 384.165 2794.295 384.495 2794.300 ;
        RECT 386.925 2794.295 387.255 2794.300 ;
        RECT 392.905 2794.295 393.235 2794.310 ;
        RECT 395.870 2794.610 396.250 2794.620 ;
        RECT 396.585 2794.610 396.915 2794.625 ;
        RECT 399.805 2794.620 400.135 2794.625 ;
        RECT 395.870 2794.310 396.915 2794.610 ;
        RECT 395.870 2794.300 396.250 2794.310 ;
        RECT 396.585 2794.295 396.915 2794.310 ;
        RECT 399.550 2794.610 400.135 2794.620 ;
        RECT 403.230 2794.610 403.610 2794.620 ;
        RECT 403.945 2794.610 404.275 2794.625 ;
        RECT 406.245 2794.620 406.575 2794.625 ;
        RECT 409.925 2794.620 410.255 2794.625 ;
        RECT 413.605 2794.620 413.935 2794.625 ;
        RECT 419.125 2794.620 419.455 2794.625 ;
        RECT 420.965 2794.620 421.295 2794.625 ;
        RECT 405.990 2794.610 406.575 2794.620 ;
        RECT 409.670 2794.610 410.255 2794.620 ;
        RECT 399.550 2794.310 400.360 2794.610 ;
        RECT 403.230 2794.310 404.275 2794.610 ;
        RECT 405.790 2794.310 406.575 2794.610 ;
        RECT 409.470 2794.310 410.255 2794.610 ;
        RECT 399.550 2794.300 400.135 2794.310 ;
        RECT 403.230 2794.300 403.610 2794.310 ;
        RECT 399.805 2794.295 400.135 2794.300 ;
        RECT 403.945 2794.295 404.275 2794.310 ;
        RECT 405.990 2794.300 406.575 2794.310 ;
        RECT 409.670 2794.300 410.255 2794.310 ;
        RECT 413.350 2794.610 413.935 2794.620 ;
        RECT 418.870 2794.610 419.455 2794.620 ;
        RECT 413.350 2794.310 414.160 2794.610 ;
        RECT 418.670 2794.310 419.455 2794.610 ;
        RECT 413.350 2794.300 413.935 2794.310 ;
        RECT 418.870 2794.300 419.455 2794.310 ;
        RECT 420.710 2794.610 421.295 2794.620 ;
        RECT 425.310 2794.610 425.690 2794.620 ;
        RECT 427.405 2794.610 427.735 2794.625 ;
        RECT 433.845 2794.620 434.175 2794.625 ;
        RECT 439.365 2794.620 439.695 2794.625 ;
        RECT 441.205 2794.620 441.535 2794.625 ;
        RECT 420.710 2794.310 421.520 2794.610 ;
        RECT 425.310 2794.310 427.735 2794.610 ;
        RECT 420.710 2794.300 421.295 2794.310 ;
        RECT 425.310 2794.300 425.690 2794.310 ;
        RECT 406.245 2794.295 406.575 2794.300 ;
        RECT 409.925 2794.295 410.255 2794.300 ;
        RECT 413.605 2794.295 413.935 2794.300 ;
        RECT 419.125 2794.295 419.455 2794.300 ;
        RECT 420.965 2794.295 421.295 2794.300 ;
        RECT 427.405 2794.295 427.735 2794.310 ;
        RECT 433.590 2794.610 434.175 2794.620 ;
        RECT 439.110 2794.610 439.695 2794.620 ;
        RECT 433.590 2794.310 434.400 2794.610 ;
        RECT 438.910 2794.310 439.695 2794.610 ;
        RECT 433.590 2794.300 434.175 2794.310 ;
        RECT 439.110 2794.300 439.695 2794.310 ;
        RECT 440.950 2794.610 441.535 2794.620 ;
        RECT 444.425 2794.620 444.755 2794.625 ;
        RECT 444.425 2794.610 445.010 2794.620 ;
        RECT 445.550 2794.610 445.930 2794.620 ;
        RECT 446.725 2794.610 447.055 2794.625 ;
        RECT 440.950 2794.310 441.760 2794.610 ;
        RECT 444.425 2794.310 445.210 2794.610 ;
        RECT 445.550 2794.310 447.055 2794.610 ;
        RECT 440.950 2794.300 441.535 2794.310 ;
        RECT 433.845 2794.295 434.175 2794.300 ;
        RECT 439.365 2794.295 439.695 2794.300 ;
        RECT 441.205 2794.295 441.535 2794.300 ;
        RECT 444.425 2794.300 445.010 2794.310 ;
        RECT 445.550 2794.300 445.930 2794.310 ;
        RECT 444.425 2794.295 444.755 2794.300 ;
        RECT 446.725 2794.295 447.055 2794.310 ;
        RECT 449.025 2794.620 449.355 2794.625 ;
        RECT 455.005 2794.620 455.335 2794.625 ;
        RECT 449.025 2794.610 449.610 2794.620 ;
        RECT 454.750 2794.610 455.335 2794.620 ;
        RECT 460.270 2794.610 460.650 2794.620 ;
        RECT 461.445 2794.610 461.775 2794.625 ;
        RECT 462.365 2794.620 462.695 2794.625 ;
        RECT 449.025 2794.310 449.810 2794.610 ;
        RECT 454.750 2794.310 455.560 2794.610 ;
        RECT 460.270 2794.310 461.775 2794.610 ;
        RECT 449.025 2794.300 449.610 2794.310 ;
        RECT 454.750 2794.300 455.335 2794.310 ;
        RECT 460.270 2794.300 460.650 2794.310 ;
        RECT 449.025 2794.295 449.355 2794.300 ;
        RECT 455.005 2794.295 455.335 2794.300 ;
        RECT 461.445 2794.295 461.775 2794.310 ;
        RECT 462.110 2794.610 462.695 2794.620 ;
        RECT 465.790 2794.610 466.170 2794.620 ;
        RECT 468.345 2794.610 468.675 2794.625 ;
        RECT 474.325 2794.620 474.655 2794.625 ;
        RECT 475.245 2794.620 475.575 2794.625 ;
        RECT 474.070 2794.610 474.655 2794.620 ;
        RECT 462.110 2794.310 462.920 2794.610 ;
        RECT 465.790 2794.310 468.675 2794.610 ;
        RECT 473.870 2794.310 474.655 2794.610 ;
        RECT 462.110 2794.300 462.695 2794.310 ;
        RECT 465.790 2794.300 466.170 2794.310 ;
        RECT 462.365 2794.295 462.695 2794.300 ;
        RECT 468.345 2794.295 468.675 2794.310 ;
        RECT 474.070 2794.300 474.655 2794.310 ;
        RECT 474.990 2794.610 475.575 2794.620 ;
        RECT 478.465 2794.620 478.795 2794.625 ;
        RECT 482.605 2794.620 482.935 2794.625 ;
        RECT 485.365 2794.620 485.695 2794.625 ;
        RECT 488.125 2794.620 488.455 2794.625 ;
        RECT 478.465 2794.610 479.050 2794.620 ;
        RECT 482.350 2794.610 482.935 2794.620 ;
        RECT 485.110 2794.610 485.695 2794.620 ;
        RECT 487.870 2794.610 488.455 2794.620 ;
        RECT 474.990 2794.310 475.800 2794.610 ;
        RECT 478.465 2794.310 479.250 2794.610 ;
        RECT 482.350 2794.310 483.160 2794.610 ;
        RECT 484.910 2794.310 485.695 2794.610 ;
        RECT 487.670 2794.310 488.455 2794.610 ;
        RECT 474.990 2794.300 475.575 2794.310 ;
        RECT 474.325 2794.295 474.655 2794.300 ;
        RECT 475.245 2794.295 475.575 2794.300 ;
        RECT 478.465 2794.300 479.050 2794.310 ;
        RECT 482.350 2794.300 482.935 2794.310 ;
        RECT 485.110 2794.300 485.695 2794.310 ;
        RECT 487.870 2794.300 488.455 2794.310 ;
        RECT 491.550 2794.610 491.930 2794.620 ;
        RECT 492.725 2794.610 493.055 2794.625 ;
        RECT 491.550 2794.310 493.055 2794.610 ;
        RECT 491.550 2794.300 491.930 2794.310 ;
        RECT 478.465 2794.295 478.795 2794.300 ;
        RECT 482.605 2794.295 482.935 2794.300 ;
        RECT 485.365 2794.295 485.695 2794.300 ;
        RECT 488.125 2794.295 488.455 2794.300 ;
        RECT 492.725 2794.295 493.055 2794.310 ;
        RECT 495.230 2794.610 495.610 2794.620 ;
        RECT 496.405 2794.610 496.735 2794.625 ;
        RECT 495.230 2794.310 496.735 2794.610 ;
        RECT 495.230 2794.300 495.610 2794.310 ;
        RECT 496.405 2794.295 496.735 2794.310 ;
        RECT 500.750 2794.610 501.130 2794.620 ;
        RECT 502.845 2794.610 503.175 2794.625 ;
        RECT 510.205 2794.620 510.535 2794.625 ;
        RECT 524.005 2794.620 524.335 2794.625 ;
        RECT 509.950 2794.610 510.535 2794.620 ;
        RECT 523.750 2794.610 524.335 2794.620 ;
        RECT 500.750 2794.310 503.175 2794.610 ;
        RECT 509.750 2794.310 510.535 2794.610 ;
        RECT 523.550 2794.310 524.335 2794.610 ;
        RECT 500.750 2794.300 501.130 2794.310 ;
        RECT 502.845 2794.295 503.175 2794.310 ;
        RECT 509.950 2794.300 510.535 2794.310 ;
        RECT 523.750 2794.300 524.335 2794.310 ;
        RECT 535.710 2794.610 536.090 2794.620 ;
        RECT 537.345 2794.610 537.675 2794.625 ;
        RECT 542.405 2794.620 542.735 2794.625 ;
        RECT 542.150 2794.610 542.735 2794.620 ;
        RECT 535.710 2794.310 537.675 2794.610 ;
        RECT 541.950 2794.310 542.735 2794.610 ;
        RECT 535.710 2794.300 536.090 2794.310 ;
        RECT 510.205 2794.295 510.535 2794.300 ;
        RECT 524.005 2794.295 524.335 2794.300 ;
        RECT 537.345 2794.295 537.675 2794.310 ;
        RECT 542.150 2794.300 542.735 2794.310 ;
        RECT 542.405 2794.295 542.735 2794.300 ;
        RECT 979.865 2794.610 980.195 2794.625 ;
        RECT 1001.025 2794.620 1001.355 2794.625 ;
        RECT 1007.465 2794.620 1007.795 2794.625 ;
        RECT 980.990 2794.610 981.370 2794.620 ;
        RECT 1001.025 2794.610 1001.610 2794.620 ;
        RECT 1007.465 2794.610 1008.050 2794.620 ;
        RECT 979.865 2794.310 981.370 2794.610 ;
        RECT 1000.800 2794.310 1001.610 2794.610 ;
        RECT 1007.240 2794.310 1008.050 2794.610 ;
        RECT 979.865 2794.295 980.195 2794.310 ;
        RECT 980.990 2794.300 981.370 2794.310 ;
        RECT 1001.025 2794.300 1001.610 2794.310 ;
        RECT 1007.465 2794.300 1008.050 2794.310 ;
        RECT 1013.190 2794.610 1013.570 2794.620 ;
        RECT 1013.905 2794.610 1014.235 2794.625 ;
        RECT 1018.965 2794.620 1019.295 2794.625 ;
        RECT 1018.710 2794.610 1019.295 2794.620 ;
        RECT 1013.190 2794.310 1014.235 2794.610 ;
        RECT 1018.510 2794.310 1019.295 2794.610 ;
        RECT 1013.190 2794.300 1013.570 2794.310 ;
        RECT 1001.025 2794.295 1001.355 2794.300 ;
        RECT 1007.465 2794.295 1007.795 2794.300 ;
        RECT 1013.905 2794.295 1014.235 2794.310 ;
        RECT 1018.710 2794.300 1019.295 2794.310 ;
        RECT 1019.630 2794.610 1020.010 2794.620 ;
        RECT 1020.805 2794.610 1021.135 2794.625 ;
        RECT 1019.630 2794.310 1021.135 2794.610 ;
        RECT 1019.630 2794.300 1020.010 2794.310 ;
        RECT 1018.965 2794.295 1019.295 2794.300 ;
        RECT 1020.805 2794.295 1021.135 2794.310 ;
        RECT 1026.990 2794.610 1027.370 2794.620 ;
        RECT 1027.705 2794.610 1028.035 2794.625 ;
        RECT 1026.990 2794.310 1028.035 2794.610 ;
        RECT 1026.990 2794.300 1027.370 2794.310 ;
        RECT 1027.705 2794.295 1028.035 2794.310 ;
        RECT 1030.670 2794.610 1031.050 2794.620 ;
        RECT 1031.845 2794.610 1032.175 2794.625 ;
        RECT 1030.670 2794.310 1032.175 2794.610 ;
        RECT 1030.670 2794.300 1031.050 2794.310 ;
        RECT 1031.845 2794.295 1032.175 2794.310 ;
        RECT 1041.710 2794.610 1042.090 2794.620 ;
        RECT 1042.425 2794.610 1042.755 2794.625 ;
        RECT 1059.445 2794.620 1059.775 2794.625 ;
        RECT 1059.190 2794.610 1059.775 2794.620 ;
        RECT 1041.710 2794.310 1042.755 2794.610 ;
        RECT 1058.990 2794.310 1059.775 2794.610 ;
        RECT 1041.710 2794.300 1042.090 2794.310 ;
        RECT 1042.425 2794.295 1042.755 2794.310 ;
        RECT 1059.190 2794.300 1059.775 2794.310 ;
        RECT 1059.445 2794.295 1059.775 2794.300 ;
        RECT 1065.425 2794.620 1065.755 2794.625 ;
        RECT 1065.425 2794.610 1066.010 2794.620 ;
        RECT 1069.565 2794.610 1069.895 2794.625 ;
        RECT 1076.465 2794.620 1076.795 2794.625 ;
        RECT 1093.945 2794.620 1094.275 2794.625 ;
        RECT 1100.385 2794.620 1100.715 2794.625 ;
        RECT 1105.445 2794.620 1105.775 2794.625 ;
        RECT 1070.230 2794.610 1070.610 2794.620 ;
        RECT 1065.425 2794.310 1066.210 2794.610 ;
        RECT 1069.565 2794.310 1070.610 2794.610 ;
        RECT 1065.425 2794.300 1066.010 2794.310 ;
        RECT 1065.425 2794.295 1065.755 2794.300 ;
        RECT 1069.565 2794.295 1069.895 2794.310 ;
        RECT 1070.230 2794.300 1070.610 2794.310 ;
        RECT 1076.465 2794.610 1077.050 2794.620 ;
        RECT 1093.945 2794.610 1094.530 2794.620 ;
        RECT 1100.385 2794.610 1100.970 2794.620 ;
        RECT 1105.190 2794.610 1105.775 2794.620 ;
        RECT 1076.465 2794.310 1077.250 2794.610 ;
        RECT 1093.945 2794.310 1094.730 2794.610 ;
        RECT 1100.385 2794.310 1101.170 2794.610 ;
        RECT 1104.990 2794.310 1105.775 2794.610 ;
        RECT 1076.465 2794.300 1077.050 2794.310 ;
        RECT 1093.945 2794.300 1094.530 2794.310 ;
        RECT 1100.385 2794.300 1100.970 2794.310 ;
        RECT 1105.190 2794.300 1105.775 2794.310 ;
        RECT 1076.465 2794.295 1076.795 2794.300 ;
        RECT 1093.945 2794.295 1094.275 2794.300 ;
        RECT 1100.385 2794.295 1100.715 2794.300 ;
        RECT 1105.445 2794.295 1105.775 2794.300 ;
        RECT 1111.425 2794.620 1111.755 2794.625 ;
        RECT 1117.865 2794.620 1118.195 2794.625 ;
        RECT 1111.425 2794.610 1112.010 2794.620 ;
        RECT 1117.865 2794.610 1118.450 2794.620 ;
        RECT 1119.705 2794.610 1120.035 2794.625 ;
        RECT 1140.405 2794.620 1140.735 2794.625 ;
        RECT 1122.670 2794.610 1123.050 2794.620 ;
        RECT 1140.150 2794.610 1140.735 2794.620 ;
        RECT 1111.425 2794.310 1112.210 2794.610 ;
        RECT 1117.865 2794.310 1118.650 2794.610 ;
        RECT 1119.705 2794.310 1123.050 2794.610 ;
        RECT 1139.950 2794.310 1140.735 2794.610 ;
        RECT 1111.425 2794.300 1112.010 2794.310 ;
        RECT 1117.865 2794.300 1118.450 2794.310 ;
        RECT 1111.425 2794.295 1111.755 2794.300 ;
        RECT 1117.865 2794.295 1118.195 2794.300 ;
        RECT 1119.705 2794.295 1120.035 2794.310 ;
        RECT 1122.670 2794.300 1123.050 2794.310 ;
        RECT 1140.150 2794.300 1140.735 2794.310 ;
        RECT 1178.790 2794.610 1179.170 2794.620 ;
        RECT 1179.505 2794.610 1179.835 2794.625 ;
        RECT 1186.405 2794.620 1186.735 2794.625 ;
        RECT 1178.790 2794.310 1179.835 2794.610 ;
        RECT 1178.790 2794.300 1179.170 2794.310 ;
        RECT 1140.405 2794.295 1140.735 2794.300 ;
        RECT 1179.505 2794.295 1179.835 2794.310 ;
        RECT 1186.150 2794.610 1186.735 2794.620 ;
        RECT 1198.110 2794.610 1198.490 2794.620 ;
        RECT 1200.205 2794.610 1200.535 2794.625 ;
        RECT 1186.150 2794.310 1186.960 2794.610 ;
        RECT 1198.110 2794.310 1200.535 2794.610 ;
        RECT 1186.150 2794.300 1186.735 2794.310 ;
        RECT 1198.110 2794.300 1198.490 2794.310 ;
        RECT 1186.405 2794.295 1186.735 2794.300 ;
        RECT 1200.205 2794.295 1200.535 2794.310 ;
        RECT 1580.165 2794.610 1580.495 2794.625 ;
        RECT 1587.065 2794.620 1587.395 2794.625 ;
        RECT 1580.830 2794.610 1581.210 2794.620 ;
        RECT 1587.065 2794.610 1587.650 2794.620 ;
        RECT 1580.165 2794.310 1581.210 2794.610 ;
        RECT 1586.840 2794.310 1587.650 2794.610 ;
        RECT 1580.165 2794.295 1580.495 2794.310 ;
        RECT 1580.830 2794.300 1581.210 2794.310 ;
        RECT 1587.065 2794.300 1587.650 2794.310 ;
        RECT 1601.325 2794.610 1601.655 2794.625 ;
        RECT 1604.750 2794.610 1605.130 2794.620 ;
        RECT 1601.325 2794.310 1605.130 2794.610 ;
        RECT 1587.065 2794.295 1587.395 2794.300 ;
        RECT 1601.325 2794.295 1601.655 2794.310 ;
        RECT 1604.750 2794.300 1605.130 2794.310 ;
        RECT 1613.030 2794.610 1613.410 2794.620 ;
        RECT 1614.205 2794.610 1614.535 2794.625 ;
        RECT 1613.030 2794.310 1614.535 2794.610 ;
        RECT 1613.030 2794.300 1613.410 2794.310 ;
        RECT 1614.205 2794.295 1614.535 2794.310 ;
        RECT 1617.425 2794.620 1617.755 2794.625 ;
        RECT 1642.725 2794.620 1643.055 2794.625 ;
        RECT 1617.425 2794.610 1618.010 2794.620 ;
        RECT 1642.470 2794.610 1643.055 2794.620 ;
        RECT 1617.425 2794.310 1618.210 2794.610 ;
        RECT 1642.270 2794.310 1643.055 2794.610 ;
        RECT 1617.425 2794.300 1618.010 2794.310 ;
        RECT 1642.470 2794.300 1643.055 2794.310 ;
        RECT 1617.425 2794.295 1617.755 2794.300 ;
        RECT 1642.725 2794.295 1643.055 2794.300 ;
        RECT 1647.785 2794.620 1648.115 2794.625 ;
        RECT 1652.385 2794.620 1652.715 2794.625 ;
        RECT 1647.785 2794.610 1648.370 2794.620 ;
        RECT 1652.385 2794.610 1652.970 2794.620 ;
        RECT 1659.030 2794.610 1659.410 2794.620 ;
        RECT 1662.505 2794.610 1662.835 2794.625 ;
        RECT 1665.725 2794.620 1666.055 2794.625 ;
        RECT 1665.470 2794.610 1666.055 2794.620 ;
        RECT 1647.785 2794.310 1648.570 2794.610 ;
        RECT 1652.385 2794.310 1653.170 2794.610 ;
        RECT 1659.030 2794.310 1662.835 2794.610 ;
        RECT 1665.270 2794.310 1666.055 2794.610 ;
        RECT 1647.785 2794.300 1648.370 2794.310 ;
        RECT 1652.385 2794.300 1652.970 2794.310 ;
        RECT 1659.030 2794.300 1659.410 2794.310 ;
        RECT 1647.785 2794.295 1648.115 2794.300 ;
        RECT 1652.385 2794.295 1652.715 2794.300 ;
        RECT 1662.505 2794.295 1662.835 2794.310 ;
        RECT 1665.470 2794.300 1666.055 2794.310 ;
        RECT 1670.070 2794.610 1670.450 2794.620 ;
        RECT 1671.245 2794.610 1671.575 2794.625 ;
        RECT 1670.070 2794.310 1671.575 2794.610 ;
        RECT 1670.070 2794.300 1670.450 2794.310 ;
        RECT 1665.725 2794.295 1666.055 2794.300 ;
        RECT 1671.245 2794.295 1671.575 2794.310 ;
        RECT 1677.430 2794.610 1677.810 2794.620 ;
        RECT 1679.525 2794.610 1679.855 2794.625 ;
        RECT 1677.430 2794.310 1679.855 2794.610 ;
        RECT 1677.430 2794.300 1677.810 2794.310 ;
        RECT 1679.525 2794.295 1679.855 2794.310 ;
        RECT 1681.365 2794.610 1681.695 2794.625 ;
        RECT 1688.725 2794.620 1689.055 2794.625 ;
        RECT 1695.165 2794.620 1695.495 2794.625 ;
        RECT 1682.030 2794.610 1682.410 2794.620 ;
        RECT 1688.470 2794.610 1689.055 2794.620 ;
        RECT 1694.910 2794.610 1695.495 2794.620 ;
        RECT 1681.365 2794.310 1682.410 2794.610 ;
        RECT 1688.270 2794.310 1689.055 2794.610 ;
        RECT 1694.710 2794.310 1695.495 2794.610 ;
        RECT 1681.365 2794.295 1681.695 2794.310 ;
        RECT 1682.030 2794.300 1682.410 2794.310 ;
        RECT 1688.470 2794.300 1689.055 2794.310 ;
        RECT 1694.910 2794.300 1695.495 2794.310 ;
        RECT 1688.725 2794.295 1689.055 2794.300 ;
        RECT 1695.165 2794.295 1695.495 2794.300 ;
        RECT 1699.305 2794.620 1699.635 2794.625 ;
        RECT 1706.205 2794.620 1706.535 2794.625 ;
        RECT 1712.645 2794.620 1712.975 2794.625 ;
        RECT 1718.165 2794.620 1718.495 2794.625 ;
        RECT 1699.305 2794.610 1699.890 2794.620 ;
        RECT 1705.950 2794.610 1706.535 2794.620 ;
        RECT 1712.390 2794.610 1712.975 2794.620 ;
        RECT 1717.910 2794.610 1718.495 2794.620 ;
        RECT 1699.305 2794.310 1700.090 2794.610 ;
        RECT 1705.750 2794.310 1706.535 2794.610 ;
        RECT 1712.190 2794.310 1712.975 2794.610 ;
        RECT 1717.710 2794.310 1718.495 2794.610 ;
        RECT 1699.305 2794.300 1699.890 2794.310 ;
        RECT 1705.950 2794.300 1706.535 2794.310 ;
        RECT 1712.390 2794.300 1712.975 2794.310 ;
        RECT 1717.910 2794.300 1718.495 2794.310 ;
        RECT 1723.430 2794.610 1723.810 2794.620 ;
        RECT 1724.145 2794.610 1724.475 2794.625 ;
        RECT 1723.430 2794.310 1724.475 2794.610 ;
        RECT 1723.430 2794.300 1723.810 2794.310 ;
        RECT 1699.305 2794.295 1699.635 2794.300 ;
        RECT 1706.205 2794.295 1706.535 2794.300 ;
        RECT 1712.645 2794.295 1712.975 2794.300 ;
        RECT 1718.165 2794.295 1718.495 2794.300 ;
        RECT 1724.145 2794.295 1724.475 2794.310 ;
        RECT 1728.745 2794.620 1729.075 2794.625 ;
        RECT 1732.425 2794.620 1732.755 2794.625 ;
        RECT 1741.165 2794.620 1741.495 2794.625 ;
        RECT 1728.745 2794.610 1729.330 2794.620 ;
        RECT 1732.425 2794.610 1733.010 2794.620 ;
        RECT 1740.910 2794.610 1741.495 2794.620 ;
        RECT 1728.745 2794.310 1729.530 2794.610 ;
        RECT 1732.425 2794.310 1733.210 2794.610 ;
        RECT 1740.710 2794.310 1741.495 2794.610 ;
        RECT 1728.745 2794.300 1729.330 2794.310 ;
        RECT 1732.425 2794.300 1733.010 2794.310 ;
        RECT 1740.910 2794.300 1741.495 2794.310 ;
        RECT 1728.745 2794.295 1729.075 2794.300 ;
        RECT 1732.425 2794.295 1732.755 2794.300 ;
        RECT 1741.165 2794.295 1741.495 2794.300 ;
        RECT 1746.685 2794.610 1747.015 2794.625 ;
        RECT 1752.665 2794.620 1752.995 2794.625 ;
        RECT 1747.350 2794.610 1747.730 2794.620 ;
        RECT 1746.685 2794.310 1747.730 2794.610 ;
        RECT 1746.685 2794.295 1747.015 2794.310 ;
        RECT 1747.350 2794.300 1747.730 2794.310 ;
        RECT 1752.665 2794.610 1753.250 2794.620 ;
        RECT 1760.025 2794.610 1760.355 2794.625 ;
        RECT 1762.070 2794.610 1762.450 2794.620 ;
        RECT 1752.665 2794.310 1753.450 2794.610 ;
        RECT 1760.025 2794.310 1762.450 2794.610 ;
        RECT 1752.665 2794.300 1753.250 2794.310 ;
        RECT 1752.665 2794.295 1752.995 2794.300 ;
        RECT 1760.025 2794.295 1760.355 2794.310 ;
        RECT 1762.070 2794.300 1762.450 2794.310 ;
        RECT 1766.465 2794.610 1766.795 2794.625 ;
        RECT 1767.590 2794.610 1767.970 2794.620 ;
        RECT 1766.465 2794.310 1767.970 2794.610 ;
        RECT 1766.465 2794.295 1766.795 2794.310 ;
        RECT 1767.590 2794.300 1767.970 2794.310 ;
        RECT 2228.765 2794.610 2229.095 2794.625 ;
        RECT 2231.270 2794.610 2231.650 2794.620 ;
        RECT 2228.765 2794.310 2231.650 2794.610 ;
        RECT 2228.765 2794.295 2229.095 2794.310 ;
        RECT 2231.270 2794.300 2231.650 2794.310 ;
        RECT 2237.965 2794.610 2238.295 2794.625 ;
        RECT 2268.325 2794.620 2268.655 2794.625 ;
        RECT 2238.630 2794.610 2239.010 2794.620 ;
        RECT 2268.070 2794.610 2268.655 2794.620 ;
        RECT 2237.965 2794.310 2239.010 2794.610 ;
        RECT 2267.870 2794.310 2268.655 2794.610 ;
        RECT 2237.965 2794.295 2238.295 2794.310 ;
        RECT 2238.630 2794.300 2239.010 2794.310 ;
        RECT 2268.070 2794.300 2268.655 2794.310 ;
        RECT 2268.325 2794.295 2268.655 2794.300 ;
        RECT 2273.385 2794.620 2273.715 2794.625 ;
        RECT 2279.825 2794.620 2280.155 2794.625 ;
        RECT 2286.725 2794.620 2287.055 2794.625 ;
        RECT 2291.325 2794.620 2291.655 2794.625 ;
        RECT 2304.205 2794.620 2304.535 2794.625 ;
        RECT 2273.385 2794.610 2273.970 2794.620 ;
        RECT 2279.825 2794.610 2280.410 2794.620 ;
        RECT 2286.470 2794.610 2287.055 2794.620 ;
        RECT 2291.070 2794.610 2291.655 2794.620 ;
        RECT 2303.950 2794.610 2304.535 2794.620 ;
        RECT 2273.385 2794.310 2274.170 2794.610 ;
        RECT 2279.825 2794.310 2280.610 2794.610 ;
        RECT 2286.270 2794.310 2287.055 2794.610 ;
        RECT 2290.870 2794.310 2291.655 2794.610 ;
        RECT 2303.750 2794.310 2304.535 2794.610 ;
        RECT 2273.385 2794.300 2273.970 2794.310 ;
        RECT 2279.825 2794.300 2280.410 2794.310 ;
        RECT 2286.470 2794.300 2287.055 2794.310 ;
        RECT 2291.070 2794.300 2291.655 2794.310 ;
        RECT 2303.950 2794.300 2304.535 2794.310 ;
        RECT 2273.385 2794.295 2273.715 2794.300 ;
        RECT 2279.825 2794.295 2280.155 2794.300 ;
        RECT 2286.725 2794.295 2287.055 2794.300 ;
        RECT 2291.325 2794.295 2291.655 2794.300 ;
        RECT 2304.205 2794.295 2304.535 2794.300 ;
        RECT 2308.345 2794.620 2308.675 2794.625 ;
        RECT 2312.945 2794.620 2313.275 2794.625 ;
        RECT 2321.225 2794.620 2321.555 2794.625 ;
        RECT 2326.285 2794.620 2326.615 2794.625 ;
        RECT 2308.345 2794.610 2308.930 2794.620 ;
        RECT 2312.945 2794.610 2313.530 2794.620 ;
        RECT 2321.225 2794.610 2321.810 2794.620 ;
        RECT 2326.030 2794.610 2326.615 2794.620 ;
        RECT 2308.345 2794.310 2309.130 2794.610 ;
        RECT 2312.945 2794.310 2313.730 2794.610 ;
        RECT 2321.225 2794.310 2322.010 2794.610 ;
        RECT 2325.830 2794.310 2326.615 2794.610 ;
        RECT 2308.345 2794.300 2308.930 2794.310 ;
        RECT 2312.945 2794.300 2313.530 2794.310 ;
        RECT 2321.225 2794.300 2321.810 2794.310 ;
        RECT 2326.030 2794.300 2326.615 2794.310 ;
        RECT 2308.345 2794.295 2308.675 2794.300 ;
        RECT 2312.945 2794.295 2313.275 2794.300 ;
        RECT 2321.225 2794.295 2321.555 2794.300 ;
        RECT 2326.285 2794.295 2326.615 2794.300 ;
        RECT 2332.265 2794.610 2332.595 2794.625 ;
        RECT 2334.310 2794.610 2334.690 2794.620 ;
        RECT 2332.265 2794.310 2334.690 2794.610 ;
        RECT 2332.265 2794.295 2332.595 2794.310 ;
        RECT 2334.310 2794.300 2334.690 2794.310 ;
        RECT 2339.165 2794.610 2339.495 2794.625 ;
        RECT 2343.305 2794.620 2343.635 2794.625 ;
        RECT 2339.830 2794.610 2340.210 2794.620 ;
        RECT 2339.165 2794.310 2340.210 2794.610 ;
        RECT 2339.165 2794.295 2339.495 2794.310 ;
        RECT 2339.830 2794.300 2340.210 2794.310 ;
        RECT 2343.305 2794.610 2343.890 2794.620 ;
        RECT 2346.065 2794.610 2346.395 2794.625 ;
        RECT 2351.790 2794.610 2352.170 2794.620 ;
        RECT 2343.305 2794.310 2344.090 2794.610 ;
        RECT 2346.065 2794.310 2352.170 2794.610 ;
        RECT 2343.305 2794.300 2343.890 2794.310 ;
        RECT 2343.305 2794.295 2343.635 2794.300 ;
        RECT 2346.065 2794.295 2346.395 2794.310 ;
        RECT 2351.790 2794.300 2352.170 2794.310 ;
        RECT 2352.965 2794.610 2353.295 2794.625 ;
        RECT 2357.310 2794.610 2357.690 2794.620 ;
        RECT 2352.965 2794.310 2357.690 2794.610 ;
        RECT 2352.965 2794.295 2353.295 2794.310 ;
        RECT 2357.310 2794.300 2357.690 2794.310 ;
        RECT 2359.865 2794.610 2360.195 2794.625 ;
        RECT 2363.750 2794.610 2364.130 2794.620 ;
        RECT 2359.865 2794.310 2364.130 2794.610 ;
        RECT 2359.865 2794.295 2360.195 2794.310 ;
        RECT 2363.750 2794.300 2364.130 2794.310 ;
        RECT 2366.765 2794.610 2367.095 2794.625 ;
        RECT 2374.125 2794.620 2374.455 2794.625 ;
        RECT 2370.190 2794.610 2370.570 2794.620 ;
        RECT 2373.870 2794.610 2374.455 2794.620 ;
        RECT 2366.765 2794.310 2370.570 2794.610 ;
        RECT 2373.670 2794.310 2374.455 2794.610 ;
        RECT 2366.765 2794.295 2367.095 2794.310 ;
        RECT 2370.190 2794.300 2370.570 2794.310 ;
        RECT 2373.870 2794.300 2374.455 2794.310 ;
        RECT 2374.125 2794.295 2374.455 2794.300 ;
        RECT 2377.345 2794.620 2377.675 2794.625 ;
        RECT 2385.625 2794.620 2385.955 2794.625 ;
        RECT 2391.145 2794.620 2391.475 2794.625 ;
        RECT 2394.825 2794.620 2395.155 2794.625 ;
        RECT 2377.345 2794.610 2377.930 2794.620 ;
        RECT 2385.625 2794.610 2386.210 2794.620 ;
        RECT 2391.145 2794.610 2391.730 2794.620 ;
        RECT 2394.825 2794.610 2395.410 2794.620 ;
        RECT 2402.645 2794.610 2402.975 2794.625 ;
        RECT 2404.230 2794.610 2404.610 2794.620 ;
        RECT 2377.345 2794.310 2378.130 2794.610 ;
        RECT 2385.625 2794.310 2386.410 2794.610 ;
        RECT 2391.145 2794.310 2391.930 2794.610 ;
        RECT 2394.825 2794.310 2395.610 2794.610 ;
        RECT 2402.645 2794.310 2404.610 2794.610 ;
        RECT 2377.345 2794.300 2377.930 2794.310 ;
        RECT 2385.625 2794.300 2386.210 2794.310 ;
        RECT 2391.145 2794.300 2391.730 2794.310 ;
        RECT 2394.825 2794.300 2395.410 2794.310 ;
        RECT 2377.345 2794.295 2377.675 2794.300 ;
        RECT 2385.625 2794.295 2385.955 2794.300 ;
        RECT 2391.145 2794.295 2391.475 2794.300 ;
        RECT 2394.825 2794.295 2395.155 2794.300 ;
        RECT 2402.645 2794.295 2402.975 2794.310 ;
        RECT 2404.230 2794.300 2404.610 2794.310 ;
        RECT 2415.065 2794.610 2415.395 2794.625 ;
        RECT 2418.030 2794.610 2418.410 2794.620 ;
        RECT 2415.065 2794.310 2418.410 2794.610 ;
        RECT 2415.065 2794.295 2415.395 2794.310 ;
        RECT 2418.030 2794.300 2418.410 2794.310 ;
        RECT 348.950 2793.930 349.330 2793.940 ;
        RECT 351.505 2793.930 351.835 2793.945 ;
        RECT 379.565 2793.940 379.895 2793.945 ;
        RECT 392.445 2793.940 392.775 2793.945 ;
        RECT 379.310 2793.930 379.895 2793.940 ;
        RECT 392.190 2793.930 392.775 2793.940 ;
        RECT 348.950 2793.630 351.835 2793.930 ;
        RECT 379.110 2793.630 379.895 2793.930 ;
        RECT 391.990 2793.630 392.775 2793.930 ;
        RECT 348.950 2793.620 349.330 2793.630 ;
        RECT 351.505 2793.615 351.835 2793.630 ;
        RECT 379.310 2793.620 379.895 2793.630 ;
        RECT 392.190 2793.620 392.775 2793.630 ;
        RECT 396.790 2793.930 397.170 2793.940 ;
        RECT 397.505 2793.930 397.835 2793.945 ;
        RECT 414.525 2793.940 414.855 2793.945 ;
        RECT 414.270 2793.930 414.855 2793.940 ;
        RECT 396.790 2793.630 397.835 2793.930 ;
        RECT 414.070 2793.630 414.855 2793.930 ;
        RECT 396.790 2793.620 397.170 2793.630 ;
        RECT 379.565 2793.615 379.895 2793.620 ;
        RECT 392.445 2793.615 392.775 2793.620 ;
        RECT 397.505 2793.615 397.835 2793.630 ;
        RECT 414.270 2793.620 414.855 2793.630 ;
        RECT 414.525 2793.615 414.855 2793.620 ;
        RECT 426.945 2793.940 427.275 2793.945 ;
        RECT 426.945 2793.930 427.530 2793.940 ;
        RECT 430.830 2793.930 431.210 2793.940 ;
        RECT 434.305 2793.930 434.635 2793.945 ;
        RECT 426.945 2793.630 427.730 2793.930 ;
        RECT 430.830 2793.630 434.635 2793.930 ;
        RECT 426.945 2793.620 427.530 2793.630 ;
        RECT 430.830 2793.620 431.210 2793.630 ;
        RECT 426.945 2793.615 427.275 2793.620 ;
        RECT 434.305 2793.615 434.635 2793.630 ;
        RECT 455.465 2793.940 455.795 2793.945 ;
        RECT 468.805 2793.940 469.135 2793.945 ;
        RECT 455.465 2793.930 456.050 2793.940 ;
        RECT 468.550 2793.930 469.135 2793.940 ;
        RECT 455.465 2793.630 456.250 2793.930 ;
        RECT 468.350 2793.630 469.135 2793.930 ;
        RECT 455.465 2793.620 456.050 2793.630 ;
        RECT 468.550 2793.620 469.135 2793.630 ;
        RECT 455.465 2793.615 455.795 2793.620 ;
        RECT 468.805 2793.615 469.135 2793.620 ;
        RECT 524.465 2793.930 524.795 2793.945 ;
        RECT 526.510 2793.930 526.890 2793.940 ;
        RECT 524.465 2793.630 526.890 2793.930 ;
        RECT 524.465 2793.615 524.795 2793.630 ;
        RECT 526.510 2793.620 526.890 2793.630 ;
        RECT 1010.685 2793.930 1011.015 2793.945 ;
        RECT 1012.270 2793.930 1012.650 2793.940 ;
        RECT 1010.685 2793.630 1012.650 2793.930 ;
        RECT 1010.685 2793.615 1011.015 2793.630 ;
        RECT 1012.270 2793.620 1012.650 2793.630 ;
        RECT 1083.110 2793.930 1083.490 2793.940 ;
        RECT 1089.805 2793.930 1090.135 2793.945 ;
        RECT 1083.110 2793.630 1090.135 2793.930 ;
        RECT 1083.110 2793.620 1083.490 2793.630 ;
        RECT 1089.805 2793.615 1090.135 2793.630 ;
        RECT 1159.725 2793.930 1160.055 2793.945 ;
        RECT 1164.070 2793.930 1164.450 2793.940 ;
        RECT 1159.725 2793.630 1164.450 2793.930 ;
        RECT 1159.725 2793.615 1160.055 2793.630 ;
        RECT 1164.070 2793.620 1164.450 2793.630 ;
        RECT 1166.165 2793.930 1166.495 2793.945 ;
        RECT 1173.065 2793.940 1173.395 2793.945 ;
        RECT 1167.750 2793.930 1168.130 2793.940 ;
        RECT 1173.065 2793.930 1173.650 2793.940 ;
        RECT 1166.165 2793.630 1168.130 2793.930 ;
        RECT 1172.840 2793.630 1173.650 2793.930 ;
        RECT 1166.165 2793.615 1166.495 2793.630 ;
        RECT 1167.750 2793.620 1168.130 2793.630 ;
        RECT 1173.065 2793.620 1173.650 2793.630 ;
        RECT 1179.965 2793.930 1180.295 2793.945 ;
        RECT 1600.865 2793.940 1601.195 2793.945 ;
        RECT 1180.630 2793.930 1181.010 2793.940 ;
        RECT 1600.865 2793.930 1601.450 2793.940 ;
        RECT 1179.965 2793.630 1181.010 2793.930 ;
        RECT 1600.640 2793.630 1601.450 2793.930 ;
        RECT 1173.065 2793.615 1173.395 2793.620 ;
        RECT 1179.965 2793.615 1180.295 2793.630 ;
        RECT 1180.630 2793.620 1181.010 2793.630 ;
        RECT 1600.865 2793.620 1601.450 2793.630 ;
        RECT 1773.365 2793.930 1773.695 2793.945 ;
        RECT 1780.265 2793.940 1780.595 2793.945 ;
        RECT 1774.030 2793.930 1774.410 2793.940 ;
        RECT 1780.265 2793.930 1780.850 2793.940 ;
        RECT 1773.365 2793.630 1774.410 2793.930 ;
        RECT 1780.040 2793.630 1780.850 2793.930 ;
        RECT 1600.865 2793.615 1601.195 2793.620 ;
        RECT 1773.365 2793.615 1773.695 2793.630 ;
        RECT 1774.030 2793.620 1774.410 2793.630 ;
        RECT 1780.265 2793.620 1780.850 2793.630 ;
        RECT 2263.265 2793.930 2263.595 2793.945 ;
        RECT 2332.725 2793.940 2333.055 2793.945 ;
        RECT 2268.990 2793.930 2269.370 2793.940 ;
        RECT 2332.470 2793.930 2333.055 2793.940 ;
        RECT 2263.265 2793.630 2269.370 2793.930 ;
        RECT 2332.270 2793.630 2333.055 2793.930 ;
        RECT 1780.265 2793.615 1780.595 2793.620 ;
        RECT 2263.265 2793.615 2263.595 2793.630 ;
        RECT 2268.990 2793.620 2269.370 2793.630 ;
        RECT 2332.470 2793.620 2333.055 2793.630 ;
        RECT 2332.725 2793.615 2333.055 2793.620 ;
        RECT 2339.625 2793.930 2339.955 2793.945 ;
        RECT 2350.205 2793.940 2350.535 2793.945 ;
        RECT 2356.645 2793.940 2356.975 2793.945 ;
        RECT 2345.350 2793.930 2345.730 2793.940 ;
        RECT 2349.950 2793.930 2350.535 2793.940 ;
        RECT 2356.390 2793.930 2356.975 2793.940 ;
        RECT 2339.625 2793.630 2345.730 2793.930 ;
        RECT 2349.750 2793.630 2350.535 2793.930 ;
        RECT 2356.190 2793.630 2356.975 2793.930 ;
        RECT 2339.625 2793.615 2339.955 2793.630 ;
        RECT 2345.350 2793.620 2345.730 2793.630 ;
        RECT 2349.950 2793.620 2350.535 2793.630 ;
        RECT 2356.390 2793.620 2356.975 2793.630 ;
        RECT 2350.205 2793.615 2350.535 2793.620 ;
        RECT 2356.645 2793.615 2356.975 2793.620 ;
        RECT 2360.785 2793.940 2361.115 2793.945 ;
        RECT 2360.785 2793.930 2361.370 2793.940 ;
        RECT 2401.725 2793.930 2402.055 2793.945 ;
        RECT 2408.165 2793.940 2408.495 2793.945 ;
        RECT 2402.390 2793.930 2402.770 2793.940 ;
        RECT 2360.785 2793.630 2361.570 2793.930 ;
        RECT 2401.725 2793.630 2402.770 2793.930 ;
        RECT 2360.785 2793.620 2361.370 2793.630 ;
        RECT 2360.785 2793.615 2361.115 2793.620 ;
        RECT 2401.725 2793.615 2402.055 2793.630 ;
        RECT 2402.390 2793.620 2402.770 2793.630 ;
        RECT 2407.910 2793.930 2408.495 2793.940 ;
        RECT 2407.910 2793.630 2408.720 2793.930 ;
        RECT 2407.910 2793.620 2408.495 2793.630 ;
        RECT 2408.165 2793.615 2408.495 2793.620 ;
        RECT 431.750 2793.250 432.130 2793.260 ;
        RECT 433.385 2793.250 433.715 2793.265 ;
        RECT 467.885 2793.260 468.215 2793.265 ;
        RECT 1024.485 2793.260 1024.815 2793.265 ;
        RECT 467.630 2793.250 468.215 2793.260 ;
        RECT 1024.230 2793.250 1024.815 2793.260 ;
        RECT 431.750 2792.950 433.715 2793.250 ;
        RECT 467.430 2792.950 468.215 2793.250 ;
        RECT 1024.030 2792.950 1024.815 2793.250 ;
        RECT 431.750 2792.940 432.130 2792.950 ;
        RECT 433.385 2792.935 433.715 2792.950 ;
        RECT 467.630 2792.940 468.215 2792.950 ;
        RECT 1024.230 2792.940 1024.815 2792.950 ;
        RECT 467.885 2792.935 468.215 2792.940 ;
        RECT 1024.485 2792.935 1024.815 2792.940 ;
        RECT 1052.545 2793.260 1052.875 2793.265 ;
        RECT 1052.545 2793.250 1053.130 2793.260 ;
        RECT 1055.765 2793.250 1056.095 2793.265 ;
        RECT 1087.710 2793.250 1088.090 2793.260 ;
        RECT 1103.605 2793.250 1103.935 2793.265 ;
        RECT 1159.265 2793.260 1159.595 2793.265 ;
        RECT 1186.865 2793.260 1187.195 2793.265 ;
        RECT 1159.265 2793.250 1159.850 2793.260 ;
        RECT 1186.865 2793.250 1187.450 2793.260 ;
        RECT 1052.545 2792.950 1053.330 2793.250 ;
        RECT 1055.765 2792.950 1103.935 2793.250 ;
        RECT 1159.040 2792.950 1159.850 2793.250 ;
        RECT 1186.640 2792.950 1187.450 2793.250 ;
        RECT 1052.545 2792.940 1053.130 2792.950 ;
        RECT 1052.545 2792.935 1052.875 2792.940 ;
        RECT 1055.765 2792.935 1056.095 2792.950 ;
        RECT 1087.710 2792.940 1088.090 2792.950 ;
        RECT 1103.605 2792.935 1103.935 2792.950 ;
        RECT 1159.265 2792.940 1159.850 2792.950 ;
        RECT 1186.865 2792.940 1187.450 2792.950 ;
        RECT 1462.865 2793.250 1463.195 2793.265 ;
        RECT 1510.705 2793.250 1511.035 2793.265 ;
        RECT 1462.865 2792.950 1511.035 2793.250 ;
        RECT 1159.265 2792.935 1159.595 2792.940 ;
        RECT 1186.865 2792.935 1187.195 2792.940 ;
        RECT 1462.865 2792.935 1463.195 2792.950 ;
        RECT 1510.705 2792.935 1511.035 2792.950 ;
        RECT 1593.965 2793.250 1594.295 2793.265 ;
        RECT 1594.630 2793.250 1595.010 2793.260 ;
        RECT 1593.965 2792.950 1595.010 2793.250 ;
        RECT 1593.965 2792.935 1594.295 2792.950 ;
        RECT 1594.630 2792.940 1595.010 2792.950 ;
        RECT 2263.470 2793.250 2263.850 2793.260 ;
        RECT 2266.485 2793.250 2266.815 2793.265 ;
        RECT 2269.705 2793.250 2270.035 2793.265 ;
        RECT 2263.470 2792.950 2270.035 2793.250 ;
        RECT 2263.470 2792.940 2263.850 2792.950 ;
        RECT 2266.485 2792.935 2266.815 2792.950 ;
        RECT 2269.705 2792.935 2270.035 2792.950 ;
        RECT 2297.510 2793.250 2297.890 2793.260 ;
        RECT 2298.225 2793.250 2298.555 2793.265 ;
        RECT 2314.785 2793.250 2315.115 2793.265 ;
        RECT 2297.510 2792.950 2315.115 2793.250 ;
        RECT 2297.510 2792.940 2297.890 2792.950 ;
        RECT 2298.225 2792.935 2298.555 2792.950 ;
        RECT 2314.785 2792.935 2315.115 2792.950 ;
        RECT 2338.910 2793.250 2339.290 2793.260 ;
        RECT 2340.085 2793.250 2340.415 2793.265 ;
        RECT 2338.910 2792.950 2340.415 2793.250 ;
        RECT 2338.910 2792.940 2339.290 2792.950 ;
        RECT 2340.085 2792.935 2340.415 2792.950 ;
        RECT 2367.225 2793.260 2367.555 2793.265 ;
        RECT 2367.225 2793.250 2367.810 2793.260 ;
        RECT 2421.965 2793.250 2422.295 2793.265 ;
        RECT 2442.665 2793.260 2442.995 2793.265 ;
        RECT 2423.550 2793.250 2423.930 2793.260 ;
        RECT 2442.665 2793.250 2443.250 2793.260 ;
        RECT 2367.225 2792.950 2368.010 2793.250 ;
        RECT 2421.965 2792.950 2423.930 2793.250 ;
        RECT 2442.440 2792.950 2443.250 2793.250 ;
        RECT 2367.225 2792.940 2367.810 2792.950 ;
        RECT 2367.225 2792.935 2367.555 2792.940 ;
        RECT 2421.965 2792.935 2422.295 2792.950 ;
        RECT 2423.550 2792.940 2423.930 2792.950 ;
        RECT 2442.665 2792.940 2443.250 2792.950 ;
        RECT 2442.665 2792.935 2442.995 2792.940 ;
        RECT 496.865 2792.580 497.195 2792.585 ;
        RECT 496.865 2792.570 497.450 2792.580 ;
        RECT 541.485 2792.570 541.815 2792.585 ;
        RECT 543.070 2792.570 543.450 2792.580 ;
        RECT 496.865 2792.270 497.650 2792.570 ;
        RECT 541.485 2792.270 543.450 2792.570 ;
        RECT 496.865 2792.260 497.450 2792.270 ;
        RECT 496.865 2792.255 497.195 2792.260 ;
        RECT 541.485 2792.255 541.815 2792.270 ;
        RECT 543.070 2792.260 543.450 2792.270 ;
        RECT 1152.365 2792.570 1152.695 2792.585 ;
        RECT 1153.030 2792.570 1153.410 2792.580 ;
        RECT 1152.365 2792.270 1153.410 2792.570 ;
        RECT 1152.365 2792.255 1152.695 2792.270 ;
        RECT 1153.030 2792.260 1153.410 2792.270 ;
        RECT 1787.165 2792.570 1787.495 2792.585 ;
        RECT 2249.465 2792.580 2249.795 2792.585 ;
        RECT 1787.830 2792.570 1788.210 2792.580 ;
        RECT 2249.465 2792.570 2250.050 2792.580 ;
        RECT 1787.165 2792.270 1788.210 2792.570 ;
        RECT 2249.240 2792.270 2250.050 2792.570 ;
        RECT 1787.165 2792.255 1787.495 2792.270 ;
        RECT 1787.830 2792.260 1788.210 2792.270 ;
        RECT 2249.465 2792.260 2250.050 2792.270 ;
        RECT 2380.565 2792.570 2380.895 2792.585 ;
        RECT 2386.750 2792.570 2387.130 2792.580 ;
        RECT 2380.565 2792.270 2387.130 2792.570 ;
        RECT 2249.465 2792.255 2249.795 2792.260 ;
        RECT 2380.565 2792.255 2380.895 2792.270 ;
        RECT 2386.750 2792.260 2387.130 2792.270 ;
        RECT 2408.165 2792.570 2408.495 2792.585 ;
        RECT 2410.670 2792.570 2411.050 2792.580 ;
        RECT 2408.165 2792.270 2411.050 2792.570 ;
        RECT 2408.165 2792.255 2408.495 2792.270 ;
        RECT 2410.670 2792.260 2411.050 2792.270 ;
        RECT 2428.865 2792.570 2429.195 2792.585 ;
        RECT 2429.990 2792.570 2430.370 2792.580 ;
        RECT 2428.865 2792.270 2430.370 2792.570 ;
        RECT 2428.865 2792.255 2429.195 2792.270 ;
        RECT 2429.990 2792.260 2430.370 2792.270 ;
        RECT 2435.765 2792.570 2436.095 2792.585 ;
        RECT 2436.430 2792.570 2436.810 2792.580 ;
        RECT 2435.765 2792.270 2436.810 2792.570 ;
        RECT 2435.765 2792.255 2436.095 2792.270 ;
        RECT 2436.430 2792.260 2436.810 2792.270 ;
        RECT 310.105 2791.890 310.435 2791.905 ;
        RECT 1193.765 2791.900 1194.095 2791.905 ;
        RECT 986.510 2791.890 986.890 2791.900 ;
        RECT 310.105 2791.590 986.890 2791.890 ;
        RECT 310.105 2791.575 310.435 2791.590 ;
        RECT 986.510 2791.580 986.890 2791.590 ;
        RECT 1193.510 2791.890 1194.095 2791.900 ;
        RECT 1783.485 2791.890 1783.815 2791.905 ;
        RECT 2381.025 2791.900 2381.355 2791.905 ;
        RECT 2374.790 2791.890 2375.170 2791.900 ;
        RECT 2381.025 2791.890 2381.610 2791.900 ;
        RECT 1193.510 2791.590 1194.320 2791.890 ;
        RECT 1783.485 2791.590 2375.170 2791.890 ;
        RECT 2380.800 2791.590 2381.610 2791.890 ;
        RECT 1193.510 2791.580 1194.095 2791.590 ;
        RECT 1193.765 2791.575 1194.095 2791.580 ;
        RECT 1783.485 2791.575 1783.815 2791.590 ;
        RECT 2374.790 2791.580 2375.170 2791.590 ;
        RECT 2381.025 2791.580 2381.610 2791.590 ;
        RECT 2387.465 2791.890 2387.795 2791.905 ;
        RECT 2392.270 2791.890 2392.650 2791.900 ;
        RECT 2387.465 2791.590 2392.650 2791.890 ;
        RECT 2381.025 2791.575 2381.355 2791.580 ;
        RECT 2387.465 2791.575 2387.795 2791.590 ;
        RECT 2392.270 2791.580 2392.650 2791.590 ;
        RECT 317.005 2791.210 317.335 2791.225 ;
        RECT 993.870 2791.210 994.250 2791.220 ;
        RECT 317.005 2790.910 994.250 2791.210 ;
        RECT 317.005 2790.895 317.335 2790.910 ;
        RECT 993.870 2790.900 994.250 2790.910 ;
        RECT 1418.245 2791.210 1418.575 2791.225 ;
        RECT 2242.310 2791.210 2242.690 2791.220 ;
        RECT 1418.245 2790.910 2242.690 2791.210 ;
        RECT 1418.245 2790.895 1418.575 2790.910 ;
        RECT 2242.310 2790.900 2242.690 2790.910 ;
        RECT 2394.365 2791.210 2394.695 2791.225 ;
        RECT 2398.710 2791.210 2399.090 2791.220 ;
        RECT 2394.365 2790.910 2399.090 2791.210 ;
        RECT 2394.365 2790.895 2394.695 2790.910 ;
        RECT 2398.710 2790.900 2399.090 2790.910 ;
        RECT 2415.065 2791.210 2415.395 2791.225 ;
        RECT 2417.110 2791.210 2417.490 2791.220 ;
        RECT 2415.065 2790.910 2417.490 2791.210 ;
        RECT 2415.065 2790.895 2415.395 2790.910 ;
        RECT 2417.110 2790.900 2417.490 2790.910 ;
        RECT 2421.965 2791.210 2422.295 2791.225 ;
        RECT 2428.150 2791.210 2428.530 2791.220 ;
        RECT 2421.965 2790.910 2428.530 2791.210 ;
        RECT 2421.965 2790.895 2422.295 2790.910 ;
        RECT 2428.150 2790.900 2428.530 2790.910 ;
        RECT 2428.865 2791.210 2429.195 2791.225 ;
        RECT 2434.590 2791.210 2434.970 2791.220 ;
        RECT 2428.865 2790.910 2434.970 2791.210 ;
        RECT 2428.865 2790.895 2429.195 2790.910 ;
        RECT 2434.590 2790.900 2434.970 2790.910 ;
        RECT 1191.670 2790.530 1192.050 2790.540 ;
        RECT 1193.305 2790.530 1193.635 2790.545 ;
        RECT 1191.670 2790.230 1193.635 2790.530 ;
        RECT 1191.670 2790.220 1192.050 2790.230 ;
        RECT 1193.305 2790.215 1193.635 2790.230 ;
        RECT 2256.365 2790.530 2256.695 2790.545 ;
        RECT 2257.030 2790.530 2257.410 2790.540 ;
        RECT 2256.365 2790.230 2257.410 2790.530 ;
        RECT 2256.365 2790.215 2256.695 2790.230 ;
        RECT 2257.030 2790.220 2257.410 2790.230 ;
        RECT 2415.525 2790.530 2415.855 2790.545 ;
        RECT 2420.790 2790.530 2421.170 2790.540 ;
        RECT 2415.525 2790.230 2421.170 2790.530 ;
        RECT 2415.525 2790.215 2415.855 2790.230 ;
        RECT 2420.790 2790.220 2421.170 2790.230 ;
        RECT 2442.665 2790.530 2442.995 2790.545 ;
        RECT 2445.630 2790.530 2446.010 2790.540 ;
        RECT 2442.665 2790.230 2446.010 2790.530 ;
        RECT 2442.665 2790.215 2442.995 2790.230 ;
        RECT 2445.630 2790.220 2446.010 2790.230 ;
        RECT 2435.765 2789.850 2436.095 2789.865 ;
        RECT 2439.190 2789.850 2439.570 2789.860 ;
        RECT 2435.765 2789.550 2439.570 2789.850 ;
        RECT 2435.765 2789.535 2436.095 2789.550 ;
        RECT 2439.190 2789.540 2439.570 2789.550 ;
        RECT 500.085 2789.170 500.415 2789.185 ;
        RECT 501.670 2789.170 502.050 2789.180 ;
        RECT 500.085 2788.870 502.050 2789.170 ;
        RECT 500.085 2788.855 500.415 2788.870 ;
        RECT 501.670 2788.860 502.050 2788.870 ;
        RECT 504.225 2788.490 504.555 2788.505 ;
        RECT 506.985 2788.490 507.315 2788.505 ;
        RECT 531.365 2788.500 531.695 2788.505 ;
        RECT 508.110 2788.490 508.490 2788.500 ;
        RECT 531.110 2788.490 531.695 2788.500 ;
        RECT 534.585 2788.490 534.915 2788.505 ;
        RECT 504.225 2788.190 508.490 2788.490 ;
        RECT 530.730 2788.190 534.915 2788.490 ;
        RECT 504.225 2788.175 504.555 2788.190 ;
        RECT 506.985 2788.175 507.315 2788.190 ;
        RECT 508.110 2788.180 508.490 2788.190 ;
        RECT 531.110 2788.180 531.695 2788.190 ;
        RECT 531.365 2788.175 531.695 2788.180 ;
        RECT 534.585 2788.175 534.915 2788.190 ;
        RECT 1035.270 2788.490 1035.650 2788.500 ;
        RECT 1038.285 2788.490 1038.615 2788.505 ;
        RECT 1035.270 2788.190 1038.615 2788.490 ;
        RECT 1035.270 2788.180 1035.650 2788.190 ;
        RECT 1038.285 2788.175 1038.615 2788.190 ;
        RECT 1045.185 2788.490 1045.515 2788.505 ;
        RECT 1048.150 2788.490 1048.530 2788.500 ;
        RECT 1045.185 2788.190 1048.530 2788.490 ;
        RECT 1045.185 2788.175 1045.515 2788.190 ;
        RECT 1048.150 2788.180 1048.530 2788.190 ;
        RECT 1051.830 2788.490 1052.210 2788.500 ;
        RECT 1054.845 2788.490 1055.175 2788.505 ;
        RECT 1051.830 2788.190 1055.175 2788.490 ;
        RECT 1051.830 2788.180 1052.210 2788.190 ;
        RECT 1054.845 2788.175 1055.175 2788.190 ;
        RECT 1086.790 2788.490 1087.170 2788.500 ;
        RECT 1089.345 2788.490 1089.675 2788.505 ;
        RECT 1086.790 2788.190 1089.675 2788.490 ;
        RECT 1086.790 2788.180 1087.170 2788.190 ;
        RECT 1089.345 2788.175 1089.675 2788.190 ;
        RECT 1128.190 2788.490 1128.570 2788.500 ;
        RECT 1131.205 2788.490 1131.535 2788.505 ;
        RECT 1128.190 2788.190 1131.535 2788.490 ;
        RECT 1128.190 2788.180 1128.570 2788.190 ;
        RECT 1131.205 2788.175 1131.535 2788.190 ;
        RECT 1163.150 2788.490 1163.530 2788.500 ;
        RECT 1165.705 2788.490 1166.035 2788.505 ;
        RECT 1163.150 2788.190 1166.035 2788.490 ;
        RECT 1163.150 2788.180 1163.530 2788.190 ;
        RECT 1165.705 2788.175 1166.035 2788.190 ;
        RECT 1624.070 2788.490 1624.450 2788.500 ;
        RECT 1624.785 2788.490 1625.115 2788.505 ;
        RECT 1624.070 2788.190 1625.115 2788.490 ;
        RECT 1624.070 2788.180 1624.450 2788.190 ;
        RECT 1624.785 2788.175 1625.115 2788.190 ;
        RECT 1630.510 2788.490 1630.890 2788.500 ;
        RECT 1631.685 2788.490 1632.015 2788.505 ;
        RECT 1630.510 2788.190 1632.015 2788.490 ;
        RECT 1630.510 2788.180 1630.890 2788.190 ;
        RECT 1631.685 2788.175 1632.015 2788.190 ;
        RECT 1635.110 2788.490 1635.490 2788.500 ;
        RECT 1638.585 2788.490 1638.915 2788.505 ;
        RECT 1635.110 2788.190 1638.915 2788.490 ;
        RECT 1635.110 2788.180 1635.490 2788.190 ;
        RECT 1638.585 2788.175 1638.915 2788.190 ;
        RECT 1649.625 2788.490 1649.955 2788.505 ;
        RECT 1655.350 2788.490 1655.730 2788.500 ;
        RECT 1649.625 2788.190 1655.730 2788.490 ;
        RECT 1649.625 2788.175 1649.955 2788.190 ;
        RECT 1655.350 2788.180 1655.730 2788.190 ;
        RECT 1684.125 2788.490 1684.455 2788.505 ;
        RECT 1689.390 2788.490 1689.770 2788.500 ;
        RECT 1684.125 2788.190 1689.770 2788.490 ;
        RECT 1684.125 2788.175 1684.455 2788.190 ;
        RECT 1689.390 2788.180 1689.770 2788.190 ;
        RECT 1718.625 2788.490 1718.955 2788.505 ;
        RECT 1724.350 2788.490 1724.730 2788.500 ;
        RECT 1718.625 2788.190 1724.730 2788.490 ;
        RECT 1718.625 2788.175 1718.955 2788.190 ;
        RECT 1724.350 2788.180 1724.730 2788.190 ;
        RECT 1760.025 2788.490 1760.355 2788.505 ;
        RECT 1765.750 2788.490 1766.130 2788.500 ;
        RECT 1760.025 2788.190 1766.130 2788.490 ;
        RECT 1760.025 2788.175 1760.355 2788.190 ;
        RECT 1765.750 2788.180 1766.130 2788.190 ;
        RECT 2305.125 2788.490 2305.455 2788.505 ;
        RECT 2415.065 2788.500 2415.395 2788.505 ;
        RECT 2310.390 2788.490 2310.770 2788.500 ;
        RECT 2415.065 2788.490 2415.650 2788.500 ;
        RECT 2305.125 2788.190 2310.770 2788.490 ;
        RECT 2414.840 2788.190 2415.650 2788.490 ;
        RECT 2305.125 2788.175 2305.455 2788.190 ;
        RECT 2310.390 2788.180 2310.770 2788.190 ;
        RECT 2415.065 2788.180 2415.650 2788.190 ;
        RECT 2415.065 2788.175 2415.395 2788.180 ;
        RECT 507.190 2787.810 507.570 2787.820 ;
        RECT 510.205 2787.810 510.535 2787.825 ;
        RECT 513.885 2787.820 514.215 2787.825 ;
        RECT 513.630 2787.810 514.215 2787.820 ;
        RECT 507.190 2787.510 510.535 2787.810 ;
        RECT 513.430 2787.510 514.215 2787.810 ;
        RECT 507.190 2787.500 507.570 2787.510 ;
        RECT 510.205 2787.495 510.535 2787.510 ;
        RECT 513.630 2787.500 514.215 2787.510 ;
        RECT 516.390 2787.810 516.770 2787.820 ;
        RECT 517.105 2787.810 517.435 2787.825 ;
        RECT 516.390 2787.510 517.435 2787.810 ;
        RECT 516.390 2787.500 516.770 2787.510 ;
        RECT 513.885 2787.495 514.215 2787.500 ;
        RECT 517.105 2787.495 517.435 2787.510 ;
        RECT 520.070 2787.810 520.450 2787.820 ;
        RECT 520.785 2787.810 521.115 2787.825 ;
        RECT 520.070 2787.510 521.115 2787.810 ;
        RECT 520.070 2787.500 520.450 2787.510 ;
        RECT 520.785 2787.495 521.115 2787.510 ;
        RECT 526.510 2787.810 526.890 2787.820 ;
        RECT 527.685 2787.810 528.015 2787.825 ;
        RECT 526.510 2787.510 528.015 2787.810 ;
        RECT 526.510 2787.500 526.890 2787.510 ;
        RECT 527.685 2787.495 528.015 2787.510 ;
        RECT 530.190 2787.810 530.570 2787.820 ;
        RECT 530.905 2787.810 531.235 2787.825 ;
        RECT 538.265 2787.820 538.595 2787.825 ;
        RECT 538.265 2787.810 538.850 2787.820 ;
        RECT 542.405 2787.810 542.735 2787.825 ;
        RECT 530.190 2787.510 531.235 2787.810 ;
        RECT 537.860 2787.510 542.735 2787.810 ;
        RECT 530.190 2787.500 530.570 2787.510 ;
        RECT 530.905 2787.495 531.235 2787.510 ;
        RECT 538.265 2787.500 538.850 2787.510 ;
        RECT 538.265 2787.495 538.595 2787.500 ;
        RECT 542.405 2787.495 542.735 2787.510 ;
        RECT 544.910 2787.810 545.290 2787.820 ;
        RECT 551.605 2787.810 551.935 2787.825 ;
        RECT 1034.605 2787.820 1034.935 2787.825 ;
        RECT 544.910 2787.510 551.935 2787.810 ;
        RECT 544.910 2787.500 545.290 2787.510 ;
        RECT 551.605 2787.495 551.935 2787.510 ;
        RECT 1034.350 2787.810 1034.935 2787.820 ;
        RECT 1039.870 2787.810 1040.250 2787.820 ;
        RECT 1041.505 2787.810 1041.835 2787.825 ;
        RECT 1034.350 2787.510 1035.160 2787.810 ;
        RECT 1039.870 2787.510 1041.835 2787.810 ;
        RECT 1034.350 2787.500 1034.935 2787.510 ;
        RECT 1039.870 2787.500 1040.250 2787.510 ;
        RECT 1034.605 2787.495 1034.935 2787.500 ;
        RECT 1041.505 2787.495 1041.835 2787.510 ;
        RECT 1046.310 2787.810 1046.690 2787.820 ;
        RECT 1048.405 2787.810 1048.735 2787.825 ;
        RECT 1046.310 2787.510 1048.735 2787.810 ;
        RECT 1046.310 2787.500 1046.690 2787.510 ;
        RECT 1048.405 2787.495 1048.735 2787.510 ;
        RECT 1054.590 2787.810 1054.970 2787.820 ;
        RECT 1055.305 2787.810 1055.635 2787.825 ;
        RECT 1062.205 2787.820 1062.535 2787.825 ;
        RECT 1054.590 2787.510 1055.635 2787.810 ;
        RECT 1054.590 2787.500 1054.970 2787.510 ;
        RECT 1055.305 2787.495 1055.635 2787.510 ;
        RECT 1061.950 2787.810 1062.535 2787.820 ;
        RECT 1067.470 2787.810 1067.850 2787.820 ;
        RECT 1069.105 2787.810 1069.435 2787.825 ;
        RECT 1061.950 2787.510 1062.760 2787.810 ;
        RECT 1067.470 2787.510 1069.435 2787.810 ;
        RECT 1061.950 2787.500 1062.535 2787.510 ;
        RECT 1067.470 2787.500 1067.850 2787.510 ;
        RECT 1062.205 2787.495 1062.535 2787.500 ;
        RECT 1069.105 2787.495 1069.435 2787.510 ;
        RECT 1073.910 2787.810 1074.290 2787.820 ;
        RECT 1076.005 2787.810 1076.335 2787.825 ;
        RECT 1073.910 2787.510 1076.335 2787.810 ;
        RECT 1073.910 2787.500 1074.290 2787.510 ;
        RECT 1076.005 2787.495 1076.335 2787.510 ;
        RECT 1081.270 2787.810 1081.650 2787.820 ;
        RECT 1082.905 2787.810 1083.235 2787.825 ;
        RECT 1089.805 2787.820 1090.135 2787.825 ;
        RECT 1081.270 2787.510 1083.235 2787.810 ;
        RECT 1081.270 2787.500 1081.650 2787.510 ;
        RECT 1082.905 2787.495 1083.235 2787.510 ;
        RECT 1089.550 2787.810 1090.135 2787.820 ;
        RECT 1095.990 2787.810 1096.370 2787.820 ;
        RECT 1096.705 2787.810 1097.035 2787.825 ;
        RECT 1103.605 2787.820 1103.935 2787.825 ;
        RECT 1089.550 2787.510 1090.360 2787.810 ;
        RECT 1095.990 2787.510 1097.035 2787.810 ;
        RECT 1089.550 2787.500 1090.135 2787.510 ;
        RECT 1095.990 2787.500 1096.370 2787.510 ;
        RECT 1089.805 2787.495 1090.135 2787.500 ;
        RECT 1096.705 2787.495 1097.035 2787.510 ;
        RECT 1103.350 2787.810 1103.935 2787.820 ;
        RECT 1109.790 2787.810 1110.170 2787.820 ;
        RECT 1110.505 2787.810 1110.835 2787.825 ;
        RECT 1103.350 2787.510 1104.160 2787.810 ;
        RECT 1109.790 2787.510 1110.835 2787.810 ;
        RECT 1103.350 2787.500 1103.935 2787.510 ;
        RECT 1109.790 2787.500 1110.170 2787.510 ;
        RECT 1103.605 2787.495 1103.935 2787.500 ;
        RECT 1110.505 2787.495 1110.835 2787.510 ;
        RECT 1116.230 2787.810 1116.610 2787.820 ;
        RECT 1117.405 2787.810 1117.735 2787.825 ;
        RECT 1116.230 2787.510 1117.735 2787.810 ;
        RECT 1116.230 2787.500 1116.610 2787.510 ;
        RECT 1117.405 2787.495 1117.735 2787.510 ;
        RECT 1121.750 2787.810 1122.130 2787.820 ;
        RECT 1124.305 2787.810 1124.635 2787.825 ;
        RECT 1130.745 2787.820 1131.075 2787.825 ;
        RECT 1130.745 2787.810 1131.330 2787.820 ;
        RECT 1121.750 2787.510 1124.635 2787.810 ;
        RECT 1130.520 2787.510 1131.330 2787.810 ;
        RECT 1121.750 2787.500 1122.130 2787.510 ;
        RECT 1124.305 2787.495 1124.635 2787.510 ;
        RECT 1130.745 2787.500 1131.330 2787.510 ;
        RECT 1137.390 2787.810 1137.770 2787.820 ;
        RECT 1138.105 2787.810 1138.435 2787.825 ;
        RECT 1137.390 2787.510 1138.435 2787.810 ;
        RECT 1137.390 2787.500 1137.770 2787.510 ;
        RECT 1130.745 2787.495 1131.075 2787.500 ;
        RECT 1138.105 2787.495 1138.435 2787.510 ;
        RECT 1143.830 2787.810 1144.210 2787.820 ;
        RECT 1145.005 2787.810 1145.335 2787.825 ;
        RECT 1143.830 2787.510 1145.335 2787.810 ;
        RECT 1143.830 2787.500 1144.210 2787.510 ;
        RECT 1145.005 2787.495 1145.335 2787.510 ;
        RECT 1151.190 2787.810 1151.570 2787.820 ;
        RECT 1151.905 2787.810 1152.235 2787.825 ;
        RECT 1151.190 2787.510 1152.235 2787.810 ;
        RECT 1151.190 2787.500 1151.570 2787.510 ;
        RECT 1151.905 2787.495 1152.235 2787.510 ;
        RECT 1153.950 2787.810 1154.330 2787.820 ;
        RECT 1158.805 2787.810 1159.135 2787.825 ;
        RECT 1165.245 2787.820 1165.575 2787.825 ;
        RECT 1172.605 2787.820 1172.935 2787.825 ;
        RECT 1153.950 2787.510 1159.135 2787.810 ;
        RECT 1153.950 2787.500 1154.330 2787.510 ;
        RECT 1158.805 2787.495 1159.135 2787.510 ;
        RECT 1164.990 2787.810 1165.575 2787.820 ;
        RECT 1172.350 2787.810 1172.935 2787.820 ;
        RECT 1164.990 2787.510 1165.800 2787.810 ;
        RECT 1172.150 2787.510 1172.935 2787.810 ;
        RECT 1164.990 2787.500 1165.575 2787.510 ;
        RECT 1172.350 2787.500 1172.935 2787.510 ;
        RECT 1165.245 2787.495 1165.575 2787.500 ;
        RECT 1172.605 2787.495 1172.935 2787.500 ;
        RECT 1607.765 2787.810 1608.095 2787.825 ;
        RECT 1613.950 2787.810 1614.330 2787.820 ;
        RECT 1607.765 2787.510 1614.330 2787.810 ;
        RECT 1607.765 2787.495 1608.095 2787.510 ;
        RECT 1613.950 2787.500 1614.330 2787.510 ;
        RECT 1614.665 2787.810 1614.995 2787.825 ;
        RECT 1620.390 2787.810 1620.770 2787.820 ;
        RECT 1614.665 2787.510 1620.770 2787.810 ;
        RECT 1614.665 2787.495 1614.995 2787.510 ;
        RECT 1620.390 2787.500 1620.770 2787.510 ;
        RECT 1621.565 2787.810 1621.895 2787.825 ;
        RECT 1626.830 2787.810 1627.210 2787.820 ;
        RECT 1621.565 2787.510 1627.210 2787.810 ;
        RECT 1621.565 2787.495 1621.895 2787.510 ;
        RECT 1626.830 2787.500 1627.210 2787.510 ;
        RECT 1628.465 2787.810 1628.795 2787.825 ;
        RECT 1631.430 2787.810 1631.810 2787.820 ;
        RECT 1628.465 2787.510 1631.810 2787.810 ;
        RECT 1628.465 2787.495 1628.795 2787.510 ;
        RECT 1631.430 2787.500 1631.810 2787.510 ;
        RECT 1635.365 2787.810 1635.695 2787.825 ;
        RECT 1637.870 2787.810 1638.250 2787.820 ;
        RECT 1635.365 2787.510 1638.250 2787.810 ;
        RECT 1635.365 2787.495 1635.695 2787.510 ;
        RECT 1637.870 2787.500 1638.250 2787.510 ;
        RECT 1642.265 2787.810 1642.595 2787.825 ;
        RECT 1649.165 2787.820 1649.495 2787.825 ;
        RECT 1644.310 2787.810 1644.690 2787.820 ;
        RECT 1642.265 2787.510 1644.690 2787.810 ;
        RECT 1642.265 2787.495 1642.595 2787.510 ;
        RECT 1644.310 2787.500 1644.690 2787.510 ;
        RECT 1648.910 2787.810 1649.495 2787.820 ;
        RECT 1656.065 2787.810 1656.395 2787.825 ;
        RECT 1661.790 2787.810 1662.170 2787.820 ;
        RECT 1648.910 2787.510 1649.720 2787.810 ;
        RECT 1656.065 2787.510 1662.170 2787.810 ;
        RECT 1648.910 2787.500 1649.495 2787.510 ;
        RECT 1649.165 2787.495 1649.495 2787.500 ;
        RECT 1656.065 2787.495 1656.395 2787.510 ;
        RECT 1661.790 2787.500 1662.170 2787.510 ;
        RECT 1662.965 2787.810 1663.295 2787.825 ;
        RECT 1666.390 2787.810 1666.770 2787.820 ;
        RECT 1662.965 2787.510 1666.770 2787.810 ;
        RECT 1662.965 2787.495 1663.295 2787.510 ;
        RECT 1666.390 2787.500 1666.770 2787.510 ;
        RECT 1669.865 2787.810 1670.195 2787.825 ;
        RECT 1672.830 2787.810 1673.210 2787.820 ;
        RECT 1669.865 2787.510 1673.210 2787.810 ;
        RECT 1669.865 2787.495 1670.195 2787.510 ;
        RECT 1672.830 2787.500 1673.210 2787.510 ;
        RECT 1676.765 2787.810 1677.095 2787.825 ;
        RECT 1683.665 2787.820 1683.995 2787.825 ;
        RECT 1679.270 2787.810 1679.650 2787.820 ;
        RECT 1683.665 2787.810 1684.250 2787.820 ;
        RECT 1676.765 2787.510 1679.650 2787.810 ;
        RECT 1683.440 2787.510 1684.250 2787.810 ;
        RECT 1676.765 2787.495 1677.095 2787.510 ;
        RECT 1679.270 2787.500 1679.650 2787.510 ;
        RECT 1683.665 2787.500 1684.250 2787.510 ;
        RECT 1690.565 2787.810 1690.895 2787.825 ;
        RECT 1695.830 2787.810 1696.210 2787.820 ;
        RECT 1690.565 2787.510 1696.210 2787.810 ;
        RECT 1683.665 2787.495 1683.995 2787.500 ;
        RECT 1690.565 2787.495 1690.895 2787.510 ;
        RECT 1695.830 2787.500 1696.210 2787.510 ;
        RECT 1697.465 2787.810 1697.795 2787.825 ;
        RECT 1702.270 2787.810 1702.650 2787.820 ;
        RECT 1697.465 2787.510 1702.650 2787.810 ;
        RECT 1697.465 2787.495 1697.795 2787.510 ;
        RECT 1702.270 2787.500 1702.650 2787.510 ;
        RECT 1704.365 2787.810 1704.695 2787.825 ;
        RECT 1708.710 2787.810 1709.090 2787.820 ;
        RECT 1704.365 2787.510 1709.090 2787.810 ;
        RECT 1704.365 2787.495 1704.695 2787.510 ;
        RECT 1708.710 2787.500 1709.090 2787.510 ;
        RECT 1711.265 2787.810 1711.595 2787.825 ;
        RECT 1713.310 2787.810 1713.690 2787.820 ;
        RECT 1711.265 2787.510 1713.690 2787.810 ;
        RECT 1711.265 2787.495 1711.595 2787.510 ;
        RECT 1713.310 2787.500 1713.690 2787.510 ;
        RECT 1718.165 2787.810 1718.495 2787.825 ;
        RECT 1719.750 2787.810 1720.130 2787.820 ;
        RECT 1718.165 2787.510 1720.130 2787.810 ;
        RECT 1718.165 2787.495 1718.495 2787.510 ;
        RECT 1719.750 2787.500 1720.130 2787.510 ;
        RECT 1725.065 2787.810 1725.395 2787.825 ;
        RECT 1730.790 2787.810 1731.170 2787.820 ;
        RECT 1725.065 2787.510 1731.170 2787.810 ;
        RECT 1725.065 2787.495 1725.395 2787.510 ;
        RECT 1730.790 2787.500 1731.170 2787.510 ;
        RECT 1731.965 2787.810 1732.295 2787.825 ;
        RECT 1737.230 2787.810 1737.610 2787.820 ;
        RECT 1731.965 2787.510 1737.610 2787.810 ;
        RECT 1731.965 2787.495 1732.295 2787.510 ;
        RECT 1737.230 2787.500 1737.610 2787.510 ;
        RECT 1738.865 2787.810 1739.195 2787.825 ;
        RECT 1743.670 2787.810 1744.050 2787.820 ;
        RECT 1738.865 2787.510 1744.050 2787.810 ;
        RECT 1738.865 2787.495 1739.195 2787.510 ;
        RECT 1743.670 2787.500 1744.050 2787.510 ;
        RECT 1745.765 2787.810 1746.095 2787.825 ;
        RECT 1748.270 2787.810 1748.650 2787.820 ;
        RECT 1745.765 2787.510 1748.650 2787.810 ;
        RECT 1745.765 2787.495 1746.095 2787.510 ;
        RECT 1748.270 2787.500 1748.650 2787.510 ;
        RECT 1752.665 2787.810 1752.995 2787.825 ;
        RECT 1754.710 2787.810 1755.090 2787.820 ;
        RECT 1752.665 2787.510 1755.090 2787.810 ;
        RECT 1752.665 2787.495 1752.995 2787.510 ;
        RECT 1754.710 2787.500 1755.090 2787.510 ;
        RECT 1766.465 2787.810 1766.795 2787.825 ;
        RECT 1772.190 2787.810 1772.570 2787.820 ;
        RECT 1766.465 2787.510 1772.570 2787.810 ;
        RECT 1766.465 2787.495 1766.795 2787.510 ;
        RECT 1772.190 2787.500 1772.570 2787.510 ;
        RECT 1773.365 2787.810 1773.695 2787.825 ;
        RECT 1778.630 2787.810 1779.010 2787.820 ;
        RECT 1773.365 2787.510 1779.010 2787.810 ;
        RECT 1773.365 2787.495 1773.695 2787.510 ;
        RECT 1778.630 2787.500 1779.010 2787.510 ;
        RECT 1780.265 2787.810 1780.595 2787.825 ;
        RECT 1783.230 2787.810 1783.610 2787.820 ;
        RECT 1780.265 2787.510 1783.610 2787.810 ;
        RECT 1780.265 2787.495 1780.595 2787.510 ;
        RECT 1783.230 2787.500 1783.610 2787.510 ;
        RECT 1787.625 2787.810 1787.955 2787.825 ;
        RECT 1789.670 2787.810 1790.050 2787.820 ;
        RECT 1787.625 2787.510 1790.050 2787.810 ;
        RECT 1787.625 2787.495 1787.955 2787.510 ;
        RECT 1789.670 2787.500 1790.050 2787.510 ;
        RECT 2263.265 2787.810 2263.595 2787.825 ;
        RECT 2264.390 2787.810 2264.770 2787.820 ;
        RECT 2263.265 2787.510 2264.770 2787.810 ;
        RECT 2263.265 2787.495 2263.595 2787.510 ;
        RECT 2264.390 2787.500 2264.770 2787.510 ;
        RECT 2266.945 2787.810 2267.275 2787.825 ;
        RECT 2276.350 2787.810 2276.730 2787.820 ;
        RECT 2266.945 2787.510 2276.730 2787.810 ;
        RECT 2266.945 2787.495 2267.275 2787.510 ;
        RECT 2276.350 2787.500 2276.730 2787.510 ;
        RECT 2277.065 2787.810 2277.395 2787.825 ;
        RECT 2282.790 2787.810 2283.170 2787.820 ;
        RECT 2277.065 2787.510 2283.170 2787.810 ;
        RECT 2277.065 2787.495 2277.395 2787.510 ;
        RECT 2282.790 2787.500 2283.170 2787.510 ;
        RECT 2283.965 2787.810 2284.295 2787.825 ;
        RECT 2287.390 2787.810 2287.770 2787.820 ;
        RECT 2283.965 2787.510 2287.770 2787.810 ;
        RECT 2283.965 2787.495 2284.295 2787.510 ;
        RECT 2287.390 2787.500 2287.770 2787.510 ;
        RECT 2290.865 2787.810 2291.195 2787.825 ;
        RECT 2293.830 2787.810 2294.210 2787.820 ;
        RECT 2290.865 2787.510 2294.210 2787.810 ;
        RECT 2290.865 2787.495 2291.195 2787.510 ;
        RECT 2293.830 2787.500 2294.210 2787.510 ;
        RECT 2297.765 2787.810 2298.095 2787.825 ;
        RECT 2304.665 2787.820 2304.995 2787.825 ;
        RECT 2300.270 2787.810 2300.650 2787.820 ;
        RECT 2304.665 2787.810 2305.250 2787.820 ;
        RECT 2297.765 2787.510 2300.650 2787.810 ;
        RECT 2304.440 2787.510 2305.250 2787.810 ;
        RECT 2297.765 2787.495 2298.095 2787.510 ;
        RECT 2300.270 2787.500 2300.650 2787.510 ;
        RECT 2304.665 2787.500 2305.250 2787.510 ;
        RECT 2311.565 2787.810 2311.895 2787.825 ;
        RECT 2317.750 2787.810 2318.130 2787.820 ;
        RECT 2311.565 2787.510 2318.130 2787.810 ;
        RECT 2304.665 2787.495 2304.995 2787.500 ;
        RECT 2311.565 2787.495 2311.895 2787.510 ;
        RECT 2317.750 2787.500 2318.130 2787.510 ;
        RECT 2318.465 2787.810 2318.795 2787.825 ;
        RECT 2322.350 2787.810 2322.730 2787.820 ;
        RECT 2318.465 2787.510 2322.730 2787.810 ;
        RECT 2318.465 2787.495 2318.795 2787.510 ;
        RECT 2322.350 2787.500 2322.730 2787.510 ;
        RECT 2325.365 2787.810 2325.695 2787.825 ;
        RECT 2328.790 2787.810 2329.170 2787.820 ;
        RECT 2325.365 2787.510 2329.170 2787.810 ;
        RECT 2325.365 2787.495 2325.695 2787.510 ;
        RECT 2328.790 2787.500 2329.170 2787.510 ;
        RECT 2373.205 2787.810 2373.535 2787.825 ;
        RECT 2381.945 2787.810 2382.275 2787.825 ;
        RECT 2373.205 2787.510 2382.275 2787.810 ;
        RECT 2373.205 2787.495 2373.535 2787.510 ;
        RECT 2381.945 2787.495 2382.275 2787.510 ;
        RECT 1760.945 2777.620 1761.275 2777.625 ;
        RECT 1760.945 2777.610 1761.530 2777.620 ;
        RECT 1760.720 2777.310 1761.530 2777.610 ;
        RECT 1760.945 2777.300 1761.530 2777.310 ;
        RECT 1794.525 2777.610 1794.855 2777.625 ;
        RECT 1796.110 2777.610 1796.490 2777.620 ;
        RECT 1794.525 2777.310 1796.490 2777.610 ;
        RECT 1760.945 2777.295 1761.275 2777.300 ;
        RECT 1794.525 2777.295 1794.855 2777.310 ;
        RECT 1796.110 2777.300 1796.490 2777.310 ;
        RECT 700.185 2718.450 700.515 2718.465 ;
        RECT 1000.105 2718.450 1000.435 2718.465 ;
        RECT 700.185 2718.150 1000.435 2718.450 ;
        RECT 700.185 2718.135 700.515 2718.150 ;
        RECT 1000.105 2718.135 1000.435 2718.150 ;
        RECT 741.585 2717.770 741.915 2717.785 ;
        RECT 1052.085 2717.770 1052.415 2717.785 ;
        RECT 741.585 2717.470 1052.415 2717.770 ;
        RECT 741.585 2717.455 741.915 2717.470 ;
        RECT 1052.085 2717.455 1052.415 2717.470 ;
        RECT 707.085 2717.090 707.415 2717.105 ;
        RECT 1041.505 2717.090 1041.835 2717.105 ;
        RECT 707.085 2716.790 1041.835 2717.090 ;
        RECT 707.085 2716.775 707.415 2716.790 ;
        RECT 1041.505 2716.775 1041.835 2716.790 ;
        RECT 481.225 2716.410 481.555 2716.425 ;
        RECT 941.685 2716.410 942.015 2716.425 ;
        RECT 481.225 2716.110 942.015 2716.410 ;
        RECT 481.225 2716.095 481.555 2716.110 ;
        RECT 941.685 2716.095 942.015 2716.110 ;
        RECT 517.105 2715.730 517.435 2715.745 ;
        RECT 1010.225 2715.730 1010.555 2715.745 ;
        RECT 517.105 2715.430 1010.555 2715.730 ;
        RECT 517.105 2715.415 517.435 2715.430 ;
        RECT 1010.225 2715.415 1010.555 2715.430 ;
        RECT 387.845 2715.050 388.175 2715.065 ;
        RECT 944.905 2715.050 945.235 2715.065 ;
        RECT 387.845 2714.750 945.235 2715.050 ;
        RECT 387.845 2714.735 388.175 2714.750 ;
        RECT 944.905 2714.735 945.235 2714.750 ;
        RECT 1395.930 2695.330 1399.930 2695.440 ;
        RECT 1408.585 2695.330 1408.915 2695.345 ;
      LAYER met3 ;
        RECT 300.915 2694.440 1395.530 2695.305 ;
      LAYER met3 ;
        RECT 1395.930 2695.030 1408.915 2695.330 ;
        RECT 1395.930 2694.840 1399.930 2695.030 ;
        RECT 1408.585 2695.015 1408.915 2695.030 ;
      LAYER met3 ;
        RECT 300.915 2685.640 1395.930 2694.440 ;
        RECT 300.915 2684.240 1395.530 2685.640 ;
      LAYER met3 ;
        RECT 1395.930 2685.130 1399.930 2685.240 ;
        RECT 1408.585 2685.130 1408.915 2685.145 ;
        RECT 1395.930 2684.830 1408.915 2685.130 ;
        RECT 1395.930 2684.640 1399.930 2684.830 ;
        RECT 1408.585 2684.815 1408.915 2684.830 ;
      LAYER met3 ;
        RECT 300.915 2675.440 1395.930 2684.240 ;
        RECT 300.915 2674.040 1395.530 2675.440 ;
      LAYER met3 ;
        RECT 1395.930 2674.930 1399.930 2675.040 ;
        RECT 1408.585 2674.930 1408.915 2674.945 ;
        RECT 1395.930 2674.630 1408.915 2674.930 ;
        RECT 1395.930 2674.440 1399.930 2674.630 ;
        RECT 1408.585 2674.615 1408.915 2674.630 ;
      LAYER met3 ;
        RECT 300.915 2665.240 1395.930 2674.040 ;
        RECT 300.915 2663.840 1395.530 2665.240 ;
      LAYER met3 ;
        RECT 1395.930 2664.730 1399.930 2664.840 ;
        RECT 1408.585 2664.730 1408.915 2664.745 ;
        RECT 1395.930 2664.430 1408.915 2664.730 ;
        RECT 1395.930 2664.240 1399.930 2664.430 ;
        RECT 1408.585 2664.415 1408.915 2664.430 ;
      LAYER met3 ;
        RECT 300.915 2655.040 1395.930 2663.840 ;
        RECT 300.915 2653.640 1395.530 2655.040 ;
      LAYER met3 ;
        RECT 1395.930 2654.530 1399.930 2654.640 ;
        RECT 1408.585 2654.530 1408.915 2654.545 ;
        RECT 1395.930 2654.230 1408.915 2654.530 ;
        RECT 1395.930 2654.040 1399.930 2654.230 ;
        RECT 1408.585 2654.215 1408.915 2654.230 ;
      LAYER met3 ;
        RECT 300.915 2644.840 1395.930 2653.640 ;
        RECT 300.915 2643.440 1395.530 2644.840 ;
      LAYER met3 ;
        RECT 1395.930 2644.330 1399.930 2644.440 ;
        RECT 1408.585 2644.330 1408.915 2644.345 ;
        RECT 1395.930 2644.030 1408.915 2644.330 ;
        RECT 1395.930 2643.840 1399.930 2644.030 ;
        RECT 1408.585 2644.015 1408.915 2644.030 ;
      LAYER met3 ;
        RECT 300.915 2634.640 1395.930 2643.440 ;
        RECT 300.915 2633.240 1395.530 2634.640 ;
      LAYER met3 ;
        RECT 1395.930 2634.130 1399.930 2634.240 ;
        RECT 1408.585 2634.130 1408.915 2634.145 ;
        RECT 1395.930 2633.830 1408.915 2634.130 ;
        RECT 1395.930 2633.640 1399.930 2633.830 ;
        RECT 1408.585 2633.815 1408.915 2633.830 ;
      LAYER met3 ;
        RECT 300.915 2624.440 1395.930 2633.240 ;
        RECT 300.915 2623.040 1395.530 2624.440 ;
      LAYER met3 ;
        RECT 1395.930 2623.930 1399.930 2624.040 ;
        RECT 1408.585 2623.930 1408.915 2623.945 ;
        RECT 1395.930 2623.630 1408.915 2623.930 ;
        RECT 1395.930 2623.440 1399.930 2623.630 ;
        RECT 1408.585 2623.615 1408.915 2623.630 ;
      LAYER met3 ;
        RECT 300.915 2614.240 1395.930 2623.040 ;
        RECT 300.915 2612.840 1395.530 2614.240 ;
      LAYER met3 ;
        RECT 1395.930 2613.730 1399.930 2613.840 ;
        RECT 1408.585 2613.730 1408.915 2613.745 ;
        RECT 1395.930 2613.430 1408.915 2613.730 ;
        RECT 1395.930 2613.240 1399.930 2613.430 ;
        RECT 1408.585 2613.415 1408.915 2613.430 ;
      LAYER met3 ;
        RECT 300.915 2604.040 1395.930 2612.840 ;
        RECT 300.915 2602.640 1395.530 2604.040 ;
      LAYER met3 ;
        RECT 1395.930 2603.530 1399.930 2603.640 ;
        RECT 1408.585 2603.530 1408.915 2603.545 ;
        RECT 1395.930 2603.230 1408.915 2603.530 ;
        RECT 1395.930 2603.040 1399.930 2603.230 ;
        RECT 1408.585 2603.215 1408.915 2603.230 ;
      LAYER met3 ;
        RECT 300.915 2593.840 1395.930 2602.640 ;
        RECT 300.915 2592.440 1395.530 2593.840 ;
      LAYER met3 ;
        RECT 1395.930 2593.330 1399.930 2593.440 ;
        RECT 1408.585 2593.330 1408.915 2593.345 ;
        RECT 1395.930 2593.030 1408.915 2593.330 ;
        RECT 1395.930 2592.840 1399.930 2593.030 ;
        RECT 1408.585 2593.015 1408.915 2593.030 ;
      LAYER met3 ;
        RECT 300.915 2583.640 1395.930 2592.440 ;
        RECT 300.915 2582.240 1395.530 2583.640 ;
      LAYER met3 ;
        RECT 1395.930 2583.130 1399.930 2583.240 ;
        RECT 1408.585 2583.130 1408.915 2583.145 ;
        RECT 1395.930 2582.830 1408.915 2583.130 ;
        RECT 1395.930 2582.640 1399.930 2582.830 ;
        RECT 1408.585 2582.815 1408.915 2582.830 ;
      LAYER met3 ;
        RECT 300.915 2573.440 1395.930 2582.240 ;
        RECT 300.915 2572.040 1395.530 2573.440 ;
      LAYER met3 ;
        RECT 1395.930 2572.930 1399.930 2573.040 ;
        RECT 1408.585 2572.930 1408.915 2572.945 ;
        RECT 1395.930 2572.630 1408.915 2572.930 ;
        RECT 1395.930 2572.440 1399.930 2572.630 ;
        RECT 1408.585 2572.615 1408.915 2572.630 ;
      LAYER met3 ;
        RECT 300.915 2563.240 1395.930 2572.040 ;
        RECT 300.915 2561.840 1395.530 2563.240 ;
      LAYER met3 ;
        RECT 1395.930 2562.730 1399.930 2562.840 ;
        RECT 1408.585 2562.730 1408.915 2562.745 ;
        RECT 1395.930 2562.430 1408.915 2562.730 ;
        RECT 1395.930 2562.240 1399.930 2562.430 ;
        RECT 1408.585 2562.415 1408.915 2562.430 ;
      LAYER met3 ;
        RECT 300.915 2553.040 1395.930 2561.840 ;
        RECT 300.915 2551.640 1395.530 2553.040 ;
      LAYER met3 ;
        RECT 1395.930 2552.530 1399.930 2552.640 ;
        RECT 1408.585 2552.530 1408.915 2552.545 ;
        RECT 1395.930 2552.230 1408.915 2552.530 ;
        RECT 1395.930 2552.040 1399.930 2552.230 ;
        RECT 1408.585 2552.215 1408.915 2552.230 ;
      LAYER met3 ;
        RECT 300.915 2542.840 1395.930 2551.640 ;
        RECT 300.915 2541.440 1395.530 2542.840 ;
      LAYER met3 ;
        RECT 1395.930 2542.330 1399.930 2542.440 ;
        RECT 1408.585 2542.330 1408.915 2542.345 ;
        RECT 1395.930 2542.030 1408.915 2542.330 ;
        RECT 1395.930 2541.840 1399.930 2542.030 ;
        RECT 1408.585 2542.015 1408.915 2542.030 ;
      LAYER met3 ;
        RECT 300.915 2532.640 1395.930 2541.440 ;
        RECT 300.915 2531.240 1395.530 2532.640 ;
      LAYER met3 ;
        RECT 1395.930 2532.130 1399.930 2532.240 ;
        RECT 1408.585 2532.130 1408.915 2532.145 ;
        RECT 1395.930 2531.830 1408.915 2532.130 ;
        RECT 1395.930 2531.640 1399.930 2531.830 ;
        RECT 1408.585 2531.815 1408.915 2531.830 ;
      LAYER met3 ;
        RECT 300.915 2522.440 1395.930 2531.240 ;
        RECT 300.915 2521.040 1395.530 2522.440 ;
      LAYER met3 ;
        RECT 1395.930 2521.930 1399.930 2522.040 ;
        RECT 1408.585 2521.930 1408.915 2521.945 ;
        RECT 1395.930 2521.630 1408.915 2521.930 ;
        RECT 1395.930 2521.440 1399.930 2521.630 ;
        RECT 1408.585 2521.615 1408.915 2521.630 ;
      LAYER met3 ;
        RECT 300.915 2512.240 1395.930 2521.040 ;
        RECT 300.915 2510.840 1395.530 2512.240 ;
      LAYER met3 ;
        RECT 1395.930 2511.730 1399.930 2511.840 ;
        RECT 1408.585 2511.730 1408.915 2511.745 ;
        RECT 1395.930 2511.430 1408.915 2511.730 ;
        RECT 1395.930 2511.240 1399.930 2511.430 ;
        RECT 1408.585 2511.415 1408.915 2511.430 ;
      LAYER met3 ;
        RECT 300.915 2502.040 1395.930 2510.840 ;
        RECT 300.915 2500.640 1395.530 2502.040 ;
      LAYER met3 ;
        RECT 1395.930 2501.530 1399.930 2501.640 ;
        RECT 1408.585 2501.530 1408.915 2501.545 ;
        RECT 1395.930 2501.230 1408.915 2501.530 ;
        RECT 1395.930 2501.040 1399.930 2501.230 ;
        RECT 1408.585 2501.215 1408.915 2501.230 ;
      LAYER met3 ;
        RECT 300.915 2491.840 1395.930 2500.640 ;
        RECT 300.915 2490.440 1395.530 2491.840 ;
      LAYER met3 ;
        RECT 1395.930 2491.330 1399.930 2491.440 ;
        RECT 1408.585 2491.330 1408.915 2491.345 ;
        RECT 1395.930 2491.030 1408.915 2491.330 ;
        RECT 1395.930 2490.840 1399.930 2491.030 ;
        RECT 1408.585 2491.015 1408.915 2491.030 ;
      LAYER met3 ;
        RECT 300.915 2481.640 1395.930 2490.440 ;
        RECT 300.915 2480.240 1395.530 2481.640 ;
      LAYER met3 ;
        RECT 1395.930 2481.130 1399.930 2481.240 ;
        RECT 1408.585 2481.130 1408.915 2481.145 ;
        RECT 1395.930 2480.830 1408.915 2481.130 ;
        RECT 1395.930 2480.640 1399.930 2480.830 ;
        RECT 1408.585 2480.815 1408.915 2480.830 ;
      LAYER met3 ;
        RECT 300.915 2471.440 1395.930 2480.240 ;
        RECT 300.915 2470.040 1395.530 2471.440 ;
      LAYER met3 ;
        RECT 1395.930 2470.930 1399.930 2471.040 ;
        RECT 1408.585 2470.930 1408.915 2470.945 ;
        RECT 1395.930 2470.630 1408.915 2470.930 ;
        RECT 1395.930 2470.440 1399.930 2470.630 ;
        RECT 1408.585 2470.615 1408.915 2470.630 ;
      LAYER met3 ;
        RECT 300.915 2461.240 1395.930 2470.040 ;
        RECT 300.915 2459.840 1395.530 2461.240 ;
      LAYER met3 ;
        RECT 1395.930 2460.730 1399.930 2460.840 ;
        RECT 1408.585 2460.730 1408.915 2460.745 ;
        RECT 1395.930 2460.430 1408.915 2460.730 ;
        RECT 1395.930 2460.240 1399.930 2460.430 ;
        RECT 1408.585 2460.415 1408.915 2460.430 ;
      LAYER met3 ;
        RECT 300.915 2451.040 1395.930 2459.840 ;
        RECT 300.915 2449.640 1395.530 2451.040 ;
      LAYER met3 ;
        RECT 1395.930 2450.530 1399.930 2450.640 ;
        RECT 1408.585 2450.530 1408.915 2450.545 ;
        RECT 1395.930 2450.230 1408.915 2450.530 ;
        RECT 1395.930 2450.040 1399.930 2450.230 ;
        RECT 1408.585 2450.215 1408.915 2450.230 ;
      LAYER met3 ;
        RECT 300.915 2440.840 1395.930 2449.640 ;
        RECT 300.915 2439.440 1395.530 2440.840 ;
      LAYER met3 ;
        RECT 1395.930 2440.330 1399.930 2440.440 ;
        RECT 1408.585 2440.330 1408.915 2440.345 ;
        RECT 1395.930 2440.030 1408.915 2440.330 ;
        RECT 1395.930 2439.840 1399.930 2440.030 ;
        RECT 1408.585 2440.015 1408.915 2440.030 ;
      LAYER met3 ;
        RECT 300.915 2430.640 1395.930 2439.440 ;
        RECT 300.915 2429.240 1395.530 2430.640 ;
      LAYER met3 ;
        RECT 1395.930 2430.130 1399.930 2430.240 ;
        RECT 1408.585 2430.130 1408.915 2430.145 ;
        RECT 1395.930 2429.830 1408.915 2430.130 ;
        RECT 1395.930 2429.640 1399.930 2429.830 ;
        RECT 1408.585 2429.815 1408.915 2429.830 ;
      LAYER met3 ;
        RECT 300.915 2420.440 1395.930 2429.240 ;
        RECT 300.915 2419.040 1395.530 2420.440 ;
      LAYER met3 ;
        RECT 1395.930 2419.930 1399.930 2420.040 ;
        RECT 1408.585 2419.930 1408.915 2419.945 ;
        RECT 1395.930 2419.630 1408.915 2419.930 ;
        RECT 1395.930 2419.440 1399.930 2419.630 ;
        RECT 1408.585 2419.615 1408.915 2419.630 ;
      LAYER met3 ;
        RECT 300.915 2410.240 1395.930 2419.040 ;
        RECT 300.915 2408.840 1395.530 2410.240 ;
      LAYER met3 ;
        RECT 1395.930 2409.730 1399.930 2409.840 ;
        RECT 1408.585 2409.730 1408.915 2409.745 ;
        RECT 1395.930 2409.430 1408.915 2409.730 ;
        RECT 1395.930 2409.240 1399.930 2409.430 ;
        RECT 1408.585 2409.415 1408.915 2409.430 ;
      LAYER met3 ;
        RECT 300.915 2400.040 1395.930 2408.840 ;
        RECT 300.915 2398.640 1395.530 2400.040 ;
      LAYER met3 ;
        RECT 1395.930 2399.530 1399.930 2399.640 ;
        RECT 1408.585 2399.530 1408.915 2399.545 ;
        RECT 1395.930 2399.230 1408.915 2399.530 ;
        RECT 1395.930 2399.040 1399.930 2399.230 ;
        RECT 1408.585 2399.215 1408.915 2399.230 ;
      LAYER met3 ;
        RECT 300.915 2389.840 1395.930 2398.640 ;
        RECT 300.915 2388.440 1395.530 2389.840 ;
      LAYER met3 ;
        RECT 1395.930 2389.330 1399.930 2389.440 ;
        RECT 1408.585 2389.330 1408.915 2389.345 ;
        RECT 1395.930 2389.030 1408.915 2389.330 ;
        RECT 1395.930 2388.840 1399.930 2389.030 ;
        RECT 1408.585 2389.015 1408.915 2389.030 ;
      LAYER met3 ;
        RECT 300.915 2379.640 1395.930 2388.440 ;
        RECT 300.915 2378.240 1395.530 2379.640 ;
      LAYER met3 ;
        RECT 1395.930 2379.130 1399.930 2379.240 ;
        RECT 1408.585 2379.130 1408.915 2379.145 ;
        RECT 1395.930 2378.830 1408.915 2379.130 ;
        RECT 1395.930 2378.640 1399.930 2378.830 ;
        RECT 1408.585 2378.815 1408.915 2378.830 ;
      LAYER met3 ;
        RECT 300.915 2369.440 1395.930 2378.240 ;
        RECT 300.915 2368.040 1395.530 2369.440 ;
      LAYER met3 ;
        RECT 1395.930 2368.930 1399.930 2369.040 ;
        RECT 1408.585 2368.930 1408.915 2368.945 ;
        RECT 1395.930 2368.630 1408.915 2368.930 ;
        RECT 1395.930 2368.440 1399.930 2368.630 ;
        RECT 1408.585 2368.615 1408.915 2368.630 ;
      LAYER met3 ;
        RECT 300.915 2359.240 1395.930 2368.040 ;
        RECT 300.915 2357.840 1395.530 2359.240 ;
      LAYER met3 ;
        RECT 1395.930 2358.730 1399.930 2358.840 ;
        RECT 1408.585 2358.730 1408.915 2358.745 ;
        RECT 1395.930 2358.430 1408.915 2358.730 ;
        RECT 1395.930 2358.240 1399.930 2358.430 ;
        RECT 1408.585 2358.415 1408.915 2358.430 ;
      LAYER met3 ;
        RECT 300.915 2349.040 1395.930 2357.840 ;
        RECT 300.915 2347.640 1395.530 2349.040 ;
      LAYER met3 ;
        RECT 1395.930 2348.530 1399.930 2348.640 ;
        RECT 1408.585 2348.530 1408.915 2348.545 ;
        RECT 1395.930 2348.230 1408.915 2348.530 ;
        RECT 1395.930 2348.040 1399.930 2348.230 ;
        RECT 1408.585 2348.215 1408.915 2348.230 ;
      LAYER met3 ;
        RECT 300.915 2338.840 1395.930 2347.640 ;
        RECT 300.915 2337.440 1395.530 2338.840 ;
      LAYER met3 ;
        RECT 1395.930 2338.330 1399.930 2338.440 ;
        RECT 1408.585 2338.330 1408.915 2338.345 ;
        RECT 1395.930 2338.030 1408.915 2338.330 ;
        RECT 1395.930 2337.840 1399.930 2338.030 ;
        RECT 1408.585 2338.015 1408.915 2338.030 ;
      LAYER met3 ;
        RECT 300.915 2328.640 1395.930 2337.440 ;
        RECT 300.915 2327.240 1395.530 2328.640 ;
      LAYER met3 ;
        RECT 1395.930 2328.130 1399.930 2328.240 ;
        RECT 1408.585 2328.130 1408.915 2328.145 ;
        RECT 1395.930 2327.830 1408.915 2328.130 ;
        RECT 1395.930 2327.640 1399.930 2327.830 ;
        RECT 1408.585 2327.815 1408.915 2327.830 ;
      LAYER met3 ;
        RECT 300.915 2318.440 1395.930 2327.240 ;
        RECT 300.915 2317.040 1395.530 2318.440 ;
      LAYER met3 ;
        RECT 1395.930 2317.930 1399.930 2318.040 ;
        RECT 1408.585 2317.930 1408.915 2317.945 ;
        RECT 1395.930 2317.630 1408.915 2317.930 ;
        RECT 1395.930 2317.440 1399.930 2317.630 ;
        RECT 1408.585 2317.615 1408.915 2317.630 ;
      LAYER met3 ;
        RECT 300.915 2308.240 1395.930 2317.040 ;
        RECT 300.915 2306.840 1395.530 2308.240 ;
      LAYER met3 ;
        RECT 1395.930 2307.730 1399.930 2307.840 ;
        RECT 1408.585 2307.730 1408.915 2307.745 ;
        RECT 1395.930 2307.430 1408.915 2307.730 ;
        RECT 1395.930 2307.240 1399.930 2307.430 ;
        RECT 1408.585 2307.415 1408.915 2307.430 ;
      LAYER met3 ;
        RECT 300.915 2298.040 1395.930 2306.840 ;
        RECT 300.915 2296.640 1395.530 2298.040 ;
      LAYER met3 ;
        RECT 1395.930 2297.530 1399.930 2297.640 ;
        RECT 1408.585 2297.530 1408.915 2297.545 ;
        RECT 1395.930 2297.230 1408.915 2297.530 ;
        RECT 1395.930 2297.040 1399.930 2297.230 ;
        RECT 1408.585 2297.215 1408.915 2297.230 ;
      LAYER met3 ;
        RECT 300.915 2287.840 1395.930 2296.640 ;
        RECT 300.915 2286.440 1395.530 2287.840 ;
      LAYER met3 ;
        RECT 1395.930 2287.330 1399.930 2287.440 ;
        RECT 1408.585 2287.330 1408.915 2287.345 ;
        RECT 1395.930 2287.030 1408.915 2287.330 ;
        RECT 1395.930 2286.840 1399.930 2287.030 ;
        RECT 1408.585 2287.015 1408.915 2287.030 ;
      LAYER met3 ;
        RECT 300.915 2277.640 1395.930 2286.440 ;
        RECT 300.915 2276.240 1395.530 2277.640 ;
      LAYER met3 ;
        RECT 1395.930 2277.130 1399.930 2277.240 ;
        RECT 1408.585 2277.130 1408.915 2277.145 ;
        RECT 1395.930 2276.830 1408.915 2277.130 ;
        RECT 1395.930 2276.640 1399.930 2276.830 ;
        RECT 1408.585 2276.815 1408.915 2276.830 ;
      LAYER met3 ;
        RECT 300.915 2267.440 1395.930 2276.240 ;
        RECT 300.915 2266.040 1395.530 2267.440 ;
      LAYER met3 ;
        RECT 1395.930 2266.930 1399.930 2267.040 ;
        RECT 1408.585 2266.930 1408.915 2266.945 ;
        RECT 1395.930 2266.630 1408.915 2266.930 ;
        RECT 1395.930 2266.440 1399.930 2266.630 ;
        RECT 1408.585 2266.615 1408.915 2266.630 ;
      LAYER met3 ;
        RECT 300.915 2257.240 1395.930 2266.040 ;
        RECT 300.915 2255.840 1395.530 2257.240 ;
      LAYER met3 ;
        RECT 1395.930 2256.730 1399.930 2256.840 ;
        RECT 1408.585 2256.730 1408.915 2256.745 ;
        RECT 1395.930 2256.430 1408.915 2256.730 ;
        RECT 1395.930 2256.240 1399.930 2256.430 ;
        RECT 1408.585 2256.415 1408.915 2256.430 ;
      LAYER met3 ;
        RECT 300.915 2247.040 1395.930 2255.840 ;
        RECT 300.915 2245.640 1395.530 2247.040 ;
      LAYER met3 ;
        RECT 1395.930 2246.530 1399.930 2246.640 ;
        RECT 1408.585 2246.530 1408.915 2246.545 ;
        RECT 1395.930 2246.230 1408.915 2246.530 ;
        RECT 1395.930 2246.040 1399.930 2246.230 ;
        RECT 1408.585 2246.215 1408.915 2246.230 ;
      LAYER met3 ;
        RECT 300.915 2236.840 1395.930 2245.640 ;
        RECT 300.915 2235.440 1395.530 2236.840 ;
      LAYER met3 ;
        RECT 1395.930 2236.330 1399.930 2236.440 ;
        RECT 1408.585 2236.330 1408.915 2236.345 ;
        RECT 1395.930 2236.030 1408.915 2236.330 ;
        RECT 1395.930 2235.840 1399.930 2236.030 ;
        RECT 1408.585 2236.015 1408.915 2236.030 ;
      LAYER met3 ;
        RECT 300.915 2226.640 1395.930 2235.440 ;
        RECT 300.915 2225.240 1395.530 2226.640 ;
      LAYER met3 ;
        RECT 1395.930 2226.130 1399.930 2226.240 ;
        RECT 1408.585 2226.130 1408.915 2226.145 ;
        RECT 1395.930 2225.830 1408.915 2226.130 ;
        RECT 1395.930 2225.640 1399.930 2225.830 ;
        RECT 1408.585 2225.815 1408.915 2225.830 ;
      LAYER met3 ;
        RECT 300.915 2216.440 1395.930 2225.240 ;
        RECT 300.915 2215.040 1395.530 2216.440 ;
      LAYER met3 ;
        RECT 1395.930 2215.930 1399.930 2216.040 ;
        RECT 1408.585 2215.930 1408.915 2215.945 ;
        RECT 1395.930 2215.630 1408.915 2215.930 ;
        RECT 1395.930 2215.440 1399.930 2215.630 ;
        RECT 1408.585 2215.615 1408.915 2215.630 ;
      LAYER met3 ;
        RECT 300.915 2206.240 1395.930 2215.040 ;
        RECT 300.915 2204.840 1395.530 2206.240 ;
      LAYER met3 ;
        RECT 1395.930 2205.730 1399.930 2205.840 ;
        RECT 1408.585 2205.730 1408.915 2205.745 ;
        RECT 1395.930 2205.430 1408.915 2205.730 ;
        RECT 1395.930 2205.240 1399.930 2205.430 ;
        RECT 1408.585 2205.415 1408.915 2205.430 ;
      LAYER met3 ;
        RECT 300.915 2196.040 1395.930 2204.840 ;
        RECT 300.915 2194.640 1395.530 2196.040 ;
      LAYER met3 ;
        RECT 1395.930 2195.530 1399.930 2195.640 ;
        RECT 1408.585 2195.530 1408.915 2195.545 ;
        RECT 1395.930 2195.230 1408.915 2195.530 ;
        RECT 1395.930 2195.040 1399.930 2195.230 ;
        RECT 1408.585 2195.215 1408.915 2195.230 ;
      LAYER met3 ;
        RECT 300.915 2185.840 1395.930 2194.640 ;
        RECT 300.915 2184.440 1395.530 2185.840 ;
      LAYER met3 ;
        RECT 1395.930 2185.330 1399.930 2185.440 ;
        RECT 1408.585 2185.330 1408.915 2185.345 ;
        RECT 1395.930 2185.030 1408.915 2185.330 ;
        RECT 1395.930 2184.840 1399.930 2185.030 ;
        RECT 1408.585 2185.015 1408.915 2185.030 ;
      LAYER met3 ;
        RECT 300.915 2175.640 1395.930 2184.440 ;
        RECT 300.915 2174.240 1395.530 2175.640 ;
      LAYER met3 ;
        RECT 1395.930 2175.130 1399.930 2175.240 ;
        RECT 1408.585 2175.130 1408.915 2175.145 ;
        RECT 1395.930 2174.830 1408.915 2175.130 ;
        RECT 1395.930 2174.640 1399.930 2174.830 ;
        RECT 1408.585 2174.815 1408.915 2174.830 ;
      LAYER met3 ;
        RECT 300.915 2165.440 1395.930 2174.240 ;
        RECT 300.915 2164.040 1395.530 2165.440 ;
      LAYER met3 ;
        RECT 1395.930 2164.930 1399.930 2165.040 ;
        RECT 1408.585 2164.930 1408.915 2164.945 ;
        RECT 1395.930 2164.630 1408.915 2164.930 ;
        RECT 1395.930 2164.440 1399.930 2164.630 ;
        RECT 1408.585 2164.615 1408.915 2164.630 ;
      LAYER met3 ;
        RECT 300.915 2155.920 1395.930 2164.040 ;
        RECT 300.915 2154.520 1395.530 2155.920 ;
      LAYER met3 ;
        RECT 1395.930 2155.410 1399.930 2155.520 ;
        RECT 1408.585 2155.410 1408.915 2155.425 ;
        RECT 1395.930 2155.110 1408.915 2155.410 ;
        RECT 1395.930 2154.920 1399.930 2155.110 ;
        RECT 1408.585 2155.095 1408.915 2155.110 ;
      LAYER met3 ;
        RECT 300.915 2145.720 1395.930 2154.520 ;
        RECT 300.915 2144.320 1395.530 2145.720 ;
      LAYER met3 ;
        RECT 1395.930 2145.210 1399.930 2145.320 ;
        RECT 1408.585 2145.210 1408.915 2145.225 ;
        RECT 1395.930 2144.910 1408.915 2145.210 ;
        RECT 1395.930 2144.720 1399.930 2144.910 ;
        RECT 1408.585 2144.895 1408.915 2144.910 ;
      LAYER met3 ;
        RECT 300.915 2135.520 1395.930 2144.320 ;
        RECT 300.915 2134.120 1395.530 2135.520 ;
      LAYER met3 ;
        RECT 1395.930 2135.010 1399.930 2135.120 ;
        RECT 1408.585 2135.010 1408.915 2135.025 ;
        RECT 1395.930 2134.710 1408.915 2135.010 ;
        RECT 1395.930 2134.520 1399.930 2134.710 ;
        RECT 1408.585 2134.695 1408.915 2134.710 ;
      LAYER met3 ;
        RECT 300.915 2125.320 1395.930 2134.120 ;
        RECT 300.915 2123.920 1395.530 2125.320 ;
      LAYER met3 ;
        RECT 1395.930 2124.810 1399.930 2124.920 ;
        RECT 1408.585 2124.810 1408.915 2124.825 ;
        RECT 1395.930 2124.510 1408.915 2124.810 ;
        RECT 1395.930 2124.320 1399.930 2124.510 ;
        RECT 1408.585 2124.495 1408.915 2124.510 ;
      LAYER met3 ;
        RECT 300.915 2115.120 1395.930 2123.920 ;
        RECT 300.915 2113.720 1395.530 2115.120 ;
      LAYER met3 ;
        RECT 1395.930 2114.610 1399.930 2114.720 ;
        RECT 1408.585 2114.610 1408.915 2114.625 ;
        RECT 1395.930 2114.310 1408.915 2114.610 ;
        RECT 1395.930 2114.120 1399.930 2114.310 ;
        RECT 1408.585 2114.295 1408.915 2114.310 ;
      LAYER met3 ;
        RECT 300.915 2104.920 1395.930 2113.720 ;
        RECT 300.915 2103.520 1395.530 2104.920 ;
      LAYER met3 ;
        RECT 1395.930 2104.410 1399.930 2104.520 ;
        RECT 1408.585 2104.410 1408.915 2104.425 ;
        RECT 1395.930 2104.110 1408.915 2104.410 ;
        RECT 1395.930 2103.920 1399.930 2104.110 ;
        RECT 1408.585 2104.095 1408.915 2104.110 ;
      LAYER met3 ;
        RECT 300.915 2094.720 1395.930 2103.520 ;
        RECT 300.915 2093.320 1395.530 2094.720 ;
      LAYER met3 ;
        RECT 1395.930 2094.210 1399.930 2094.320 ;
        RECT 1408.585 2094.210 1408.915 2094.225 ;
        RECT 1395.930 2093.910 1408.915 2094.210 ;
        RECT 1395.930 2093.720 1399.930 2093.910 ;
        RECT 1408.585 2093.895 1408.915 2093.910 ;
      LAYER met3 ;
        RECT 300.915 2084.520 1395.930 2093.320 ;
        RECT 300.915 2083.120 1395.530 2084.520 ;
      LAYER met3 ;
        RECT 1395.930 2084.010 1399.930 2084.120 ;
        RECT 1408.585 2084.010 1408.915 2084.025 ;
        RECT 1395.930 2083.710 1408.915 2084.010 ;
        RECT 1395.930 2083.520 1399.930 2083.710 ;
        RECT 1408.585 2083.695 1408.915 2083.710 ;
      LAYER met3 ;
        RECT 300.915 2074.320 1395.930 2083.120 ;
        RECT 300.915 2072.920 1395.530 2074.320 ;
      LAYER met3 ;
        RECT 1395.930 2073.810 1399.930 2073.920 ;
        RECT 1408.585 2073.810 1408.915 2073.825 ;
        RECT 1395.930 2073.510 1408.915 2073.810 ;
        RECT 1395.930 2073.320 1399.930 2073.510 ;
        RECT 1408.585 2073.495 1408.915 2073.510 ;
      LAYER met3 ;
        RECT 300.915 2064.120 1395.930 2072.920 ;
        RECT 300.915 2062.720 1395.530 2064.120 ;
      LAYER met3 ;
        RECT 1395.930 2063.610 1399.930 2063.720 ;
        RECT 1408.585 2063.610 1408.915 2063.625 ;
        RECT 1395.930 2063.310 1408.915 2063.610 ;
        RECT 1395.930 2063.120 1399.930 2063.310 ;
        RECT 1408.585 2063.295 1408.915 2063.310 ;
      LAYER met3 ;
        RECT 300.915 2053.920 1395.930 2062.720 ;
        RECT 300.915 2052.520 1395.530 2053.920 ;
      LAYER met3 ;
        RECT 1395.930 2053.410 1399.930 2053.520 ;
        RECT 1409.965 2053.410 1410.295 2053.425 ;
        RECT 1395.930 2053.110 1410.295 2053.410 ;
        RECT 1395.930 2052.920 1399.930 2053.110 ;
        RECT 1409.965 2053.095 1410.295 2053.110 ;
      LAYER met3 ;
        RECT 300.915 2043.720 1395.930 2052.520 ;
      LAYER met3 ;
        RECT 2559.280 2051.235 2561.020 2052.140 ;
      LAYER met3 ;
        RECT 300.915 2042.320 1395.530 2043.720 ;
      LAYER met3 ;
        RECT 1395.930 2043.210 1399.930 2043.320 ;
        RECT 1409.045 2043.210 1409.375 2043.225 ;
        RECT 1395.930 2042.910 1409.375 2043.210 ;
        RECT 1395.930 2042.720 1399.930 2042.910 ;
        RECT 1409.045 2042.895 1409.375 2042.910 ;
      LAYER met3 ;
        RECT 300.915 2033.520 1395.930 2042.320 ;
        RECT 300.915 2032.120 1395.530 2033.520 ;
      LAYER met3 ;
        RECT 1395.930 2033.010 1399.930 2033.120 ;
        RECT 1409.505 2033.010 1409.835 2033.025 ;
        RECT 1395.930 2032.710 1409.835 2033.010 ;
        RECT 1395.930 2032.520 1399.930 2032.710 ;
        RECT 1409.505 2032.695 1409.835 2032.710 ;
      LAYER met3 ;
        RECT 300.915 2023.320 1395.930 2032.120 ;
        RECT 300.915 2021.920 1395.530 2023.320 ;
      LAYER met3 ;
        RECT 1395.930 2022.810 1399.930 2022.920 ;
        RECT 1408.585 2022.810 1408.915 2022.825 ;
        RECT 1395.930 2022.510 1408.915 2022.810 ;
        RECT 1395.930 2022.320 1399.930 2022.510 ;
        RECT 1408.585 2022.495 1408.915 2022.510 ;
      LAYER met3 ;
        RECT 300.915 2013.120 1395.930 2021.920 ;
        RECT 300.915 2011.720 1395.530 2013.120 ;
      LAYER met3 ;
        RECT 1395.930 2012.610 1399.930 2012.720 ;
        RECT 1407.665 2012.610 1407.995 2012.625 ;
        RECT 1395.930 2012.310 1407.995 2012.610 ;
        RECT 1395.930 2012.120 1399.930 2012.310 ;
        RECT 1407.665 2012.295 1407.995 2012.310 ;
      LAYER met3 ;
        RECT 300.915 2002.920 1395.930 2011.720 ;
        RECT 300.915 2001.520 1395.530 2002.920 ;
      LAYER met3 ;
        RECT 1395.930 2002.410 1399.930 2002.520 ;
        RECT 1408.125 2002.410 1408.455 2002.425 ;
        RECT 1395.930 2002.110 1408.455 2002.410 ;
        RECT 1395.930 2001.920 1399.930 2002.110 ;
        RECT 1408.125 2002.095 1408.455 2002.110 ;
      LAYER met3 ;
        RECT 300.915 1992.720 1395.930 2001.520 ;
        RECT 300.915 1991.320 1395.530 1992.720 ;
      LAYER met3 ;
        RECT 1395.930 1992.210 1399.930 1992.320 ;
        RECT 1408.585 1992.210 1408.915 1992.225 ;
        RECT 1395.930 1991.910 1408.915 1992.210 ;
        RECT 1395.930 1991.720 1399.930 1991.910 ;
        RECT 1408.585 1991.895 1408.915 1991.910 ;
      LAYER met3 ;
        RECT 300.915 1982.520 1395.930 1991.320 ;
        RECT 300.915 1981.120 1395.530 1982.520 ;
      LAYER met3 ;
        RECT 1395.930 1982.010 1399.930 1982.120 ;
        RECT 1407.665 1982.010 1407.995 1982.025 ;
        RECT 1395.930 1981.710 1407.995 1982.010 ;
        RECT 1395.930 1981.520 1399.930 1981.710 ;
        RECT 1407.665 1981.695 1407.995 1981.710 ;
      LAYER met3 ;
        RECT 300.915 1972.320 1395.930 1981.120 ;
        RECT 300.915 1970.920 1395.530 1972.320 ;
      LAYER met3 ;
        RECT 1395.930 1971.810 1399.930 1971.920 ;
        RECT 1410.425 1971.810 1410.755 1971.825 ;
        RECT 1395.930 1971.510 1410.755 1971.810 ;
        RECT 1395.930 1971.320 1399.930 1971.510 ;
        RECT 1410.425 1971.495 1410.755 1971.510 ;
      LAYER met3 ;
        RECT 300.915 1962.120 1395.930 1970.920 ;
        RECT 300.915 1960.720 1395.530 1962.120 ;
      LAYER met3 ;
        RECT 1395.930 1961.610 1399.930 1961.720 ;
        RECT 1414.105 1961.610 1414.435 1961.625 ;
        RECT 1395.930 1961.310 1414.435 1961.610 ;
        RECT 1395.930 1961.120 1399.930 1961.310 ;
        RECT 1414.105 1961.295 1414.435 1961.310 ;
      LAYER met3 ;
        RECT 300.915 1951.920 1395.930 1960.720 ;
        RECT 300.915 1950.520 1395.530 1951.920 ;
      LAYER met3 ;
        RECT 1395.930 1951.410 1399.930 1951.520 ;
        RECT 1550.000 1951.445 1554.600 1951.745 ;
        RECT 1413.645 1951.410 1413.975 1951.425 ;
        RECT 1395.930 1951.110 1413.975 1951.410 ;
        RECT 1395.930 1950.920 1399.930 1951.110 ;
        RECT 1413.645 1951.095 1413.975 1951.110 ;
      LAYER met3 ;
        RECT 300.915 1941.720 1395.930 1950.520 ;
      LAYER met3 ;
        RECT 1550.000 1945.805 1554.600 1946.105 ;
      LAYER met3 ;
        RECT 300.915 1940.320 1395.530 1941.720 ;
      LAYER met3 ;
        RECT 1395.930 1941.210 1399.930 1941.320 ;
        RECT 1413.185 1941.210 1413.515 1941.225 ;
        RECT 1395.930 1940.910 1413.515 1941.210 ;
        RECT 1395.930 1940.720 1399.930 1940.910 ;
        RECT 1413.185 1940.895 1413.515 1940.910 ;
      LAYER met3 ;
        RECT 300.915 1931.520 1395.930 1940.320 ;
      LAYER met3 ;
        RECT 1550.000 1937.305 1554.600 1937.605 ;
        RECT 1550.000 1931.665 1554.600 1931.965 ;
      LAYER met3 ;
        RECT 300.915 1930.120 1395.530 1931.520 ;
      LAYER met3 ;
        RECT 1395.930 1931.010 1399.930 1931.120 ;
        RECT 1412.725 1931.010 1413.055 1931.025 ;
        RECT 1395.930 1930.710 1413.055 1931.010 ;
        RECT 1395.930 1930.520 1399.930 1930.710 ;
        RECT 1412.725 1930.695 1413.055 1930.710 ;
      LAYER met3 ;
        RECT 300.915 1921.320 1395.930 1930.120 ;
      LAYER met3 ;
        RECT 1550.000 1923.165 1554.600 1923.465 ;
      LAYER met3 ;
        RECT 300.915 1919.920 1395.530 1921.320 ;
      LAYER met3 ;
        RECT 1395.930 1920.810 1399.930 1920.920 ;
        RECT 1412.265 1920.810 1412.595 1920.825 ;
        RECT 1395.930 1920.510 1412.595 1920.810 ;
        RECT 1395.930 1920.320 1399.930 1920.510 ;
        RECT 1412.265 1920.495 1412.595 1920.510 ;
      LAYER met3 ;
        RECT 300.915 1911.120 1395.930 1919.920 ;
      LAYER met3 ;
        RECT 1550.000 1917.525 1554.600 1917.825 ;
      LAYER met3 ;
        RECT 300.915 1909.720 1395.530 1911.120 ;
      LAYER met3 ;
        RECT 1395.930 1910.610 1399.930 1910.720 ;
        RECT 1411.805 1910.610 1412.135 1910.625 ;
        RECT 1395.930 1910.310 1412.135 1910.610 ;
        RECT 1395.930 1910.120 1399.930 1910.310 ;
        RECT 1411.805 1910.295 1412.135 1910.310 ;
      LAYER met3 ;
        RECT 300.915 1900.920 1395.930 1909.720 ;
      LAYER met3 ;
        RECT 1550.000 1909.025 1554.600 1909.325 ;
      LAYER met3 ;
        RECT 300.915 1899.520 1395.530 1900.920 ;
      LAYER met3 ;
        RECT 1395.930 1900.410 1399.930 1900.520 ;
        RECT 1411.345 1900.410 1411.675 1900.425 ;
        RECT 1395.930 1900.110 1411.675 1900.410 ;
        RECT 1395.930 1899.920 1399.930 1900.110 ;
        RECT 1411.345 1900.095 1411.675 1900.110 ;
      LAYER met3 ;
        RECT 300.915 1890.720 1395.930 1899.520 ;
        RECT 300.915 1889.320 1395.530 1890.720 ;
      LAYER met3 ;
        RECT 1395.930 1890.210 1399.930 1890.320 ;
        RECT 1409.505 1890.210 1409.835 1890.225 ;
        RECT 1395.930 1889.910 1409.835 1890.210 ;
        RECT 1395.930 1889.720 1399.930 1889.910 ;
        RECT 1409.505 1889.895 1409.835 1889.910 ;
      LAYER met3 ;
        RECT 300.915 1880.520 1395.930 1889.320 ;
        RECT 300.915 1879.120 1395.530 1880.520 ;
      LAYER met3 ;
        RECT 1395.930 1880.010 1399.930 1880.120 ;
        RECT 1414.105 1880.010 1414.435 1880.025 ;
        RECT 1395.930 1879.710 1414.435 1880.010 ;
        RECT 1395.930 1879.520 1399.930 1879.710 ;
        RECT 1414.105 1879.695 1414.435 1879.710 ;
      LAYER met3 ;
        RECT 300.915 1870.320 1395.930 1879.120 ;
        RECT 300.915 1868.920 1395.530 1870.320 ;
      LAYER met3 ;
        RECT 1395.930 1869.810 1399.930 1869.920 ;
        RECT 1414.105 1869.810 1414.435 1869.825 ;
        RECT 1395.930 1869.510 1414.435 1869.810 ;
        RECT 1395.930 1869.320 1399.930 1869.510 ;
        RECT 1414.105 1869.495 1414.435 1869.510 ;
      LAYER met3 ;
        RECT 300.915 1860.120 1395.930 1868.920 ;
        RECT 300.915 1858.720 1395.530 1860.120 ;
      LAYER met3 ;
        RECT 1395.930 1859.610 1399.930 1859.720 ;
        RECT 1414.105 1859.610 1414.435 1859.625 ;
        RECT 1395.930 1859.310 1414.435 1859.610 ;
        RECT 1395.930 1859.120 1399.930 1859.310 ;
        RECT 1414.105 1859.295 1414.435 1859.310 ;
      LAYER met3 ;
        RECT 300.915 1849.920 1395.930 1858.720 ;
        RECT 300.915 1848.520 1395.530 1849.920 ;
      LAYER met3 ;
        RECT 1395.930 1849.410 1399.930 1849.520 ;
        RECT 1411.805 1849.410 1412.135 1849.425 ;
        RECT 1395.930 1849.110 1412.135 1849.410 ;
        RECT 1395.930 1848.920 1399.930 1849.110 ;
        RECT 1411.805 1849.095 1412.135 1849.110 ;
      LAYER met3 ;
        RECT 300.915 1839.720 1395.930 1848.520 ;
        RECT 300.915 1838.320 1395.530 1839.720 ;
      LAYER met3 ;
        RECT 1395.930 1839.210 1399.930 1839.320 ;
        RECT 1411.345 1839.210 1411.675 1839.225 ;
        RECT 1395.930 1838.910 1411.675 1839.210 ;
        RECT 1395.930 1838.720 1399.930 1838.910 ;
        RECT 1411.345 1838.895 1411.675 1838.910 ;
      LAYER met3 ;
        RECT 300.915 1829.520 1395.930 1838.320 ;
        RECT 300.915 1828.120 1395.530 1829.520 ;
      LAYER met3 ;
        RECT 1395.930 1829.010 1399.930 1829.120 ;
        RECT 1408.585 1829.010 1408.915 1829.025 ;
        RECT 1395.930 1828.710 1408.915 1829.010 ;
        RECT 1395.930 1828.520 1399.930 1828.710 ;
        RECT 1408.585 1828.695 1408.915 1828.710 ;
      LAYER met3 ;
        RECT 300.915 1819.320 1395.930 1828.120 ;
        RECT 300.915 1817.920 1395.530 1819.320 ;
      LAYER met3 ;
        RECT 1395.930 1818.810 1399.930 1818.920 ;
        RECT 1414.105 1818.810 1414.435 1818.825 ;
        RECT 1395.930 1818.510 1414.435 1818.810 ;
        RECT 1395.930 1818.320 1399.930 1818.510 ;
        RECT 1414.105 1818.495 1414.435 1818.510 ;
      LAYER met3 ;
        RECT 300.915 1809.120 1395.930 1817.920 ;
        RECT 300.915 1807.720 1395.530 1809.120 ;
      LAYER met3 ;
        RECT 1395.930 1808.610 1399.930 1808.720 ;
        RECT 1409.505 1808.610 1409.835 1808.625 ;
        RECT 1395.930 1808.310 1409.835 1808.610 ;
        RECT 1395.930 1808.120 1399.930 1808.310 ;
        RECT 1409.505 1808.295 1409.835 1808.310 ;
      LAYER met3 ;
        RECT 300.915 1798.920 1395.930 1807.720 ;
        RECT 300.915 1797.520 1395.530 1798.920 ;
      LAYER met3 ;
        RECT 1395.930 1798.410 1399.930 1798.520 ;
        RECT 1409.505 1798.410 1409.835 1798.425 ;
        RECT 1395.930 1798.110 1409.835 1798.410 ;
        RECT 1395.930 1797.920 1399.930 1798.110 ;
        RECT 1409.505 1798.095 1409.835 1798.110 ;
      LAYER met3 ;
        RECT 300.915 1788.720 1395.930 1797.520 ;
        RECT 300.915 1787.320 1395.530 1788.720 ;
      LAYER met3 ;
        RECT 1395.930 1788.210 1399.930 1788.320 ;
        RECT 1408.585 1788.210 1408.915 1788.225 ;
        RECT 1395.930 1787.910 1408.915 1788.210 ;
        RECT 1395.930 1787.720 1399.930 1787.910 ;
        RECT 1408.585 1787.895 1408.915 1787.910 ;
      LAYER met3 ;
        RECT 300.915 1778.520 1395.930 1787.320 ;
        RECT 300.915 1777.120 1395.530 1778.520 ;
      LAYER met3 ;
        RECT 1395.930 1778.010 1399.930 1778.120 ;
        RECT 1410.425 1778.010 1410.755 1778.025 ;
        RECT 1395.930 1777.710 1410.755 1778.010 ;
        RECT 1395.930 1777.520 1399.930 1777.710 ;
        RECT 1410.425 1777.695 1410.755 1777.710 ;
      LAYER met3 ;
        RECT 300.915 1768.320 1395.930 1777.120 ;
        RECT 300.915 1766.920 1395.530 1768.320 ;
      LAYER met3 ;
        RECT 1395.930 1767.810 1399.930 1767.920 ;
        RECT 1414.105 1767.810 1414.435 1767.825 ;
        RECT 1395.930 1767.510 1414.435 1767.810 ;
        RECT 1395.930 1767.320 1399.930 1767.510 ;
        RECT 1414.105 1767.495 1414.435 1767.510 ;
      LAYER met3 ;
        RECT 300.915 1758.120 1395.930 1766.920 ;
        RECT 300.915 1756.720 1395.530 1758.120 ;
      LAYER met3 ;
        RECT 1395.930 1757.610 1399.930 1757.720 ;
        RECT 1414.105 1757.610 1414.435 1757.625 ;
        RECT 1395.930 1757.310 1414.435 1757.610 ;
        RECT 1395.930 1757.120 1399.930 1757.310 ;
        RECT 1414.105 1757.295 1414.435 1757.310 ;
      LAYER met3 ;
        RECT 300.915 1747.920 1395.930 1756.720 ;
        RECT 300.915 1746.520 1395.530 1747.920 ;
      LAYER met3 ;
        RECT 1395.930 1747.410 1399.930 1747.520 ;
        RECT 1414.105 1747.410 1414.435 1747.425 ;
        RECT 1395.930 1747.110 1414.435 1747.410 ;
        RECT 1395.930 1746.920 1399.930 1747.110 ;
        RECT 1414.105 1747.095 1414.435 1747.110 ;
      LAYER met3 ;
        RECT 300.915 1737.720 1395.930 1746.520 ;
      LAYER met3 ;
        RECT 1414.105 1738.570 1414.435 1738.585 ;
        RECT 1399.630 1738.270 1414.435 1738.570 ;
      LAYER met3 ;
        RECT 300.915 1736.320 1395.530 1737.720 ;
      LAYER met3 ;
        RECT 1399.630 1737.320 1399.930 1738.270 ;
        RECT 1414.105 1738.255 1414.435 1738.270 ;
        RECT 1395.930 1736.720 1399.930 1737.320 ;
      LAYER met3 ;
        RECT 300.915 1727.520 1395.930 1736.320 ;
        RECT 300.915 1726.120 1395.530 1727.520 ;
      LAYER met3 ;
        RECT 1395.930 1727.010 1399.930 1727.120 ;
        RECT 1407.665 1727.010 1407.995 1727.025 ;
        RECT 1395.930 1726.710 1407.995 1727.010 ;
        RECT 1395.930 1726.520 1399.930 1726.710 ;
        RECT 1407.665 1726.695 1407.995 1726.710 ;
      LAYER met3 ;
        RECT 300.915 1717.320 1395.930 1726.120 ;
        RECT 300.915 1715.920 1395.530 1717.320 ;
      LAYER met3 ;
        RECT 1395.930 1716.810 1399.930 1716.920 ;
        RECT 1414.105 1716.810 1414.435 1716.825 ;
        RECT 1395.930 1716.510 1414.435 1716.810 ;
        RECT 1395.930 1716.320 1399.930 1716.510 ;
        RECT 1414.105 1716.495 1414.435 1716.510 ;
      LAYER met3 ;
        RECT 300.915 1707.120 1395.930 1715.920 ;
        RECT 300.915 1705.720 1395.530 1707.120 ;
      LAYER met3 ;
        RECT 1395.930 1706.610 1399.930 1706.720 ;
        RECT 1407.665 1706.610 1407.995 1706.625 ;
        RECT 1395.930 1706.310 1407.995 1706.610 ;
        RECT 1395.930 1706.120 1399.930 1706.310 ;
        RECT 1407.665 1706.295 1407.995 1706.310 ;
      LAYER met3 ;
        RECT 300.915 1696.920 1395.930 1705.720 ;
        RECT 300.915 1695.520 1395.530 1696.920 ;
      LAYER met3 ;
        RECT 1395.930 1696.410 1399.930 1696.520 ;
        RECT 1408.585 1696.410 1408.915 1696.425 ;
        RECT 1395.930 1696.110 1408.915 1696.410 ;
        RECT 1395.930 1695.920 1399.930 1696.110 ;
        RECT 1408.585 1696.095 1408.915 1696.110 ;
      LAYER met3 ;
        RECT 300.915 1686.720 1395.930 1695.520 ;
        RECT 300.915 1685.320 1395.530 1686.720 ;
      LAYER met3 ;
        RECT 1395.930 1686.210 1399.930 1686.320 ;
        RECT 1407.665 1686.210 1407.995 1686.225 ;
        RECT 1395.930 1685.910 1407.995 1686.210 ;
        RECT 1395.930 1685.720 1399.930 1685.910 ;
        RECT 1407.665 1685.895 1407.995 1685.910 ;
      LAYER met3 ;
        RECT 300.915 1676.520 1395.930 1685.320 ;
        RECT 300.915 1675.120 1395.530 1676.520 ;
      LAYER met3 ;
        RECT 1395.930 1676.010 1399.930 1676.120 ;
        RECT 1408.125 1676.010 1408.455 1676.025 ;
        RECT 1395.930 1675.710 1408.455 1676.010 ;
        RECT 1395.930 1675.520 1399.930 1675.710 ;
        RECT 1408.125 1675.695 1408.455 1675.710 ;
      LAYER met3 ;
        RECT 300.915 1666.320 1395.930 1675.120 ;
        RECT 300.915 1664.920 1395.530 1666.320 ;
      LAYER met3 ;
        RECT 1395.930 1665.810 1399.930 1665.920 ;
        RECT 1407.665 1665.810 1407.995 1665.825 ;
        RECT 1395.930 1665.510 1407.995 1665.810 ;
        RECT 1395.930 1665.320 1399.930 1665.510 ;
        RECT 1407.665 1665.495 1407.995 1665.510 ;
      LAYER met3 ;
        RECT 300.915 1656.120 1395.930 1664.920 ;
        RECT 300.915 1654.720 1395.530 1656.120 ;
      LAYER met3 ;
        RECT 1395.930 1655.610 1399.930 1655.720 ;
        RECT 1407.665 1655.610 1407.995 1655.625 ;
        RECT 1395.930 1655.310 1407.995 1655.610 ;
        RECT 1395.930 1655.120 1399.930 1655.310 ;
        RECT 1407.665 1655.295 1407.995 1655.310 ;
      LAYER met3 ;
        RECT 300.915 1645.920 1395.930 1654.720 ;
        RECT 300.915 1644.520 1395.530 1645.920 ;
      LAYER met3 ;
        RECT 1395.930 1645.410 1399.930 1645.520 ;
        RECT 1407.665 1645.410 1407.995 1645.425 ;
        RECT 1395.930 1645.110 1407.995 1645.410 ;
        RECT 1395.930 1644.920 1399.930 1645.110 ;
        RECT 1407.665 1645.095 1407.995 1645.110 ;
      LAYER met3 ;
        RECT 300.915 1635.720 1395.930 1644.520 ;
        RECT 300.915 1634.320 1395.530 1635.720 ;
      LAYER met3 ;
        RECT 1395.930 1635.210 1399.930 1635.320 ;
        RECT 1407.665 1635.210 1407.995 1635.225 ;
        RECT 1395.930 1634.910 1407.995 1635.210 ;
        RECT 1395.930 1634.720 1399.930 1634.910 ;
        RECT 1407.665 1634.895 1407.995 1634.910 ;
      LAYER met3 ;
        RECT 300.915 1625.520 1395.930 1634.320 ;
        RECT 300.915 1624.120 1395.530 1625.520 ;
      LAYER met3 ;
        RECT 1395.930 1625.010 1399.930 1625.120 ;
        RECT 1407.665 1625.010 1407.995 1625.025 ;
        RECT 1395.930 1624.710 1407.995 1625.010 ;
        RECT 1395.930 1624.520 1399.930 1624.710 ;
        RECT 1407.665 1624.695 1407.995 1624.710 ;
      LAYER met3 ;
        RECT 300.915 1615.320 1395.930 1624.120 ;
        RECT 300.915 1613.920 1395.530 1615.320 ;
      LAYER met3 ;
        RECT 1395.930 1614.810 1399.930 1614.920 ;
        RECT 1411.550 1614.810 1411.930 1614.820 ;
        RECT 1395.930 1614.510 1411.930 1614.810 ;
        RECT 1395.930 1614.320 1399.930 1614.510 ;
        RECT 1411.550 1614.500 1411.930 1614.510 ;
      LAYER met3 ;
        RECT 300.915 1605.800 1395.930 1613.920 ;
      LAYER met3 ;
        RECT 1550.000 1607.670 1554.600 1607.970 ;
      LAYER met3 ;
        RECT 300.915 1604.935 1395.530 1605.800 ;
      LAYER met3 ;
        RECT 1395.930 1605.290 1399.930 1605.400 ;
        RECT 1410.885 1605.290 1411.215 1605.305 ;
        RECT 1395.930 1604.990 1411.215 1605.290 ;
      LAYER met3 ;
        RECT 1555.000 1605.000 1931.480 2051.235 ;
      LAYER met3 ;
        RECT 2200.000 2032.785 2204.600 2033.085 ;
        RECT 2200.000 2027.145 2204.600 2027.445 ;
        RECT 2200.000 2018.645 2204.600 2018.945 ;
        RECT 2200.000 2013.005 2204.600 2013.305 ;
        RECT 2200.000 2004.505 2204.600 2004.805 ;
        RECT 2200.000 1998.865 2204.600 1999.165 ;
        RECT 2200.000 1990.365 2204.600 1990.665 ;
        RECT 1931.880 1963.310 1936.480 1963.610 ;
        RECT 1931.880 1954.810 1936.480 1955.110 ;
        RECT 2200.000 1701.125 2204.600 1701.425 ;
        RECT 2200.000 1692.625 2204.600 1692.925 ;
        RECT 1931.880 1665.570 1936.480 1665.870 ;
        RECT 1931.880 1657.070 1936.480 1657.370 ;
        RECT 1931.880 1651.430 1936.480 1651.730 ;
        RECT 1931.880 1642.930 1936.480 1643.230 ;
        RECT 1931.880 1637.290 1936.480 1637.590 ;
        RECT 1931.880 1628.790 1936.480 1629.090 ;
        RECT 1931.880 1623.150 1936.480 1623.450 ;
      LAYER met3 ;
        RECT 2205.000 1605.000 2581.480 2051.235 ;
      LAYER met3 ;
        RECT 2581.880 2048.265 2586.480 2048.565 ;
        RECT 2581.880 1746.910 2586.480 1747.210 ;
        RECT 2581.880 1738.410 2586.480 1738.710 ;
        RECT 2581.880 1732.770 2586.480 1733.070 ;
        RECT 2581.880 1724.270 2586.480 1724.570 ;
        RECT 2581.880 1718.630 2586.480 1718.930 ;
        RECT 2581.880 1710.130 2586.480 1710.430 ;
        RECT 2581.880 1704.490 2586.480 1704.790 ;
        RECT 1395.930 1604.800 1399.930 1604.990 ;
        RECT 1410.885 1604.975 1411.215 1604.990 ;
        RECT 1575.460 1604.095 1577.200 1605.000 ;
      LAYER met3 ;
        RECT 1550.915 1494.440 2645.530 1495.305 ;
      LAYER met3 ;
        RECT 2645.930 1494.840 2649.930 1495.440 ;
      LAYER met3 ;
        RECT 1550.915 1485.640 2645.930 1494.440 ;
        RECT 1550.915 1484.240 2645.530 1485.640 ;
      LAYER met3 ;
        RECT 2645.930 1484.640 2649.930 1485.240 ;
      LAYER met3 ;
        RECT 1550.915 1475.440 2645.930 1484.240 ;
        RECT 1550.915 1474.040 2645.530 1475.440 ;
      LAYER met3 ;
        RECT 2645.930 1474.440 2649.930 1475.040 ;
      LAYER met3 ;
        RECT 1550.915 1465.240 2645.930 1474.040 ;
        RECT 1550.915 1463.840 2645.530 1465.240 ;
      LAYER met3 ;
        RECT 2645.930 1464.240 2649.930 1464.840 ;
      LAYER met3 ;
        RECT 1550.915 1455.040 2645.930 1463.840 ;
        RECT 1550.915 1453.640 2645.530 1455.040 ;
      LAYER met3 ;
        RECT 2645.930 1454.040 2649.930 1454.640 ;
      LAYER met3 ;
        RECT 1550.915 1444.840 2645.930 1453.640 ;
        RECT 1550.915 1443.440 2645.530 1444.840 ;
      LAYER met3 ;
        RECT 2645.930 1443.840 2649.930 1444.440 ;
      LAYER met3 ;
        RECT 1550.915 1434.640 2645.930 1443.440 ;
        RECT 1550.915 1433.240 2645.530 1434.640 ;
      LAYER met3 ;
        RECT 2645.930 1433.640 2649.930 1434.240 ;
      LAYER met3 ;
        RECT 1550.915 1424.440 2645.930 1433.240 ;
        RECT 1550.915 1423.040 2645.530 1424.440 ;
      LAYER met3 ;
        RECT 2645.930 1423.440 2649.930 1424.040 ;
      LAYER met3 ;
        RECT 1550.915 1414.240 2645.930 1423.040 ;
        RECT 1550.915 1412.840 2645.530 1414.240 ;
      LAYER met3 ;
        RECT 2645.930 1413.240 2649.930 1413.840 ;
      LAYER met3 ;
        RECT 1550.915 1404.040 2645.930 1412.840 ;
        RECT 1550.915 1402.640 2645.530 1404.040 ;
      LAYER met3 ;
        RECT 2645.930 1403.040 2649.930 1403.640 ;
      LAYER met3 ;
        RECT 1550.915 1393.840 2645.930 1402.640 ;
        RECT 1550.915 1392.440 2645.530 1393.840 ;
      LAYER met3 ;
        RECT 2645.930 1392.840 2649.930 1393.440 ;
      LAYER met3 ;
        RECT 1550.915 1383.640 2645.930 1392.440 ;
        RECT 1550.915 1382.240 2645.530 1383.640 ;
      LAYER met3 ;
        RECT 2645.930 1382.640 2649.930 1383.240 ;
      LAYER met3 ;
        RECT 1550.915 1373.440 2645.930 1382.240 ;
        RECT 1550.915 1372.040 2645.530 1373.440 ;
      LAYER met3 ;
        RECT 2645.930 1372.440 2649.930 1373.040 ;
      LAYER met3 ;
        RECT 1550.915 1363.240 2645.930 1372.040 ;
        RECT 1550.915 1361.840 2645.530 1363.240 ;
      LAYER met3 ;
        RECT 2645.930 1362.240 2649.930 1362.840 ;
      LAYER met3 ;
        RECT 1550.915 1353.040 2645.930 1361.840 ;
        RECT 1550.915 1351.640 2645.530 1353.040 ;
      LAYER met3 ;
        RECT 2645.930 1352.040 2649.930 1352.640 ;
      LAYER met3 ;
        RECT 1550.915 1342.840 2645.930 1351.640 ;
        RECT 1550.915 1341.440 2645.530 1342.840 ;
      LAYER met3 ;
        RECT 2645.930 1341.840 2649.930 1342.440 ;
      LAYER met3 ;
        RECT 1550.915 1332.640 2645.930 1341.440 ;
        RECT 1550.915 1331.240 2645.530 1332.640 ;
      LAYER met3 ;
        RECT 2645.930 1331.640 2649.930 1332.240 ;
      LAYER met3 ;
        RECT 1550.915 1322.440 2645.930 1331.240 ;
        RECT 1550.915 1321.040 2645.530 1322.440 ;
      LAYER met3 ;
        RECT 2645.930 1321.440 2649.930 1322.040 ;
      LAYER met3 ;
        RECT 1550.915 1312.240 2645.930 1321.040 ;
        RECT 1550.915 1310.840 2645.530 1312.240 ;
      LAYER met3 ;
        RECT 2645.930 1311.240 2649.930 1311.840 ;
      LAYER met3 ;
        RECT 1550.915 1302.040 2645.930 1310.840 ;
        RECT 1550.915 1300.640 2645.530 1302.040 ;
      LAYER met3 ;
        RECT 2645.930 1301.040 2649.930 1301.640 ;
      LAYER met3 ;
        RECT 1550.915 1291.840 2645.930 1300.640 ;
        RECT 1550.915 1290.440 2645.530 1291.840 ;
      LAYER met3 ;
        RECT 2645.930 1290.840 2649.930 1291.440 ;
      LAYER met3 ;
        RECT 1550.915 1281.640 2645.930 1290.440 ;
        RECT 1550.915 1280.240 2645.530 1281.640 ;
      LAYER met3 ;
        RECT 2645.930 1280.640 2649.930 1281.240 ;
      LAYER met3 ;
        RECT 1550.915 1271.440 2645.930 1280.240 ;
        RECT 1550.915 1270.040 2645.530 1271.440 ;
      LAYER met3 ;
        RECT 2645.930 1270.440 2649.930 1271.040 ;
      LAYER met3 ;
        RECT 1550.915 1261.240 2645.930 1270.040 ;
        RECT 1550.915 1259.840 2645.530 1261.240 ;
      LAYER met3 ;
        RECT 2645.930 1260.240 2649.930 1260.840 ;
      LAYER met3 ;
        RECT 1550.915 1251.040 2645.930 1259.840 ;
        RECT 1550.915 1249.640 2645.530 1251.040 ;
      LAYER met3 ;
        RECT 2645.930 1250.040 2649.930 1250.640 ;
      LAYER met3 ;
        RECT 1550.915 1240.840 2645.930 1249.640 ;
        RECT 1550.915 1239.440 2645.530 1240.840 ;
      LAYER met3 ;
        RECT 2645.930 1239.840 2649.930 1240.440 ;
      LAYER met3 ;
        RECT 1550.915 1230.640 2645.930 1239.440 ;
        RECT 1550.915 1229.240 2645.530 1230.640 ;
      LAYER met3 ;
        RECT 2645.930 1229.640 2649.930 1230.240 ;
      LAYER met3 ;
        RECT 1550.915 1220.440 2645.930 1229.240 ;
        RECT 1550.915 1219.040 2645.530 1220.440 ;
      LAYER met3 ;
        RECT 2645.930 1219.440 2649.930 1220.040 ;
      LAYER met3 ;
        RECT 1550.915 1210.240 2645.930 1219.040 ;
        RECT 1550.915 1208.840 2645.530 1210.240 ;
      LAYER met3 ;
        RECT 2645.930 1209.240 2649.930 1209.840 ;
      LAYER met3 ;
        RECT 1550.915 1200.040 2645.930 1208.840 ;
        RECT 1550.915 1198.640 2645.530 1200.040 ;
      LAYER met3 ;
        RECT 2645.930 1199.040 2649.930 1199.640 ;
      LAYER met3 ;
        RECT 1550.915 1189.840 2645.930 1198.640 ;
        RECT 1550.915 1188.440 2645.530 1189.840 ;
      LAYER met3 ;
        RECT 2645.930 1188.840 2649.930 1189.440 ;
      LAYER met3 ;
        RECT 1550.915 1179.640 2645.930 1188.440 ;
        RECT 1550.915 1178.240 2645.530 1179.640 ;
      LAYER met3 ;
        RECT 2645.930 1178.640 2649.930 1179.240 ;
      LAYER met3 ;
        RECT 1550.915 1169.440 2645.930 1178.240 ;
        RECT 1550.915 1168.040 2645.530 1169.440 ;
      LAYER met3 ;
        RECT 2645.930 1168.440 2649.930 1169.040 ;
      LAYER met3 ;
        RECT 1550.915 1159.240 2645.930 1168.040 ;
        RECT 1550.915 1157.840 2645.530 1159.240 ;
      LAYER met3 ;
        RECT 2645.930 1158.240 2649.930 1158.840 ;
      LAYER met3 ;
        RECT 1550.915 1149.040 2645.930 1157.840 ;
        RECT 1550.915 1147.640 2645.530 1149.040 ;
      LAYER met3 ;
        RECT 2645.930 1148.040 2649.930 1148.640 ;
      LAYER met3 ;
        RECT 1550.915 1138.840 2645.930 1147.640 ;
        RECT 1550.915 1137.440 2645.530 1138.840 ;
      LAYER met3 ;
        RECT 2645.930 1137.840 2649.930 1138.440 ;
      LAYER met3 ;
        RECT 1550.915 1128.640 2645.930 1137.440 ;
        RECT 1550.915 1127.240 2645.530 1128.640 ;
      LAYER met3 ;
        RECT 2645.930 1127.640 2649.930 1128.240 ;
      LAYER met3 ;
        RECT 1550.915 1118.440 2645.930 1127.240 ;
        RECT 1550.915 1117.040 2645.530 1118.440 ;
      LAYER met3 ;
        RECT 2645.930 1117.440 2649.930 1118.040 ;
      LAYER met3 ;
        RECT 1550.915 1108.240 2645.930 1117.040 ;
        RECT 1550.915 1106.840 2645.530 1108.240 ;
      LAYER met3 ;
        RECT 2645.930 1107.240 2649.930 1107.840 ;
      LAYER met3 ;
        RECT 1550.915 1098.040 2645.930 1106.840 ;
        RECT 1550.915 1096.640 2645.530 1098.040 ;
      LAYER met3 ;
        RECT 2645.930 1097.040 2649.930 1097.640 ;
      LAYER met3 ;
        RECT 1550.915 1087.840 2645.930 1096.640 ;
        RECT 1550.915 1086.440 2645.530 1087.840 ;
      LAYER met3 ;
        RECT 2645.930 1086.840 2649.930 1087.440 ;
      LAYER met3 ;
        RECT 1550.915 1077.640 2645.930 1086.440 ;
        RECT 1550.915 1076.240 2645.530 1077.640 ;
      LAYER met3 ;
        RECT 2645.930 1076.640 2649.930 1077.240 ;
      LAYER met3 ;
        RECT 1550.915 1067.440 2645.930 1076.240 ;
        RECT 1550.915 1066.040 2645.530 1067.440 ;
      LAYER met3 ;
        RECT 2645.930 1066.440 2649.930 1067.040 ;
      LAYER met3 ;
        RECT 1550.915 1057.240 2645.930 1066.040 ;
        RECT 1550.915 1055.840 2645.530 1057.240 ;
      LAYER met3 ;
        RECT 2645.930 1056.240 2649.930 1056.840 ;
      LAYER met3 ;
        RECT 1550.915 1047.040 2645.930 1055.840 ;
        RECT 1550.915 1045.640 2645.530 1047.040 ;
      LAYER met3 ;
        RECT 2645.930 1046.040 2649.930 1046.640 ;
      LAYER met3 ;
        RECT 1550.915 1036.840 2645.930 1045.640 ;
        RECT 1550.915 1035.440 2645.530 1036.840 ;
      LAYER met3 ;
        RECT 2645.930 1035.840 2649.930 1036.440 ;
      LAYER met3 ;
        RECT 1550.915 1026.640 2645.930 1035.440 ;
        RECT 1550.915 1025.240 2645.530 1026.640 ;
      LAYER met3 ;
        RECT 2645.930 1025.640 2649.930 1026.240 ;
      LAYER met3 ;
        RECT 1550.915 1016.440 2645.930 1025.240 ;
        RECT 1550.915 1015.040 2645.530 1016.440 ;
      LAYER met3 ;
        RECT 2645.930 1015.440 2649.930 1016.040 ;
      LAYER met3 ;
        RECT 1550.915 1006.240 2645.930 1015.040 ;
        RECT 1550.915 1004.840 2645.530 1006.240 ;
      LAYER met3 ;
        RECT 2645.930 1005.240 2649.930 1005.840 ;
      LAYER met3 ;
        RECT 1550.915 996.040 2645.930 1004.840 ;
        RECT 1550.915 994.640 2645.530 996.040 ;
      LAYER met3 ;
        RECT 2645.930 995.040 2649.930 995.640 ;
      LAYER met3 ;
        RECT 1550.915 985.840 2645.930 994.640 ;
        RECT 1550.915 984.440 2645.530 985.840 ;
      LAYER met3 ;
        RECT 2645.930 984.840 2649.930 985.440 ;
      LAYER met3 ;
        RECT 1550.915 975.640 2645.930 984.440 ;
        RECT 1550.915 974.240 2645.530 975.640 ;
      LAYER met3 ;
        RECT 2645.930 974.640 2649.930 975.240 ;
      LAYER met3 ;
        RECT 1550.915 965.440 2645.930 974.240 ;
        RECT 1550.915 964.040 2645.530 965.440 ;
      LAYER met3 ;
        RECT 2645.930 964.440 2649.930 965.040 ;
      LAYER met3 ;
        RECT 1550.915 955.920 2645.930 964.040 ;
        RECT 1550.915 954.520 2645.530 955.920 ;
      LAYER met3 ;
        RECT 2645.930 954.920 2649.930 955.520 ;
      LAYER met3 ;
        RECT 1550.915 945.720 2645.930 954.520 ;
        RECT 1550.915 944.320 2645.530 945.720 ;
      LAYER met3 ;
        RECT 2645.930 944.720 2649.930 945.320 ;
      LAYER met3 ;
        RECT 1550.915 935.520 2645.930 944.320 ;
        RECT 1550.915 934.120 2645.530 935.520 ;
      LAYER met3 ;
        RECT 2645.930 934.520 2649.930 935.120 ;
      LAYER met3 ;
        RECT 1550.915 925.320 2645.930 934.120 ;
        RECT 1550.915 923.920 2645.530 925.320 ;
      LAYER met3 ;
        RECT 2645.930 924.320 2649.930 924.920 ;
      LAYER met3 ;
        RECT 1550.915 915.120 2645.930 923.920 ;
        RECT 1550.915 913.720 2645.530 915.120 ;
      LAYER met3 ;
        RECT 2645.930 914.120 2649.930 914.720 ;
      LAYER met3 ;
        RECT 1550.915 904.920 2645.930 913.720 ;
        RECT 1550.915 903.520 2645.530 904.920 ;
      LAYER met3 ;
        RECT 2645.930 903.920 2649.930 904.520 ;
      LAYER met3 ;
        RECT 1550.915 894.720 2645.930 903.520 ;
        RECT 1550.915 893.320 2645.530 894.720 ;
      LAYER met3 ;
        RECT 2645.930 893.720 2649.930 894.320 ;
      LAYER met3 ;
        RECT 1550.915 884.520 2645.930 893.320 ;
        RECT 1550.915 883.120 2645.530 884.520 ;
      LAYER met3 ;
        RECT 2645.930 883.520 2649.930 884.120 ;
      LAYER met3 ;
        RECT 1550.915 874.320 2645.930 883.120 ;
        RECT 1550.915 872.920 2645.530 874.320 ;
      LAYER met3 ;
        RECT 2645.930 873.320 2649.930 873.920 ;
      LAYER met3 ;
        RECT 1550.915 864.120 2645.930 872.920 ;
        RECT 1550.915 862.720 2645.530 864.120 ;
      LAYER met3 ;
        RECT 2645.930 863.120 2649.930 863.720 ;
      LAYER met3 ;
        RECT 1550.915 853.920 2645.930 862.720 ;
        RECT 1550.915 852.520 2645.530 853.920 ;
      LAYER met3 ;
        RECT 2645.930 852.920 2649.930 853.520 ;
      LAYER met3 ;
        RECT 1550.915 843.720 2645.930 852.520 ;
        RECT 1550.915 842.320 2645.530 843.720 ;
      LAYER met3 ;
        RECT 2645.930 842.720 2649.930 843.320 ;
      LAYER met3 ;
        RECT 1550.915 833.520 2645.930 842.320 ;
        RECT 1550.915 832.120 2645.530 833.520 ;
      LAYER met3 ;
        RECT 2645.930 832.520 2649.930 833.120 ;
      LAYER met3 ;
        RECT 1550.915 823.320 2645.930 832.120 ;
        RECT 1550.915 821.920 2645.530 823.320 ;
      LAYER met3 ;
        RECT 2645.930 822.320 2649.930 822.920 ;
      LAYER met3 ;
        RECT 1550.915 813.120 2645.930 821.920 ;
        RECT 1550.915 811.720 2645.530 813.120 ;
      LAYER met3 ;
        RECT 2645.930 812.120 2649.930 812.720 ;
      LAYER met3 ;
        RECT 1550.915 802.920 2645.930 811.720 ;
        RECT 1550.915 801.520 2645.530 802.920 ;
      LAYER met3 ;
        RECT 2645.930 801.920 2649.930 802.520 ;
      LAYER met3 ;
        RECT 1550.915 792.720 2645.930 801.520 ;
        RECT 1550.915 791.320 2645.530 792.720 ;
      LAYER met3 ;
        RECT 2645.930 791.720 2649.930 792.320 ;
      LAYER met3 ;
        RECT 1550.915 782.520 2645.930 791.320 ;
        RECT 1550.915 781.120 2645.530 782.520 ;
      LAYER met3 ;
        RECT 2645.930 781.520 2649.930 782.120 ;
      LAYER met3 ;
        RECT 1550.915 772.320 2645.930 781.120 ;
        RECT 1550.915 770.920 2645.530 772.320 ;
      LAYER met3 ;
        RECT 2645.930 771.320 2649.930 771.920 ;
      LAYER met3 ;
        RECT 1550.915 762.120 2645.930 770.920 ;
        RECT 1550.915 760.720 2645.530 762.120 ;
      LAYER met3 ;
        RECT 2645.930 761.120 2649.930 761.720 ;
      LAYER met3 ;
        RECT 1550.915 751.920 2645.930 760.720 ;
        RECT 1550.915 750.520 2645.530 751.920 ;
      LAYER met3 ;
        RECT 2645.930 750.920 2649.930 751.520 ;
      LAYER met3 ;
        RECT 1550.915 741.720 2645.930 750.520 ;
        RECT 1550.915 740.320 2645.530 741.720 ;
      LAYER met3 ;
        RECT 2645.930 740.720 2649.930 741.320 ;
      LAYER met3 ;
        RECT 1550.915 731.520 2645.930 740.320 ;
        RECT 1550.915 730.120 2645.530 731.520 ;
      LAYER met3 ;
        RECT 2645.930 730.520 2649.930 731.120 ;
      LAYER met3 ;
        RECT 1550.915 721.320 2645.930 730.120 ;
        RECT 1550.915 719.920 2645.530 721.320 ;
      LAYER met3 ;
        RECT 2645.930 720.320 2649.930 720.920 ;
      LAYER met3 ;
        RECT 1550.915 711.120 2645.930 719.920 ;
        RECT 1550.915 709.720 2645.530 711.120 ;
      LAYER met3 ;
        RECT 2645.930 710.120 2649.930 710.720 ;
      LAYER met3 ;
        RECT 1550.915 700.920 2645.930 709.720 ;
        RECT 1550.915 699.520 2645.530 700.920 ;
      LAYER met3 ;
        RECT 2645.930 699.920 2649.930 700.520 ;
      LAYER met3 ;
        RECT 1550.915 690.720 2645.930 699.520 ;
        RECT 1550.915 689.320 2645.530 690.720 ;
      LAYER met3 ;
        RECT 2645.930 689.720 2649.930 690.320 ;
      LAYER met3 ;
        RECT 1550.915 680.520 2645.930 689.320 ;
        RECT 1550.915 679.120 2645.530 680.520 ;
      LAYER met3 ;
        RECT 2645.930 679.520 2649.930 680.120 ;
      LAYER met3 ;
        RECT 1550.915 670.320 2645.930 679.120 ;
        RECT 1550.915 668.920 2645.530 670.320 ;
      LAYER met3 ;
        RECT 2645.930 669.320 2649.930 669.920 ;
      LAYER met3 ;
        RECT 1550.915 660.120 2645.930 668.920 ;
        RECT 1550.915 658.720 2645.530 660.120 ;
      LAYER met3 ;
        RECT 2645.930 659.120 2649.930 659.720 ;
      LAYER met3 ;
        RECT 1550.915 649.920 2645.930 658.720 ;
        RECT 1550.915 648.520 2645.530 649.920 ;
      LAYER met3 ;
        RECT 2645.930 648.920 2649.930 649.520 ;
      LAYER met3 ;
        RECT 1550.915 639.720 2645.930 648.520 ;
        RECT 1550.915 638.320 2645.530 639.720 ;
      LAYER met3 ;
        RECT 2645.930 638.720 2649.930 639.320 ;
      LAYER met3 ;
        RECT 1550.915 629.520 2645.930 638.320 ;
        RECT 1550.915 628.120 2645.530 629.520 ;
      LAYER met3 ;
        RECT 2645.930 628.520 2649.930 629.120 ;
      LAYER met3 ;
        RECT 1550.915 619.320 2645.930 628.120 ;
        RECT 1550.915 617.920 2645.530 619.320 ;
      LAYER met3 ;
        RECT 2645.930 618.320 2649.930 618.920 ;
      LAYER met3 ;
        RECT 1550.915 609.120 2645.930 617.920 ;
        RECT 1550.915 607.720 2645.530 609.120 ;
      LAYER met3 ;
        RECT 2645.930 608.120 2649.930 608.720 ;
      LAYER met3 ;
        RECT 1550.915 598.920 2645.930 607.720 ;
        RECT 1550.915 597.520 2645.530 598.920 ;
      LAYER met3 ;
        RECT 2645.930 597.920 2649.930 598.520 ;
      LAYER met3 ;
        RECT 1550.915 588.720 2645.930 597.520 ;
        RECT 1550.915 587.320 2645.530 588.720 ;
      LAYER met3 ;
        RECT 2645.930 587.720 2649.930 588.320 ;
      LAYER met3 ;
        RECT 1550.915 578.520 2645.930 587.320 ;
        RECT 1550.915 577.120 2645.530 578.520 ;
      LAYER met3 ;
        RECT 2645.930 577.520 2649.930 578.120 ;
      LAYER met3 ;
        RECT 1550.915 568.320 2645.930 577.120 ;
        RECT 1550.915 566.920 2645.530 568.320 ;
      LAYER met3 ;
        RECT 2645.930 567.320 2649.930 567.920 ;
      LAYER met3 ;
        RECT 1550.915 558.120 2645.930 566.920 ;
        RECT 1550.915 556.720 2645.530 558.120 ;
      LAYER met3 ;
        RECT 2645.930 557.120 2649.930 557.720 ;
      LAYER met3 ;
        RECT 1550.915 547.920 2645.930 556.720 ;
        RECT 1550.915 546.520 2645.530 547.920 ;
      LAYER met3 ;
        RECT 2645.930 546.920 2649.930 547.520 ;
      LAYER met3 ;
        RECT 1550.915 537.720 2645.930 546.520 ;
        RECT 1550.915 536.320 2645.530 537.720 ;
      LAYER met3 ;
        RECT 2645.930 536.720 2649.930 537.320 ;
      LAYER met3 ;
        RECT 1550.915 527.520 2645.930 536.320 ;
        RECT 1550.915 526.120 2645.530 527.520 ;
      LAYER met3 ;
        RECT 2645.930 526.520 2649.930 527.120 ;
      LAYER met3 ;
        RECT 1550.915 517.320 2645.930 526.120 ;
        RECT 1550.915 515.920 2645.530 517.320 ;
      LAYER met3 ;
        RECT 2645.930 516.320 2649.930 516.920 ;
      LAYER met3 ;
        RECT 1550.915 507.120 2645.930 515.920 ;
        RECT 1550.915 505.720 2645.530 507.120 ;
      LAYER met3 ;
        RECT 2645.930 506.120 2649.930 506.720 ;
      LAYER met3 ;
        RECT 1550.915 496.920 2645.930 505.720 ;
        RECT 1550.915 495.520 2645.530 496.920 ;
      LAYER met3 ;
        RECT 2645.930 495.920 2649.930 496.520 ;
      LAYER met3 ;
        RECT 1550.915 486.720 2645.930 495.520 ;
        RECT 1550.915 485.320 2645.530 486.720 ;
      LAYER met3 ;
        RECT 2645.930 485.720 2649.930 486.320 ;
      LAYER met3 ;
        RECT 1550.915 476.520 2645.930 485.320 ;
        RECT 1550.915 475.120 2645.530 476.520 ;
      LAYER met3 ;
        RECT 2645.930 475.520 2649.930 476.120 ;
      LAYER met3 ;
        RECT 1550.915 466.320 2645.930 475.120 ;
        RECT 1550.915 464.920 2645.530 466.320 ;
      LAYER met3 ;
        RECT 2645.930 465.320 2649.930 465.920 ;
      LAYER met3 ;
        RECT 1550.915 456.120 2645.930 464.920 ;
        RECT 1550.915 454.720 2645.530 456.120 ;
      LAYER met3 ;
        RECT 2645.930 455.120 2649.930 455.720 ;
      LAYER met3 ;
        RECT 1550.915 445.920 2645.930 454.720 ;
        RECT 1550.915 444.520 2645.530 445.920 ;
      LAYER met3 ;
        RECT 2645.930 444.920 2649.930 445.520 ;
      LAYER met3 ;
        RECT 1550.915 435.720 2645.930 444.520 ;
        RECT 1550.915 434.320 2645.530 435.720 ;
      LAYER met3 ;
        RECT 2645.930 434.720 2649.930 435.320 ;
      LAYER met3 ;
        RECT 1550.915 425.520 2645.930 434.320 ;
        RECT 1550.915 424.120 2645.530 425.520 ;
      LAYER met3 ;
        RECT 2645.930 424.520 2649.930 425.120 ;
      LAYER met3 ;
        RECT 1550.915 415.320 2645.930 424.120 ;
        RECT 1550.915 413.920 2645.530 415.320 ;
      LAYER met3 ;
        RECT 2645.930 414.320 2649.930 414.920 ;
      LAYER met3 ;
        RECT 1550.915 405.800 2645.930 413.920 ;
        RECT 1550.915 404.935 2645.530 405.800 ;
      LAYER met3 ;
        RECT 2645.930 404.800 2649.930 405.400 ;
      LAYER via3 ;
        RECT 646.140 3264.180 646.460 3264.500 ;
        RECT 668.220 3264.180 668.540 3264.500 ;
        RECT 1295.660 3264.180 1295.980 3264.500 ;
        RECT 1317.740 3264.180 1318.060 3264.500 ;
        RECT 1890.900 3264.180 1891.220 3264.500 ;
        RECT 1917.580 3264.180 1917.900 3264.500 ;
        RECT 2542.260 3264.180 2542.580 3264.500 ;
        RECT 2567.100 3264.180 2567.420 3264.500 ;
        RECT 302.980 2894.940 303.300 2895.260 ;
        RECT 687.540 2901.740 687.860 2902.060 ;
        RECT 950.660 2894.940 950.980 2895.260 ;
        RECT 1411.580 3243.100 1411.900 3243.420 ;
        RECT 1413.420 2935.740 1413.740 2936.060 ;
        RECT 1345.340 2904.460 1345.660 2904.780 ;
        RECT 1937.820 2935.740 1938.140 2936.060 ;
        RECT 2200.020 2895.620 2200.340 2895.940 ;
        RECT 2594.700 2904.460 2595.020 2904.780 ;
        RECT 1146.620 2799.740 1146.940 2800.060 ;
        RECT 1129.140 2799.060 1129.460 2799.380 ;
        RECT 1135.580 2796.340 1135.900 2796.660 ;
        RECT 1759.340 2796.340 1759.660 2796.660 ;
        RECT 1794.300 2796.340 1794.620 2796.660 ;
        RECT 337.020 2794.300 337.340 2794.620 ;
        RECT 342.540 2794.300 342.860 2794.620 ;
        RECT 350.820 2794.300 351.140 2794.620 ;
        RECT 358.180 2794.300 358.500 2794.620 ;
        RECT 361.860 2794.300 362.180 2794.620 ;
        RECT 364.620 2794.300 364.940 2794.620 ;
        RECT 368.300 2794.300 368.620 2794.620 ;
        RECT 371.060 2794.300 371.380 2794.620 ;
        RECT 374.740 2794.300 375.060 2794.620 ;
        RECT 378.420 2794.300 378.740 2794.620 ;
        RECT 383.940 2794.300 384.260 2794.620 ;
        RECT 386.700 2794.300 387.020 2794.620 ;
        RECT 390.380 2794.300 390.700 2794.620 ;
        RECT 395.900 2794.300 396.220 2794.620 ;
        RECT 399.580 2794.300 399.900 2794.620 ;
        RECT 403.260 2794.300 403.580 2794.620 ;
        RECT 406.020 2794.300 406.340 2794.620 ;
        RECT 409.700 2794.300 410.020 2794.620 ;
        RECT 413.380 2794.300 413.700 2794.620 ;
        RECT 418.900 2794.300 419.220 2794.620 ;
        RECT 420.740 2794.300 421.060 2794.620 ;
        RECT 425.340 2794.300 425.660 2794.620 ;
        RECT 433.620 2794.300 433.940 2794.620 ;
        RECT 439.140 2794.300 439.460 2794.620 ;
        RECT 440.980 2794.300 441.300 2794.620 ;
        RECT 444.660 2794.300 444.980 2794.620 ;
        RECT 445.580 2794.300 445.900 2794.620 ;
        RECT 449.260 2794.300 449.580 2794.620 ;
        RECT 454.780 2794.300 455.100 2794.620 ;
        RECT 460.300 2794.300 460.620 2794.620 ;
        RECT 462.140 2794.300 462.460 2794.620 ;
        RECT 465.820 2794.300 466.140 2794.620 ;
        RECT 474.100 2794.300 474.420 2794.620 ;
        RECT 475.020 2794.300 475.340 2794.620 ;
        RECT 478.700 2794.300 479.020 2794.620 ;
        RECT 482.380 2794.300 482.700 2794.620 ;
        RECT 485.140 2794.300 485.460 2794.620 ;
        RECT 487.900 2794.300 488.220 2794.620 ;
        RECT 491.580 2794.300 491.900 2794.620 ;
        RECT 495.260 2794.300 495.580 2794.620 ;
        RECT 500.780 2794.300 501.100 2794.620 ;
        RECT 509.980 2794.300 510.300 2794.620 ;
        RECT 523.780 2794.300 524.100 2794.620 ;
        RECT 535.740 2794.300 536.060 2794.620 ;
        RECT 542.180 2794.300 542.500 2794.620 ;
        RECT 981.020 2794.300 981.340 2794.620 ;
        RECT 1001.260 2794.300 1001.580 2794.620 ;
        RECT 1007.700 2794.300 1008.020 2794.620 ;
        RECT 1013.220 2794.300 1013.540 2794.620 ;
        RECT 1018.740 2794.300 1019.060 2794.620 ;
        RECT 1019.660 2794.300 1019.980 2794.620 ;
        RECT 1027.020 2794.300 1027.340 2794.620 ;
        RECT 1030.700 2794.300 1031.020 2794.620 ;
        RECT 1041.740 2794.300 1042.060 2794.620 ;
        RECT 1059.220 2794.300 1059.540 2794.620 ;
        RECT 1065.660 2794.300 1065.980 2794.620 ;
        RECT 1070.260 2794.300 1070.580 2794.620 ;
        RECT 1076.700 2794.300 1077.020 2794.620 ;
        RECT 1094.180 2794.300 1094.500 2794.620 ;
        RECT 1100.620 2794.300 1100.940 2794.620 ;
        RECT 1105.220 2794.300 1105.540 2794.620 ;
        RECT 1111.660 2794.300 1111.980 2794.620 ;
        RECT 1118.100 2794.300 1118.420 2794.620 ;
        RECT 1122.700 2794.300 1123.020 2794.620 ;
        RECT 1140.180 2794.300 1140.500 2794.620 ;
        RECT 1178.820 2794.300 1179.140 2794.620 ;
        RECT 1186.180 2794.300 1186.500 2794.620 ;
        RECT 1198.140 2794.300 1198.460 2794.620 ;
        RECT 1580.860 2794.300 1581.180 2794.620 ;
        RECT 1587.300 2794.300 1587.620 2794.620 ;
        RECT 1604.780 2794.300 1605.100 2794.620 ;
        RECT 1613.060 2794.300 1613.380 2794.620 ;
        RECT 1617.660 2794.300 1617.980 2794.620 ;
        RECT 1642.500 2794.300 1642.820 2794.620 ;
        RECT 1648.020 2794.300 1648.340 2794.620 ;
        RECT 1652.620 2794.300 1652.940 2794.620 ;
        RECT 1659.060 2794.300 1659.380 2794.620 ;
        RECT 1665.500 2794.300 1665.820 2794.620 ;
        RECT 1670.100 2794.300 1670.420 2794.620 ;
        RECT 1677.460 2794.300 1677.780 2794.620 ;
        RECT 1682.060 2794.300 1682.380 2794.620 ;
        RECT 1688.500 2794.300 1688.820 2794.620 ;
        RECT 1694.940 2794.300 1695.260 2794.620 ;
        RECT 1699.540 2794.300 1699.860 2794.620 ;
        RECT 1705.980 2794.300 1706.300 2794.620 ;
        RECT 1712.420 2794.300 1712.740 2794.620 ;
        RECT 1717.940 2794.300 1718.260 2794.620 ;
        RECT 1723.460 2794.300 1723.780 2794.620 ;
        RECT 1728.980 2794.300 1729.300 2794.620 ;
        RECT 1732.660 2794.300 1732.980 2794.620 ;
        RECT 1740.940 2794.300 1741.260 2794.620 ;
        RECT 1747.380 2794.300 1747.700 2794.620 ;
        RECT 1752.900 2794.300 1753.220 2794.620 ;
        RECT 1762.100 2794.300 1762.420 2794.620 ;
        RECT 1767.620 2794.300 1767.940 2794.620 ;
        RECT 2231.300 2794.300 2231.620 2794.620 ;
        RECT 2238.660 2794.300 2238.980 2794.620 ;
        RECT 2268.100 2794.300 2268.420 2794.620 ;
        RECT 2273.620 2794.300 2273.940 2794.620 ;
        RECT 2280.060 2794.300 2280.380 2794.620 ;
        RECT 2286.500 2794.300 2286.820 2794.620 ;
        RECT 2291.100 2794.300 2291.420 2794.620 ;
        RECT 2303.980 2794.300 2304.300 2794.620 ;
        RECT 2308.580 2794.300 2308.900 2794.620 ;
        RECT 2313.180 2794.300 2313.500 2794.620 ;
        RECT 2321.460 2794.300 2321.780 2794.620 ;
        RECT 2326.060 2794.300 2326.380 2794.620 ;
        RECT 2334.340 2794.300 2334.660 2794.620 ;
        RECT 2339.860 2794.300 2340.180 2794.620 ;
        RECT 2343.540 2794.300 2343.860 2794.620 ;
        RECT 2351.820 2794.300 2352.140 2794.620 ;
        RECT 2357.340 2794.300 2357.660 2794.620 ;
        RECT 2363.780 2794.300 2364.100 2794.620 ;
        RECT 2370.220 2794.300 2370.540 2794.620 ;
        RECT 2373.900 2794.300 2374.220 2794.620 ;
        RECT 2377.580 2794.300 2377.900 2794.620 ;
        RECT 2385.860 2794.300 2386.180 2794.620 ;
        RECT 2391.380 2794.300 2391.700 2794.620 ;
        RECT 2395.060 2794.300 2395.380 2794.620 ;
        RECT 2404.260 2794.300 2404.580 2794.620 ;
        RECT 2418.060 2794.300 2418.380 2794.620 ;
        RECT 348.980 2793.620 349.300 2793.940 ;
        RECT 379.340 2793.620 379.660 2793.940 ;
        RECT 392.220 2793.620 392.540 2793.940 ;
        RECT 396.820 2793.620 397.140 2793.940 ;
        RECT 414.300 2793.620 414.620 2793.940 ;
        RECT 427.180 2793.620 427.500 2793.940 ;
        RECT 430.860 2793.620 431.180 2793.940 ;
        RECT 455.700 2793.620 456.020 2793.940 ;
        RECT 468.580 2793.620 468.900 2793.940 ;
        RECT 526.540 2793.620 526.860 2793.940 ;
        RECT 1012.300 2793.620 1012.620 2793.940 ;
        RECT 1083.140 2793.620 1083.460 2793.940 ;
        RECT 1164.100 2793.620 1164.420 2793.940 ;
        RECT 1167.780 2793.620 1168.100 2793.940 ;
        RECT 1173.300 2793.620 1173.620 2793.940 ;
        RECT 1180.660 2793.620 1180.980 2793.940 ;
        RECT 1601.100 2793.620 1601.420 2793.940 ;
        RECT 1774.060 2793.620 1774.380 2793.940 ;
        RECT 1780.500 2793.620 1780.820 2793.940 ;
        RECT 2269.020 2793.620 2269.340 2793.940 ;
        RECT 2332.500 2793.620 2332.820 2793.940 ;
        RECT 2345.380 2793.620 2345.700 2793.940 ;
        RECT 2349.980 2793.620 2350.300 2793.940 ;
        RECT 2356.420 2793.620 2356.740 2793.940 ;
        RECT 2361.020 2793.620 2361.340 2793.940 ;
        RECT 2402.420 2793.620 2402.740 2793.940 ;
        RECT 2407.940 2793.620 2408.260 2793.940 ;
        RECT 431.780 2792.940 432.100 2793.260 ;
        RECT 467.660 2792.940 467.980 2793.260 ;
        RECT 1024.260 2792.940 1024.580 2793.260 ;
        RECT 1052.780 2792.940 1053.100 2793.260 ;
        RECT 1087.740 2792.940 1088.060 2793.260 ;
        RECT 1159.500 2792.940 1159.820 2793.260 ;
        RECT 1187.100 2792.940 1187.420 2793.260 ;
        RECT 1594.660 2792.940 1594.980 2793.260 ;
        RECT 2263.500 2792.940 2263.820 2793.260 ;
        RECT 2297.540 2792.940 2297.860 2793.260 ;
        RECT 2338.940 2792.940 2339.260 2793.260 ;
        RECT 2367.460 2792.940 2367.780 2793.260 ;
        RECT 2423.580 2792.940 2423.900 2793.260 ;
        RECT 2442.900 2792.940 2443.220 2793.260 ;
        RECT 497.100 2792.260 497.420 2792.580 ;
        RECT 543.100 2792.260 543.420 2792.580 ;
        RECT 1153.060 2792.260 1153.380 2792.580 ;
        RECT 1787.860 2792.260 1788.180 2792.580 ;
        RECT 2249.700 2792.260 2250.020 2792.580 ;
        RECT 2386.780 2792.260 2387.100 2792.580 ;
        RECT 2410.700 2792.260 2411.020 2792.580 ;
        RECT 2430.020 2792.260 2430.340 2792.580 ;
        RECT 2436.460 2792.260 2436.780 2792.580 ;
        RECT 986.540 2791.580 986.860 2791.900 ;
        RECT 1193.540 2791.580 1193.860 2791.900 ;
        RECT 2374.820 2791.580 2375.140 2791.900 ;
        RECT 2381.260 2791.580 2381.580 2791.900 ;
        RECT 2392.300 2791.580 2392.620 2791.900 ;
        RECT 993.900 2790.900 994.220 2791.220 ;
        RECT 2242.340 2790.900 2242.660 2791.220 ;
        RECT 2398.740 2790.900 2399.060 2791.220 ;
        RECT 2417.140 2790.900 2417.460 2791.220 ;
        RECT 2428.180 2790.900 2428.500 2791.220 ;
        RECT 2434.620 2790.900 2434.940 2791.220 ;
        RECT 1191.700 2790.220 1192.020 2790.540 ;
        RECT 2257.060 2790.220 2257.380 2790.540 ;
        RECT 2420.820 2790.220 2421.140 2790.540 ;
        RECT 2445.660 2790.220 2445.980 2790.540 ;
        RECT 2439.220 2789.540 2439.540 2789.860 ;
        RECT 501.700 2788.860 502.020 2789.180 ;
        RECT 508.140 2788.180 508.460 2788.500 ;
        RECT 531.140 2788.180 531.460 2788.500 ;
        RECT 1035.300 2788.180 1035.620 2788.500 ;
        RECT 1048.180 2788.180 1048.500 2788.500 ;
        RECT 1051.860 2788.180 1052.180 2788.500 ;
        RECT 1086.820 2788.180 1087.140 2788.500 ;
        RECT 1128.220 2788.180 1128.540 2788.500 ;
        RECT 1163.180 2788.180 1163.500 2788.500 ;
        RECT 1624.100 2788.180 1624.420 2788.500 ;
        RECT 1630.540 2788.180 1630.860 2788.500 ;
        RECT 1635.140 2788.180 1635.460 2788.500 ;
        RECT 1655.380 2788.180 1655.700 2788.500 ;
        RECT 1689.420 2788.180 1689.740 2788.500 ;
        RECT 1724.380 2788.180 1724.700 2788.500 ;
        RECT 1765.780 2788.180 1766.100 2788.500 ;
        RECT 2310.420 2788.180 2310.740 2788.500 ;
        RECT 2415.300 2788.180 2415.620 2788.500 ;
        RECT 507.220 2787.500 507.540 2787.820 ;
        RECT 513.660 2787.500 513.980 2787.820 ;
        RECT 516.420 2787.500 516.740 2787.820 ;
        RECT 520.100 2787.500 520.420 2787.820 ;
        RECT 526.540 2787.500 526.860 2787.820 ;
        RECT 530.220 2787.500 530.540 2787.820 ;
        RECT 538.500 2787.500 538.820 2787.820 ;
        RECT 544.940 2787.500 545.260 2787.820 ;
        RECT 1034.380 2787.500 1034.700 2787.820 ;
        RECT 1039.900 2787.500 1040.220 2787.820 ;
        RECT 1046.340 2787.500 1046.660 2787.820 ;
        RECT 1054.620 2787.500 1054.940 2787.820 ;
        RECT 1061.980 2787.500 1062.300 2787.820 ;
        RECT 1067.500 2787.500 1067.820 2787.820 ;
        RECT 1073.940 2787.500 1074.260 2787.820 ;
        RECT 1081.300 2787.500 1081.620 2787.820 ;
        RECT 1089.580 2787.500 1089.900 2787.820 ;
        RECT 1096.020 2787.500 1096.340 2787.820 ;
        RECT 1103.380 2787.500 1103.700 2787.820 ;
        RECT 1109.820 2787.500 1110.140 2787.820 ;
        RECT 1116.260 2787.500 1116.580 2787.820 ;
        RECT 1121.780 2787.500 1122.100 2787.820 ;
        RECT 1130.980 2787.500 1131.300 2787.820 ;
        RECT 1137.420 2787.500 1137.740 2787.820 ;
        RECT 1143.860 2787.500 1144.180 2787.820 ;
        RECT 1151.220 2787.500 1151.540 2787.820 ;
        RECT 1153.980 2787.500 1154.300 2787.820 ;
        RECT 1165.020 2787.500 1165.340 2787.820 ;
        RECT 1172.380 2787.500 1172.700 2787.820 ;
        RECT 1613.980 2787.500 1614.300 2787.820 ;
        RECT 1620.420 2787.500 1620.740 2787.820 ;
        RECT 1626.860 2787.500 1627.180 2787.820 ;
        RECT 1631.460 2787.500 1631.780 2787.820 ;
        RECT 1637.900 2787.500 1638.220 2787.820 ;
        RECT 1644.340 2787.500 1644.660 2787.820 ;
        RECT 1648.940 2787.500 1649.260 2787.820 ;
        RECT 1661.820 2787.500 1662.140 2787.820 ;
        RECT 1666.420 2787.500 1666.740 2787.820 ;
        RECT 1672.860 2787.500 1673.180 2787.820 ;
        RECT 1679.300 2787.500 1679.620 2787.820 ;
        RECT 1683.900 2787.500 1684.220 2787.820 ;
        RECT 1695.860 2787.500 1696.180 2787.820 ;
        RECT 1702.300 2787.500 1702.620 2787.820 ;
        RECT 1708.740 2787.500 1709.060 2787.820 ;
        RECT 1713.340 2787.500 1713.660 2787.820 ;
        RECT 1719.780 2787.500 1720.100 2787.820 ;
        RECT 1730.820 2787.500 1731.140 2787.820 ;
        RECT 1737.260 2787.500 1737.580 2787.820 ;
        RECT 1743.700 2787.500 1744.020 2787.820 ;
        RECT 1748.300 2787.500 1748.620 2787.820 ;
        RECT 1754.740 2787.500 1755.060 2787.820 ;
        RECT 1772.220 2787.500 1772.540 2787.820 ;
        RECT 1778.660 2787.500 1778.980 2787.820 ;
        RECT 1783.260 2787.500 1783.580 2787.820 ;
        RECT 1789.700 2787.500 1790.020 2787.820 ;
        RECT 2264.420 2787.500 2264.740 2787.820 ;
        RECT 2276.380 2787.500 2276.700 2787.820 ;
        RECT 2282.820 2787.500 2283.140 2787.820 ;
        RECT 2287.420 2787.500 2287.740 2787.820 ;
        RECT 2293.860 2787.500 2294.180 2787.820 ;
        RECT 2300.300 2787.500 2300.620 2787.820 ;
        RECT 2304.900 2787.500 2305.220 2787.820 ;
        RECT 2317.780 2787.500 2318.100 2787.820 ;
        RECT 2322.380 2787.500 2322.700 2787.820 ;
        RECT 2328.820 2787.500 2329.140 2787.820 ;
        RECT 1761.180 2777.300 1761.500 2777.620 ;
        RECT 1796.140 2777.300 1796.460 2777.620 ;
        RECT 1411.580 1614.500 1411.900 1614.820 ;
      LAYER met4 ;
        RECT 646.135 3264.175 646.465 3264.505 ;
        RECT 668.215 3264.175 668.545 3264.505 ;
        RECT 1295.655 3264.175 1295.985 3264.505 ;
        RECT 1317.735 3264.175 1318.065 3264.505 ;
        RECT 1890.895 3264.175 1891.225 3264.505 ;
        RECT 1917.575 3264.175 1917.905 3264.505 ;
        RECT 2542.255 3264.175 2542.585 3264.505 ;
        RECT 2567.095 3264.175 2567.425 3264.505 ;
        RECT 394.025 3251.635 394.325 3256.235 ;
        RECT 400.265 3251.635 400.565 3256.235 ;
        RECT 406.505 3251.635 406.805 3256.235 ;
        RECT 412.745 3251.635 413.045 3256.235 ;
        RECT 418.985 3251.635 419.285 3256.235 ;
        RECT 425.225 3251.635 425.525 3256.235 ;
        RECT 431.465 3251.635 431.765 3256.235 ;
        RECT 437.705 3251.635 438.005 3256.235 ;
        RECT 443.945 3251.635 444.245 3256.235 ;
        RECT 450.185 3251.635 450.485 3256.235 ;
        RECT 456.425 3251.635 456.725 3256.235 ;
        RECT 462.665 3251.635 462.965 3256.235 ;
        RECT 468.905 3251.635 469.205 3256.235 ;
        RECT 475.145 3251.635 475.445 3256.235 ;
        RECT 481.385 3251.635 481.685 3256.235 ;
        RECT 487.625 3251.635 487.925 3256.235 ;
        RECT 493.865 3251.635 494.165 3256.235 ;
        RECT 500.105 3251.635 500.405 3256.235 ;
        RECT 506.345 3251.635 506.645 3256.235 ;
        RECT 512.585 3251.635 512.885 3256.235 ;
        RECT 518.825 3251.635 519.125 3256.235 ;
        RECT 525.065 3251.635 525.365 3256.235 ;
        RECT 531.305 3251.635 531.605 3256.235 ;
        RECT 537.545 3251.635 537.845 3256.235 ;
        RECT 543.785 3251.635 544.085 3256.235 ;
        RECT 550.025 3251.635 550.325 3256.235 ;
        RECT 556.265 3251.635 556.565 3256.235 ;
        RECT 562.505 3251.635 562.805 3256.235 ;
        RECT 568.745 3251.635 569.045 3256.235 ;
        RECT 574.985 3251.635 575.285 3256.235 ;
        RECT 581.225 3251.635 581.525 3256.235 ;
        RECT 587.465 3251.635 587.765 3256.235 ;
        RECT 642.890 3255.650 643.190 3256.235 ;
        RECT 646.150 3255.650 646.450 3264.175 ;
        RECT 668.230 3259.050 668.530 3264.175 ;
        RECT 642.890 3255.350 646.450 3255.650 ;
        RECT 667.865 3258.750 668.530 3259.050 ;
        RECT 642.890 3251.635 643.190 3255.350 ;
        RECT 667.865 3251.635 668.165 3258.750 ;
        RECT 1044.025 3251.635 1044.325 3256.235 ;
        RECT 1050.265 3251.635 1050.565 3256.235 ;
        RECT 1056.505 3251.635 1056.805 3256.235 ;
        RECT 1062.745 3251.635 1063.045 3256.235 ;
        RECT 1068.985 3251.635 1069.285 3256.235 ;
        RECT 1075.225 3251.635 1075.525 3256.235 ;
        RECT 1081.465 3251.635 1081.765 3256.235 ;
        RECT 1087.705 3251.635 1088.005 3256.235 ;
        RECT 1093.945 3251.635 1094.245 3256.235 ;
        RECT 1100.185 3251.635 1100.485 3256.235 ;
        RECT 1106.425 3251.635 1106.725 3256.235 ;
        RECT 1112.665 3251.635 1112.965 3256.235 ;
        RECT 1118.905 3251.635 1119.205 3256.235 ;
        RECT 1125.145 3251.635 1125.445 3256.235 ;
        RECT 1131.385 3251.635 1131.685 3256.235 ;
        RECT 1137.625 3251.635 1137.925 3256.235 ;
        RECT 1143.865 3251.635 1144.165 3256.235 ;
        RECT 1150.105 3251.635 1150.405 3256.235 ;
        RECT 1156.345 3251.635 1156.645 3256.235 ;
        RECT 1162.585 3251.635 1162.885 3256.235 ;
        RECT 1168.825 3251.635 1169.125 3256.235 ;
        RECT 1175.065 3251.635 1175.365 3256.235 ;
        RECT 1181.305 3251.635 1181.605 3256.235 ;
        RECT 1187.545 3251.635 1187.845 3256.235 ;
        RECT 1193.785 3251.635 1194.085 3256.235 ;
        RECT 1200.025 3251.635 1200.325 3256.235 ;
        RECT 1206.265 3251.635 1206.565 3256.235 ;
        RECT 1212.505 3251.635 1212.805 3256.235 ;
        RECT 1218.745 3251.635 1219.045 3256.235 ;
        RECT 1224.985 3251.635 1225.285 3256.235 ;
        RECT 1231.225 3251.635 1231.525 3256.235 ;
        RECT 1237.465 3251.635 1237.765 3256.235 ;
        RECT 1292.890 3255.650 1293.190 3256.235 ;
        RECT 1295.670 3255.650 1295.970 3264.175 ;
        RECT 1292.890 3255.350 1295.970 3255.650 ;
        RECT 1317.750 3256.235 1318.050 3264.175 ;
        RECT 1317.750 3255.350 1318.165 3256.235 ;
        RECT 1292.890 3251.635 1293.190 3255.350 ;
        RECT 1317.865 3251.635 1318.165 3255.350 ;
        RECT 1644.025 3251.635 1644.325 3256.235 ;
        RECT 1650.265 3251.635 1650.565 3256.235 ;
        RECT 1656.505 3251.635 1656.805 3256.235 ;
        RECT 1662.745 3251.635 1663.045 3256.235 ;
        RECT 1668.985 3251.635 1669.285 3256.235 ;
        RECT 1675.225 3251.635 1675.525 3256.235 ;
        RECT 1681.465 3251.635 1681.765 3256.235 ;
        RECT 1687.705 3251.635 1688.005 3256.235 ;
        RECT 1693.945 3251.635 1694.245 3256.235 ;
        RECT 1700.185 3251.635 1700.485 3256.235 ;
        RECT 1706.425 3251.635 1706.725 3256.235 ;
        RECT 1712.665 3251.635 1712.965 3256.235 ;
        RECT 1718.905 3251.635 1719.205 3256.235 ;
        RECT 1725.145 3251.635 1725.445 3256.235 ;
        RECT 1731.385 3251.635 1731.685 3256.235 ;
        RECT 1737.625 3251.635 1737.925 3256.235 ;
        RECT 1743.865 3251.635 1744.165 3256.235 ;
        RECT 1750.105 3251.635 1750.405 3256.235 ;
        RECT 1756.345 3251.635 1756.645 3256.235 ;
        RECT 1762.585 3251.635 1762.885 3256.235 ;
        RECT 1768.825 3251.635 1769.125 3256.235 ;
        RECT 1775.065 3251.635 1775.365 3256.235 ;
        RECT 1781.305 3251.635 1781.605 3256.235 ;
        RECT 1787.545 3251.635 1787.845 3256.235 ;
        RECT 1793.785 3251.635 1794.085 3256.235 ;
        RECT 1800.025 3251.635 1800.325 3256.235 ;
        RECT 1806.265 3251.635 1806.565 3256.235 ;
        RECT 1812.505 3251.635 1812.805 3256.235 ;
        RECT 1818.745 3251.635 1819.045 3256.235 ;
        RECT 1824.985 3251.635 1825.285 3256.235 ;
        RECT 1831.225 3251.635 1831.525 3256.235 ;
        RECT 1837.465 3251.635 1837.765 3256.235 ;
        RECT 1890.910 3255.650 1891.210 3264.175 ;
        RECT 1917.590 3256.235 1917.890 3264.175 ;
        RECT 1892.890 3255.650 1893.190 3256.235 ;
        RECT 1890.910 3255.350 1893.190 3255.650 ;
        RECT 1917.590 3255.350 1918.165 3256.235 ;
        RECT 1892.890 3251.635 1893.190 3255.350 ;
        RECT 1917.865 3251.635 1918.165 3255.350 ;
        RECT 2294.025 3251.635 2294.325 3256.235 ;
        RECT 2300.265 3251.635 2300.565 3256.235 ;
        RECT 2306.505 3251.635 2306.805 3256.235 ;
        RECT 2312.745 3251.635 2313.045 3256.235 ;
        RECT 2318.985 3251.635 2319.285 3256.235 ;
        RECT 2325.225 3251.635 2325.525 3256.235 ;
        RECT 2331.465 3251.635 2331.765 3256.235 ;
        RECT 2337.705 3251.635 2338.005 3256.235 ;
        RECT 2343.945 3251.635 2344.245 3256.235 ;
        RECT 2350.185 3251.635 2350.485 3256.235 ;
        RECT 2356.425 3251.635 2356.725 3256.235 ;
        RECT 2362.665 3251.635 2362.965 3256.235 ;
        RECT 2368.905 3251.635 2369.205 3256.235 ;
        RECT 2375.145 3251.635 2375.445 3256.235 ;
        RECT 2381.385 3251.635 2381.685 3256.235 ;
        RECT 2387.625 3251.635 2387.925 3256.235 ;
        RECT 2393.865 3251.635 2394.165 3256.235 ;
        RECT 2400.105 3251.635 2400.405 3256.235 ;
        RECT 2406.345 3251.635 2406.645 3256.235 ;
        RECT 2412.585 3251.635 2412.885 3256.235 ;
        RECT 2418.825 3251.635 2419.125 3256.235 ;
        RECT 2425.065 3251.635 2425.365 3256.235 ;
        RECT 2431.305 3251.635 2431.605 3256.235 ;
        RECT 2437.545 3251.635 2437.845 3256.235 ;
        RECT 2443.785 3251.635 2444.085 3256.235 ;
        RECT 2450.025 3251.635 2450.325 3256.235 ;
        RECT 2456.265 3251.635 2456.565 3256.235 ;
        RECT 2462.505 3251.635 2462.805 3256.235 ;
        RECT 2468.745 3251.635 2469.045 3256.235 ;
        RECT 2474.985 3251.635 2475.285 3256.235 ;
        RECT 2481.225 3251.635 2481.525 3256.235 ;
        RECT 2487.465 3251.635 2487.765 3256.235 ;
        RECT 2542.270 3255.650 2542.570 3264.175 ;
        RECT 2542.890 3255.650 2543.190 3256.235 ;
        RECT 2542.270 3255.350 2543.190 3255.650 ;
        RECT 2567.110 3255.650 2567.410 3264.175 ;
        RECT 2567.865 3255.650 2568.165 3256.235 ;
        RECT 2567.110 3255.350 2568.165 3255.650 ;
        RECT 2542.890 3251.635 2543.190 3255.350 ;
        RECT 2567.865 3251.635 2568.165 3255.350 ;
        RECT 302.550 2894.510 303.730 2895.690 ;
      LAYER met4 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met4 ;
        RECT 687.535 2901.735 687.865 2902.065 ;
        RECT 687.550 2895.690 687.850 2901.735 ;
        RECT 687.110 2894.510 688.290 2895.690 ;
        RECT 950.230 2894.510 951.410 2895.690 ;
      LAYER met4 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met4 ;
        RECT 1411.575 3243.095 1411.905 3243.425 ;
        RECT 1345.335 2904.455 1345.665 2904.785 ;
        RECT 1345.350 2895.690 1345.650 2904.455 ;
        RECT 1344.910 2894.510 1346.090 2895.690 ;
        RECT 334.010 2801.750 334.310 2804.600 ;
        RECT 339.850 2801.750 340.150 2804.600 ;
        RECT 345.690 2801.750 345.990 2804.600 ;
        RECT 351.530 2801.750 351.830 2804.600 ;
        RECT 334.010 2801.450 337.330 2801.750 ;
        RECT 334.010 2800.000 334.310 2801.450 ;
        RECT 337.030 2794.625 337.330 2801.450 ;
        RECT 339.850 2801.450 342.850 2801.750 ;
        RECT 339.850 2800.000 340.150 2801.450 ;
        RECT 342.550 2794.625 342.850 2801.450 ;
        RECT 345.690 2801.450 349.290 2801.750 ;
        RECT 345.690 2800.000 345.990 2801.450 ;
        RECT 337.015 2794.295 337.345 2794.625 ;
        RECT 342.535 2794.295 342.865 2794.625 ;
        RECT 348.990 2793.945 349.290 2801.450 ;
        RECT 350.830 2801.450 351.830 2801.750 ;
        RECT 350.830 2794.625 351.130 2801.450 ;
        RECT 351.530 2800.000 351.830 2801.450 ;
        RECT 357.370 2801.750 357.670 2804.600 ;
        RECT 363.210 2802.450 363.510 2804.600 ;
        RECT 361.870 2802.150 363.510 2802.450 ;
        RECT 357.370 2801.450 358.490 2801.750 ;
        RECT 357.370 2800.000 357.670 2801.450 ;
        RECT 358.190 2794.625 358.490 2801.450 ;
        RECT 361.870 2794.625 362.170 2802.150 ;
        RECT 363.210 2800.000 363.510 2802.150 ;
        RECT 363.830 2801.750 364.130 2804.600 ;
        RECT 369.050 2801.750 369.350 2804.600 ;
        RECT 363.830 2801.450 364.930 2801.750 ;
        RECT 363.830 2800.000 364.130 2801.450 ;
        RECT 364.630 2794.625 364.930 2801.450 ;
        RECT 368.310 2801.450 369.350 2801.750 ;
        RECT 368.310 2794.625 368.610 2801.450 ;
        RECT 369.050 2800.000 369.350 2801.450 ;
        RECT 369.670 2801.750 369.970 2804.600 ;
        RECT 374.890 2801.750 375.190 2804.600 ;
        RECT 369.670 2801.450 371.370 2801.750 ;
        RECT 369.670 2800.000 369.970 2801.450 ;
        RECT 371.070 2794.625 371.370 2801.450 ;
        RECT 374.750 2800.000 375.190 2801.750 ;
        RECT 375.510 2801.750 375.810 2804.600 ;
        RECT 380.730 2801.750 381.030 2804.600 ;
        RECT 375.510 2801.450 378.730 2801.750 ;
        RECT 375.510 2800.000 375.810 2801.450 ;
        RECT 374.750 2794.625 375.050 2800.000 ;
        RECT 378.430 2794.625 378.730 2801.450 ;
        RECT 379.350 2801.450 381.030 2801.750 ;
        RECT 350.815 2794.295 351.145 2794.625 ;
        RECT 358.175 2794.295 358.505 2794.625 ;
        RECT 361.855 2794.295 362.185 2794.625 ;
        RECT 364.615 2794.295 364.945 2794.625 ;
        RECT 368.295 2794.295 368.625 2794.625 ;
        RECT 371.055 2794.295 371.385 2794.625 ;
        RECT 374.735 2794.295 375.065 2794.625 ;
        RECT 378.415 2794.295 378.745 2794.625 ;
        RECT 379.350 2793.945 379.650 2801.450 ;
        RECT 380.730 2800.000 381.030 2801.450 ;
        RECT 381.350 2801.750 381.650 2804.600 ;
        RECT 381.350 2801.450 384.250 2801.750 ;
        RECT 381.350 2800.000 381.650 2801.450 ;
        RECT 383.950 2794.625 384.250 2801.450 ;
        RECT 386.570 2796.650 386.870 2804.600 ;
        RECT 387.190 2801.750 387.490 2804.600 ;
        RECT 392.410 2801.750 392.710 2804.600 ;
        RECT 387.190 2801.450 390.690 2801.750 ;
        RECT 387.190 2800.000 387.490 2801.450 ;
        RECT 386.570 2796.350 387.010 2796.650 ;
        RECT 386.710 2794.625 387.010 2796.350 ;
        RECT 390.390 2794.625 390.690 2801.450 ;
        RECT 392.230 2800.000 392.710 2801.750 ;
        RECT 393.030 2801.750 393.330 2804.600 ;
        RECT 398.250 2802.450 398.550 2804.600 ;
        RECT 396.830 2802.150 398.550 2802.450 ;
        RECT 393.030 2801.450 396.210 2801.750 ;
        RECT 393.030 2800.000 393.330 2801.450 ;
        RECT 383.935 2794.295 384.265 2794.625 ;
        RECT 386.695 2794.295 387.025 2794.625 ;
        RECT 390.375 2794.295 390.705 2794.625 ;
        RECT 392.230 2793.945 392.530 2800.000 ;
        RECT 395.910 2794.625 396.210 2801.450 ;
        RECT 395.895 2794.295 396.225 2794.625 ;
        RECT 396.830 2793.945 397.130 2802.150 ;
        RECT 398.250 2800.000 398.550 2802.150 ;
        RECT 398.870 2801.750 399.170 2804.600 ;
        RECT 404.090 2801.750 404.390 2804.600 ;
        RECT 398.870 2801.450 399.890 2801.750 ;
        RECT 398.870 2800.000 399.170 2801.450 ;
        RECT 399.590 2794.625 399.890 2801.450 ;
        RECT 403.270 2801.450 404.390 2801.750 ;
        RECT 403.270 2794.625 403.570 2801.450 ;
        RECT 404.090 2800.000 404.390 2801.450 ;
        RECT 404.710 2801.750 405.010 2804.600 ;
        RECT 409.930 2801.750 410.230 2804.600 ;
        RECT 404.710 2801.450 406.330 2801.750 ;
        RECT 404.710 2800.000 405.010 2801.450 ;
        RECT 406.030 2794.625 406.330 2801.450 ;
        RECT 409.710 2800.000 410.230 2801.750 ;
        RECT 410.550 2801.750 410.850 2804.600 ;
        RECT 415.770 2802.450 416.070 2804.600 ;
        RECT 414.310 2802.150 416.070 2802.450 ;
        RECT 410.550 2801.450 413.690 2801.750 ;
        RECT 410.550 2800.000 410.850 2801.450 ;
        RECT 409.710 2794.625 410.010 2800.000 ;
        RECT 413.390 2794.625 413.690 2801.450 ;
        RECT 399.575 2794.295 399.905 2794.625 ;
        RECT 403.255 2794.295 403.585 2794.625 ;
        RECT 406.015 2794.295 406.345 2794.625 ;
        RECT 409.695 2794.295 410.025 2794.625 ;
        RECT 413.375 2794.295 413.705 2794.625 ;
        RECT 414.310 2793.945 414.610 2802.150 ;
        RECT 415.770 2800.000 416.070 2802.150 ;
        RECT 416.390 2801.750 416.690 2804.600 ;
        RECT 421.610 2801.750 421.910 2804.600 ;
        RECT 416.390 2801.450 419.210 2801.750 ;
        RECT 416.390 2800.000 416.690 2801.450 ;
        RECT 418.910 2794.625 419.210 2801.450 ;
        RECT 420.750 2801.450 421.910 2801.750 ;
        RECT 420.750 2794.625 421.050 2801.450 ;
        RECT 421.610 2800.000 421.910 2801.450 ;
        RECT 422.230 2801.750 422.530 2804.600 ;
        RECT 427.450 2801.750 427.750 2804.600 ;
        RECT 422.230 2801.450 425.650 2801.750 ;
        RECT 422.230 2800.000 422.530 2801.450 ;
        RECT 425.350 2794.625 425.650 2801.450 ;
        RECT 427.190 2800.000 427.750 2801.750 ;
        RECT 428.070 2801.750 428.370 2804.600 ;
        RECT 433.290 2802.450 433.590 2804.600 ;
        RECT 431.790 2802.150 433.590 2802.450 ;
        RECT 428.070 2801.450 431.170 2801.750 ;
        RECT 428.070 2800.000 428.370 2801.450 ;
        RECT 418.895 2794.295 419.225 2794.625 ;
        RECT 420.735 2794.295 421.065 2794.625 ;
        RECT 425.335 2794.295 425.665 2794.625 ;
        RECT 427.190 2793.945 427.490 2800.000 ;
        RECT 430.870 2793.945 431.170 2801.450 ;
        RECT 348.975 2793.615 349.305 2793.945 ;
        RECT 379.335 2793.615 379.665 2793.945 ;
        RECT 392.215 2793.615 392.545 2793.945 ;
        RECT 396.815 2793.615 397.145 2793.945 ;
        RECT 414.295 2793.615 414.625 2793.945 ;
        RECT 427.175 2793.615 427.505 2793.945 ;
        RECT 430.855 2793.615 431.185 2793.945 ;
        RECT 431.790 2793.265 432.090 2802.150 ;
        RECT 433.290 2800.000 433.590 2802.150 ;
        RECT 433.910 2796.650 434.210 2804.600 ;
        RECT 439.130 2800.050 439.430 2804.600 ;
        RECT 439.750 2801.750 440.050 2804.600 ;
        RECT 444.970 2801.750 445.270 2804.600 ;
        RECT 439.750 2801.450 441.290 2801.750 ;
        RECT 439.130 2799.750 439.450 2800.050 ;
        RECT 439.750 2800.000 440.050 2801.450 ;
        RECT 433.630 2796.350 434.210 2796.650 ;
        RECT 433.630 2794.625 433.930 2796.350 ;
        RECT 439.150 2794.625 439.450 2799.750 ;
        RECT 440.990 2794.625 441.290 2801.450 ;
        RECT 444.670 2800.000 445.270 2801.750 ;
        RECT 444.670 2794.625 444.970 2800.000 ;
        RECT 445.590 2794.625 445.890 2804.600 ;
        RECT 450.810 2801.750 451.110 2804.600 ;
        RECT 449.270 2801.450 451.110 2801.750 ;
        RECT 449.270 2794.625 449.570 2801.450 ;
        RECT 450.810 2800.000 451.110 2801.450 ;
        RECT 451.430 2801.750 451.730 2804.600 ;
        RECT 456.650 2801.750 456.950 2804.600 ;
        RECT 451.430 2801.450 455.090 2801.750 ;
        RECT 451.430 2800.000 451.730 2801.450 ;
        RECT 454.790 2794.625 455.090 2801.450 ;
        RECT 455.710 2801.450 456.950 2801.750 ;
        RECT 433.615 2794.295 433.945 2794.625 ;
        RECT 439.135 2794.295 439.465 2794.625 ;
        RECT 440.975 2794.295 441.305 2794.625 ;
        RECT 444.655 2794.295 444.985 2794.625 ;
        RECT 445.575 2794.295 445.905 2794.625 ;
        RECT 449.255 2794.295 449.585 2794.625 ;
        RECT 454.775 2794.295 455.105 2794.625 ;
        RECT 455.710 2793.945 456.010 2801.450 ;
        RECT 456.650 2800.000 456.950 2801.450 ;
        RECT 457.270 2801.750 457.570 2804.600 ;
        RECT 457.270 2801.450 460.610 2801.750 ;
        RECT 457.270 2800.000 457.570 2801.450 ;
        RECT 460.310 2794.625 460.610 2801.450 ;
        RECT 462.490 2800.050 462.790 2804.600 ;
        RECT 462.150 2799.750 462.790 2800.050 ;
        RECT 463.110 2801.750 463.410 2804.600 ;
        RECT 468.330 2801.750 468.630 2804.600 ;
        RECT 463.110 2801.450 466.130 2801.750 ;
        RECT 463.110 2800.000 463.410 2801.450 ;
        RECT 462.150 2794.625 462.450 2799.750 ;
        RECT 465.830 2794.625 466.130 2801.450 ;
        RECT 467.670 2801.450 468.630 2801.750 ;
        RECT 460.295 2794.295 460.625 2794.625 ;
        RECT 462.135 2794.295 462.465 2794.625 ;
        RECT 465.815 2794.295 466.145 2794.625 ;
        RECT 455.695 2793.615 456.025 2793.945 ;
        RECT 467.670 2793.265 467.970 2801.450 ;
        RECT 468.330 2800.000 468.630 2801.450 ;
        RECT 468.950 2796.650 469.250 2804.600 ;
        RECT 474.170 2801.750 474.470 2804.600 ;
        RECT 468.590 2796.350 469.250 2796.650 ;
        RECT 474.110 2800.000 474.470 2801.750 ;
        RECT 474.790 2801.750 475.090 2804.600 ;
        RECT 480.010 2801.750 480.310 2804.600 ;
        RECT 474.790 2800.000 475.330 2801.750 ;
        RECT 468.590 2793.945 468.890 2796.350 ;
        RECT 474.110 2794.625 474.410 2800.000 ;
        RECT 475.030 2794.625 475.330 2800.000 ;
        RECT 478.710 2801.450 480.310 2801.750 ;
        RECT 478.710 2794.625 479.010 2801.450 ;
        RECT 480.010 2800.000 480.310 2801.450 ;
        RECT 480.630 2801.750 480.930 2804.600 ;
        RECT 485.850 2801.750 486.150 2804.600 ;
        RECT 480.630 2801.450 482.690 2801.750 ;
        RECT 480.630 2800.000 480.930 2801.450 ;
        RECT 482.390 2794.625 482.690 2801.450 ;
        RECT 485.150 2801.450 486.150 2801.750 ;
        RECT 485.150 2794.625 485.450 2801.450 ;
        RECT 485.850 2800.000 486.150 2801.450 ;
        RECT 486.470 2801.750 486.770 2804.600 ;
        RECT 491.690 2801.750 491.990 2804.600 ;
        RECT 486.470 2801.450 488.210 2801.750 ;
        RECT 486.470 2800.000 486.770 2801.450 ;
        RECT 487.910 2794.625 488.210 2801.450 ;
        RECT 491.590 2800.000 491.990 2801.750 ;
        RECT 492.310 2801.750 492.610 2804.600 ;
        RECT 492.310 2801.450 495.570 2801.750 ;
        RECT 492.310 2800.000 492.610 2801.450 ;
        RECT 491.590 2794.625 491.890 2800.000 ;
        RECT 495.270 2794.625 495.570 2801.450 ;
        RECT 497.530 2800.050 497.830 2804.600 ;
        RECT 497.110 2799.750 497.830 2800.050 ;
        RECT 498.150 2801.750 498.450 2804.600 ;
        RECT 503.370 2801.750 503.670 2804.600 ;
        RECT 498.150 2801.450 501.090 2801.750 ;
        RECT 498.150 2800.000 498.450 2801.450 ;
        RECT 474.095 2794.295 474.425 2794.625 ;
        RECT 475.015 2794.295 475.345 2794.625 ;
        RECT 478.695 2794.295 479.025 2794.625 ;
        RECT 482.375 2794.295 482.705 2794.625 ;
        RECT 485.135 2794.295 485.465 2794.625 ;
        RECT 487.895 2794.295 488.225 2794.625 ;
        RECT 491.575 2794.295 491.905 2794.625 ;
        RECT 495.255 2794.295 495.585 2794.625 ;
        RECT 468.575 2793.615 468.905 2793.945 ;
        RECT 431.775 2792.935 432.105 2793.265 ;
        RECT 467.655 2792.935 467.985 2793.265 ;
        RECT 497.110 2792.585 497.410 2799.750 ;
        RECT 500.790 2794.625 501.090 2801.450 ;
        RECT 501.710 2801.450 503.670 2801.750 ;
        RECT 500.775 2794.295 501.105 2794.625 ;
        RECT 497.095 2792.255 497.425 2792.585 ;
        RECT 501.710 2789.185 502.010 2801.450 ;
        RECT 503.370 2800.000 503.670 2801.450 ;
        RECT 503.990 2801.750 504.290 2804.600 ;
        RECT 509.210 2801.750 509.510 2804.600 ;
        RECT 503.990 2801.450 507.530 2801.750 ;
        RECT 503.990 2800.000 504.290 2801.450 ;
        RECT 501.695 2788.855 502.025 2789.185 ;
        RECT 507.230 2787.825 507.530 2801.450 ;
        RECT 508.150 2801.450 509.510 2801.750 ;
        RECT 508.150 2788.505 508.450 2801.450 ;
        RECT 509.210 2800.000 509.510 2801.450 ;
        RECT 509.830 2801.750 510.130 2804.600 ;
        RECT 515.050 2802.450 515.350 2804.600 ;
        RECT 513.670 2802.150 515.350 2802.450 ;
        RECT 509.830 2800.000 510.290 2801.750 ;
        RECT 509.990 2794.625 510.290 2800.000 ;
        RECT 509.975 2794.295 510.305 2794.625 ;
        RECT 508.135 2788.175 508.465 2788.505 ;
        RECT 513.670 2787.825 513.970 2802.150 ;
        RECT 515.050 2800.000 515.350 2802.150 ;
        RECT 515.670 2801.750 515.970 2804.600 ;
        RECT 520.890 2801.750 521.190 2804.600 ;
        RECT 515.670 2801.450 516.730 2801.750 ;
        RECT 515.670 2800.000 515.970 2801.450 ;
        RECT 516.430 2787.825 516.730 2801.450 ;
        RECT 520.110 2801.450 521.190 2801.750 ;
        RECT 520.110 2787.825 520.410 2801.450 ;
        RECT 520.890 2800.000 521.190 2801.450 ;
        RECT 521.510 2801.750 521.810 2804.600 ;
        RECT 526.730 2801.750 527.030 2804.600 ;
        RECT 521.510 2801.450 524.090 2801.750 ;
        RECT 521.510 2800.000 521.810 2801.450 ;
        RECT 523.790 2794.625 524.090 2801.450 ;
        RECT 526.550 2800.000 527.030 2801.750 ;
        RECT 527.350 2801.750 527.650 2804.600 ;
        RECT 532.570 2802.450 532.870 2804.600 ;
        RECT 531.150 2802.150 532.870 2802.450 ;
        RECT 527.350 2801.450 530.530 2801.750 ;
        RECT 527.350 2800.000 527.650 2801.450 ;
        RECT 523.775 2794.295 524.105 2794.625 ;
        RECT 526.550 2793.945 526.850 2800.000 ;
        RECT 526.535 2793.615 526.865 2793.945 ;
        RECT 526.550 2787.825 526.850 2793.615 ;
        RECT 530.230 2787.825 530.530 2801.450 ;
        RECT 531.150 2788.505 531.450 2802.150 ;
        RECT 532.570 2800.000 532.870 2802.150 ;
        RECT 533.190 2801.750 533.490 2804.600 ;
        RECT 533.190 2801.450 536.050 2801.750 ;
        RECT 533.190 2800.000 533.490 2801.450 ;
        RECT 535.750 2794.625 536.050 2801.450 ;
        RECT 538.410 2796.650 538.710 2804.600 ;
        RECT 539.030 2801.750 539.330 2804.600 ;
        RECT 544.250 2801.750 544.550 2804.600 ;
        RECT 539.030 2801.450 542.490 2801.750 ;
        RECT 539.030 2800.000 539.330 2801.450 ;
        RECT 538.410 2796.350 538.810 2796.650 ;
        RECT 535.735 2794.295 536.065 2794.625 ;
        RECT 531.135 2788.175 531.465 2788.505 ;
        RECT 538.510 2787.825 538.810 2796.350 ;
        RECT 542.190 2794.625 542.490 2801.450 ;
        RECT 543.110 2801.450 544.550 2801.750 ;
        RECT 542.175 2794.295 542.505 2794.625 ;
        RECT 543.110 2792.585 543.410 2801.450 ;
        RECT 544.250 2800.000 544.550 2801.450 ;
        RECT 544.870 2801.750 545.170 2804.600 ;
        RECT 984.010 2801.750 984.310 2804.600 ;
        RECT 989.850 2801.750 990.150 2804.600 ;
        RECT 995.690 2801.750 995.990 2804.600 ;
        RECT 1001.530 2801.750 1001.830 2804.600 ;
        RECT 544.870 2800.000 545.250 2801.750 ;
        RECT 543.095 2792.255 543.425 2792.585 ;
        RECT 544.950 2787.825 545.250 2800.000 ;
        RECT 981.030 2801.450 984.310 2801.750 ;
        RECT 981.030 2794.625 981.330 2801.450 ;
        RECT 984.010 2800.000 984.310 2801.450 ;
        RECT 986.550 2801.450 990.150 2801.750 ;
        RECT 981.015 2794.295 981.345 2794.625 ;
        RECT 986.550 2791.905 986.850 2801.450 ;
        RECT 989.850 2800.000 990.150 2801.450 ;
        RECT 993.910 2801.450 995.990 2801.750 ;
        RECT 986.535 2791.575 986.865 2791.905 ;
        RECT 993.910 2791.225 994.210 2801.450 ;
        RECT 995.690 2800.000 995.990 2801.450 ;
        RECT 1001.270 2800.000 1001.830 2801.750 ;
        RECT 1007.370 2800.050 1007.670 2804.600 ;
        RECT 1013.210 2801.750 1013.510 2804.600 ;
        RECT 1012.310 2801.450 1013.510 2801.750 ;
        RECT 1001.270 2794.625 1001.570 2800.000 ;
        RECT 1007.370 2799.750 1008.010 2800.050 ;
        RECT 1007.710 2794.625 1008.010 2799.750 ;
        RECT 1001.255 2794.295 1001.585 2794.625 ;
        RECT 1007.695 2794.295 1008.025 2794.625 ;
        RECT 1012.310 2793.945 1012.610 2801.450 ;
        RECT 1013.210 2800.000 1013.510 2801.450 ;
        RECT 1013.830 2796.650 1014.130 2804.600 ;
        RECT 1019.050 2801.750 1019.350 2804.600 ;
        RECT 1013.230 2796.350 1014.130 2796.650 ;
        RECT 1018.750 2800.000 1019.350 2801.750 ;
        RECT 1013.230 2794.625 1013.530 2796.350 ;
        RECT 1018.750 2794.625 1019.050 2800.000 ;
        RECT 1019.670 2794.625 1019.970 2804.600 ;
        RECT 1024.890 2801.750 1025.190 2804.600 ;
        RECT 1024.270 2801.450 1025.190 2801.750 ;
        RECT 1013.215 2794.295 1013.545 2794.625 ;
        RECT 1018.735 2794.295 1019.065 2794.625 ;
        RECT 1019.655 2794.295 1019.985 2794.625 ;
        RECT 1012.295 2793.615 1012.625 2793.945 ;
        RECT 1024.270 2793.265 1024.570 2801.450 ;
        RECT 1024.890 2800.000 1025.190 2801.450 ;
        RECT 1025.510 2801.750 1025.810 2804.600 ;
        RECT 1030.730 2801.750 1031.030 2804.600 ;
        RECT 1025.510 2801.450 1027.330 2801.750 ;
        RECT 1025.510 2800.000 1025.810 2801.450 ;
        RECT 1027.030 2794.625 1027.330 2801.450 ;
        RECT 1030.710 2800.000 1031.030 2801.750 ;
        RECT 1031.350 2801.750 1031.650 2804.600 ;
        RECT 1036.570 2802.450 1036.870 2804.600 ;
        RECT 1035.310 2802.150 1036.870 2802.450 ;
        RECT 1031.350 2801.450 1034.690 2801.750 ;
        RECT 1031.350 2800.000 1031.650 2801.450 ;
        RECT 1030.710 2794.625 1031.010 2800.000 ;
        RECT 1027.015 2794.295 1027.345 2794.625 ;
        RECT 1030.695 2794.295 1031.025 2794.625 ;
        RECT 1024.255 2792.935 1024.585 2793.265 ;
        RECT 993.895 2790.895 994.225 2791.225 ;
        RECT 1034.390 2787.825 1034.690 2801.450 ;
        RECT 1035.310 2788.505 1035.610 2802.150 ;
        RECT 1036.570 2800.000 1036.870 2802.150 ;
        RECT 1037.190 2801.750 1037.490 2804.600 ;
        RECT 1042.410 2801.750 1042.710 2804.600 ;
        RECT 1037.190 2801.450 1040.210 2801.750 ;
        RECT 1037.190 2800.000 1037.490 2801.450 ;
        RECT 1035.295 2788.175 1035.625 2788.505 ;
        RECT 1039.910 2787.825 1040.210 2801.450 ;
        RECT 1041.750 2801.450 1042.710 2801.750 ;
        RECT 1041.750 2794.625 1042.050 2801.450 ;
        RECT 1042.410 2800.000 1042.710 2801.450 ;
        RECT 1043.030 2801.750 1043.330 2804.600 ;
        RECT 1048.250 2801.750 1048.550 2804.600 ;
        RECT 1043.030 2801.450 1046.650 2801.750 ;
        RECT 1043.030 2800.000 1043.330 2801.450 ;
        RECT 1041.735 2794.295 1042.065 2794.625 ;
        RECT 1046.350 2787.825 1046.650 2801.450 ;
        RECT 1048.190 2800.000 1048.550 2801.750 ;
        RECT 1048.870 2801.750 1049.170 2804.600 ;
        RECT 1054.090 2801.750 1054.390 2804.600 ;
        RECT 1048.870 2801.450 1052.170 2801.750 ;
        RECT 1048.870 2800.000 1049.170 2801.450 ;
        RECT 1048.190 2788.505 1048.490 2800.000 ;
        RECT 1051.870 2788.505 1052.170 2801.450 ;
        RECT 1052.790 2801.450 1054.390 2801.750 ;
        RECT 1052.790 2793.265 1053.090 2801.450 ;
        RECT 1054.090 2800.000 1054.390 2801.450 ;
        RECT 1054.710 2796.650 1055.010 2804.600 ;
        RECT 1059.930 2801.750 1060.230 2804.600 ;
        RECT 1054.630 2796.350 1055.010 2796.650 ;
        RECT 1059.230 2801.450 1060.230 2801.750 ;
        RECT 1052.775 2792.935 1053.105 2793.265 ;
        RECT 1048.175 2788.175 1048.505 2788.505 ;
        RECT 1051.855 2788.175 1052.185 2788.505 ;
        RECT 1054.630 2787.825 1054.930 2796.350 ;
        RECT 1059.230 2794.625 1059.530 2801.450 ;
        RECT 1059.930 2800.000 1060.230 2801.450 ;
        RECT 1060.550 2801.750 1060.850 2804.600 ;
        RECT 1065.770 2801.750 1066.070 2804.600 ;
        RECT 1060.550 2801.450 1062.290 2801.750 ;
        RECT 1060.550 2800.000 1060.850 2801.450 ;
        RECT 1059.215 2794.295 1059.545 2794.625 ;
        RECT 1061.990 2787.825 1062.290 2801.450 ;
        RECT 1065.670 2800.000 1066.070 2801.750 ;
        RECT 1066.390 2801.750 1066.690 2804.600 ;
        RECT 1071.610 2801.750 1071.910 2804.600 ;
        RECT 1066.390 2801.450 1067.810 2801.750 ;
        RECT 1066.390 2800.000 1066.690 2801.450 ;
        RECT 1065.670 2794.625 1065.970 2800.000 ;
        RECT 1065.655 2794.295 1065.985 2794.625 ;
        RECT 1067.510 2787.825 1067.810 2801.450 ;
        RECT 1070.270 2801.450 1071.910 2801.750 ;
        RECT 1070.270 2794.625 1070.570 2801.450 ;
        RECT 1071.610 2800.000 1071.910 2801.450 ;
        RECT 1072.230 2801.750 1072.530 2804.600 ;
        RECT 1077.450 2801.750 1077.750 2804.600 ;
        RECT 1072.230 2801.450 1074.250 2801.750 ;
        RECT 1072.230 2800.000 1072.530 2801.450 ;
        RECT 1070.255 2794.295 1070.585 2794.625 ;
        RECT 1073.950 2787.825 1074.250 2801.450 ;
        RECT 1076.710 2801.450 1077.750 2801.750 ;
        RECT 1076.710 2794.625 1077.010 2801.450 ;
        RECT 1077.450 2800.000 1077.750 2801.450 ;
        RECT 1078.070 2801.750 1078.370 2804.600 ;
        RECT 1083.290 2801.750 1083.590 2804.600 ;
        RECT 1078.070 2801.450 1081.610 2801.750 ;
        RECT 1078.070 2800.000 1078.370 2801.450 ;
        RECT 1076.695 2794.295 1077.025 2794.625 ;
        RECT 1081.310 2787.825 1081.610 2801.450 ;
        RECT 1083.150 2800.000 1083.590 2801.750 ;
        RECT 1083.910 2801.750 1084.210 2804.600 ;
        RECT 1089.130 2801.750 1089.430 2804.600 ;
        RECT 1083.910 2801.450 1087.130 2801.750 ;
        RECT 1083.910 2800.000 1084.210 2801.450 ;
        RECT 1083.150 2793.945 1083.450 2800.000 ;
        RECT 1083.135 2793.615 1083.465 2793.945 ;
        RECT 1086.830 2788.505 1087.130 2801.450 ;
        RECT 1087.750 2801.450 1089.430 2801.750 ;
        RECT 1087.750 2793.265 1088.050 2801.450 ;
        RECT 1089.130 2800.000 1089.430 2801.450 ;
        RECT 1089.750 2796.650 1090.050 2804.600 ;
        RECT 1094.970 2801.750 1095.270 2804.600 ;
        RECT 1089.590 2796.350 1090.050 2796.650 ;
        RECT 1094.190 2801.450 1095.270 2801.750 ;
        RECT 1087.735 2792.935 1088.065 2793.265 ;
        RECT 1086.815 2788.175 1087.145 2788.505 ;
        RECT 1089.590 2787.825 1089.890 2796.350 ;
        RECT 1094.190 2794.625 1094.490 2801.450 ;
        RECT 1094.970 2800.000 1095.270 2801.450 ;
        RECT 1095.590 2800.050 1095.890 2804.600 ;
        RECT 1100.810 2801.750 1101.110 2804.600 ;
        RECT 1095.590 2799.750 1096.330 2800.050 ;
        RECT 1094.175 2794.295 1094.505 2794.625 ;
        RECT 1096.030 2787.825 1096.330 2799.750 ;
        RECT 1100.630 2800.000 1101.110 2801.750 ;
        RECT 1101.430 2801.750 1101.730 2804.600 ;
        RECT 1106.650 2802.450 1106.950 2804.600 ;
        RECT 1105.230 2802.150 1106.950 2802.450 ;
        RECT 1101.430 2801.450 1103.690 2801.750 ;
        RECT 1101.430 2800.000 1101.730 2801.450 ;
        RECT 1100.630 2794.625 1100.930 2800.000 ;
        RECT 1100.615 2794.295 1100.945 2794.625 ;
        RECT 1103.390 2787.825 1103.690 2801.450 ;
        RECT 1105.230 2794.625 1105.530 2802.150 ;
        RECT 1106.650 2800.000 1106.950 2802.150 ;
        RECT 1107.270 2801.750 1107.570 2804.600 ;
        RECT 1112.490 2801.750 1112.790 2804.600 ;
        RECT 1107.270 2801.450 1110.130 2801.750 ;
        RECT 1107.270 2800.000 1107.570 2801.450 ;
        RECT 1105.215 2794.295 1105.545 2794.625 ;
        RECT 1109.830 2787.825 1110.130 2801.450 ;
        RECT 1111.670 2801.450 1112.790 2801.750 ;
        RECT 1111.670 2794.625 1111.970 2801.450 ;
        RECT 1112.490 2800.000 1112.790 2801.450 ;
        RECT 1113.110 2801.750 1113.410 2804.600 ;
        RECT 1118.330 2801.750 1118.630 2804.600 ;
        RECT 1113.110 2801.450 1116.570 2801.750 ;
        RECT 1113.110 2800.000 1113.410 2801.450 ;
        RECT 1111.655 2794.295 1111.985 2794.625 ;
        RECT 1116.270 2787.825 1116.570 2801.450 ;
        RECT 1118.110 2800.000 1118.630 2801.750 ;
        RECT 1118.950 2801.750 1119.250 2804.600 ;
        RECT 1124.170 2801.750 1124.470 2804.600 ;
        RECT 1118.950 2801.450 1122.090 2801.750 ;
        RECT 1118.950 2800.000 1119.250 2801.450 ;
        RECT 1118.110 2794.625 1118.410 2800.000 ;
        RECT 1118.095 2794.295 1118.425 2794.625 ;
        RECT 1121.790 2787.825 1122.090 2801.450 ;
        RECT 1122.710 2801.450 1124.470 2801.750 ;
        RECT 1122.710 2794.625 1123.010 2801.450 ;
        RECT 1124.170 2800.000 1124.470 2801.450 ;
        RECT 1124.790 2801.750 1125.090 2804.600 ;
        RECT 1130.010 2801.750 1130.310 2804.600 ;
        RECT 1124.790 2801.450 1128.530 2801.750 ;
        RECT 1124.790 2800.000 1125.090 2801.450 ;
        RECT 1122.695 2794.295 1123.025 2794.625 ;
        RECT 1128.230 2788.505 1128.530 2801.450 ;
        RECT 1129.150 2801.450 1130.310 2801.750 ;
        RECT 1129.150 2799.385 1129.450 2801.450 ;
        RECT 1130.010 2800.000 1130.310 2801.450 ;
        RECT 1130.630 2800.050 1130.930 2804.600 ;
        RECT 1135.850 2801.750 1136.150 2804.600 ;
        RECT 1130.630 2799.750 1131.290 2800.050 ;
        RECT 1129.135 2799.055 1129.465 2799.385 ;
        RECT 1128.215 2788.175 1128.545 2788.505 ;
        RECT 1130.990 2787.825 1131.290 2799.750 ;
        RECT 1135.590 2800.000 1136.150 2801.750 ;
        RECT 1136.470 2801.750 1136.770 2804.600 ;
        RECT 1141.690 2802.450 1141.990 2804.600 ;
        RECT 1140.190 2802.150 1141.990 2802.450 ;
        RECT 1136.470 2801.450 1137.730 2801.750 ;
        RECT 1136.470 2800.000 1136.770 2801.450 ;
        RECT 1135.590 2796.665 1135.890 2800.000 ;
        RECT 1135.575 2796.335 1135.905 2796.665 ;
        RECT 1137.430 2787.825 1137.730 2801.450 ;
        RECT 1140.190 2794.625 1140.490 2802.150 ;
        RECT 1141.690 2800.000 1141.990 2802.150 ;
        RECT 1142.310 2801.750 1142.610 2804.600 ;
        RECT 1142.310 2801.450 1144.170 2801.750 ;
        RECT 1142.310 2800.000 1142.610 2801.450 ;
        RECT 1140.175 2794.295 1140.505 2794.625 ;
        RECT 1143.870 2787.825 1144.170 2801.450 ;
        RECT 1146.615 2800.050 1146.945 2800.065 ;
        RECT 1147.530 2800.050 1147.830 2804.600 ;
        RECT 1146.615 2799.750 1147.830 2800.050 ;
        RECT 1148.150 2801.750 1148.450 2804.600 ;
        RECT 1153.370 2801.750 1153.670 2804.600 ;
        RECT 1148.150 2801.450 1151.530 2801.750 ;
        RECT 1148.150 2800.000 1148.450 2801.450 ;
        RECT 1146.615 2799.735 1146.945 2799.750 ;
        RECT 1151.230 2787.825 1151.530 2801.450 ;
        RECT 1153.070 2800.000 1153.670 2801.750 ;
        RECT 1153.070 2792.585 1153.370 2800.000 ;
        RECT 1153.055 2792.255 1153.385 2792.585 ;
        RECT 1153.990 2787.825 1154.290 2804.600 ;
        RECT 1159.210 2796.650 1159.510 2804.600 ;
        RECT 1159.830 2801.750 1160.130 2804.600 ;
        RECT 1165.050 2801.750 1165.350 2804.600 ;
        RECT 1159.830 2801.450 1163.490 2801.750 ;
        RECT 1159.830 2800.000 1160.130 2801.450 ;
        RECT 1159.210 2796.350 1159.810 2796.650 ;
        RECT 1159.510 2793.265 1159.810 2796.350 ;
        RECT 1159.495 2792.935 1159.825 2793.265 ;
        RECT 1163.190 2788.505 1163.490 2801.450 ;
        RECT 1164.110 2801.450 1165.350 2801.750 ;
        RECT 1164.110 2793.945 1164.410 2801.450 ;
        RECT 1165.050 2800.000 1165.350 2801.450 ;
        RECT 1165.670 2796.650 1165.970 2804.600 ;
        RECT 1170.890 2801.750 1171.190 2804.600 ;
        RECT 1165.030 2796.350 1165.970 2796.650 ;
        RECT 1167.790 2801.450 1171.190 2801.750 ;
        RECT 1164.095 2793.615 1164.425 2793.945 ;
        RECT 1163.175 2788.175 1163.505 2788.505 ;
        RECT 1165.030 2787.825 1165.330 2796.350 ;
        RECT 1167.790 2793.945 1168.090 2801.450 ;
        RECT 1170.890 2800.000 1171.190 2801.450 ;
        RECT 1171.510 2801.750 1171.810 2804.600 ;
        RECT 1176.730 2801.750 1177.030 2804.600 ;
        RECT 1171.510 2801.450 1172.690 2801.750 ;
        RECT 1171.510 2800.000 1171.810 2801.450 ;
        RECT 1167.775 2793.615 1168.105 2793.945 ;
        RECT 1172.390 2787.825 1172.690 2801.450 ;
        RECT 1173.310 2801.450 1177.030 2801.750 ;
        RECT 1173.310 2793.945 1173.610 2801.450 ;
        RECT 1176.730 2800.000 1177.030 2801.450 ;
        RECT 1177.350 2801.750 1177.650 2804.600 ;
        RECT 1182.570 2801.750 1182.870 2804.600 ;
        RECT 1177.350 2801.450 1179.130 2801.750 ;
        RECT 1177.350 2800.000 1177.650 2801.450 ;
        RECT 1178.830 2794.625 1179.130 2801.450 ;
        RECT 1180.670 2801.450 1182.870 2801.750 ;
        RECT 1178.815 2794.295 1179.145 2794.625 ;
        RECT 1180.670 2793.945 1180.970 2801.450 ;
        RECT 1182.570 2800.000 1182.870 2801.450 ;
        RECT 1183.190 2801.750 1183.490 2804.600 ;
        RECT 1188.410 2801.750 1188.710 2804.600 ;
        RECT 1183.190 2801.450 1186.490 2801.750 ;
        RECT 1183.190 2800.000 1183.490 2801.450 ;
        RECT 1186.190 2794.625 1186.490 2801.450 ;
        RECT 1187.110 2801.450 1188.710 2801.750 ;
        RECT 1186.175 2794.295 1186.505 2794.625 ;
        RECT 1173.295 2793.615 1173.625 2793.945 ;
        RECT 1180.655 2793.615 1180.985 2793.945 ;
        RECT 1187.110 2793.265 1187.410 2801.450 ;
        RECT 1188.410 2800.000 1188.710 2801.450 ;
        RECT 1189.030 2801.750 1189.330 2804.600 ;
        RECT 1194.250 2801.750 1194.550 2804.600 ;
        RECT 1189.030 2801.450 1192.010 2801.750 ;
        RECT 1189.030 2800.000 1189.330 2801.450 ;
        RECT 1187.095 2792.935 1187.425 2793.265 ;
        RECT 1191.710 2790.545 1192.010 2801.450 ;
        RECT 1193.550 2801.450 1194.550 2801.750 ;
        RECT 1193.550 2791.905 1193.850 2801.450 ;
        RECT 1194.250 2800.000 1194.550 2801.450 ;
        RECT 1194.870 2801.750 1195.170 2804.600 ;
        RECT 1194.870 2801.450 1198.450 2801.750 ;
        RECT 1194.870 2800.000 1195.170 2801.450 ;
        RECT 1198.150 2794.625 1198.450 2801.450 ;
        RECT 1198.135 2794.295 1198.465 2794.625 ;
        RECT 1193.535 2791.575 1193.865 2791.905 ;
        RECT 1191.695 2790.215 1192.025 2790.545 ;
        RECT 507.215 2787.495 507.545 2787.825 ;
        RECT 513.655 2787.495 513.985 2787.825 ;
        RECT 516.415 2787.495 516.745 2787.825 ;
        RECT 520.095 2787.495 520.425 2787.825 ;
        RECT 526.535 2787.495 526.865 2787.825 ;
        RECT 530.215 2787.495 530.545 2787.825 ;
        RECT 538.495 2787.495 538.825 2787.825 ;
        RECT 544.935 2787.495 545.265 2787.825 ;
        RECT 1034.375 2787.495 1034.705 2787.825 ;
        RECT 1039.895 2787.495 1040.225 2787.825 ;
        RECT 1046.335 2787.495 1046.665 2787.825 ;
        RECT 1054.615 2787.495 1054.945 2787.825 ;
        RECT 1061.975 2787.495 1062.305 2787.825 ;
        RECT 1067.495 2787.495 1067.825 2787.825 ;
        RECT 1073.935 2787.495 1074.265 2787.825 ;
        RECT 1081.295 2787.495 1081.625 2787.825 ;
        RECT 1089.575 2787.495 1089.905 2787.825 ;
        RECT 1096.015 2787.495 1096.345 2787.825 ;
        RECT 1103.375 2787.495 1103.705 2787.825 ;
        RECT 1109.815 2787.495 1110.145 2787.825 ;
        RECT 1116.255 2787.495 1116.585 2787.825 ;
        RECT 1121.775 2787.495 1122.105 2787.825 ;
        RECT 1130.975 2787.495 1131.305 2787.825 ;
        RECT 1137.415 2787.495 1137.745 2787.825 ;
        RECT 1143.855 2787.495 1144.185 2787.825 ;
        RECT 1151.215 2787.495 1151.545 2787.825 ;
        RECT 1153.975 2787.495 1154.305 2787.825 ;
        RECT 1165.015 2787.495 1165.345 2787.825 ;
        RECT 1172.375 2787.495 1172.705 2787.825 ;
        RECT 292.020 2715.000 295.020 2785.000 ;
        RECT 310.020 2715.000 313.020 2785.000 ;
        RECT 328.020 2715.000 331.020 2785.000 ;
        RECT 364.020 2715.000 367.020 2785.000 ;
        RECT 454.020 2715.000 457.020 2785.000 ;
        RECT 472.020 2715.000 475.020 2785.000 ;
        RECT 490.020 2715.000 493.020 2785.000 ;
        RECT 508.020 2715.000 511.020 2785.000 ;
        RECT 544.020 2715.000 547.020 2785.000 ;
        RECT 634.020 2715.000 637.020 2785.000 ;
        RECT 652.020 2715.000 655.020 2785.000 ;
        RECT 670.020 2715.000 673.020 2785.000 ;
        RECT 688.020 2715.000 691.020 2785.000 ;
        RECT 994.020 2715.000 997.020 2785.000 ;
        RECT 1012.020 2715.000 1015.020 2785.000 ;
        RECT 1030.020 2715.000 1033.020 2785.000 ;
        RECT 1048.020 2715.000 1051.020 2785.000 ;
        RECT 1084.020 2715.000 1087.020 2785.000 ;
        RECT 1174.020 2715.000 1177.020 2785.000 ;
        RECT 1192.020 2715.000 1195.020 2785.000 ;
        RECT 1210.020 2715.000 1213.020 2785.000 ;
        RECT 1228.020 2715.000 1231.020 2785.000 ;
        RECT 1264.020 2715.000 1267.020 2785.000 ;
      LAYER met4 ;
        RECT 366.465 1610.640 397.370 2688.240 ;
        RECT 399.770 1610.640 1387.995 2688.240 ;
      LAYER met4 ;
        RECT 1411.590 1614.825 1411.890 3243.095 ;
        RECT 1412.990 2935.310 1414.170 2936.490 ;
      LAYER met4 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met4 ;
        RECT 1937.390 2935.310 1938.570 2936.490 ;
        RECT 2199.590 2897.910 2200.770 2899.090 ;
        RECT 2200.030 2895.945 2200.330 2897.910 ;
        RECT 2200.015 2895.615 2200.345 2895.945 ;
      LAYER met4 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met4 ;
        RECT 2594.695 2904.455 2595.025 2904.785 ;
        RECT 2594.710 2899.090 2595.010 2904.455 ;
        RECT 2594.270 2897.910 2595.450 2899.090 ;
        RECT 1584.010 2801.750 1584.310 2804.600 ;
        RECT 1589.850 2801.750 1590.150 2804.600 ;
        RECT 1595.690 2801.750 1595.990 2804.600 ;
        RECT 1580.870 2801.450 1584.310 2801.750 ;
        RECT 1580.870 2794.625 1581.170 2801.450 ;
        RECT 1584.010 2800.000 1584.310 2801.450 ;
        RECT 1587.310 2801.450 1590.150 2801.750 ;
        RECT 1587.310 2794.625 1587.610 2801.450 ;
        RECT 1589.850 2800.000 1590.150 2801.450 ;
        RECT 1594.670 2801.450 1595.990 2801.750 ;
        RECT 1580.855 2794.295 1581.185 2794.625 ;
        RECT 1587.295 2794.295 1587.625 2794.625 ;
        RECT 1594.670 2793.265 1594.970 2801.450 ;
        RECT 1595.690 2800.000 1595.990 2801.450 ;
        RECT 1601.530 2800.050 1601.830 2804.600 ;
        RECT 1607.370 2801.750 1607.670 2804.600 ;
        RECT 1613.210 2801.750 1613.510 2804.600 ;
        RECT 1601.110 2799.750 1601.830 2800.050 ;
        RECT 1604.790 2801.450 1607.670 2801.750 ;
        RECT 1601.110 2793.945 1601.410 2799.750 ;
        RECT 1604.790 2794.625 1605.090 2801.450 ;
        RECT 1607.370 2800.000 1607.670 2801.450 ;
        RECT 1613.070 2800.000 1613.510 2801.750 ;
        RECT 1613.830 2801.750 1614.130 2804.600 ;
        RECT 1619.050 2802.450 1619.350 2804.600 ;
        RECT 1617.670 2802.150 1619.350 2802.450 ;
        RECT 1613.830 2800.000 1614.290 2801.750 ;
        RECT 1613.070 2794.625 1613.370 2800.000 ;
        RECT 1604.775 2794.295 1605.105 2794.625 ;
        RECT 1613.055 2794.295 1613.385 2794.625 ;
        RECT 1601.095 2793.615 1601.425 2793.945 ;
        RECT 1594.655 2792.935 1594.985 2793.265 ;
        RECT 1613.990 2787.825 1614.290 2800.000 ;
        RECT 1617.670 2794.625 1617.970 2802.150 ;
        RECT 1619.050 2800.000 1619.350 2802.150 ;
        RECT 1619.670 2801.750 1619.970 2804.600 ;
        RECT 1624.890 2801.750 1625.190 2804.600 ;
        RECT 1619.670 2801.450 1620.730 2801.750 ;
        RECT 1619.670 2800.000 1619.970 2801.450 ;
        RECT 1617.655 2794.295 1617.985 2794.625 ;
        RECT 1620.430 2787.825 1620.730 2801.450 ;
        RECT 1624.110 2801.450 1625.190 2801.750 ;
        RECT 1624.110 2788.505 1624.410 2801.450 ;
        RECT 1624.890 2800.000 1625.190 2801.450 ;
        RECT 1625.510 2802.450 1625.810 2804.600 ;
        RECT 1625.510 2802.150 1627.170 2802.450 ;
        RECT 1625.510 2800.000 1625.810 2802.150 ;
        RECT 1624.095 2788.175 1624.425 2788.505 ;
        RECT 1626.870 2787.825 1627.170 2802.150 ;
        RECT 1630.730 2801.750 1631.030 2804.600 ;
        RECT 1630.550 2800.000 1631.030 2801.750 ;
        RECT 1631.350 2801.750 1631.650 2804.600 ;
        RECT 1636.570 2802.450 1636.870 2804.600 ;
        RECT 1635.150 2802.150 1636.870 2802.450 ;
        RECT 1631.350 2800.000 1631.770 2801.750 ;
        RECT 1630.550 2788.505 1630.850 2800.000 ;
        RECT 1630.535 2788.175 1630.865 2788.505 ;
        RECT 1631.470 2787.825 1631.770 2800.000 ;
        RECT 1635.150 2788.505 1635.450 2802.150 ;
        RECT 1636.570 2800.000 1636.870 2802.150 ;
        RECT 1637.190 2801.750 1637.490 2804.600 ;
        RECT 1637.190 2801.450 1638.210 2801.750 ;
        RECT 1637.190 2800.000 1637.490 2801.450 ;
        RECT 1635.135 2788.175 1635.465 2788.505 ;
        RECT 1637.910 2787.825 1638.210 2801.450 ;
        RECT 1642.410 2796.650 1642.710 2804.600 ;
        RECT 1643.030 2802.450 1643.330 2804.600 ;
        RECT 1643.030 2802.150 1644.650 2802.450 ;
        RECT 1643.030 2800.000 1643.330 2802.150 ;
        RECT 1642.410 2796.350 1642.810 2796.650 ;
        RECT 1642.510 2794.625 1642.810 2796.350 ;
        RECT 1642.495 2794.295 1642.825 2794.625 ;
        RECT 1644.350 2787.825 1644.650 2802.150 ;
        RECT 1648.250 2801.750 1648.550 2804.600 ;
        RECT 1648.030 2800.000 1648.550 2801.750 ;
        RECT 1648.870 2801.750 1649.170 2804.600 ;
        RECT 1654.090 2802.450 1654.390 2804.600 ;
        RECT 1652.630 2802.150 1654.390 2802.450 ;
        RECT 1648.870 2800.000 1649.250 2801.750 ;
        RECT 1648.030 2794.625 1648.330 2800.000 ;
        RECT 1648.015 2794.295 1648.345 2794.625 ;
        RECT 1648.950 2787.825 1649.250 2800.000 ;
        RECT 1652.630 2794.625 1652.930 2802.150 ;
        RECT 1654.090 2800.000 1654.390 2802.150 ;
        RECT 1654.710 2801.750 1655.010 2804.600 ;
        RECT 1659.930 2801.750 1660.230 2804.600 ;
        RECT 1654.710 2801.450 1655.690 2801.750 ;
        RECT 1654.710 2800.000 1655.010 2801.450 ;
        RECT 1652.615 2794.295 1652.945 2794.625 ;
        RECT 1655.390 2788.505 1655.690 2801.450 ;
        RECT 1659.070 2801.450 1660.230 2801.750 ;
        RECT 1659.070 2794.625 1659.370 2801.450 ;
        RECT 1659.930 2800.000 1660.230 2801.450 ;
        RECT 1660.550 2802.450 1660.850 2804.600 ;
        RECT 1660.550 2802.150 1662.130 2802.450 ;
        RECT 1660.550 2800.000 1660.850 2802.150 ;
        RECT 1659.055 2794.295 1659.385 2794.625 ;
        RECT 1655.375 2788.175 1655.705 2788.505 ;
        RECT 1661.830 2787.825 1662.130 2802.150 ;
        RECT 1665.770 2801.750 1666.070 2804.600 ;
        RECT 1665.510 2800.000 1666.070 2801.750 ;
        RECT 1666.390 2801.750 1666.690 2804.600 ;
        RECT 1671.610 2802.450 1671.910 2804.600 ;
        RECT 1670.110 2802.150 1671.910 2802.450 ;
        RECT 1666.390 2800.000 1666.730 2801.750 ;
        RECT 1665.510 2794.625 1665.810 2800.000 ;
        RECT 1665.495 2794.295 1665.825 2794.625 ;
        RECT 1666.430 2787.825 1666.730 2800.000 ;
        RECT 1670.110 2794.625 1670.410 2802.150 ;
        RECT 1671.610 2800.000 1671.910 2802.150 ;
        RECT 1672.230 2801.750 1672.530 2804.600 ;
        RECT 1672.230 2801.450 1673.170 2801.750 ;
        RECT 1672.230 2800.000 1672.530 2801.450 ;
        RECT 1670.095 2794.295 1670.425 2794.625 ;
        RECT 1672.870 2787.825 1673.170 2801.450 ;
        RECT 1677.450 2800.050 1677.750 2804.600 ;
        RECT 1678.070 2802.450 1678.370 2804.600 ;
        RECT 1678.070 2802.150 1679.610 2802.450 ;
        RECT 1677.450 2799.750 1677.770 2800.050 ;
        RECT 1678.070 2800.000 1678.370 2802.150 ;
        RECT 1677.470 2794.625 1677.770 2799.750 ;
        RECT 1677.455 2794.295 1677.785 2794.625 ;
        RECT 1679.310 2787.825 1679.610 2802.150 ;
        RECT 1683.290 2801.750 1683.590 2804.600 ;
        RECT 1682.070 2801.450 1683.590 2801.750 ;
        RECT 1682.070 2794.625 1682.370 2801.450 ;
        RECT 1683.290 2800.000 1683.590 2801.450 ;
        RECT 1682.055 2794.295 1682.385 2794.625 ;
        RECT 1683.910 2787.825 1684.210 2804.600 ;
        RECT 1689.130 2801.750 1689.430 2804.600 ;
        RECT 1688.510 2801.450 1689.430 2801.750 ;
        RECT 1688.510 2794.625 1688.810 2801.450 ;
        RECT 1689.130 2800.000 1689.430 2801.450 ;
        RECT 1689.750 2796.650 1690.050 2804.600 ;
        RECT 1694.970 2801.750 1695.270 2804.600 ;
        RECT 1689.430 2796.350 1690.050 2796.650 ;
        RECT 1694.950 2800.000 1695.270 2801.750 ;
        RECT 1695.590 2801.750 1695.890 2804.600 ;
        RECT 1700.810 2802.450 1701.110 2804.600 ;
        RECT 1699.550 2802.150 1701.110 2802.450 ;
        RECT 1695.590 2800.000 1696.170 2801.750 ;
        RECT 1688.495 2794.295 1688.825 2794.625 ;
        RECT 1689.430 2788.505 1689.730 2796.350 ;
        RECT 1694.950 2794.625 1695.250 2800.000 ;
        RECT 1694.935 2794.295 1695.265 2794.625 ;
        RECT 1689.415 2788.175 1689.745 2788.505 ;
        RECT 1695.870 2787.825 1696.170 2800.000 ;
        RECT 1699.550 2794.625 1699.850 2802.150 ;
        RECT 1700.810 2800.000 1701.110 2802.150 ;
        RECT 1701.430 2801.750 1701.730 2804.600 ;
        RECT 1706.650 2801.750 1706.950 2804.600 ;
        RECT 1701.430 2801.450 1702.610 2801.750 ;
        RECT 1701.430 2800.000 1701.730 2801.450 ;
        RECT 1699.535 2794.295 1699.865 2794.625 ;
        RECT 1702.310 2787.825 1702.610 2801.450 ;
        RECT 1705.990 2801.450 1706.950 2801.750 ;
        RECT 1705.990 2794.625 1706.290 2801.450 ;
        RECT 1706.650 2800.000 1706.950 2801.450 ;
        RECT 1707.270 2802.450 1707.570 2804.600 ;
        RECT 1707.270 2802.150 1709.050 2802.450 ;
        RECT 1707.270 2800.000 1707.570 2802.150 ;
        RECT 1705.975 2794.295 1706.305 2794.625 ;
        RECT 1708.750 2787.825 1709.050 2802.150 ;
        RECT 1712.490 2801.750 1712.790 2804.600 ;
        RECT 1712.430 2800.000 1712.790 2801.750 ;
        RECT 1713.110 2801.750 1713.410 2804.600 ;
        RECT 1713.110 2800.000 1713.650 2801.750 ;
        RECT 1718.330 2800.050 1718.630 2804.600 ;
        RECT 1712.430 2794.625 1712.730 2800.000 ;
        RECT 1712.415 2794.295 1712.745 2794.625 ;
        RECT 1713.350 2787.825 1713.650 2800.000 ;
        RECT 1717.950 2799.750 1718.630 2800.050 ;
        RECT 1718.950 2801.750 1719.250 2804.600 ;
        RECT 1724.170 2801.750 1724.470 2804.600 ;
        RECT 1718.950 2801.450 1720.090 2801.750 ;
        RECT 1718.950 2800.000 1719.250 2801.450 ;
        RECT 1717.950 2794.625 1718.250 2799.750 ;
        RECT 1717.935 2794.295 1718.265 2794.625 ;
        RECT 1719.790 2787.825 1720.090 2801.450 ;
        RECT 1723.470 2801.450 1724.470 2801.750 ;
        RECT 1723.470 2794.625 1723.770 2801.450 ;
        RECT 1724.170 2800.000 1724.470 2801.450 ;
        RECT 1724.790 2796.650 1725.090 2804.600 ;
        RECT 1730.010 2801.750 1730.310 2804.600 ;
        RECT 1724.390 2796.350 1725.090 2796.650 ;
        RECT 1728.990 2801.450 1730.310 2801.750 ;
        RECT 1723.455 2794.295 1723.785 2794.625 ;
        RECT 1724.390 2788.505 1724.690 2796.350 ;
        RECT 1728.990 2794.625 1729.290 2801.450 ;
        RECT 1730.010 2800.000 1730.310 2801.450 ;
        RECT 1730.630 2801.750 1730.930 2804.600 ;
        RECT 1735.850 2801.750 1736.150 2804.600 ;
        RECT 1730.630 2800.000 1731.130 2801.750 ;
        RECT 1728.975 2794.295 1729.305 2794.625 ;
        RECT 1724.375 2788.175 1724.705 2788.505 ;
        RECT 1730.830 2787.825 1731.130 2800.000 ;
        RECT 1732.670 2801.450 1736.150 2801.750 ;
        RECT 1732.670 2794.625 1732.970 2801.450 ;
        RECT 1735.850 2800.000 1736.150 2801.450 ;
        RECT 1736.470 2801.750 1736.770 2804.600 ;
        RECT 1741.690 2801.750 1741.990 2804.600 ;
        RECT 1736.470 2801.450 1737.570 2801.750 ;
        RECT 1736.470 2800.000 1736.770 2801.450 ;
        RECT 1732.655 2794.295 1732.985 2794.625 ;
        RECT 1737.270 2787.825 1737.570 2801.450 ;
        RECT 1740.950 2801.450 1741.990 2801.750 ;
        RECT 1740.950 2794.625 1741.250 2801.450 ;
        RECT 1741.690 2800.000 1741.990 2801.450 ;
        RECT 1742.310 2802.450 1742.610 2804.600 ;
        RECT 1742.310 2802.150 1744.010 2802.450 ;
        RECT 1742.310 2800.000 1742.610 2802.150 ;
        RECT 1740.935 2794.295 1741.265 2794.625 ;
        RECT 1743.710 2787.825 1744.010 2802.150 ;
        RECT 1747.530 2801.750 1747.830 2804.600 ;
        RECT 1747.390 2800.000 1747.830 2801.750 ;
        RECT 1748.150 2801.750 1748.450 2804.600 ;
        RECT 1748.150 2800.000 1748.610 2801.750 ;
        RECT 1753.370 2800.050 1753.670 2804.600 ;
        RECT 1747.390 2794.625 1747.690 2800.000 ;
        RECT 1747.375 2794.295 1747.705 2794.625 ;
        RECT 1748.310 2787.825 1748.610 2800.000 ;
        RECT 1752.910 2799.750 1753.670 2800.050 ;
        RECT 1753.990 2801.750 1754.290 2804.600 ;
        RECT 1753.990 2801.450 1755.050 2801.750 ;
        RECT 1753.990 2800.000 1754.290 2801.450 ;
        RECT 1752.910 2794.625 1753.210 2799.750 ;
        RECT 1752.895 2794.295 1753.225 2794.625 ;
        RECT 1754.750 2787.825 1755.050 2801.450 ;
        RECT 1759.210 2796.665 1759.510 2804.600 ;
        RECT 1759.830 2802.450 1760.130 2804.600 ;
        RECT 1759.830 2802.150 1761.490 2802.450 ;
        RECT 1759.830 2800.000 1760.130 2802.150 ;
        RECT 1759.210 2796.350 1759.665 2796.665 ;
        RECT 1759.335 2796.335 1759.665 2796.350 ;
        RECT 1613.975 2787.495 1614.305 2787.825 ;
        RECT 1620.415 2787.495 1620.745 2787.825 ;
        RECT 1626.855 2787.495 1627.185 2787.825 ;
        RECT 1631.455 2787.495 1631.785 2787.825 ;
        RECT 1637.895 2787.495 1638.225 2787.825 ;
        RECT 1644.335 2787.495 1644.665 2787.825 ;
        RECT 1648.935 2787.495 1649.265 2787.825 ;
        RECT 1661.815 2787.495 1662.145 2787.825 ;
        RECT 1666.415 2787.495 1666.745 2787.825 ;
        RECT 1672.855 2787.495 1673.185 2787.825 ;
        RECT 1679.295 2787.495 1679.625 2787.825 ;
        RECT 1683.895 2787.495 1684.225 2787.825 ;
        RECT 1695.855 2787.495 1696.185 2787.825 ;
        RECT 1702.295 2787.495 1702.625 2787.825 ;
        RECT 1708.735 2787.495 1709.065 2787.825 ;
        RECT 1713.335 2787.495 1713.665 2787.825 ;
        RECT 1719.775 2787.495 1720.105 2787.825 ;
        RECT 1730.815 2787.495 1731.145 2787.825 ;
        RECT 1737.255 2787.495 1737.585 2787.825 ;
        RECT 1743.695 2787.495 1744.025 2787.825 ;
        RECT 1748.295 2787.495 1748.625 2787.825 ;
        RECT 1754.735 2787.495 1755.065 2787.825 ;
        RECT 1761.190 2777.625 1761.490 2802.150 ;
        RECT 1765.050 2801.750 1765.350 2804.600 ;
        RECT 1762.110 2801.450 1765.350 2801.750 ;
        RECT 1762.110 2794.625 1762.410 2801.450 ;
        RECT 1765.050 2800.000 1765.350 2801.450 ;
        RECT 1765.670 2801.750 1765.970 2804.600 ;
        RECT 1770.890 2801.750 1771.190 2804.600 ;
        RECT 1765.670 2800.000 1766.090 2801.750 ;
        RECT 1762.095 2794.295 1762.425 2794.625 ;
        RECT 1765.790 2788.505 1766.090 2800.000 ;
        RECT 1767.630 2801.450 1771.190 2801.750 ;
        RECT 1767.630 2794.625 1767.930 2801.450 ;
        RECT 1770.890 2800.000 1771.190 2801.450 ;
        RECT 1771.510 2801.750 1771.810 2804.600 ;
        RECT 1776.730 2801.750 1777.030 2804.600 ;
        RECT 1771.510 2801.450 1772.530 2801.750 ;
        RECT 1771.510 2800.000 1771.810 2801.450 ;
        RECT 1767.615 2794.295 1767.945 2794.625 ;
        RECT 1765.775 2788.175 1766.105 2788.505 ;
        RECT 1772.230 2787.825 1772.530 2801.450 ;
        RECT 1774.070 2801.450 1777.030 2801.750 ;
        RECT 1774.070 2793.945 1774.370 2801.450 ;
        RECT 1776.730 2800.000 1777.030 2801.450 ;
        RECT 1777.350 2802.450 1777.650 2804.600 ;
        RECT 1777.350 2802.150 1778.970 2802.450 ;
        RECT 1777.350 2800.000 1777.650 2802.150 ;
        RECT 1774.055 2793.615 1774.385 2793.945 ;
        RECT 1778.670 2787.825 1778.970 2802.150 ;
        RECT 1782.570 2801.750 1782.870 2804.600 ;
        RECT 1780.510 2801.450 1782.870 2801.750 ;
        RECT 1780.510 2793.945 1780.810 2801.450 ;
        RECT 1782.570 2800.000 1782.870 2801.450 ;
        RECT 1783.190 2801.750 1783.490 2804.600 ;
        RECT 1783.190 2800.000 1783.570 2801.750 ;
        RECT 1788.410 2800.050 1788.710 2804.600 ;
        RECT 1780.495 2793.615 1780.825 2793.945 ;
        RECT 1783.270 2787.825 1783.570 2800.000 ;
        RECT 1787.870 2799.750 1788.710 2800.050 ;
        RECT 1789.030 2801.750 1789.330 2804.600 ;
        RECT 1789.030 2801.450 1790.010 2801.750 ;
        RECT 1789.030 2800.000 1789.330 2801.450 ;
        RECT 1787.870 2792.585 1788.170 2799.750 ;
        RECT 1787.855 2792.255 1788.185 2792.585 ;
        RECT 1789.710 2787.825 1790.010 2801.450 ;
        RECT 1794.250 2796.665 1794.550 2804.600 ;
        RECT 1794.870 2802.450 1795.170 2804.600 ;
        RECT 1794.870 2802.150 1796.450 2802.450 ;
        RECT 1794.870 2800.000 1795.170 2802.150 ;
        RECT 1794.250 2796.350 1794.625 2796.665 ;
        RECT 1794.295 2796.335 1794.625 2796.350 ;
        RECT 1772.215 2787.495 1772.545 2787.825 ;
        RECT 1778.655 2787.495 1778.985 2787.825 ;
        RECT 1783.255 2787.495 1783.585 2787.825 ;
        RECT 1789.695 2787.495 1790.025 2787.825 ;
        RECT 1796.150 2777.625 1796.450 2802.150 ;
        RECT 2234.010 2801.750 2234.310 2804.600 ;
        RECT 2239.850 2801.750 2240.150 2804.600 ;
        RECT 2245.690 2801.750 2245.990 2804.600 ;
        RECT 2251.530 2801.750 2251.830 2804.600 ;
        RECT 2257.370 2801.750 2257.670 2804.600 ;
        RECT 2231.310 2801.450 2234.310 2801.750 ;
        RECT 2231.310 2794.625 2231.610 2801.450 ;
        RECT 2234.010 2800.000 2234.310 2801.450 ;
        RECT 2238.670 2801.450 2240.150 2801.750 ;
        RECT 2238.670 2794.625 2238.970 2801.450 ;
        RECT 2239.850 2800.000 2240.150 2801.450 ;
        RECT 2242.350 2801.450 2245.990 2801.750 ;
        RECT 2231.295 2794.295 2231.625 2794.625 ;
        RECT 2238.655 2794.295 2238.985 2794.625 ;
        RECT 2242.350 2791.225 2242.650 2801.450 ;
        RECT 2245.690 2800.000 2245.990 2801.450 ;
        RECT 2249.710 2801.450 2251.830 2801.750 ;
        RECT 2249.710 2792.585 2250.010 2801.450 ;
        RECT 2251.530 2800.000 2251.830 2801.450 ;
        RECT 2257.070 2800.000 2257.670 2801.750 ;
        RECT 2249.695 2792.255 2250.025 2792.585 ;
        RECT 2242.335 2790.895 2242.665 2791.225 ;
        RECT 2257.070 2790.545 2257.370 2800.000 ;
        RECT 2263.210 2796.650 2263.510 2804.600 ;
        RECT 2263.830 2801.750 2264.130 2804.600 ;
        RECT 2269.050 2801.750 2269.350 2804.600 ;
        RECT 2263.830 2801.450 2264.730 2801.750 ;
        RECT 2263.830 2800.000 2264.130 2801.450 ;
        RECT 2263.210 2796.350 2263.810 2796.650 ;
        RECT 2263.510 2793.265 2263.810 2796.350 ;
        RECT 2263.495 2792.935 2263.825 2793.265 ;
        RECT 2257.055 2790.215 2257.385 2790.545 ;
        RECT 2264.430 2787.825 2264.730 2801.450 ;
        RECT 2268.110 2801.450 2269.350 2801.750 ;
        RECT 2268.110 2794.625 2268.410 2801.450 ;
        RECT 2269.050 2800.000 2269.350 2801.450 ;
        RECT 2269.670 2796.650 2269.970 2804.600 ;
        RECT 2274.890 2802.450 2275.190 2804.600 ;
        RECT 2269.030 2796.350 2269.970 2796.650 ;
        RECT 2273.630 2802.150 2275.190 2802.450 ;
        RECT 2268.095 2794.295 2268.425 2794.625 ;
        RECT 2269.030 2793.945 2269.330 2796.350 ;
        RECT 2273.630 2794.625 2273.930 2802.150 ;
        RECT 2274.890 2800.000 2275.190 2802.150 ;
        RECT 2275.510 2801.750 2275.810 2804.600 ;
        RECT 2280.730 2801.750 2281.030 2804.600 ;
        RECT 2275.510 2801.450 2276.690 2801.750 ;
        RECT 2275.510 2800.000 2275.810 2801.450 ;
        RECT 2273.615 2794.295 2273.945 2794.625 ;
        RECT 2269.015 2793.615 2269.345 2793.945 ;
        RECT 2276.390 2787.825 2276.690 2801.450 ;
        RECT 2280.070 2801.450 2281.030 2801.750 ;
        RECT 2280.070 2794.625 2280.370 2801.450 ;
        RECT 2280.730 2800.000 2281.030 2801.450 ;
        RECT 2281.350 2802.450 2281.650 2804.600 ;
        RECT 2281.350 2802.150 2283.130 2802.450 ;
        RECT 2281.350 2800.000 2281.650 2802.150 ;
        RECT 2280.055 2794.295 2280.385 2794.625 ;
        RECT 2282.830 2787.825 2283.130 2802.150 ;
        RECT 2286.570 2801.750 2286.870 2804.600 ;
        RECT 2286.510 2800.000 2286.870 2801.750 ;
        RECT 2287.190 2801.750 2287.490 2804.600 ;
        RECT 2292.410 2802.450 2292.710 2804.600 ;
        RECT 2291.110 2802.150 2292.710 2802.450 ;
        RECT 2287.190 2800.000 2287.730 2801.750 ;
        RECT 2286.510 2794.625 2286.810 2800.000 ;
        RECT 2286.495 2794.295 2286.825 2794.625 ;
        RECT 2287.430 2787.825 2287.730 2800.000 ;
        RECT 2291.110 2794.625 2291.410 2802.150 ;
        RECT 2292.410 2800.000 2292.710 2802.150 ;
        RECT 2293.030 2801.750 2293.330 2804.600 ;
        RECT 2298.250 2801.750 2298.550 2804.600 ;
        RECT 2293.030 2801.450 2294.170 2801.750 ;
        RECT 2293.030 2800.000 2293.330 2801.450 ;
        RECT 2291.095 2794.295 2291.425 2794.625 ;
        RECT 2293.870 2787.825 2294.170 2801.450 ;
        RECT 2297.550 2801.450 2298.550 2801.750 ;
        RECT 2297.550 2793.265 2297.850 2801.450 ;
        RECT 2298.250 2800.000 2298.550 2801.450 ;
        RECT 2298.870 2802.450 2299.170 2804.600 ;
        RECT 2298.870 2802.150 2300.610 2802.450 ;
        RECT 2298.870 2800.000 2299.170 2802.150 ;
        RECT 2297.535 2792.935 2297.865 2793.265 ;
        RECT 2300.310 2787.825 2300.610 2802.150 ;
        RECT 2304.090 2801.750 2304.390 2804.600 ;
        RECT 2303.990 2800.000 2304.390 2801.750 ;
        RECT 2304.710 2801.750 2305.010 2804.600 ;
        RECT 2309.930 2801.750 2310.230 2804.600 ;
        RECT 2304.710 2800.000 2305.210 2801.750 ;
        RECT 2303.990 2794.625 2304.290 2800.000 ;
        RECT 2303.975 2794.295 2304.305 2794.625 ;
        RECT 2304.910 2787.825 2305.210 2800.000 ;
        RECT 2308.590 2801.450 2310.230 2801.750 ;
        RECT 2308.590 2794.625 2308.890 2801.450 ;
        RECT 2309.930 2800.000 2310.230 2801.450 ;
        RECT 2310.550 2796.650 2310.850 2804.600 ;
        RECT 2315.770 2801.750 2316.070 2804.600 ;
        RECT 2310.430 2796.350 2310.850 2796.650 ;
        RECT 2313.190 2801.450 2316.070 2801.750 ;
        RECT 2308.575 2794.295 2308.905 2794.625 ;
        RECT 2310.430 2788.505 2310.730 2796.350 ;
        RECT 2313.190 2794.625 2313.490 2801.450 ;
        RECT 2315.770 2800.000 2316.070 2801.450 ;
        RECT 2316.390 2802.450 2316.690 2804.600 ;
        RECT 2316.390 2802.150 2318.090 2802.450 ;
        RECT 2316.390 2800.000 2316.690 2802.150 ;
        RECT 2313.175 2794.295 2313.505 2794.625 ;
        RECT 2310.415 2788.175 2310.745 2788.505 ;
        RECT 2317.790 2787.825 2318.090 2802.150 ;
        RECT 2321.610 2801.750 2321.910 2804.600 ;
        RECT 2321.470 2800.000 2321.910 2801.750 ;
        RECT 2322.230 2801.750 2322.530 2804.600 ;
        RECT 2327.450 2802.450 2327.750 2804.600 ;
        RECT 2326.070 2802.150 2327.750 2802.450 ;
        RECT 2322.230 2800.000 2322.690 2801.750 ;
        RECT 2321.470 2794.625 2321.770 2800.000 ;
        RECT 2321.455 2794.295 2321.785 2794.625 ;
        RECT 2322.390 2787.825 2322.690 2800.000 ;
        RECT 2326.070 2794.625 2326.370 2802.150 ;
        RECT 2327.450 2800.000 2327.750 2802.150 ;
        RECT 2328.070 2801.750 2328.370 2804.600 ;
        RECT 2333.290 2801.750 2333.590 2804.600 ;
        RECT 2328.070 2801.450 2329.130 2801.750 ;
        RECT 2328.070 2800.000 2328.370 2801.450 ;
        RECT 2326.055 2794.295 2326.385 2794.625 ;
        RECT 2328.830 2787.825 2329.130 2801.450 ;
        RECT 2332.510 2801.450 2333.590 2801.750 ;
        RECT 2332.510 2793.945 2332.810 2801.450 ;
        RECT 2333.290 2800.000 2333.590 2801.450 ;
        RECT 2333.910 2800.050 2334.210 2804.600 ;
        RECT 2339.130 2801.750 2339.430 2804.600 ;
        RECT 2333.910 2799.750 2334.650 2800.050 ;
        RECT 2334.350 2794.625 2334.650 2799.750 ;
        RECT 2338.950 2800.000 2339.430 2801.750 ;
        RECT 2339.750 2801.750 2340.050 2804.600 ;
        RECT 2344.970 2802.450 2345.270 2804.600 ;
        RECT 2343.550 2802.150 2345.270 2802.450 ;
        RECT 2339.750 2800.000 2340.170 2801.750 ;
        RECT 2334.335 2794.295 2334.665 2794.625 ;
        RECT 2332.495 2793.615 2332.825 2793.945 ;
        RECT 2338.950 2793.265 2339.250 2800.000 ;
        RECT 2339.870 2794.625 2340.170 2800.000 ;
        RECT 2343.550 2794.625 2343.850 2802.150 ;
        RECT 2344.970 2800.000 2345.270 2802.150 ;
        RECT 2345.590 2796.650 2345.890 2804.600 ;
        RECT 2350.810 2801.750 2351.110 2804.600 ;
        RECT 2345.390 2796.350 2345.890 2796.650 ;
        RECT 2349.990 2801.450 2351.110 2801.750 ;
        RECT 2339.855 2794.295 2340.185 2794.625 ;
        RECT 2343.535 2794.295 2343.865 2794.625 ;
        RECT 2345.390 2793.945 2345.690 2796.350 ;
        RECT 2349.990 2793.945 2350.290 2801.450 ;
        RECT 2350.810 2800.000 2351.110 2801.450 ;
        RECT 2351.430 2800.050 2351.730 2804.600 ;
        RECT 2356.650 2801.750 2356.950 2804.600 ;
        RECT 2351.430 2799.750 2352.130 2800.050 ;
        RECT 2351.830 2794.625 2352.130 2799.750 ;
        RECT 2356.430 2800.000 2356.950 2801.750 ;
        RECT 2357.270 2801.750 2357.570 2804.600 ;
        RECT 2362.490 2802.450 2362.790 2804.600 ;
        RECT 2361.030 2802.150 2362.790 2802.450 ;
        RECT 2357.270 2800.000 2357.650 2801.750 ;
        RECT 2351.815 2794.295 2352.145 2794.625 ;
        RECT 2356.430 2793.945 2356.730 2800.000 ;
        RECT 2357.350 2794.625 2357.650 2800.000 ;
        RECT 2357.335 2794.295 2357.665 2794.625 ;
        RECT 2361.030 2793.945 2361.330 2802.150 ;
        RECT 2362.490 2800.000 2362.790 2802.150 ;
        RECT 2363.110 2801.750 2363.410 2804.600 ;
        RECT 2368.330 2801.750 2368.630 2804.600 ;
        RECT 2363.110 2801.450 2364.090 2801.750 ;
        RECT 2363.110 2800.000 2363.410 2801.450 ;
        RECT 2363.790 2794.625 2364.090 2801.450 ;
        RECT 2367.470 2801.450 2368.630 2801.750 ;
        RECT 2363.775 2794.295 2364.105 2794.625 ;
        RECT 2345.375 2793.615 2345.705 2793.945 ;
        RECT 2349.975 2793.615 2350.305 2793.945 ;
        RECT 2356.415 2793.615 2356.745 2793.945 ;
        RECT 2361.015 2793.615 2361.345 2793.945 ;
        RECT 2367.470 2793.265 2367.770 2801.450 ;
        RECT 2368.330 2800.000 2368.630 2801.450 ;
        RECT 2368.950 2802.450 2369.250 2804.600 ;
        RECT 2368.950 2802.150 2370.530 2802.450 ;
        RECT 2368.950 2800.000 2369.250 2802.150 ;
        RECT 2370.230 2794.625 2370.530 2802.150 ;
        RECT 2374.170 2801.750 2374.470 2804.600 ;
        RECT 2373.910 2800.000 2374.470 2801.750 ;
        RECT 2374.790 2801.750 2375.090 2804.600 ;
        RECT 2380.010 2801.750 2380.310 2804.600 ;
        RECT 2374.790 2800.000 2375.130 2801.750 ;
        RECT 2373.910 2794.625 2374.210 2800.000 ;
        RECT 2370.215 2794.295 2370.545 2794.625 ;
        RECT 2373.895 2794.295 2374.225 2794.625 ;
        RECT 2338.935 2792.935 2339.265 2793.265 ;
        RECT 2367.455 2792.935 2367.785 2793.265 ;
        RECT 2374.830 2791.905 2375.130 2800.000 ;
        RECT 2377.590 2801.450 2380.310 2801.750 ;
        RECT 2377.590 2794.625 2377.890 2801.450 ;
        RECT 2380.010 2800.000 2380.310 2801.450 ;
        RECT 2380.630 2801.750 2380.930 2804.600 ;
        RECT 2380.630 2801.450 2381.570 2801.750 ;
        RECT 2380.630 2800.000 2380.930 2801.450 ;
        RECT 2377.575 2794.295 2377.905 2794.625 ;
        RECT 2381.270 2791.905 2381.570 2801.450 ;
        RECT 2385.850 2800.050 2386.150 2804.600 ;
        RECT 2386.470 2800.050 2386.770 2804.600 ;
        RECT 2391.690 2801.750 2391.990 2804.600 ;
        RECT 2385.850 2799.750 2386.170 2800.050 ;
        RECT 2386.470 2799.750 2387.090 2800.050 ;
        RECT 2385.870 2794.625 2386.170 2799.750 ;
        RECT 2385.855 2794.295 2386.185 2794.625 ;
        RECT 2386.790 2792.585 2387.090 2799.750 ;
        RECT 2391.390 2800.000 2391.990 2801.750 ;
        RECT 2391.390 2794.625 2391.690 2800.000 ;
        RECT 2391.375 2794.295 2391.705 2794.625 ;
        RECT 2386.775 2792.255 2387.105 2792.585 ;
        RECT 2392.310 2791.905 2392.610 2804.600 ;
        RECT 2397.530 2801.750 2397.830 2804.600 ;
        RECT 2395.070 2801.450 2397.830 2801.750 ;
        RECT 2395.070 2794.625 2395.370 2801.450 ;
        RECT 2397.530 2800.000 2397.830 2801.450 ;
        RECT 2398.150 2801.750 2398.450 2804.600 ;
        RECT 2403.370 2801.750 2403.670 2804.600 ;
        RECT 2398.150 2801.450 2399.050 2801.750 ;
        RECT 2398.150 2800.000 2398.450 2801.450 ;
        RECT 2395.055 2794.295 2395.385 2794.625 ;
        RECT 2374.815 2791.575 2375.145 2791.905 ;
        RECT 2381.255 2791.575 2381.585 2791.905 ;
        RECT 2392.295 2791.575 2392.625 2791.905 ;
        RECT 2398.750 2791.225 2399.050 2801.450 ;
        RECT 2402.430 2801.450 2403.670 2801.750 ;
        RECT 2402.430 2793.945 2402.730 2801.450 ;
        RECT 2403.370 2800.000 2403.670 2801.450 ;
        RECT 2403.990 2801.750 2404.290 2804.600 ;
        RECT 2409.210 2802.450 2409.510 2804.600 ;
        RECT 2407.950 2802.150 2409.510 2802.450 ;
        RECT 2403.990 2800.000 2404.570 2801.750 ;
        RECT 2404.270 2794.625 2404.570 2800.000 ;
        RECT 2404.255 2794.295 2404.585 2794.625 ;
        RECT 2407.950 2793.945 2408.250 2802.150 ;
        RECT 2409.210 2800.000 2409.510 2802.150 ;
        RECT 2409.830 2801.750 2410.130 2804.600 ;
        RECT 2409.830 2801.450 2411.010 2801.750 ;
        RECT 2409.830 2800.000 2410.130 2801.450 ;
        RECT 2402.415 2793.615 2402.745 2793.945 ;
        RECT 2407.935 2793.615 2408.265 2793.945 ;
        RECT 2410.710 2792.585 2411.010 2801.450 ;
        RECT 2415.050 2796.650 2415.350 2804.600 ;
        RECT 2415.670 2802.450 2415.970 2804.600 ;
        RECT 2415.670 2802.150 2417.450 2802.450 ;
        RECT 2415.670 2800.000 2415.970 2802.150 ;
        RECT 2415.050 2796.350 2415.610 2796.650 ;
        RECT 2410.695 2792.255 2411.025 2792.585 ;
        RECT 2398.735 2790.895 2399.065 2791.225 ;
        RECT 2415.310 2788.505 2415.610 2796.350 ;
        RECT 2417.150 2791.225 2417.450 2802.150 ;
        RECT 2420.890 2801.750 2421.190 2804.600 ;
        RECT 2418.070 2801.450 2421.190 2801.750 ;
        RECT 2418.070 2794.625 2418.370 2801.450 ;
        RECT 2420.890 2800.000 2421.190 2801.450 ;
        RECT 2421.510 2796.650 2421.810 2804.600 ;
        RECT 2426.730 2801.750 2427.030 2804.600 ;
        RECT 2420.830 2796.350 2421.810 2796.650 ;
        RECT 2423.590 2801.450 2427.030 2801.750 ;
        RECT 2418.055 2794.295 2418.385 2794.625 ;
        RECT 2417.135 2790.895 2417.465 2791.225 ;
        RECT 2420.830 2790.545 2421.130 2796.350 ;
        RECT 2423.590 2793.265 2423.890 2801.450 ;
        RECT 2426.730 2800.000 2427.030 2801.450 ;
        RECT 2427.350 2801.750 2427.650 2804.600 ;
        RECT 2432.570 2801.750 2432.870 2804.600 ;
        RECT 2427.350 2801.450 2428.490 2801.750 ;
        RECT 2427.350 2800.000 2427.650 2801.450 ;
        RECT 2423.575 2792.935 2423.905 2793.265 ;
        RECT 2428.190 2791.225 2428.490 2801.450 ;
        RECT 2430.030 2801.450 2432.870 2801.750 ;
        RECT 2430.030 2792.585 2430.330 2801.450 ;
        RECT 2432.570 2800.000 2432.870 2801.450 ;
        RECT 2433.190 2802.450 2433.490 2804.600 ;
        RECT 2433.190 2802.150 2434.930 2802.450 ;
        RECT 2433.190 2800.000 2433.490 2802.150 ;
        RECT 2430.015 2792.255 2430.345 2792.585 ;
        RECT 2434.630 2791.225 2434.930 2802.150 ;
        RECT 2438.410 2801.750 2438.710 2804.600 ;
        RECT 2436.470 2801.450 2438.710 2801.750 ;
        RECT 2436.470 2792.585 2436.770 2801.450 ;
        RECT 2438.410 2800.000 2438.710 2801.450 ;
        RECT 2439.030 2801.750 2439.330 2804.600 ;
        RECT 2444.250 2801.750 2444.550 2804.600 ;
        RECT 2439.030 2800.000 2439.530 2801.750 ;
        RECT 2436.455 2792.255 2436.785 2792.585 ;
        RECT 2428.175 2790.895 2428.505 2791.225 ;
        RECT 2434.615 2790.895 2434.945 2791.225 ;
        RECT 2420.815 2790.215 2421.145 2790.545 ;
        RECT 2439.230 2789.865 2439.530 2800.000 ;
        RECT 2442.910 2801.450 2444.550 2801.750 ;
        RECT 2442.910 2793.265 2443.210 2801.450 ;
        RECT 2444.250 2800.000 2444.550 2801.450 ;
        RECT 2444.870 2801.750 2445.170 2804.600 ;
        RECT 2444.870 2801.450 2445.970 2801.750 ;
        RECT 2444.870 2800.000 2445.170 2801.450 ;
        RECT 2442.895 2792.935 2443.225 2793.265 ;
        RECT 2445.670 2790.545 2445.970 2801.450 ;
        RECT 2445.655 2790.215 2445.985 2790.545 ;
        RECT 2439.215 2789.535 2439.545 2789.865 ;
        RECT 2415.295 2788.175 2415.625 2788.505 ;
        RECT 2264.415 2787.495 2264.745 2787.825 ;
        RECT 2276.375 2787.495 2276.705 2787.825 ;
        RECT 2282.815 2787.495 2283.145 2787.825 ;
        RECT 2287.415 2787.495 2287.745 2787.825 ;
        RECT 2293.855 2787.495 2294.185 2787.825 ;
        RECT 2300.295 2787.495 2300.625 2787.825 ;
        RECT 2304.895 2787.495 2305.225 2787.825 ;
        RECT 2317.775 2787.495 2318.105 2787.825 ;
        RECT 2322.375 2787.495 2322.705 2787.825 ;
        RECT 2328.815 2787.495 2329.145 2787.825 ;
        RECT 1761.175 2777.295 1761.505 2777.625 ;
        RECT 1796.135 2777.295 1796.465 2777.625 ;
        RECT 1691.310 2051.635 1691.610 2056.235 ;
        RECT 1691.930 2051.635 1692.230 2056.235 ;
        RECT 1697.150 2051.635 1697.450 2056.235 ;
        RECT 1697.770 2051.635 1698.070 2056.235 ;
        RECT 1702.990 2051.635 1703.290 2056.235 ;
        RECT 1703.610 2051.635 1703.910 2056.235 ;
        RECT 1708.830 2051.635 1709.130 2056.235 ;
        RECT 1709.450 2051.635 1709.750 2056.235 ;
        RECT 1714.670 2051.635 1714.970 2056.235 ;
        RECT 1715.290 2051.635 1715.590 2056.235 ;
        RECT 1720.510 2051.635 1720.810 2056.235 ;
        RECT 1721.130 2051.635 1721.430 2056.235 ;
        RECT 1726.350 2051.635 1726.650 2056.235 ;
        RECT 1726.970 2051.635 1727.270 2056.235 ;
        RECT 1732.190 2051.635 1732.490 2056.235 ;
        RECT 1732.810 2051.635 1733.110 2056.235 ;
        RECT 1738.030 2051.635 1738.330 2056.235 ;
        RECT 1738.650 2051.635 1738.950 2056.235 ;
        RECT 1743.870 2051.635 1744.170 2056.235 ;
        RECT 1744.490 2051.635 1744.790 2056.235 ;
        RECT 1749.710 2051.635 1750.010 2056.235 ;
        RECT 1750.330 2051.635 1750.630 2056.235 ;
        RECT 1755.550 2051.635 1755.850 2056.235 ;
        RECT 1756.170 2051.635 1756.470 2056.235 ;
        RECT 1761.390 2051.635 1761.690 2056.235 ;
        RECT 1762.010 2051.635 1762.310 2056.235 ;
        RECT 1767.230 2051.635 1767.530 2056.235 ;
        RECT 1767.850 2051.635 1768.150 2056.235 ;
        RECT 1773.070 2051.635 1773.370 2056.235 ;
        RECT 1773.690 2051.635 1773.990 2056.235 ;
        RECT 1778.910 2051.635 1779.210 2056.235 ;
        RECT 1779.530 2051.635 1779.830 2056.235 ;
        RECT 1784.750 2051.635 1785.050 2056.235 ;
        RECT 1785.370 2051.635 1785.670 2056.235 ;
        RECT 1790.590 2051.635 1790.890 2056.235 ;
        RECT 1791.210 2051.635 1791.510 2056.235 ;
        RECT 1796.430 2051.635 1796.730 2056.235 ;
        RECT 1797.050 2051.635 1797.350 2056.235 ;
        RECT 1802.270 2051.635 1802.570 2056.235 ;
        RECT 1802.890 2051.635 1803.190 2056.235 ;
        RECT 1808.110 2051.635 1808.410 2056.235 ;
        RECT 1808.730 2051.635 1809.030 2056.235 ;
        RECT 1813.950 2051.635 1814.250 2056.235 ;
        RECT 1814.570 2051.635 1814.870 2056.235 ;
        RECT 1819.790 2051.635 1820.090 2056.235 ;
        RECT 1820.410 2051.635 1820.710 2056.235 ;
        RECT 1825.630 2051.635 1825.930 2056.235 ;
        RECT 1826.250 2051.635 1826.550 2056.235 ;
        RECT 1831.470 2051.635 1831.770 2056.235 ;
        RECT 1832.090 2051.635 1832.390 2056.235 ;
        RECT 1837.310 2051.635 1837.610 2056.235 ;
        RECT 1837.930 2051.635 1838.230 2056.235 ;
        RECT 1843.150 2051.635 1843.450 2056.235 ;
        RECT 1843.770 2051.635 1844.070 2056.235 ;
        RECT 1848.990 2051.635 1849.290 2056.235 ;
        RECT 1849.610 2051.635 1849.910 2056.235 ;
        RECT 1854.830 2051.635 1855.130 2056.235 ;
        RECT 1855.450 2051.635 1855.750 2056.235 ;
        RECT 1860.670 2051.635 1860.970 2056.235 ;
        RECT 1861.290 2051.635 1861.590 2056.235 ;
        RECT 1866.510 2051.635 1866.810 2056.235 ;
        RECT 1867.130 2051.635 1867.430 2056.235 ;
        RECT 1872.350 2051.635 1872.650 2056.235 ;
        RECT 1872.970 2051.635 1873.270 2056.235 ;
        RECT 1878.810 2051.635 1879.110 2056.235 ;
        RECT 1884.650 2051.635 1884.950 2056.235 ;
        RECT 1890.490 2051.635 1890.790 2056.235 ;
        RECT 1896.330 2051.635 1896.630 2056.235 ;
        RECT 1902.170 2051.635 1902.470 2056.235 ;
        RECT 2294.025 2051.635 2294.325 2056.235 ;
        RECT 2300.265 2051.635 2300.565 2056.235 ;
        RECT 2306.505 2051.635 2306.805 2056.235 ;
        RECT 2312.745 2051.635 2313.045 2056.235 ;
        RECT 2318.985 2051.635 2319.285 2056.235 ;
        RECT 2325.225 2051.635 2325.525 2056.235 ;
        RECT 2331.465 2051.635 2331.765 2056.235 ;
        RECT 2337.705 2051.635 2338.005 2056.235 ;
        RECT 2343.945 2051.635 2344.245 2056.235 ;
        RECT 2350.185 2051.635 2350.485 2056.235 ;
        RECT 2356.425 2051.635 2356.725 2056.235 ;
        RECT 2362.665 2051.635 2362.965 2056.235 ;
        RECT 2368.905 2051.635 2369.205 2056.235 ;
        RECT 2375.145 2051.635 2375.445 2056.235 ;
        RECT 2381.385 2051.635 2381.685 2056.235 ;
        RECT 2387.625 2051.635 2387.925 2056.235 ;
        RECT 2393.865 2051.635 2394.165 2056.235 ;
        RECT 2400.105 2051.635 2400.405 2056.235 ;
        RECT 2406.345 2051.635 2406.645 2056.235 ;
        RECT 2412.585 2051.635 2412.885 2056.235 ;
        RECT 2418.825 2051.635 2419.125 2056.235 ;
        RECT 2425.065 2051.635 2425.365 2056.235 ;
        RECT 2431.305 2051.635 2431.605 2056.235 ;
        RECT 2437.545 2051.635 2437.845 2056.235 ;
        RECT 2443.785 2051.635 2444.085 2056.235 ;
        RECT 2450.025 2051.635 2450.325 2056.235 ;
        RECT 2456.265 2051.635 2456.565 2056.235 ;
        RECT 2462.505 2051.635 2462.805 2056.235 ;
        RECT 2468.745 2051.635 2469.045 2056.235 ;
        RECT 2474.985 2051.635 2475.285 2056.235 ;
        RECT 2481.225 2051.635 2481.525 2056.235 ;
        RECT 2487.465 2051.635 2487.765 2056.235 ;
        RECT 2542.890 2051.635 2543.190 2056.235 ;
        RECT 1411.575 1614.495 1411.905 1614.825 ;
      LAYER met4 ;
        RECT 1555.000 1605.000 1931.480 2051.235 ;
        RECT 2205.000 1605.000 2581.480 2051.235 ;
      LAYER met4 ;
        RECT 1593.290 1600.000 1593.590 1604.600 ;
        RECT 1648.715 1600.000 1649.015 1604.600 ;
        RECT 1654.955 1600.000 1655.255 1604.600 ;
        RECT 1661.195 1600.000 1661.495 1604.600 ;
        RECT 1667.435 1600.000 1667.735 1604.600 ;
        RECT 1673.675 1600.000 1673.975 1604.600 ;
        RECT 1679.915 1600.000 1680.215 1604.600 ;
        RECT 1686.155 1600.000 1686.455 1604.600 ;
        RECT 1692.395 1600.000 1692.695 1604.600 ;
        RECT 1698.635 1600.000 1698.935 1604.600 ;
        RECT 1704.875 1600.000 1705.175 1604.600 ;
        RECT 1711.115 1600.000 1711.415 1604.600 ;
        RECT 1717.355 1600.000 1717.655 1604.600 ;
        RECT 1723.595 1600.000 1723.895 1604.600 ;
        RECT 1729.835 1600.000 1730.135 1604.600 ;
        RECT 1736.075 1600.000 1736.375 1604.600 ;
        RECT 1742.315 1600.000 1742.615 1604.600 ;
        RECT 1748.555 1600.000 1748.855 1604.600 ;
        RECT 1754.795 1600.000 1755.095 1604.600 ;
        RECT 1761.035 1600.000 1761.335 1604.600 ;
        RECT 1767.275 1600.000 1767.575 1604.600 ;
        RECT 1773.515 1600.000 1773.815 1604.600 ;
        RECT 1779.755 1600.000 1780.055 1604.600 ;
        RECT 1785.995 1600.000 1786.295 1604.600 ;
        RECT 1792.235 1600.000 1792.535 1604.600 ;
        RECT 1798.475 1600.000 1798.775 1604.600 ;
        RECT 1804.715 1600.000 1805.015 1604.600 ;
        RECT 1810.955 1600.000 1811.255 1604.600 ;
        RECT 1817.195 1600.000 1817.495 1604.600 ;
        RECT 1823.435 1600.000 1823.735 1604.600 ;
        RECT 1829.675 1600.000 1829.975 1604.600 ;
        RECT 1835.915 1600.000 1836.215 1604.600 ;
        RECT 1842.155 1600.000 1842.455 1604.600 ;
        RECT 2234.010 1600.000 2234.310 1604.600 ;
        RECT 2239.850 1600.000 2240.150 1604.600 ;
        RECT 2245.690 1600.000 2245.990 1604.600 ;
        RECT 2251.530 1600.000 2251.830 1604.600 ;
        RECT 2257.370 1600.000 2257.670 1604.600 ;
        RECT 2263.210 1600.000 2263.510 1604.600 ;
        RECT 2263.830 1600.000 2264.130 1604.600 ;
        RECT 2269.050 1600.000 2269.350 1604.600 ;
        RECT 2269.670 1600.000 2269.970 1604.600 ;
        RECT 2274.890 1600.000 2275.190 1604.600 ;
        RECT 2275.510 1600.000 2275.810 1604.600 ;
        RECT 2280.730 1600.000 2281.030 1604.600 ;
        RECT 2281.350 1600.000 2281.650 1604.600 ;
        RECT 2286.570 1600.000 2286.870 1604.600 ;
        RECT 2287.190 1600.000 2287.490 1604.600 ;
        RECT 2292.410 1600.000 2292.710 1604.600 ;
        RECT 2293.030 1600.000 2293.330 1604.600 ;
        RECT 2298.250 1600.000 2298.550 1604.600 ;
        RECT 2298.870 1600.000 2299.170 1604.600 ;
        RECT 2304.090 1600.000 2304.390 1604.600 ;
        RECT 2304.710 1600.000 2305.010 1604.600 ;
        RECT 2309.930 1600.000 2310.230 1604.600 ;
        RECT 2310.550 1600.000 2310.850 1604.600 ;
        RECT 2315.770 1600.000 2316.070 1604.600 ;
        RECT 2316.390 1600.000 2316.690 1604.600 ;
        RECT 2321.610 1600.000 2321.910 1604.600 ;
        RECT 2322.230 1600.000 2322.530 1604.600 ;
        RECT 2327.450 1600.000 2327.750 1604.600 ;
        RECT 2328.070 1600.000 2328.370 1604.600 ;
        RECT 2333.290 1600.000 2333.590 1604.600 ;
        RECT 2333.910 1600.000 2334.210 1604.600 ;
        RECT 2339.130 1600.000 2339.430 1604.600 ;
        RECT 2339.750 1600.000 2340.050 1604.600 ;
        RECT 2344.970 1600.000 2345.270 1604.600 ;
        RECT 2345.590 1600.000 2345.890 1604.600 ;
        RECT 2350.810 1600.000 2351.110 1604.600 ;
        RECT 2351.430 1600.000 2351.730 1604.600 ;
        RECT 2356.650 1600.000 2356.950 1604.600 ;
        RECT 2357.270 1600.000 2357.570 1604.600 ;
        RECT 2362.490 1600.000 2362.790 1604.600 ;
        RECT 2363.110 1600.000 2363.410 1604.600 ;
        RECT 2368.330 1600.000 2368.630 1604.600 ;
        RECT 2368.950 1600.000 2369.250 1604.600 ;
        RECT 2374.170 1600.000 2374.470 1604.600 ;
        RECT 2374.790 1600.000 2375.090 1604.600 ;
        RECT 2380.010 1600.000 2380.310 1604.600 ;
        RECT 2380.630 1600.000 2380.930 1604.600 ;
        RECT 2385.850 1600.000 2386.150 1604.600 ;
        RECT 2386.470 1600.000 2386.770 1604.600 ;
        RECT 2391.690 1600.000 2391.990 1604.600 ;
        RECT 2392.310 1600.000 2392.610 1604.600 ;
        RECT 2397.530 1600.000 2397.830 1604.600 ;
        RECT 2398.150 1600.000 2398.450 1604.600 ;
        RECT 2403.370 1600.000 2403.670 1604.600 ;
        RECT 2403.990 1600.000 2404.290 1604.600 ;
        RECT 2409.210 1600.000 2409.510 1604.600 ;
        RECT 2409.830 1600.000 2410.130 1604.600 ;
        RECT 2415.050 1600.000 2415.350 1604.600 ;
        RECT 2415.670 1600.000 2415.970 1604.600 ;
        RECT 2420.890 1600.000 2421.190 1604.600 ;
        RECT 2421.510 1600.000 2421.810 1604.600 ;
        RECT 2426.730 1600.000 2427.030 1604.600 ;
        RECT 2427.350 1600.000 2427.650 1604.600 ;
        RECT 2432.570 1600.000 2432.870 1604.600 ;
        RECT 2433.190 1600.000 2433.490 1604.600 ;
        RECT 2438.410 1600.000 2438.710 1604.600 ;
        RECT 2439.030 1600.000 2439.330 1604.600 ;
        RECT 2444.250 1600.000 2444.550 1604.600 ;
        RECT 2444.870 1600.000 2445.170 1604.600 ;
        RECT 1588.020 1515.000 1591.020 1585.000 ;
        RECT 1624.020 1515.000 1627.020 1585.000 ;
        RECT 1642.020 1515.000 1645.020 1585.000 ;
        RECT 1660.020 1515.000 1663.020 1585.000 ;
        RECT 1678.020 1515.000 1681.020 1585.000 ;
        RECT 1768.020 1515.000 1771.020 1585.000 ;
        RECT 1804.020 1515.000 1807.020 1585.000 ;
        RECT 1822.020 1515.000 1825.020 1585.000 ;
        RECT 1840.020 1515.000 1843.020 1585.000 ;
        RECT 1858.020 1515.000 1861.020 1585.000 ;
        RECT 1948.020 1515.000 1951.020 1585.000 ;
        RECT 2182.020 1515.000 2185.020 1585.000 ;
        RECT 2200.020 1515.000 2203.020 1585.000 ;
        RECT 2218.020 1515.000 2221.020 1585.000 ;
        RECT 2308.020 1515.000 2311.020 1585.000 ;
        RECT 2344.020 1515.000 2347.020 1585.000 ;
        RECT 2362.020 1515.000 2365.020 1585.000 ;
        RECT 2380.020 1515.000 2383.020 1585.000 ;
        RECT 2398.020 1515.000 2401.020 1585.000 ;
        RECT 2488.020 1515.000 2491.020 1585.000 ;
        RECT 2524.020 1515.000 2527.020 1585.000 ;
        RECT 2542.020 1515.000 2545.020 1585.000 ;
        RECT 2560.020 1515.000 2563.020 1585.000 ;
        RECT 2578.020 1515.000 2581.020 1585.000 ;
      LAYER met4 ;
        RECT 1616.465 410.640 1647.370 1488.240 ;
        RECT 1649.770 410.640 2637.995 1488.240 ;
      LAYER met5 ;
        RECT 1412.780 2935.100 1938.780 2936.700 ;
        RECT 2199.380 2897.700 2595.660 2899.300 ;
        RECT 302.340 2894.300 688.500 2895.900 ;
        RECT 950.020 2894.300 1346.300 2895.900 ;
  END
END user_project_wrapper
END LIBRARY

