VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2433.460 2924.800 2434.660 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2903.340 2924.800 2904.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3410.620 2.400 3411.820 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 2.400 3124.860 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2836.020 2.400 2837.220 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 2.400 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 2.400 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1974.460 2.400 1975.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 2.400 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 2.400 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 2.400 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 2.400 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 2.400 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 2.400 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 2.400 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 2.400 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1964.260 2924.800 1965.460 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2198.860 2924.800 2200.060 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 2.400 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 2.400 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 2.400 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 2.400 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 2.400 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 2.400 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 2.400 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 2.400 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 2.400 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 2.400 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 2.400 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 2.400 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.220 2.400 3340.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 2.400 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 2.400 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2476.980 2.400 2478.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 2.400 2190.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 2.400 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 2.400 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 2.400 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 2.400 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 2.400 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 2.400 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 2.400 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 2.400 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 616.085 17.765 618.095 17.935 ;
      LAYER mcon ;
        RECT 617.925 17.765 618.095 17.935 ;
      LAYER met1 ;
        RECT 569.550 1590.420 569.870 1590.480 ;
        RECT 571.850 1590.420 572.170 1590.480 ;
        RECT 569.550 1590.280 572.170 1590.420 ;
        RECT 569.550 1590.220 569.870 1590.280 ;
        RECT 571.850 1590.220 572.170 1590.280 ;
        RECT 616.025 17.920 616.315 17.965 ;
        RECT 591.720 17.780 616.315 17.920 ;
        RECT 571.850 16.900 572.170 16.960 ;
        RECT 591.720 16.900 591.860 17.780 ;
        RECT 616.025 17.735 616.315 17.780 ;
        RECT 617.865 17.920 618.155 17.965 ;
        RECT 633.030 17.920 633.350 17.980 ;
        RECT 617.865 17.780 633.350 17.920 ;
        RECT 617.865 17.735 618.155 17.780 ;
        RECT 633.030 17.720 633.350 17.780 ;
        RECT 571.850 16.760 591.860 16.900 ;
        RECT 571.850 16.700 572.170 16.760 ;
      LAYER via ;
        RECT 569.580 1590.220 569.840 1590.480 ;
        RECT 571.880 1590.220 572.140 1590.480 ;
        RECT 571.880 16.700 572.140 16.960 ;
        RECT 633.060 17.720 633.320 17.980 ;
      LAYER met2 ;
        RECT 569.440 1600.380 569.720 1604.000 ;
        RECT 569.440 1600.000 569.780 1600.380 ;
        RECT 569.640 1590.510 569.780 1600.000 ;
        RECT 569.580 1590.190 569.840 1590.510 ;
        RECT 571.880 1590.190 572.140 1590.510 ;
        RECT 571.940 16.990 572.080 1590.190 ;
        RECT 633.060 17.690 633.320 18.010 ;
        RECT 571.880 16.670 572.140 16.990 ;
        RECT 633.120 2.400 633.260 17.690 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.870 1535.340 1187.190 1535.400 ;
        RECT 1193.310 1535.340 1193.630 1535.400 ;
        RECT 1186.870 1535.200 1193.630 1535.340 ;
        RECT 1186.870 1535.140 1187.190 1535.200 ;
        RECT 1193.310 1535.140 1193.630 1535.200 ;
        RECT 1193.310 62.800 1193.630 62.860 ;
        RECT 2415.070 62.800 2415.390 62.860 ;
        RECT 1193.310 62.660 2415.390 62.800 ;
        RECT 1193.310 62.600 1193.630 62.660 ;
        RECT 2415.070 62.600 2415.390 62.660 ;
      LAYER via ;
        RECT 1186.900 1535.140 1187.160 1535.400 ;
        RECT 1193.340 1535.140 1193.600 1535.400 ;
        RECT 1193.340 62.600 1193.600 62.860 ;
        RECT 2415.100 62.600 2415.360 62.860 ;
      LAYER met2 ;
        RECT 1187.680 1600.450 1187.960 1604.000 ;
        RECT 1186.960 1600.310 1187.960 1600.450 ;
        RECT 1186.960 1535.430 1187.100 1600.310 ;
        RECT 1187.680 1600.000 1187.960 1600.310 ;
        RECT 1186.900 1535.110 1187.160 1535.430 ;
        RECT 1193.340 1535.110 1193.600 1535.430 ;
        RECT 1193.400 62.890 1193.540 1535.110 ;
        RECT 1193.340 62.570 1193.600 62.890 ;
        RECT 2415.100 62.570 2415.360 62.890 ;
        RECT 2415.160 17.410 2415.300 62.570 ;
        RECT 2415.160 17.270 2417.600 17.410 ;
        RECT 2417.460 2.400 2417.600 17.270 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1194.230 1580.900 1194.550 1580.960 ;
        RECT 1199.750 1580.900 1200.070 1580.960 ;
        RECT 1194.230 1580.760 1200.070 1580.900 ;
        RECT 1194.230 1580.700 1194.550 1580.760 ;
        RECT 1199.750 1580.700 1200.070 1580.760 ;
        RECT 1199.750 63.140 1200.070 63.200 ;
        RECT 2429.330 63.140 2429.650 63.200 ;
        RECT 1199.750 63.000 2429.650 63.140 ;
        RECT 1199.750 62.940 1200.070 63.000 ;
        RECT 2429.330 62.940 2429.650 63.000 ;
      LAYER via ;
        RECT 1194.260 1580.700 1194.520 1580.960 ;
        RECT 1199.780 1580.700 1200.040 1580.960 ;
        RECT 1199.780 62.940 1200.040 63.200 ;
        RECT 2429.360 62.940 2429.620 63.200 ;
      LAYER met2 ;
        RECT 1193.660 1600.450 1193.940 1604.000 ;
        RECT 1193.660 1600.310 1194.460 1600.450 ;
        RECT 1193.660 1600.000 1193.940 1600.310 ;
        RECT 1194.320 1580.990 1194.460 1600.310 ;
        RECT 1194.260 1580.670 1194.520 1580.990 ;
        RECT 1199.780 1580.670 1200.040 1580.990 ;
        RECT 1199.840 63.230 1199.980 1580.670 ;
        RECT 1199.780 62.910 1200.040 63.230 ;
        RECT 2429.360 62.910 2429.620 63.230 ;
        RECT 2429.420 17.410 2429.560 62.910 ;
        RECT 2429.420 17.270 2435.080 17.410 ;
        RECT 2434.940 2.400 2435.080 17.270 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1194.230 1580.220 1194.550 1580.280 ;
        RECT 1198.830 1580.220 1199.150 1580.280 ;
        RECT 1194.230 1580.080 1199.150 1580.220 ;
        RECT 1194.230 1580.020 1194.550 1580.080 ;
        RECT 1198.830 1580.020 1199.150 1580.080 ;
        RECT 1194.230 1535.340 1194.550 1535.400 ;
        RECT 1199.290 1535.340 1199.610 1535.400 ;
        RECT 1194.230 1535.200 1199.610 1535.340 ;
        RECT 1194.230 1535.140 1194.550 1535.200 ;
        RECT 1199.290 1535.140 1199.610 1535.200 ;
        RECT 2449.570 2.960 2449.890 3.020 ;
        RECT 2452.790 2.960 2453.110 3.020 ;
        RECT 2449.570 2.820 2453.110 2.960 ;
        RECT 2449.570 2.760 2449.890 2.820 ;
        RECT 2452.790 2.760 2453.110 2.820 ;
      LAYER via ;
        RECT 1194.260 1580.020 1194.520 1580.280 ;
        RECT 1198.860 1580.020 1199.120 1580.280 ;
        RECT 1194.260 1535.140 1194.520 1535.400 ;
        RECT 1199.320 1535.140 1199.580 1535.400 ;
        RECT 2449.600 2.760 2449.860 3.020 ;
        RECT 2452.820 2.760 2453.080 3.020 ;
      LAYER met2 ;
        RECT 1200.100 1600.450 1200.380 1604.000 ;
        RECT 1198.920 1600.310 1200.380 1600.450 ;
        RECT 1198.920 1580.310 1199.060 1600.310 ;
        RECT 1200.100 1600.000 1200.380 1600.310 ;
        RECT 1194.260 1579.990 1194.520 1580.310 ;
        RECT 1198.860 1579.990 1199.120 1580.310 ;
        RECT 1194.320 1535.430 1194.460 1579.990 ;
        RECT 1194.260 1535.110 1194.520 1535.430 ;
        RECT 1199.320 1535.110 1199.580 1535.430 ;
        RECT 1199.380 76.005 1199.520 1535.110 ;
        RECT 1199.310 75.635 1199.590 76.005 ;
        RECT 1283.490 75.635 1283.770 76.005 ;
        RECT 2449.590 75.635 2449.870 76.005 ;
        RECT 1283.560 73.965 1283.700 75.635 ;
        RECT 1283.490 73.595 1283.770 73.965 ;
        RECT 2449.660 3.050 2449.800 75.635 ;
        RECT 2449.600 2.730 2449.860 3.050 ;
        RECT 2452.820 2.730 2453.080 3.050 ;
        RECT 2452.880 2.400 2453.020 2.730 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
      LAYER via2 ;
        RECT 1199.310 75.680 1199.590 75.960 ;
        RECT 1283.490 75.680 1283.770 75.960 ;
        RECT 2449.590 75.680 2449.870 75.960 ;
        RECT 1283.490 73.640 1283.770 73.920 ;
      LAYER met3 ;
        RECT 1199.285 75.970 1199.615 75.985 ;
        RECT 1283.465 75.970 1283.795 75.985 ;
        RECT 1199.285 75.670 1283.795 75.970 ;
        RECT 1199.285 75.655 1199.615 75.670 ;
        RECT 1283.465 75.655 1283.795 75.670 ;
        RECT 1331.280 75.970 1331.660 75.980 ;
        RECT 2449.565 75.970 2449.895 75.985 ;
        RECT 1331.280 75.670 2449.895 75.970 ;
        RECT 1331.280 75.660 1331.660 75.670 ;
        RECT 2449.565 75.655 2449.895 75.670 ;
        RECT 1283.465 73.930 1283.795 73.945 ;
        RECT 1331.280 73.930 1331.660 73.940 ;
        RECT 1283.465 73.630 1331.660 73.930 ;
        RECT 1283.465 73.615 1283.795 73.630 ;
        RECT 1331.280 73.620 1331.660 73.630 ;
      LAYER via3 ;
        RECT 1331.310 75.660 1331.630 75.980 ;
        RECT 1331.310 73.620 1331.630 73.940 ;
      LAYER met4 ;
        RECT 1331.305 75.655 1331.635 75.985 ;
        RECT 1331.320 73.945 1331.620 75.655 ;
        RECT 1331.305 73.615 1331.635 73.945 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1207.185 20.825 1207.355 34.595 ;
      LAYER mcon ;
        RECT 1207.185 34.425 1207.355 34.595 ;
      LAYER met1 ;
        RECT 1200.670 1579.880 1200.990 1579.940 ;
        RECT 1204.810 1579.880 1205.130 1579.940 ;
        RECT 1200.670 1579.740 1205.130 1579.880 ;
        RECT 1200.670 1579.680 1200.990 1579.740 ;
        RECT 1204.810 1579.680 1205.130 1579.740 ;
        RECT 1200.670 1535.340 1200.990 1535.400 ;
        RECT 1207.110 1535.340 1207.430 1535.400 ;
        RECT 1200.670 1535.200 1207.430 1535.340 ;
        RECT 1200.670 1535.140 1200.990 1535.200 ;
        RECT 1207.110 1535.140 1207.430 1535.200 ;
        RECT 1207.110 34.580 1207.430 34.640 ;
        RECT 1206.915 34.440 1207.430 34.580 ;
        RECT 1207.110 34.380 1207.430 34.440 ;
        RECT 1207.125 20.980 1207.415 21.025 ;
        RECT 2470.730 20.980 2471.050 21.040 ;
        RECT 1207.125 20.840 2471.050 20.980 ;
        RECT 1207.125 20.795 1207.415 20.840 ;
        RECT 2470.730 20.780 2471.050 20.840 ;
      LAYER via ;
        RECT 1200.700 1579.680 1200.960 1579.940 ;
        RECT 1204.840 1579.680 1205.100 1579.940 ;
        RECT 1200.700 1535.140 1200.960 1535.400 ;
        RECT 1207.140 1535.140 1207.400 1535.400 ;
        RECT 1207.140 34.380 1207.400 34.640 ;
        RECT 2470.760 20.780 2471.020 21.040 ;
      LAYER met2 ;
        RECT 1206.080 1600.450 1206.360 1604.000 ;
        RECT 1204.900 1600.310 1206.360 1600.450 ;
        RECT 1204.900 1579.970 1205.040 1600.310 ;
        RECT 1206.080 1600.000 1206.360 1600.310 ;
        RECT 1200.700 1579.650 1200.960 1579.970 ;
        RECT 1204.840 1579.650 1205.100 1579.970 ;
        RECT 1200.760 1535.430 1200.900 1579.650 ;
        RECT 1200.700 1535.110 1200.960 1535.430 ;
        RECT 1207.140 1535.110 1207.400 1535.430 ;
        RECT 1207.200 34.670 1207.340 1535.110 ;
        RECT 1207.140 34.350 1207.400 34.670 ;
        RECT 2470.760 20.750 2471.020 21.070 ;
        RECT 2470.820 2.400 2470.960 20.750 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1244.445 21.165 1244.615 25.415 ;
      LAYER mcon ;
        RECT 1244.445 25.245 1244.615 25.415 ;
      LAYER met1 ;
        RECT 1207.570 1579.880 1207.890 1579.940 ;
        RECT 1210.790 1579.880 1211.110 1579.940 ;
        RECT 1207.570 1579.740 1211.110 1579.880 ;
        RECT 1207.570 1579.680 1207.890 1579.740 ;
        RECT 1210.790 1579.680 1211.110 1579.740 ;
        RECT 1207.570 1535.340 1207.890 1535.400 ;
        RECT 1214.010 1535.340 1214.330 1535.400 ;
        RECT 1207.570 1535.200 1214.330 1535.340 ;
        RECT 1207.570 1535.140 1207.890 1535.200 ;
        RECT 1214.010 1535.140 1214.330 1535.200 ;
        RECT 1214.010 25.400 1214.330 25.460 ;
        RECT 1244.385 25.400 1244.675 25.445 ;
        RECT 1214.010 25.260 1244.675 25.400 ;
        RECT 1214.010 25.200 1214.330 25.260 ;
        RECT 1244.385 25.215 1244.675 25.260 ;
        RECT 1244.385 21.320 1244.675 21.365 ;
        RECT 2488.670 21.320 2488.990 21.380 ;
        RECT 1244.385 21.180 2488.990 21.320 ;
        RECT 1244.385 21.135 1244.675 21.180 ;
        RECT 2488.670 21.120 2488.990 21.180 ;
      LAYER via ;
        RECT 1207.600 1579.680 1207.860 1579.940 ;
        RECT 1210.820 1579.680 1211.080 1579.940 ;
        RECT 1207.600 1535.140 1207.860 1535.400 ;
        RECT 1214.040 1535.140 1214.300 1535.400 ;
        RECT 1214.040 25.200 1214.300 25.460 ;
        RECT 2488.700 21.120 2488.960 21.380 ;
      LAYER met2 ;
        RECT 1212.520 1600.450 1212.800 1604.000 ;
        RECT 1210.880 1600.310 1212.800 1600.450 ;
        RECT 1210.880 1579.970 1211.020 1600.310 ;
        RECT 1212.520 1600.000 1212.800 1600.310 ;
        RECT 1207.600 1579.650 1207.860 1579.970 ;
        RECT 1210.820 1579.650 1211.080 1579.970 ;
        RECT 1207.660 1535.430 1207.800 1579.650 ;
        RECT 1207.600 1535.110 1207.860 1535.430 ;
        RECT 1214.040 1535.110 1214.300 1535.430 ;
        RECT 1214.100 25.490 1214.240 1535.110 ;
        RECT 1214.040 25.170 1214.300 25.490 ;
        RECT 2488.700 21.090 2488.960 21.410 ;
        RECT 2488.760 2.400 2488.900 21.090 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1246.745 21.505 1246.915 25.075 ;
      LAYER mcon ;
        RECT 1246.745 24.905 1246.915 25.075 ;
      LAYER met1 ;
        RECT 1220.910 25.060 1221.230 25.120 ;
        RECT 1246.685 25.060 1246.975 25.105 ;
        RECT 1220.910 24.920 1246.975 25.060 ;
        RECT 1220.910 24.860 1221.230 24.920 ;
        RECT 1246.685 24.875 1246.975 24.920 ;
        RECT 1246.685 21.660 1246.975 21.705 ;
        RECT 2506.150 21.660 2506.470 21.720 ;
        RECT 1246.685 21.520 2506.470 21.660 ;
        RECT 1246.685 21.475 1246.975 21.520 ;
        RECT 2506.150 21.460 2506.470 21.520 ;
      LAYER via ;
        RECT 1220.940 24.860 1221.200 25.120 ;
        RECT 2506.180 21.460 2506.440 21.720 ;
      LAYER met2 ;
        RECT 1218.500 1600.450 1218.780 1604.000 ;
        RECT 1218.500 1600.310 1220.220 1600.450 ;
        RECT 1218.500 1600.000 1218.780 1600.310 ;
        RECT 1220.080 1580.050 1220.220 1600.310 ;
        RECT 1220.080 1579.910 1221.140 1580.050 ;
        RECT 1221.000 25.150 1221.140 1579.910 ;
        RECT 1220.940 24.830 1221.200 25.150 ;
        RECT 2506.180 21.430 2506.440 21.750 ;
        RECT 2506.240 2.400 2506.380 21.430 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1227.885 1497.445 1228.055 1545.555 ;
        RECT 1247.205 21.845 1247.375 27.455 ;
      LAYER mcon ;
        RECT 1227.885 1545.385 1228.055 1545.555 ;
        RECT 1247.205 27.285 1247.375 27.455 ;
      LAYER met1 ;
        RECT 1225.050 1594.160 1225.370 1594.220 ;
        RECT 1227.810 1594.160 1228.130 1594.220 ;
        RECT 1225.050 1594.020 1228.130 1594.160 ;
        RECT 1225.050 1593.960 1225.370 1594.020 ;
        RECT 1227.810 1593.960 1228.130 1594.020 ;
        RECT 1227.810 1545.540 1228.130 1545.600 ;
        RECT 1227.615 1545.400 1228.130 1545.540 ;
        RECT 1227.810 1545.340 1228.130 1545.400 ;
        RECT 1227.810 1497.600 1228.130 1497.660 ;
        RECT 1227.615 1497.460 1228.130 1497.600 ;
        RECT 1227.810 1497.400 1228.130 1497.460 ;
        RECT 1226.430 96.460 1226.750 96.520 ;
        RECT 1227.810 96.460 1228.130 96.520 ;
        RECT 1226.430 96.320 1228.130 96.460 ;
        RECT 1226.430 96.260 1226.750 96.320 ;
        RECT 1227.810 96.260 1228.130 96.320 ;
        RECT 1226.890 27.440 1227.210 27.500 ;
        RECT 1247.145 27.440 1247.435 27.485 ;
        RECT 1226.890 27.300 1247.435 27.440 ;
        RECT 1226.890 27.240 1227.210 27.300 ;
        RECT 1247.145 27.255 1247.435 27.300 ;
        RECT 1247.145 22.000 1247.435 22.045 ;
        RECT 2524.090 22.000 2524.410 22.060 ;
        RECT 1247.145 21.860 2524.410 22.000 ;
        RECT 1247.145 21.815 1247.435 21.860 ;
        RECT 2524.090 21.800 2524.410 21.860 ;
      LAYER via ;
        RECT 1225.080 1593.960 1225.340 1594.220 ;
        RECT 1227.840 1593.960 1228.100 1594.220 ;
        RECT 1227.840 1545.340 1228.100 1545.600 ;
        RECT 1227.840 1497.400 1228.100 1497.660 ;
        RECT 1226.460 96.260 1226.720 96.520 ;
        RECT 1227.840 96.260 1228.100 96.520 ;
        RECT 1226.920 27.240 1227.180 27.500 ;
        RECT 2524.120 21.800 2524.380 22.060 ;
      LAYER met2 ;
        RECT 1224.940 1600.380 1225.220 1604.000 ;
        RECT 1224.940 1600.000 1225.280 1600.380 ;
        RECT 1225.140 1594.250 1225.280 1600.000 ;
        RECT 1225.080 1593.930 1225.340 1594.250 ;
        RECT 1227.840 1593.930 1228.100 1594.250 ;
        RECT 1227.900 1545.630 1228.040 1593.930 ;
        RECT 1227.840 1545.310 1228.100 1545.630 ;
        RECT 1227.840 1497.370 1228.100 1497.690 ;
        RECT 1227.900 96.550 1228.040 1497.370 ;
        RECT 1226.460 96.230 1226.720 96.550 ;
        RECT 1227.840 96.230 1228.100 96.550 ;
        RECT 1226.520 64.330 1226.660 96.230 ;
        RECT 1226.520 64.190 1227.120 64.330 ;
        RECT 1226.980 27.530 1227.120 64.190 ;
        RECT 1226.920 27.210 1227.180 27.530 ;
        RECT 2524.120 21.770 2524.380 22.090 ;
        RECT 2524.180 2.400 2524.320 21.770 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1234.785 1442.025 1234.955 1490.475 ;
        RECT 1234.785 476.085 1234.955 524.195 ;
        RECT 1234.785 379.525 1234.955 427.635 ;
        RECT 1234.785 282.965 1234.955 331.075 ;
        RECT 1234.785 186.405 1234.955 234.515 ;
      LAYER mcon ;
        RECT 1234.785 1490.305 1234.955 1490.475 ;
        RECT 1234.785 524.025 1234.955 524.195 ;
        RECT 1234.785 427.465 1234.955 427.635 ;
        RECT 1234.785 330.905 1234.955 331.075 ;
        RECT 1234.785 234.345 1234.955 234.515 ;
      LAYER met1 ;
        RECT 1232.410 1576.140 1232.730 1576.200 ;
        RECT 1234.710 1576.140 1235.030 1576.200 ;
        RECT 1232.410 1576.000 1235.030 1576.140 ;
        RECT 1232.410 1575.940 1232.730 1576.000 ;
        RECT 1234.710 1575.940 1235.030 1576.000 ;
        RECT 1234.710 1490.460 1235.030 1490.520 ;
        RECT 1234.515 1490.320 1235.030 1490.460 ;
        RECT 1234.710 1490.260 1235.030 1490.320 ;
        RECT 1234.710 1442.180 1235.030 1442.240 ;
        RECT 1234.515 1442.040 1235.030 1442.180 ;
        RECT 1234.710 1441.980 1235.030 1442.040 ;
        RECT 1234.710 1249.060 1235.030 1249.120 ;
        RECT 1235.630 1249.060 1235.950 1249.120 ;
        RECT 1234.710 1248.920 1235.950 1249.060 ;
        RECT 1234.710 1248.860 1235.030 1248.920 ;
        RECT 1235.630 1248.860 1235.950 1248.920 ;
        RECT 1234.710 1152.500 1235.030 1152.560 ;
        RECT 1235.630 1152.500 1235.950 1152.560 ;
        RECT 1234.710 1152.360 1235.950 1152.500 ;
        RECT 1234.710 1152.300 1235.030 1152.360 ;
        RECT 1235.630 1152.300 1235.950 1152.360 ;
        RECT 1234.710 1007.320 1235.030 1007.380 ;
        RECT 1235.630 1007.320 1235.950 1007.380 ;
        RECT 1234.710 1007.180 1235.950 1007.320 ;
        RECT 1234.710 1007.120 1235.030 1007.180 ;
        RECT 1235.630 1007.120 1235.950 1007.180 ;
        RECT 1234.710 910.760 1235.030 910.820 ;
        RECT 1235.630 910.760 1235.950 910.820 ;
        RECT 1234.710 910.620 1235.950 910.760 ;
        RECT 1234.710 910.560 1235.030 910.620 ;
        RECT 1235.630 910.560 1235.950 910.620 ;
        RECT 1234.710 717.640 1235.030 717.700 ;
        RECT 1235.630 717.640 1235.950 717.700 ;
        RECT 1234.710 717.500 1235.950 717.640 ;
        RECT 1234.710 717.440 1235.030 717.500 ;
        RECT 1235.630 717.440 1235.950 717.500 ;
        RECT 1234.710 524.180 1235.030 524.240 ;
        RECT 1234.515 524.040 1235.030 524.180 ;
        RECT 1234.710 523.980 1235.030 524.040 ;
        RECT 1234.710 476.240 1235.030 476.300 ;
        RECT 1234.515 476.100 1235.030 476.240 ;
        RECT 1234.710 476.040 1235.030 476.100 ;
        RECT 1234.710 427.620 1235.030 427.680 ;
        RECT 1234.515 427.480 1235.030 427.620 ;
        RECT 1234.710 427.420 1235.030 427.480 ;
        RECT 1234.710 379.680 1235.030 379.740 ;
        RECT 1234.515 379.540 1235.030 379.680 ;
        RECT 1234.710 379.480 1235.030 379.540 ;
        RECT 1234.710 331.060 1235.030 331.120 ;
        RECT 1234.515 330.920 1235.030 331.060 ;
        RECT 1234.710 330.860 1235.030 330.920 ;
        RECT 1234.710 283.120 1235.030 283.180 ;
        RECT 1234.515 282.980 1235.030 283.120 ;
        RECT 1234.710 282.920 1235.030 282.980 ;
        RECT 1234.710 234.500 1235.030 234.560 ;
        RECT 1234.515 234.360 1235.030 234.500 ;
        RECT 1234.710 234.300 1235.030 234.360 ;
        RECT 1234.710 186.560 1235.030 186.620 ;
        RECT 1234.515 186.420 1235.030 186.560 ;
        RECT 1234.710 186.360 1235.030 186.420 ;
        RECT 1246.210 22.340 1246.530 22.400 ;
        RECT 2542.030 22.340 2542.350 22.400 ;
        RECT 1246.210 22.200 2542.350 22.340 ;
        RECT 1246.210 22.140 1246.530 22.200 ;
        RECT 2542.030 22.140 2542.350 22.200 ;
      LAYER via ;
        RECT 1232.440 1575.940 1232.700 1576.200 ;
        RECT 1234.740 1575.940 1235.000 1576.200 ;
        RECT 1234.740 1490.260 1235.000 1490.520 ;
        RECT 1234.740 1441.980 1235.000 1442.240 ;
        RECT 1234.740 1248.860 1235.000 1249.120 ;
        RECT 1235.660 1248.860 1235.920 1249.120 ;
        RECT 1234.740 1152.300 1235.000 1152.560 ;
        RECT 1235.660 1152.300 1235.920 1152.560 ;
        RECT 1234.740 1007.120 1235.000 1007.380 ;
        RECT 1235.660 1007.120 1235.920 1007.380 ;
        RECT 1234.740 910.560 1235.000 910.820 ;
        RECT 1235.660 910.560 1235.920 910.820 ;
        RECT 1234.740 717.440 1235.000 717.700 ;
        RECT 1235.660 717.440 1235.920 717.700 ;
        RECT 1234.740 523.980 1235.000 524.240 ;
        RECT 1234.740 476.040 1235.000 476.300 ;
        RECT 1234.740 427.420 1235.000 427.680 ;
        RECT 1234.740 379.480 1235.000 379.740 ;
        RECT 1234.740 330.860 1235.000 331.120 ;
        RECT 1234.740 282.920 1235.000 283.180 ;
        RECT 1234.740 234.300 1235.000 234.560 ;
        RECT 1234.740 186.360 1235.000 186.620 ;
        RECT 1246.240 22.140 1246.500 22.400 ;
        RECT 2542.060 22.140 2542.320 22.400 ;
      LAYER met2 ;
        RECT 1230.920 1600.450 1231.200 1604.000 ;
        RECT 1230.920 1600.310 1232.640 1600.450 ;
        RECT 1230.920 1600.000 1231.200 1600.310 ;
        RECT 1232.500 1576.230 1232.640 1600.310 ;
        RECT 1232.440 1575.910 1232.700 1576.230 ;
        RECT 1234.740 1575.910 1235.000 1576.230 ;
        RECT 1234.800 1490.550 1234.940 1575.910 ;
        RECT 1234.740 1490.230 1235.000 1490.550 ;
        RECT 1234.740 1441.950 1235.000 1442.270 ;
        RECT 1234.800 1297.285 1234.940 1441.950 ;
        RECT 1234.730 1296.915 1235.010 1297.285 ;
        RECT 1235.650 1296.915 1235.930 1297.285 ;
        RECT 1235.720 1249.150 1235.860 1296.915 ;
        RECT 1234.740 1248.830 1235.000 1249.150 ;
        RECT 1235.660 1248.830 1235.920 1249.150 ;
        RECT 1234.800 1200.725 1234.940 1248.830 ;
        RECT 1234.730 1200.355 1235.010 1200.725 ;
        RECT 1235.650 1200.355 1235.930 1200.725 ;
        RECT 1235.720 1152.590 1235.860 1200.355 ;
        RECT 1234.740 1152.270 1235.000 1152.590 ;
        RECT 1235.660 1152.270 1235.920 1152.590 ;
        RECT 1234.800 1104.165 1234.940 1152.270 ;
        RECT 1234.730 1103.795 1235.010 1104.165 ;
        RECT 1235.650 1103.795 1235.930 1104.165 ;
        RECT 1235.720 1055.885 1235.860 1103.795 ;
        RECT 1234.730 1055.515 1235.010 1055.885 ;
        RECT 1235.650 1055.515 1235.930 1055.885 ;
        RECT 1234.800 1007.410 1234.940 1055.515 ;
        RECT 1234.740 1007.090 1235.000 1007.410 ;
        RECT 1235.660 1007.090 1235.920 1007.410 ;
        RECT 1235.720 959.325 1235.860 1007.090 ;
        RECT 1234.730 958.955 1235.010 959.325 ;
        RECT 1235.650 958.955 1235.930 959.325 ;
        RECT 1234.800 910.850 1234.940 958.955 ;
        RECT 1234.740 910.530 1235.000 910.850 ;
        RECT 1235.660 910.530 1235.920 910.850 ;
        RECT 1235.720 862.765 1235.860 910.530 ;
        RECT 1234.730 862.395 1235.010 862.765 ;
        RECT 1235.650 862.395 1235.930 862.765 ;
        RECT 1234.800 717.730 1234.940 862.395 ;
        RECT 1234.740 717.410 1235.000 717.730 ;
        RECT 1235.660 717.410 1235.920 717.730 ;
        RECT 1235.720 669.645 1235.860 717.410 ;
        RECT 1234.730 669.275 1235.010 669.645 ;
        RECT 1235.650 669.275 1235.930 669.645 ;
        RECT 1234.800 524.270 1234.940 669.275 ;
        RECT 1234.740 523.950 1235.000 524.270 ;
        RECT 1234.740 476.010 1235.000 476.330 ;
        RECT 1234.800 427.710 1234.940 476.010 ;
        RECT 1234.740 427.390 1235.000 427.710 ;
        RECT 1234.740 379.450 1235.000 379.770 ;
        RECT 1234.800 331.150 1234.940 379.450 ;
        RECT 1234.740 330.830 1235.000 331.150 ;
        RECT 1234.740 282.890 1235.000 283.210 ;
        RECT 1234.800 234.590 1234.940 282.890 ;
        RECT 1234.740 234.270 1235.000 234.590 ;
        RECT 1234.740 186.330 1235.000 186.650 ;
        RECT 1234.800 49.485 1234.940 186.330 ;
        RECT 1234.730 49.115 1235.010 49.485 ;
        RECT 1246.230 47.075 1246.510 47.445 ;
        RECT 1246.300 22.430 1246.440 47.075 ;
        RECT 1246.240 22.110 1246.500 22.430 ;
        RECT 2542.060 22.110 2542.320 22.430 ;
        RECT 2542.120 2.400 2542.260 22.110 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
      LAYER via2 ;
        RECT 1234.730 1296.960 1235.010 1297.240 ;
        RECT 1235.650 1296.960 1235.930 1297.240 ;
        RECT 1234.730 1200.400 1235.010 1200.680 ;
        RECT 1235.650 1200.400 1235.930 1200.680 ;
        RECT 1234.730 1103.840 1235.010 1104.120 ;
        RECT 1235.650 1103.840 1235.930 1104.120 ;
        RECT 1234.730 1055.560 1235.010 1055.840 ;
        RECT 1235.650 1055.560 1235.930 1055.840 ;
        RECT 1234.730 959.000 1235.010 959.280 ;
        RECT 1235.650 959.000 1235.930 959.280 ;
        RECT 1234.730 862.440 1235.010 862.720 ;
        RECT 1235.650 862.440 1235.930 862.720 ;
        RECT 1234.730 669.320 1235.010 669.600 ;
        RECT 1235.650 669.320 1235.930 669.600 ;
        RECT 1234.730 49.160 1235.010 49.440 ;
        RECT 1246.230 47.120 1246.510 47.400 ;
      LAYER met3 ;
        RECT 1234.705 1297.250 1235.035 1297.265 ;
        RECT 1235.625 1297.250 1235.955 1297.265 ;
        RECT 1234.705 1296.950 1235.955 1297.250 ;
        RECT 1234.705 1296.935 1235.035 1296.950 ;
        RECT 1235.625 1296.935 1235.955 1296.950 ;
        RECT 1234.705 1200.690 1235.035 1200.705 ;
        RECT 1235.625 1200.690 1235.955 1200.705 ;
        RECT 1234.705 1200.390 1235.955 1200.690 ;
        RECT 1234.705 1200.375 1235.035 1200.390 ;
        RECT 1235.625 1200.375 1235.955 1200.390 ;
        RECT 1234.705 1104.130 1235.035 1104.145 ;
        RECT 1235.625 1104.130 1235.955 1104.145 ;
        RECT 1234.705 1103.830 1235.955 1104.130 ;
        RECT 1234.705 1103.815 1235.035 1103.830 ;
        RECT 1235.625 1103.815 1235.955 1103.830 ;
        RECT 1234.705 1055.850 1235.035 1055.865 ;
        RECT 1235.625 1055.850 1235.955 1055.865 ;
        RECT 1234.705 1055.550 1235.955 1055.850 ;
        RECT 1234.705 1055.535 1235.035 1055.550 ;
        RECT 1235.625 1055.535 1235.955 1055.550 ;
        RECT 1234.705 959.290 1235.035 959.305 ;
        RECT 1235.625 959.290 1235.955 959.305 ;
        RECT 1234.705 958.990 1235.955 959.290 ;
        RECT 1234.705 958.975 1235.035 958.990 ;
        RECT 1235.625 958.975 1235.955 958.990 ;
        RECT 1234.705 862.730 1235.035 862.745 ;
        RECT 1235.625 862.730 1235.955 862.745 ;
        RECT 1234.705 862.430 1235.955 862.730 ;
        RECT 1234.705 862.415 1235.035 862.430 ;
        RECT 1235.625 862.415 1235.955 862.430 ;
        RECT 1234.705 669.610 1235.035 669.625 ;
        RECT 1235.625 669.610 1235.955 669.625 ;
        RECT 1234.705 669.310 1235.955 669.610 ;
        RECT 1234.705 669.295 1235.035 669.310 ;
        RECT 1235.625 669.295 1235.955 669.310 ;
        RECT 1234.705 49.450 1235.035 49.465 ;
        RECT 1234.030 49.150 1235.035 49.450 ;
        RECT 1234.030 47.410 1234.330 49.150 ;
        RECT 1234.705 49.135 1235.035 49.150 ;
        RECT 1246.205 47.410 1246.535 47.425 ;
        RECT 1234.030 47.110 1246.535 47.410 ;
        RECT 1246.205 47.095 1246.535 47.110 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1248.125 22.525 1248.295 34.595 ;
      LAYER mcon ;
        RECT 1248.125 34.425 1248.295 34.595 ;
      LAYER met1 ;
        RECT 1236.090 1548.940 1236.410 1549.000 ;
        RECT 1241.610 1548.940 1241.930 1549.000 ;
        RECT 1236.090 1548.800 1241.930 1548.940 ;
        RECT 1236.090 1548.740 1236.410 1548.800 ;
        RECT 1241.610 1548.740 1241.930 1548.800 ;
        RECT 1241.610 34.580 1241.930 34.640 ;
        RECT 1248.065 34.580 1248.355 34.625 ;
        RECT 1241.610 34.440 1248.355 34.580 ;
        RECT 1241.610 34.380 1241.930 34.440 ;
        RECT 1248.065 34.395 1248.355 34.440 ;
        RECT 1248.065 22.680 1248.355 22.725 ;
        RECT 2559.970 22.680 2560.290 22.740 ;
        RECT 1248.065 22.540 2560.290 22.680 ;
        RECT 1248.065 22.495 1248.355 22.540 ;
        RECT 2559.970 22.480 2560.290 22.540 ;
      LAYER via ;
        RECT 1236.120 1548.740 1236.380 1549.000 ;
        RECT 1241.640 1548.740 1241.900 1549.000 ;
        RECT 1241.640 34.380 1241.900 34.640 ;
        RECT 2560.000 22.480 2560.260 22.740 ;
      LAYER met2 ;
        RECT 1237.360 1600.450 1237.640 1604.000 ;
        RECT 1236.180 1600.310 1237.640 1600.450 ;
        RECT 1236.180 1549.030 1236.320 1600.310 ;
        RECT 1237.360 1600.000 1237.640 1600.310 ;
        RECT 1236.120 1548.710 1236.380 1549.030 ;
        RECT 1241.640 1548.710 1241.900 1549.030 ;
        RECT 1241.700 34.670 1241.840 1548.710 ;
        RECT 1241.640 34.350 1241.900 34.670 ;
        RECT 2560.000 22.450 2560.260 22.770 ;
        RECT 2560.060 2.400 2560.200 22.450 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1293.665 22.865 1293.835 26.775 ;
      LAYER mcon ;
        RECT 1293.665 26.605 1293.835 26.775 ;
      LAYER met1 ;
        RECT 1242.070 1535.340 1242.390 1535.400 ;
        RECT 1248.510 1535.340 1248.830 1535.400 ;
        RECT 1242.070 1535.200 1248.830 1535.340 ;
        RECT 1242.070 1535.140 1242.390 1535.200 ;
        RECT 1248.510 1535.140 1248.830 1535.200 ;
        RECT 1248.510 26.760 1248.830 26.820 ;
        RECT 1293.605 26.760 1293.895 26.805 ;
        RECT 1248.510 26.620 1293.895 26.760 ;
        RECT 1248.510 26.560 1248.830 26.620 ;
        RECT 1293.605 26.575 1293.895 26.620 ;
        RECT 1293.605 23.020 1293.895 23.065 ;
        RECT 2577.910 23.020 2578.230 23.080 ;
        RECT 1293.605 22.880 2578.230 23.020 ;
        RECT 1293.605 22.835 1293.895 22.880 ;
        RECT 2577.910 22.820 2578.230 22.880 ;
      LAYER via ;
        RECT 1242.100 1535.140 1242.360 1535.400 ;
        RECT 1248.540 1535.140 1248.800 1535.400 ;
        RECT 1248.540 26.560 1248.800 26.820 ;
        RECT 2577.940 22.820 2578.200 23.080 ;
      LAYER met2 ;
        RECT 1243.340 1600.450 1243.620 1604.000 ;
        RECT 1242.160 1600.310 1243.620 1600.450 ;
        RECT 1242.160 1535.430 1242.300 1600.310 ;
        RECT 1243.340 1600.000 1243.620 1600.310 ;
        RECT 1242.100 1535.110 1242.360 1535.430 ;
        RECT 1248.540 1535.110 1248.800 1535.430 ;
        RECT 1248.600 26.850 1248.740 1535.110 ;
        RECT 1248.540 26.530 1248.800 26.850 ;
        RECT 2577.940 22.790 2578.200 23.110 ;
        RECT 2578.000 2.400 2578.140 22.790 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 631.190 1589.740 631.510 1589.800 ;
        RECT 634.410 1589.740 634.730 1589.800 ;
        RECT 631.190 1589.600 634.730 1589.740 ;
        RECT 631.190 1589.540 631.510 1589.600 ;
        RECT 634.410 1589.540 634.730 1589.600 ;
        RECT 634.410 17.920 634.730 17.980 ;
        RECT 811.510 17.920 811.830 17.980 ;
        RECT 634.410 17.780 811.830 17.920 ;
        RECT 634.410 17.720 634.730 17.780 ;
        RECT 811.510 17.720 811.830 17.780 ;
      LAYER via ;
        RECT 631.220 1589.540 631.480 1589.800 ;
        RECT 634.440 1589.540 634.700 1589.800 ;
        RECT 634.440 17.720 634.700 17.980 ;
        RECT 811.540 17.720 811.800 17.980 ;
      LAYER met2 ;
        RECT 631.080 1600.380 631.360 1604.000 ;
        RECT 631.080 1600.000 631.420 1600.380 ;
        RECT 631.280 1589.830 631.420 1600.000 ;
        RECT 631.220 1589.510 631.480 1589.830 ;
        RECT 634.440 1589.510 634.700 1589.830 ;
        RECT 634.500 18.010 634.640 1589.510 ;
        RECT 634.440 17.690 634.700 18.010 ;
        RECT 811.540 17.690 811.800 18.010 ;
        RECT 811.600 2.400 811.740 17.690 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.970 1535.340 1249.290 1535.400 ;
        RECT 1255.410 1535.340 1255.730 1535.400 ;
        RECT 1248.970 1535.200 1255.730 1535.340 ;
        RECT 1248.970 1535.140 1249.290 1535.200 ;
        RECT 1255.410 1535.140 1255.730 1535.200 ;
        RECT 1255.410 23.360 1255.730 23.420 ;
        RECT 2595.390 23.360 2595.710 23.420 ;
        RECT 1255.410 23.220 2595.710 23.360 ;
        RECT 1255.410 23.160 1255.730 23.220 ;
        RECT 2595.390 23.160 2595.710 23.220 ;
      LAYER via ;
        RECT 1249.000 1535.140 1249.260 1535.400 ;
        RECT 1255.440 1535.140 1255.700 1535.400 ;
        RECT 1255.440 23.160 1255.700 23.420 ;
        RECT 2595.420 23.160 2595.680 23.420 ;
      LAYER met2 ;
        RECT 1249.320 1600.380 1249.600 1604.000 ;
        RECT 1249.320 1600.000 1249.660 1600.380 ;
        RECT 1249.520 1597.220 1249.660 1600.000 ;
        RECT 1249.060 1597.080 1249.660 1597.220 ;
        RECT 1249.060 1535.430 1249.200 1597.080 ;
        RECT 1249.000 1535.110 1249.260 1535.430 ;
        RECT 1255.440 1535.110 1255.700 1535.430 ;
        RECT 1255.500 23.450 1255.640 1535.110 ;
        RECT 1255.440 23.130 1255.700 23.450 ;
        RECT 2595.420 23.130 2595.680 23.450 ;
        RECT 2595.480 2.400 2595.620 23.130 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1275.265 23.545 1275.435 25.075 ;
      LAYER mcon ;
        RECT 1275.265 24.905 1275.435 25.075 ;
      LAYER met1 ;
        RECT 1256.790 1580.900 1257.110 1580.960 ;
        RECT 1262.310 1580.900 1262.630 1580.960 ;
        RECT 1256.790 1580.760 1262.630 1580.900 ;
        RECT 1256.790 1580.700 1257.110 1580.760 ;
        RECT 1262.310 1580.700 1262.630 1580.760 ;
        RECT 1262.310 25.060 1262.630 25.120 ;
        RECT 1275.205 25.060 1275.495 25.105 ;
        RECT 1262.310 24.920 1275.495 25.060 ;
        RECT 1262.310 24.860 1262.630 24.920 ;
        RECT 1275.205 24.875 1275.495 24.920 ;
        RECT 1275.205 23.700 1275.495 23.745 ;
        RECT 2613.330 23.700 2613.650 23.760 ;
        RECT 1275.205 23.560 2613.650 23.700 ;
        RECT 1275.205 23.515 1275.495 23.560 ;
        RECT 2613.330 23.500 2613.650 23.560 ;
      LAYER via ;
        RECT 1256.820 1580.700 1257.080 1580.960 ;
        RECT 1262.340 1580.700 1262.600 1580.960 ;
        RECT 1262.340 24.860 1262.600 25.120 ;
        RECT 2613.360 23.500 2613.620 23.760 ;
      LAYER met2 ;
        RECT 1255.760 1600.450 1256.040 1604.000 ;
        RECT 1255.760 1600.310 1257.020 1600.450 ;
        RECT 1255.760 1600.000 1256.040 1600.310 ;
        RECT 1256.880 1580.990 1257.020 1600.310 ;
        RECT 1256.820 1580.670 1257.080 1580.990 ;
        RECT 1262.340 1580.670 1262.600 1580.990 ;
        RECT 1262.400 25.150 1262.540 1580.670 ;
        RECT 1262.340 24.830 1262.600 25.150 ;
        RECT 2613.360 23.470 2613.620 23.790 ;
        RECT 2613.420 2.400 2613.560 23.470 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1261.850 27.440 1262.170 27.500 ;
        RECT 2631.270 27.440 2631.590 27.500 ;
        RECT 1261.850 27.300 2631.590 27.440 ;
        RECT 1261.850 27.240 1262.170 27.300 ;
        RECT 2631.270 27.240 2631.590 27.300 ;
      LAYER via ;
        RECT 1261.880 27.240 1262.140 27.500 ;
        RECT 2631.300 27.240 2631.560 27.500 ;
      LAYER met2 ;
        RECT 1261.740 1600.380 1262.020 1604.000 ;
        RECT 1261.740 1600.000 1262.080 1600.380 ;
        RECT 1261.940 27.530 1262.080 1600.000 ;
        RECT 1261.880 27.210 1262.140 27.530 ;
        RECT 2631.300 27.210 2631.560 27.530 ;
        RECT 2631.360 2.400 2631.500 27.210 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.770 1579.880 1263.090 1579.940 ;
        RECT 1266.910 1579.880 1267.230 1579.940 ;
        RECT 1262.770 1579.740 1267.230 1579.880 ;
        RECT 1262.770 1579.680 1263.090 1579.740 ;
        RECT 1266.910 1579.680 1267.230 1579.740 ;
        RECT 1262.770 1535.340 1263.090 1535.400 ;
        RECT 1269.210 1535.340 1269.530 1535.400 ;
        RECT 1262.770 1535.200 1269.530 1535.340 ;
        RECT 1262.770 1535.140 1263.090 1535.200 ;
        RECT 1269.210 1535.140 1269.530 1535.200 ;
        RECT 1268.290 55.320 1268.610 55.380 ;
        RECT 1269.210 55.320 1269.530 55.380 ;
        RECT 1268.290 55.180 1269.530 55.320 ;
        RECT 1268.290 55.120 1268.610 55.180 ;
        RECT 1269.210 55.120 1269.530 55.180 ;
        RECT 1268.290 27.100 1268.610 27.160 ;
        RECT 2649.210 27.100 2649.530 27.160 ;
        RECT 1268.290 26.960 2649.530 27.100 ;
        RECT 1268.290 26.900 1268.610 26.960 ;
        RECT 2649.210 26.900 2649.530 26.960 ;
      LAYER via ;
        RECT 1262.800 1579.680 1263.060 1579.940 ;
        RECT 1266.940 1579.680 1267.200 1579.940 ;
        RECT 1262.800 1535.140 1263.060 1535.400 ;
        RECT 1269.240 1535.140 1269.500 1535.400 ;
        RECT 1268.320 55.120 1268.580 55.380 ;
        RECT 1269.240 55.120 1269.500 55.380 ;
        RECT 1268.320 26.900 1268.580 27.160 ;
        RECT 2649.240 26.900 2649.500 27.160 ;
      LAYER met2 ;
        RECT 1268.180 1600.450 1268.460 1604.000 ;
        RECT 1267.000 1600.310 1268.460 1600.450 ;
        RECT 1267.000 1579.970 1267.140 1600.310 ;
        RECT 1268.180 1600.000 1268.460 1600.310 ;
        RECT 1262.800 1579.650 1263.060 1579.970 ;
        RECT 1266.940 1579.650 1267.200 1579.970 ;
        RECT 1262.860 1535.430 1263.000 1579.650 ;
        RECT 1262.800 1535.110 1263.060 1535.430 ;
        RECT 1269.240 1535.110 1269.500 1535.430 ;
        RECT 1269.300 55.410 1269.440 1535.110 ;
        RECT 1268.320 55.090 1268.580 55.410 ;
        RECT 1269.240 55.090 1269.500 55.410 ;
        RECT 1268.380 27.190 1268.520 55.090 ;
        RECT 1268.320 26.870 1268.580 27.190 ;
        RECT 2649.240 26.870 2649.500 27.190 ;
        RECT 2649.300 2.400 2649.440 26.870 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1276.185 1490.645 1276.355 1497.615 ;
        RECT 1276.185 1442.025 1276.355 1490.135 ;
        RECT 1276.185 531.505 1276.355 620.755 ;
        RECT 1276.185 434.945 1276.355 524.195 ;
        RECT 1276.185 379.525 1276.355 427.635 ;
        RECT 1276.185 282.965 1276.355 331.075 ;
        RECT 1276.185 186.405 1276.355 234.515 ;
        RECT 1276.185 89.845 1276.355 137.955 ;
        RECT 1294.125 25.585 1294.295 26.775 ;
      LAYER mcon ;
        RECT 1276.185 1497.445 1276.355 1497.615 ;
        RECT 1276.185 1489.965 1276.355 1490.135 ;
        RECT 1276.185 620.585 1276.355 620.755 ;
        RECT 1276.185 524.025 1276.355 524.195 ;
        RECT 1276.185 427.465 1276.355 427.635 ;
        RECT 1276.185 330.905 1276.355 331.075 ;
        RECT 1276.185 234.345 1276.355 234.515 ;
        RECT 1276.185 137.785 1276.355 137.955 ;
        RECT 1294.125 26.605 1294.295 26.775 ;
      LAYER met1 ;
        RECT 1276.110 1497.600 1276.430 1497.660 ;
        RECT 1275.915 1497.460 1276.430 1497.600 ;
        RECT 1276.110 1497.400 1276.430 1497.460 ;
        RECT 1276.110 1490.800 1276.430 1490.860 ;
        RECT 1275.915 1490.660 1276.430 1490.800 ;
        RECT 1276.110 1490.600 1276.430 1490.660 ;
        RECT 1276.110 1490.120 1276.430 1490.180 ;
        RECT 1275.915 1489.980 1276.430 1490.120 ;
        RECT 1276.110 1489.920 1276.430 1489.980 ;
        RECT 1276.110 1442.180 1276.430 1442.240 ;
        RECT 1275.915 1442.040 1276.430 1442.180 ;
        RECT 1276.110 1441.980 1276.430 1442.040 ;
        RECT 1276.110 1345.620 1276.430 1345.680 ;
        RECT 1276.570 1345.620 1276.890 1345.680 ;
        RECT 1276.110 1345.480 1276.890 1345.620 ;
        RECT 1276.110 1345.420 1276.430 1345.480 ;
        RECT 1276.570 1345.420 1276.890 1345.480 ;
        RECT 1276.110 1200.780 1276.430 1200.840 ;
        RECT 1276.570 1200.780 1276.890 1200.840 ;
        RECT 1276.110 1200.640 1276.890 1200.780 ;
        RECT 1276.110 1200.580 1276.430 1200.640 ;
        RECT 1276.570 1200.580 1276.890 1200.640 ;
        RECT 1276.110 1152.500 1276.430 1152.560 ;
        RECT 1276.570 1152.500 1276.890 1152.560 ;
        RECT 1276.110 1152.360 1276.890 1152.500 ;
        RECT 1276.110 1152.300 1276.430 1152.360 ;
        RECT 1276.570 1152.300 1276.890 1152.360 ;
        RECT 1276.110 1145.360 1276.430 1145.420 ;
        RECT 1277.490 1145.360 1277.810 1145.420 ;
        RECT 1276.110 1145.220 1277.810 1145.360 ;
        RECT 1276.110 1145.160 1276.430 1145.220 ;
        RECT 1277.490 1145.160 1277.810 1145.220 ;
        RECT 1276.570 1055.740 1276.890 1056.000 ;
        RECT 1276.660 1055.260 1276.800 1055.740 ;
        RECT 1277.950 1055.260 1278.270 1055.320 ;
        RECT 1276.660 1055.120 1278.270 1055.260 ;
        RECT 1277.950 1055.060 1278.270 1055.120 ;
        RECT 1277.030 1031.120 1277.350 1031.180 ;
        RECT 1277.950 1031.120 1278.270 1031.180 ;
        RECT 1277.030 1030.980 1278.270 1031.120 ;
        RECT 1277.030 1030.920 1277.350 1030.980 ;
        RECT 1277.950 1030.920 1278.270 1030.980 ;
        RECT 1276.570 952.580 1276.890 952.640 ;
        RECT 1277.030 952.580 1277.350 952.640 ;
        RECT 1276.570 952.440 1277.350 952.580 ;
        RECT 1276.570 952.380 1276.890 952.440 ;
        RECT 1277.030 952.380 1277.350 952.440 ;
        RECT 1276.570 855.680 1276.890 855.740 ;
        RECT 1277.030 855.680 1277.350 855.740 ;
        RECT 1276.570 855.540 1277.350 855.680 ;
        RECT 1276.570 855.480 1276.890 855.540 ;
        RECT 1277.030 855.480 1277.350 855.540 ;
        RECT 1276.110 620.740 1276.430 620.800 ;
        RECT 1275.915 620.600 1276.430 620.740 ;
        RECT 1276.110 620.540 1276.430 620.600 ;
        RECT 1276.110 531.660 1276.430 531.720 ;
        RECT 1275.915 531.520 1276.430 531.660 ;
        RECT 1276.110 531.460 1276.430 531.520 ;
        RECT 1276.110 524.180 1276.430 524.240 ;
        RECT 1275.915 524.040 1276.430 524.180 ;
        RECT 1276.110 523.980 1276.430 524.040 ;
        RECT 1276.110 435.100 1276.430 435.160 ;
        RECT 1275.915 434.960 1276.430 435.100 ;
        RECT 1276.110 434.900 1276.430 434.960 ;
        RECT 1276.110 427.620 1276.430 427.680 ;
        RECT 1275.915 427.480 1276.430 427.620 ;
        RECT 1276.110 427.420 1276.430 427.480 ;
        RECT 1276.110 379.680 1276.430 379.740 ;
        RECT 1275.915 379.540 1276.430 379.680 ;
        RECT 1276.110 379.480 1276.430 379.540 ;
        RECT 1276.110 331.060 1276.430 331.120 ;
        RECT 1275.915 330.920 1276.430 331.060 ;
        RECT 1276.110 330.860 1276.430 330.920 ;
        RECT 1276.110 283.120 1276.430 283.180 ;
        RECT 1275.915 282.980 1276.430 283.120 ;
        RECT 1276.110 282.920 1276.430 282.980 ;
        RECT 1276.110 234.500 1276.430 234.560 ;
        RECT 1275.915 234.360 1276.430 234.500 ;
        RECT 1276.110 234.300 1276.430 234.360 ;
        RECT 1276.110 186.560 1276.430 186.620 ;
        RECT 1275.915 186.420 1276.430 186.560 ;
        RECT 1276.110 186.360 1276.430 186.420 ;
        RECT 1276.110 137.940 1276.430 138.000 ;
        RECT 1275.915 137.800 1276.430 137.940 ;
        RECT 1276.110 137.740 1276.430 137.800 ;
        RECT 1276.110 90.000 1276.430 90.060 ;
        RECT 1275.915 89.860 1276.430 90.000 ;
        RECT 1276.110 89.800 1276.430 89.860 ;
        RECT 1294.065 26.760 1294.355 26.805 ;
        RECT 2667.150 26.760 2667.470 26.820 ;
        RECT 1294.065 26.620 2667.470 26.760 ;
        RECT 1294.065 26.575 1294.355 26.620 ;
        RECT 2667.150 26.560 2667.470 26.620 ;
        RECT 1275.650 25.740 1275.970 25.800 ;
        RECT 1294.065 25.740 1294.355 25.785 ;
        RECT 1275.650 25.600 1294.355 25.740 ;
        RECT 1275.650 25.540 1275.970 25.600 ;
        RECT 1294.065 25.555 1294.355 25.600 ;
      LAYER via ;
        RECT 1276.140 1497.400 1276.400 1497.660 ;
        RECT 1276.140 1490.600 1276.400 1490.860 ;
        RECT 1276.140 1489.920 1276.400 1490.180 ;
        RECT 1276.140 1441.980 1276.400 1442.240 ;
        RECT 1276.140 1345.420 1276.400 1345.680 ;
        RECT 1276.600 1345.420 1276.860 1345.680 ;
        RECT 1276.140 1200.580 1276.400 1200.840 ;
        RECT 1276.600 1200.580 1276.860 1200.840 ;
        RECT 1276.140 1152.300 1276.400 1152.560 ;
        RECT 1276.600 1152.300 1276.860 1152.560 ;
        RECT 1276.140 1145.160 1276.400 1145.420 ;
        RECT 1277.520 1145.160 1277.780 1145.420 ;
        RECT 1276.600 1055.740 1276.860 1056.000 ;
        RECT 1277.980 1055.060 1278.240 1055.320 ;
        RECT 1277.060 1030.920 1277.320 1031.180 ;
        RECT 1277.980 1030.920 1278.240 1031.180 ;
        RECT 1276.600 952.380 1276.860 952.640 ;
        RECT 1277.060 952.380 1277.320 952.640 ;
        RECT 1276.600 855.480 1276.860 855.740 ;
        RECT 1277.060 855.480 1277.320 855.740 ;
        RECT 1276.140 620.540 1276.400 620.800 ;
        RECT 1276.140 531.460 1276.400 531.720 ;
        RECT 1276.140 523.980 1276.400 524.240 ;
        RECT 1276.140 434.900 1276.400 435.160 ;
        RECT 1276.140 427.420 1276.400 427.680 ;
        RECT 1276.140 379.480 1276.400 379.740 ;
        RECT 1276.140 330.860 1276.400 331.120 ;
        RECT 1276.140 282.920 1276.400 283.180 ;
        RECT 1276.140 234.300 1276.400 234.560 ;
        RECT 1276.140 186.360 1276.400 186.620 ;
        RECT 1276.140 137.740 1276.400 138.000 ;
        RECT 1276.140 89.800 1276.400 90.060 ;
        RECT 2667.180 26.560 2667.440 26.820 ;
        RECT 1275.680 25.540 1275.940 25.800 ;
      LAYER met2 ;
        RECT 1274.160 1600.450 1274.440 1604.000 ;
        RECT 1274.160 1600.310 1275.880 1600.450 ;
        RECT 1274.160 1600.000 1274.440 1600.310 ;
        RECT 1275.740 1580.050 1275.880 1600.310 ;
        RECT 1275.740 1579.910 1276.340 1580.050 ;
        RECT 1276.200 1497.690 1276.340 1579.910 ;
        RECT 1276.140 1497.370 1276.400 1497.690 ;
        RECT 1276.140 1490.570 1276.400 1490.890 ;
        RECT 1276.200 1490.210 1276.340 1490.570 ;
        RECT 1276.140 1489.890 1276.400 1490.210 ;
        RECT 1276.140 1441.950 1276.400 1442.270 ;
        RECT 1276.200 1393.845 1276.340 1441.950 ;
        RECT 1276.130 1393.475 1276.410 1393.845 ;
        RECT 1276.590 1392.795 1276.870 1393.165 ;
        RECT 1276.660 1345.710 1276.800 1392.795 ;
        RECT 1276.140 1345.390 1276.400 1345.710 ;
        RECT 1276.600 1345.390 1276.860 1345.710 ;
        RECT 1276.200 1200.870 1276.340 1345.390 ;
        RECT 1276.140 1200.550 1276.400 1200.870 ;
        RECT 1276.600 1200.550 1276.860 1200.870 ;
        RECT 1276.660 1152.590 1276.800 1200.550 ;
        RECT 1276.140 1152.270 1276.400 1152.590 ;
        RECT 1276.600 1152.270 1276.860 1152.590 ;
        RECT 1276.200 1145.450 1276.340 1152.270 ;
        RECT 1276.140 1145.130 1276.400 1145.450 ;
        RECT 1277.520 1145.130 1277.780 1145.450 ;
        RECT 1277.580 1097.365 1277.720 1145.130 ;
        RECT 1276.590 1096.995 1276.870 1097.365 ;
        RECT 1277.510 1096.995 1277.790 1097.365 ;
        RECT 1276.660 1056.030 1276.800 1096.995 ;
        RECT 1276.600 1055.710 1276.860 1056.030 ;
        RECT 1277.980 1055.030 1278.240 1055.350 ;
        RECT 1278.040 1031.210 1278.180 1055.030 ;
        RECT 1277.060 1030.890 1277.320 1031.210 ;
        RECT 1277.980 1030.890 1278.240 1031.210 ;
        RECT 1277.120 952.670 1277.260 1030.890 ;
        RECT 1276.600 952.350 1276.860 952.670 ;
        RECT 1277.060 952.350 1277.320 952.670 ;
        RECT 1276.660 910.930 1276.800 952.350 ;
        RECT 1276.660 910.790 1277.260 910.930 ;
        RECT 1277.120 855.770 1277.260 910.790 ;
        RECT 1276.600 855.450 1276.860 855.770 ;
        RECT 1277.060 855.450 1277.320 855.770 ;
        RECT 1276.660 814.370 1276.800 855.450 ;
        RECT 1276.660 814.230 1277.260 814.370 ;
        RECT 1277.120 766.205 1277.260 814.230 ;
        RECT 1276.130 765.835 1276.410 766.205 ;
        RECT 1277.050 765.835 1277.330 766.205 ;
        RECT 1276.200 717.245 1276.340 765.835 ;
        RECT 1276.130 716.875 1276.410 717.245 ;
        RECT 1277.050 669.275 1277.330 669.645 ;
        RECT 1277.120 628.165 1277.260 669.275 ;
        RECT 1276.130 627.795 1276.410 628.165 ;
        RECT 1277.050 627.795 1277.330 628.165 ;
        RECT 1276.200 620.830 1276.340 627.795 ;
        RECT 1276.140 620.510 1276.400 620.830 ;
        RECT 1276.140 531.430 1276.400 531.750 ;
        RECT 1276.200 524.270 1276.340 531.430 ;
        RECT 1276.140 523.950 1276.400 524.270 ;
        RECT 1276.140 434.870 1276.400 435.190 ;
        RECT 1276.200 427.710 1276.340 434.870 ;
        RECT 1276.140 427.390 1276.400 427.710 ;
        RECT 1276.140 379.450 1276.400 379.770 ;
        RECT 1276.200 331.150 1276.340 379.450 ;
        RECT 1276.140 330.830 1276.400 331.150 ;
        RECT 1276.140 282.890 1276.400 283.210 ;
        RECT 1276.200 234.590 1276.340 282.890 ;
        RECT 1276.140 234.270 1276.400 234.590 ;
        RECT 1276.140 186.330 1276.400 186.650 ;
        RECT 1276.200 138.030 1276.340 186.330 ;
        RECT 1276.140 137.710 1276.400 138.030 ;
        RECT 1276.140 89.770 1276.400 90.090 ;
        RECT 1276.200 62.290 1276.340 89.770 ;
        RECT 1276.200 62.150 1276.800 62.290 ;
        RECT 1276.660 61.610 1276.800 62.150 ;
        RECT 1275.280 61.470 1276.800 61.610 ;
        RECT 1275.280 45.290 1275.420 61.470 ;
        RECT 1275.280 45.150 1275.880 45.290 ;
        RECT 1275.740 25.830 1275.880 45.150 ;
        RECT 2667.180 26.530 2667.440 26.850 ;
        RECT 1275.680 25.510 1275.940 25.830 ;
        RECT 2667.240 2.400 2667.380 26.530 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
      LAYER via2 ;
        RECT 1276.130 1393.520 1276.410 1393.800 ;
        RECT 1276.590 1392.840 1276.870 1393.120 ;
        RECT 1276.590 1097.040 1276.870 1097.320 ;
        RECT 1277.510 1097.040 1277.790 1097.320 ;
        RECT 1276.130 765.880 1276.410 766.160 ;
        RECT 1277.050 765.880 1277.330 766.160 ;
        RECT 1276.130 716.920 1276.410 717.200 ;
        RECT 1277.050 669.320 1277.330 669.600 ;
        RECT 1276.130 627.840 1276.410 628.120 ;
        RECT 1277.050 627.840 1277.330 628.120 ;
      LAYER met3 ;
        RECT 1276.105 1393.810 1276.435 1393.825 ;
        RECT 1275.430 1393.510 1276.435 1393.810 ;
        RECT 1275.430 1393.130 1275.730 1393.510 ;
        RECT 1276.105 1393.495 1276.435 1393.510 ;
        RECT 1276.565 1393.130 1276.895 1393.145 ;
        RECT 1275.430 1392.830 1276.895 1393.130 ;
        RECT 1276.565 1392.815 1276.895 1392.830 ;
        RECT 1276.565 1097.330 1276.895 1097.345 ;
        RECT 1277.485 1097.330 1277.815 1097.345 ;
        RECT 1276.565 1097.030 1277.815 1097.330 ;
        RECT 1276.565 1097.015 1276.895 1097.030 ;
        RECT 1277.485 1097.015 1277.815 1097.030 ;
        RECT 1276.105 766.170 1276.435 766.185 ;
        RECT 1277.025 766.170 1277.355 766.185 ;
        RECT 1276.105 765.870 1277.355 766.170 ;
        RECT 1276.105 765.855 1276.435 765.870 ;
        RECT 1277.025 765.855 1277.355 765.870 ;
        RECT 1276.105 717.220 1276.435 717.225 ;
        RECT 1276.105 717.210 1276.690 717.220 ;
        RECT 1275.880 716.910 1276.690 717.210 ;
        RECT 1276.105 716.900 1276.690 716.910 ;
        RECT 1276.105 716.895 1276.435 716.900 ;
        RECT 1276.310 669.610 1276.690 669.620 ;
        RECT 1277.025 669.610 1277.355 669.625 ;
        RECT 1276.310 669.310 1277.355 669.610 ;
        RECT 1276.310 669.300 1276.690 669.310 ;
        RECT 1277.025 669.295 1277.355 669.310 ;
        RECT 1276.105 628.130 1276.435 628.145 ;
        RECT 1277.025 628.130 1277.355 628.145 ;
        RECT 1276.105 627.830 1277.355 628.130 ;
        RECT 1276.105 627.815 1276.435 627.830 ;
        RECT 1277.025 627.815 1277.355 627.830 ;
      LAYER via3 ;
        RECT 1276.340 716.900 1276.660 717.220 ;
        RECT 1276.340 669.300 1276.660 669.620 ;
      LAYER met4 ;
        RECT 1276.335 716.895 1276.665 717.225 ;
        RECT 1276.350 669.625 1276.650 716.895 ;
        RECT 1276.335 669.295 1276.665 669.625 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1277.490 1535.000 1277.810 1535.060 ;
        RECT 1283.010 1535.000 1283.330 1535.060 ;
        RECT 1277.490 1534.860 1283.330 1535.000 ;
        RECT 1277.490 1534.800 1277.810 1534.860 ;
        RECT 1283.010 1534.800 1283.330 1534.860 ;
        RECT 1283.010 26.420 1283.330 26.480 ;
        RECT 2684.630 26.420 2684.950 26.480 ;
        RECT 1283.010 26.280 2684.950 26.420 ;
        RECT 1283.010 26.220 1283.330 26.280 ;
        RECT 2684.630 26.220 2684.950 26.280 ;
      LAYER via ;
        RECT 1277.520 1534.800 1277.780 1535.060 ;
        RECT 1283.040 1534.800 1283.300 1535.060 ;
        RECT 1283.040 26.220 1283.300 26.480 ;
        RECT 2684.660 26.220 2684.920 26.480 ;
      LAYER met2 ;
        RECT 1280.600 1600.450 1280.880 1604.000 ;
        RECT 1278.960 1600.310 1280.880 1600.450 ;
        RECT 1278.960 1580.050 1279.100 1600.310 ;
        RECT 1280.600 1600.000 1280.880 1600.310 ;
        RECT 1277.580 1579.910 1279.100 1580.050 ;
        RECT 1277.580 1535.090 1277.720 1579.910 ;
        RECT 1277.520 1534.770 1277.780 1535.090 ;
        RECT 1283.040 1534.770 1283.300 1535.090 ;
        RECT 1283.100 26.510 1283.240 1534.770 ;
        RECT 1283.040 26.190 1283.300 26.510 ;
        RECT 2684.660 26.190 2684.920 26.510 ;
        RECT 2684.720 2.400 2684.860 26.190 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1283.470 1535.340 1283.790 1535.400 ;
        RECT 1289.910 1535.340 1290.230 1535.400 ;
        RECT 1283.470 1535.200 1290.230 1535.340 ;
        RECT 1283.470 1535.140 1283.790 1535.200 ;
        RECT 1289.910 1535.140 1290.230 1535.200 ;
        RECT 1289.910 26.080 1290.230 26.140 ;
        RECT 2702.570 26.080 2702.890 26.140 ;
        RECT 1289.910 25.940 2702.890 26.080 ;
        RECT 1289.910 25.880 1290.230 25.940 ;
        RECT 2702.570 25.880 2702.890 25.940 ;
      LAYER via ;
        RECT 1283.500 1535.140 1283.760 1535.400 ;
        RECT 1289.940 1535.140 1290.200 1535.400 ;
        RECT 1289.940 25.880 1290.200 26.140 ;
        RECT 2702.600 25.880 2702.860 26.140 ;
      LAYER met2 ;
        RECT 1286.580 1600.450 1286.860 1604.000 ;
        RECT 1285.400 1600.310 1286.860 1600.450 ;
        RECT 1285.400 1580.050 1285.540 1600.310 ;
        RECT 1286.580 1600.000 1286.860 1600.310 ;
        RECT 1283.560 1579.910 1285.540 1580.050 ;
        RECT 1283.560 1535.430 1283.700 1579.910 ;
        RECT 1283.500 1535.110 1283.760 1535.430 ;
        RECT 1289.940 1535.110 1290.200 1535.430 ;
        RECT 1290.000 26.170 1290.140 1535.110 ;
        RECT 1289.940 25.850 1290.200 26.170 ;
        RECT 2702.600 25.850 2702.860 26.170 ;
        RECT 2702.660 2.400 2702.800 25.850 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1342.425 24.225 1342.595 25.755 ;
      LAYER mcon ;
        RECT 1342.425 25.585 1342.595 25.755 ;
      LAYER met1 ;
        RECT 1294.050 1579.880 1294.370 1579.940 ;
        RECT 1296.810 1579.880 1297.130 1579.940 ;
        RECT 1294.050 1579.740 1297.130 1579.880 ;
        RECT 1294.050 1579.680 1294.370 1579.740 ;
        RECT 1296.810 1579.680 1297.130 1579.740 ;
        RECT 1342.365 25.740 1342.655 25.785 ;
        RECT 2720.510 25.740 2720.830 25.800 ;
        RECT 1342.365 25.600 2720.830 25.740 ;
        RECT 1342.365 25.555 1342.655 25.600 ;
        RECT 2720.510 25.540 2720.830 25.600 ;
        RECT 1296.350 24.380 1296.670 24.440 ;
        RECT 1342.365 24.380 1342.655 24.425 ;
        RECT 1296.350 24.240 1342.655 24.380 ;
        RECT 1296.350 24.180 1296.670 24.240 ;
        RECT 1342.365 24.195 1342.655 24.240 ;
      LAYER via ;
        RECT 1294.080 1579.680 1294.340 1579.940 ;
        RECT 1296.840 1579.680 1297.100 1579.940 ;
        RECT 2720.540 25.540 2720.800 25.800 ;
        RECT 1296.380 24.180 1296.640 24.440 ;
      LAYER met2 ;
        RECT 1293.020 1600.450 1293.300 1604.000 ;
        RECT 1293.020 1600.310 1294.280 1600.450 ;
        RECT 1293.020 1600.000 1293.300 1600.310 ;
        RECT 1294.140 1579.970 1294.280 1600.310 ;
        RECT 1294.080 1579.650 1294.340 1579.970 ;
        RECT 1296.840 1579.650 1297.100 1579.970 ;
        RECT 1296.900 61.610 1297.040 1579.650 ;
        RECT 1296.440 61.470 1297.040 61.610 ;
        RECT 1296.440 24.470 1296.580 61.470 ;
        RECT 2720.540 25.510 2720.800 25.830 ;
        RECT 1296.380 24.150 1296.640 24.470 ;
        RECT 2720.600 2.400 2720.740 25.510 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1298.190 1535.340 1298.510 1535.400 ;
        RECT 1303.710 1535.340 1304.030 1535.400 ;
        RECT 1298.190 1535.200 1304.030 1535.340 ;
        RECT 1298.190 1535.140 1298.510 1535.200 ;
        RECT 1303.710 1535.140 1304.030 1535.200 ;
        RECT 1303.710 25.740 1304.030 25.800 ;
        RECT 1303.710 25.600 1342.120 25.740 ;
        RECT 1303.710 25.540 1304.030 25.600 ;
        RECT 1341.980 25.400 1342.120 25.600 ;
        RECT 2738.450 25.400 2738.770 25.460 ;
        RECT 1341.980 25.260 2738.770 25.400 ;
        RECT 2738.450 25.200 2738.770 25.260 ;
      LAYER via ;
        RECT 1298.220 1535.140 1298.480 1535.400 ;
        RECT 1303.740 1535.140 1304.000 1535.400 ;
        RECT 1303.740 25.540 1304.000 25.800 ;
        RECT 2738.480 25.200 2738.740 25.460 ;
      LAYER met2 ;
        RECT 1299.000 1600.450 1299.280 1604.000 ;
        RECT 1298.280 1600.310 1299.280 1600.450 ;
        RECT 1298.280 1535.430 1298.420 1600.310 ;
        RECT 1299.000 1600.000 1299.280 1600.310 ;
        RECT 1298.220 1535.110 1298.480 1535.430 ;
        RECT 1303.740 1535.110 1304.000 1535.430 ;
        RECT 1303.800 25.830 1303.940 1535.110 ;
        RECT 1303.740 25.510 1304.000 25.830 ;
        RECT 2738.480 25.170 2738.740 25.490 ;
        RECT 2738.540 2.400 2738.680 25.170 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1340.125 24.905 1341.675 25.075 ;
      LAYER mcon ;
        RECT 1341.505 24.905 1341.675 25.075 ;
      LAYER met1 ;
        RECT 1306.470 1579.880 1306.790 1579.940 ;
        RECT 1310.610 1579.880 1310.930 1579.940 ;
        RECT 1306.470 1579.740 1310.930 1579.880 ;
        RECT 1306.470 1579.680 1306.790 1579.740 ;
        RECT 1310.610 1579.680 1310.930 1579.740 ;
        RECT 1310.610 25.060 1310.930 25.120 ;
        RECT 1340.065 25.060 1340.355 25.105 ;
        RECT 1310.610 24.920 1340.355 25.060 ;
        RECT 1310.610 24.860 1310.930 24.920 ;
        RECT 1340.065 24.875 1340.355 24.920 ;
        RECT 1341.445 25.060 1341.735 25.105 ;
        RECT 2755.930 25.060 2756.250 25.120 ;
        RECT 1341.445 24.920 2756.250 25.060 ;
        RECT 1341.445 24.875 1341.735 24.920 ;
        RECT 2755.930 24.860 2756.250 24.920 ;
      LAYER via ;
        RECT 1306.500 1579.680 1306.760 1579.940 ;
        RECT 1310.640 1579.680 1310.900 1579.940 ;
        RECT 1310.640 24.860 1310.900 25.120 ;
        RECT 2755.960 24.860 2756.220 25.120 ;
      LAYER met2 ;
        RECT 1304.980 1600.450 1305.260 1604.000 ;
        RECT 1304.980 1600.310 1306.700 1600.450 ;
        RECT 1304.980 1600.000 1305.260 1600.310 ;
        RECT 1306.560 1579.970 1306.700 1600.310 ;
        RECT 1306.500 1579.650 1306.760 1579.970 ;
        RECT 1310.640 1579.650 1310.900 1579.970 ;
        RECT 1310.700 25.150 1310.840 1579.650 ;
        RECT 1310.640 24.830 1310.900 25.150 ;
        RECT 2755.960 24.830 2756.220 25.150 ;
        RECT 2756.020 2.400 2756.160 24.830 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 637.170 1589.740 637.490 1589.800 ;
        RECT 641.310 1589.740 641.630 1589.800 ;
        RECT 637.170 1589.600 641.630 1589.740 ;
        RECT 637.170 1589.540 637.490 1589.600 ;
        RECT 641.310 1589.540 641.630 1589.600 ;
      LAYER via ;
        RECT 637.200 1589.540 637.460 1589.800 ;
        RECT 641.340 1589.540 641.600 1589.800 ;
      LAYER met2 ;
        RECT 637.060 1600.380 637.340 1604.000 ;
        RECT 637.060 1600.000 637.400 1600.380 ;
        RECT 637.260 1589.830 637.400 1600.000 ;
        RECT 637.200 1589.510 637.460 1589.830 ;
        RECT 641.340 1589.510 641.600 1589.830 ;
        RECT 641.400 17.525 641.540 1589.510 ;
        RECT 641.330 17.155 641.610 17.525 ;
        RECT 829.470 17.155 829.750 17.525 ;
        RECT 829.540 2.400 829.680 17.155 ;
        RECT 829.330 -4.800 829.890 2.400 ;
      LAYER via2 ;
        RECT 641.330 17.200 641.610 17.480 ;
        RECT 829.470 17.200 829.750 17.480 ;
      LAYER met3 ;
        RECT 641.305 17.490 641.635 17.505 ;
        RECT 829.445 17.490 829.775 17.505 ;
        RECT 641.305 17.190 829.775 17.490 ;
        RECT 641.305 17.175 641.635 17.190 ;
        RECT 829.445 17.175 829.775 17.190 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.530 1579.880 1311.850 1579.940 ;
        RECT 1311.530 1579.740 1312.220 1579.880 ;
        RECT 1311.530 1579.680 1311.850 1579.740 ;
        RECT 1312.080 1578.920 1312.220 1579.740 ;
        RECT 1311.990 1578.660 1312.310 1578.920 ;
        RECT 1311.990 1535.000 1312.310 1535.060 ;
        RECT 1317.510 1535.000 1317.830 1535.060 ;
        RECT 1311.990 1534.860 1317.830 1535.000 ;
        RECT 1311.990 1534.800 1312.310 1534.860 ;
        RECT 1317.510 1534.800 1317.830 1534.860 ;
      LAYER via ;
        RECT 1311.560 1579.680 1311.820 1579.940 ;
        RECT 1312.020 1578.660 1312.280 1578.920 ;
        RECT 1312.020 1534.800 1312.280 1535.060 ;
        RECT 1317.540 1534.800 1317.800 1535.060 ;
      LAYER met2 ;
        RECT 1311.420 1600.380 1311.700 1604.000 ;
        RECT 1311.420 1600.000 1311.760 1600.380 ;
        RECT 1311.620 1579.970 1311.760 1600.000 ;
        RECT 1311.560 1579.650 1311.820 1579.970 ;
        RECT 1312.020 1578.630 1312.280 1578.950 ;
        RECT 1312.080 1535.090 1312.220 1578.630 ;
        RECT 1312.020 1534.770 1312.280 1535.090 ;
        RECT 1317.540 1534.770 1317.800 1535.090 ;
        RECT 1317.600 27.045 1317.740 1534.770 ;
        RECT 1317.530 26.675 1317.810 27.045 ;
        RECT 2773.890 26.675 2774.170 27.045 ;
        RECT 2773.960 2.400 2774.100 26.675 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
      LAYER via2 ;
        RECT 1317.530 26.720 1317.810 27.000 ;
        RECT 2773.890 26.720 2774.170 27.000 ;
      LAYER met3 ;
        RECT 1317.505 27.010 1317.835 27.025 ;
        RECT 2773.865 27.010 2774.195 27.025 ;
        RECT 1317.505 26.710 2774.195 27.010 ;
        RECT 1317.505 26.695 1317.835 26.710 ;
        RECT 2773.865 26.695 2774.195 26.710 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1317.400 1601.130 1317.680 1604.000 ;
        RECT 1316.680 1600.990 1317.680 1601.130 ;
        RECT 1316.680 1597.050 1316.820 1600.990 ;
        RECT 1317.400 1600.000 1317.680 1600.990 ;
        RECT 1316.680 1596.910 1317.280 1597.050 ;
        RECT 1317.140 43.930 1317.280 1596.910 ;
        RECT 1316.220 43.790 1317.280 43.930 ;
        RECT 1316.220 26.365 1316.360 43.790 ;
        RECT 1316.150 25.995 1316.430 26.365 ;
        RECT 2791.830 25.995 2792.110 26.365 ;
        RECT 2791.900 2.400 2792.040 25.995 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
      LAYER via2 ;
        RECT 1316.150 26.040 1316.430 26.320 ;
        RECT 2791.830 26.040 2792.110 26.320 ;
      LAYER met3 ;
        RECT 1316.125 26.330 1316.455 26.345 ;
        RECT 2791.805 26.330 2792.135 26.345 ;
        RECT 1316.125 26.030 2792.135 26.330 ;
        RECT 1316.125 26.015 1316.455 26.030 ;
        RECT 2791.805 26.015 2792.135 26.030 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1324.410 25.400 1324.730 25.460 ;
        RECT 1324.410 25.260 1341.200 25.400 ;
        RECT 1324.410 25.200 1324.730 25.260 ;
        RECT 1341.060 24.720 1341.200 25.260 ;
        RECT 2809.750 24.720 2810.070 24.780 ;
        RECT 1341.060 24.580 2810.070 24.720 ;
        RECT 2809.750 24.520 2810.070 24.580 ;
      LAYER via ;
        RECT 1324.440 25.200 1324.700 25.460 ;
        RECT 2809.780 24.520 2810.040 24.780 ;
      LAYER met2 ;
        RECT 1323.840 1600.450 1324.120 1604.000 ;
        RECT 1323.840 1600.310 1324.640 1600.450 ;
        RECT 1323.840 1600.000 1324.120 1600.310 ;
        RECT 1324.500 25.490 1324.640 1600.310 ;
        RECT 1324.440 25.170 1324.700 25.490 ;
        RECT 2809.780 24.490 2810.040 24.810 ;
        RECT 2809.840 2.400 2809.980 24.490 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1329.820 1600.450 1330.100 1604.000 ;
        RECT 1329.820 1600.310 1331.540 1600.450 ;
        RECT 1329.820 1600.000 1330.100 1600.310 ;
        RECT 1331.400 25.685 1331.540 1600.310 ;
        RECT 1331.330 25.315 1331.610 25.685 ;
        RECT 2827.710 25.315 2827.990 25.685 ;
        RECT 2827.780 2.400 2827.920 25.315 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
      LAYER via2 ;
        RECT 1331.330 25.360 1331.610 25.640 ;
        RECT 2827.710 25.360 2827.990 25.640 ;
      LAYER met3 ;
        RECT 1331.305 25.650 1331.635 25.665 ;
        RECT 2827.685 25.650 2828.015 25.665 ;
        RECT 1331.305 25.350 2828.015 25.650 ;
        RECT 1331.305 25.335 1331.635 25.350 ;
        RECT 2827.685 25.335 2828.015 25.350 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1334.530 1587.020 1334.850 1587.080 ;
        RECT 1338.210 1587.020 1338.530 1587.080 ;
        RECT 1334.530 1586.880 1338.530 1587.020 ;
        RECT 1334.530 1586.820 1334.850 1586.880 ;
        RECT 1338.210 1586.820 1338.530 1586.880 ;
      LAYER via ;
        RECT 1334.560 1586.820 1334.820 1587.080 ;
        RECT 1338.240 1586.820 1338.500 1587.080 ;
      LAYER met2 ;
        RECT 1336.260 1600.450 1336.540 1604.000 ;
        RECT 1334.620 1600.310 1336.540 1600.450 ;
        RECT 1334.620 1587.110 1334.760 1600.310 ;
        RECT 1336.260 1600.000 1336.540 1600.310 ;
        RECT 1334.560 1586.790 1334.820 1587.110 ;
        RECT 1338.240 1586.790 1338.500 1587.110 ;
        RECT 1338.300 25.005 1338.440 1586.790 ;
        RECT 1338.230 24.635 1338.510 25.005 ;
        RECT 2845.190 24.635 2845.470 25.005 ;
        RECT 2845.260 2.400 2845.400 24.635 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
      LAYER via2 ;
        RECT 1338.230 24.680 1338.510 24.960 ;
        RECT 2845.190 24.680 2845.470 24.960 ;
      LAYER met3 ;
        RECT 1338.205 24.970 1338.535 24.985 ;
        RECT 2845.165 24.970 2845.495 24.985 ;
        RECT 1338.205 24.670 2845.495 24.970 ;
        RECT 1338.205 24.655 1338.535 24.670 ;
        RECT 2845.165 24.655 2845.495 24.670 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1344.190 1487.060 1344.510 1487.120 ;
        RECT 1345.110 1487.060 1345.430 1487.120 ;
        RECT 1344.190 1486.920 1345.430 1487.060 ;
        RECT 1344.190 1486.860 1344.510 1486.920 ;
        RECT 1345.110 1486.860 1345.430 1486.920 ;
        RECT 1344.190 1438.780 1344.510 1438.840 ;
        RECT 1345.110 1438.780 1345.430 1438.840 ;
        RECT 1344.190 1438.640 1345.430 1438.780 ;
        RECT 1344.190 1438.580 1344.510 1438.640 ;
        RECT 1345.110 1438.580 1345.430 1438.640 ;
        RECT 1344.190 1390.500 1344.510 1390.560 ;
        RECT 1345.110 1390.500 1345.430 1390.560 ;
        RECT 1344.190 1390.360 1345.430 1390.500 ;
        RECT 1344.190 1390.300 1344.510 1390.360 ;
        RECT 1345.110 1390.300 1345.430 1390.360 ;
        RECT 1343.730 1341.200 1344.050 1341.260 ;
        RECT 1345.110 1341.200 1345.430 1341.260 ;
        RECT 1343.730 1341.060 1345.430 1341.200 ;
        RECT 1343.730 1341.000 1344.050 1341.060 ;
        RECT 1345.110 1341.000 1345.430 1341.060 ;
        RECT 1343.730 1293.940 1344.050 1294.000 ;
        RECT 1345.110 1293.940 1345.430 1294.000 ;
        RECT 1343.730 1293.800 1345.430 1293.940 ;
        RECT 1343.730 1293.740 1344.050 1293.800 ;
        RECT 1345.110 1293.740 1345.430 1293.800 ;
        RECT 1343.730 1223.560 1344.050 1223.620 ;
        RECT 1345.110 1223.560 1345.430 1223.620 ;
        RECT 1343.730 1223.420 1345.430 1223.560 ;
        RECT 1343.730 1223.360 1344.050 1223.420 ;
        RECT 1345.110 1223.360 1345.430 1223.420 ;
        RECT 1343.730 1197.380 1344.050 1197.440 ;
        RECT 1345.110 1197.380 1345.430 1197.440 ;
        RECT 1343.730 1197.240 1345.430 1197.380 ;
        RECT 1343.730 1197.180 1344.050 1197.240 ;
        RECT 1345.110 1197.180 1345.430 1197.240 ;
        RECT 1343.730 1148.760 1344.050 1148.820 ;
        RECT 1345.110 1148.760 1345.430 1148.820 ;
        RECT 1343.730 1148.620 1345.430 1148.760 ;
        RECT 1343.730 1148.560 1344.050 1148.620 ;
        RECT 1345.110 1148.560 1345.430 1148.620 ;
        RECT 1343.730 1122.580 1344.050 1122.640 ;
        RECT 1345.110 1122.580 1345.430 1122.640 ;
        RECT 1343.730 1122.440 1345.430 1122.580 ;
        RECT 1343.730 1122.380 1344.050 1122.440 ;
        RECT 1345.110 1122.380 1345.430 1122.440 ;
        RECT 1343.730 1052.200 1344.050 1052.260 ;
        RECT 1345.110 1052.200 1345.430 1052.260 ;
        RECT 1343.730 1052.060 1345.430 1052.200 ;
        RECT 1343.730 1052.000 1344.050 1052.060 ;
        RECT 1345.110 1052.000 1345.430 1052.060 ;
        RECT 1343.730 1004.940 1344.050 1005.000 ;
        RECT 1345.110 1004.940 1345.430 1005.000 ;
        RECT 1343.730 1004.800 1345.430 1004.940 ;
        RECT 1343.730 1004.740 1344.050 1004.800 ;
        RECT 1345.110 1004.740 1345.430 1004.800 ;
        RECT 1343.730 955.640 1344.050 955.700 ;
        RECT 1345.110 955.640 1345.430 955.700 ;
        RECT 1343.730 955.500 1345.430 955.640 ;
        RECT 1343.730 955.440 1344.050 955.500 ;
        RECT 1345.110 955.440 1345.430 955.500 ;
        RECT 1343.730 907.360 1344.050 907.420 ;
        RECT 1345.110 907.360 1345.430 907.420 ;
        RECT 1343.730 907.220 1345.430 907.360 ;
        RECT 1343.730 907.160 1344.050 907.220 ;
        RECT 1345.110 907.160 1345.430 907.220 ;
        RECT 1343.730 858.060 1344.050 858.120 ;
        RECT 1345.110 858.060 1345.430 858.120 ;
        RECT 1343.730 857.920 1345.430 858.060 ;
        RECT 1343.730 857.860 1344.050 857.920 ;
        RECT 1345.110 857.860 1345.430 857.920 ;
        RECT 1343.730 811.820 1344.050 811.880 ;
        RECT 1345.110 811.820 1345.430 811.880 ;
        RECT 1343.730 811.680 1345.430 811.820 ;
        RECT 1343.730 811.620 1344.050 811.680 ;
        RECT 1345.110 811.620 1345.430 811.680 ;
        RECT 1343.730 762.520 1344.050 762.580 ;
        RECT 1345.110 762.520 1345.430 762.580 ;
        RECT 1343.730 762.380 1345.430 762.520 ;
        RECT 1343.730 762.320 1344.050 762.380 ;
        RECT 1345.110 762.320 1345.430 762.380 ;
        RECT 1343.730 714.240 1344.050 714.300 ;
        RECT 1345.110 714.240 1345.430 714.300 ;
        RECT 1343.730 714.100 1345.430 714.240 ;
        RECT 1343.730 714.040 1344.050 714.100 ;
        RECT 1345.110 714.040 1345.430 714.100 ;
        RECT 1343.730 665.960 1344.050 666.020 ;
        RECT 1345.110 665.960 1345.430 666.020 ;
        RECT 1343.730 665.820 1345.430 665.960 ;
        RECT 1343.730 665.760 1344.050 665.820 ;
        RECT 1345.110 665.760 1345.430 665.820 ;
        RECT 1343.730 617.680 1344.050 617.740 ;
        RECT 1345.110 617.680 1345.430 617.740 ;
        RECT 1343.730 617.540 1345.430 617.680 ;
        RECT 1343.730 617.480 1344.050 617.540 ;
        RECT 1345.110 617.480 1345.430 617.540 ;
        RECT 1343.730 569.400 1344.050 569.460 ;
        RECT 1345.110 569.400 1345.430 569.460 ;
        RECT 1343.730 569.260 1345.430 569.400 ;
        RECT 1343.730 569.200 1344.050 569.260 ;
        RECT 1345.110 569.200 1345.430 569.260 ;
        RECT 1343.730 542.880 1344.050 542.940 ;
        RECT 1345.110 542.880 1345.430 542.940 ;
        RECT 1343.730 542.740 1345.430 542.880 ;
        RECT 1343.730 542.680 1344.050 542.740 ;
        RECT 1345.110 542.680 1345.430 542.740 ;
        RECT 1343.730 471.820 1344.050 471.880 ;
        RECT 1345.110 471.820 1345.430 471.880 ;
        RECT 1343.730 471.680 1345.430 471.820 ;
        RECT 1343.730 471.620 1344.050 471.680 ;
        RECT 1345.110 471.620 1345.430 471.680 ;
        RECT 1343.730 424.560 1344.050 424.620 ;
        RECT 1345.110 424.560 1345.430 424.620 ;
        RECT 1343.730 424.420 1345.430 424.560 ;
        RECT 1343.730 424.360 1344.050 424.420 ;
        RECT 1345.110 424.360 1345.430 424.420 ;
        RECT 1343.730 375.600 1344.050 375.660 ;
        RECT 1345.110 375.600 1345.430 375.660 ;
        RECT 1343.730 375.460 1345.430 375.600 ;
        RECT 1343.730 375.400 1344.050 375.460 ;
        RECT 1345.110 375.400 1345.430 375.460 ;
        RECT 1343.730 327.660 1344.050 327.720 ;
        RECT 1345.110 327.660 1345.430 327.720 ;
        RECT 1343.730 327.520 1345.430 327.660 ;
        RECT 1343.730 327.460 1344.050 327.520 ;
        RECT 1345.110 327.460 1345.430 327.520 ;
        RECT 1343.730 279.380 1344.050 279.440 ;
        RECT 1345.110 279.380 1345.430 279.440 ;
        RECT 1343.730 279.240 1345.430 279.380 ;
        RECT 1343.730 279.180 1344.050 279.240 ;
        RECT 1345.110 279.180 1345.430 279.240 ;
        RECT 1343.730 231.100 1344.050 231.160 ;
        RECT 1345.110 231.100 1345.430 231.160 ;
        RECT 1343.730 230.960 1345.430 231.100 ;
        RECT 1343.730 230.900 1344.050 230.960 ;
        RECT 1345.110 230.900 1345.430 230.960 ;
        RECT 1343.730 161.060 1344.050 161.120 ;
        RECT 1345.110 161.060 1345.430 161.120 ;
        RECT 1343.730 160.920 1345.430 161.060 ;
        RECT 1343.730 160.860 1344.050 160.920 ;
        RECT 1345.110 160.860 1345.430 160.920 ;
        RECT 1343.730 134.540 1344.050 134.600 ;
        RECT 1345.110 134.540 1345.430 134.600 ;
        RECT 1343.730 134.400 1345.430 134.540 ;
        RECT 1343.730 134.340 1344.050 134.400 ;
        RECT 1345.110 134.340 1345.430 134.400 ;
        RECT 1343.730 86.260 1344.050 86.320 ;
        RECT 1345.110 86.260 1345.430 86.320 ;
        RECT 1343.730 86.120 1345.430 86.260 ;
        RECT 1343.730 86.060 1344.050 86.120 ;
        RECT 1345.110 86.060 1345.430 86.120 ;
        RECT 1343.730 24.380 1344.050 24.440 ;
        RECT 2863.110 24.380 2863.430 24.440 ;
        RECT 1343.730 24.240 2863.430 24.380 ;
        RECT 1343.730 24.180 1344.050 24.240 ;
        RECT 2863.110 24.180 2863.430 24.240 ;
      LAYER via ;
        RECT 1344.220 1486.860 1344.480 1487.120 ;
        RECT 1345.140 1486.860 1345.400 1487.120 ;
        RECT 1344.220 1438.580 1344.480 1438.840 ;
        RECT 1345.140 1438.580 1345.400 1438.840 ;
        RECT 1344.220 1390.300 1344.480 1390.560 ;
        RECT 1345.140 1390.300 1345.400 1390.560 ;
        RECT 1343.760 1341.000 1344.020 1341.260 ;
        RECT 1345.140 1341.000 1345.400 1341.260 ;
        RECT 1343.760 1293.740 1344.020 1294.000 ;
        RECT 1345.140 1293.740 1345.400 1294.000 ;
        RECT 1343.760 1223.360 1344.020 1223.620 ;
        RECT 1345.140 1223.360 1345.400 1223.620 ;
        RECT 1343.760 1197.180 1344.020 1197.440 ;
        RECT 1345.140 1197.180 1345.400 1197.440 ;
        RECT 1343.760 1148.560 1344.020 1148.820 ;
        RECT 1345.140 1148.560 1345.400 1148.820 ;
        RECT 1343.760 1122.380 1344.020 1122.640 ;
        RECT 1345.140 1122.380 1345.400 1122.640 ;
        RECT 1343.760 1052.000 1344.020 1052.260 ;
        RECT 1345.140 1052.000 1345.400 1052.260 ;
        RECT 1343.760 1004.740 1344.020 1005.000 ;
        RECT 1345.140 1004.740 1345.400 1005.000 ;
        RECT 1343.760 955.440 1344.020 955.700 ;
        RECT 1345.140 955.440 1345.400 955.700 ;
        RECT 1343.760 907.160 1344.020 907.420 ;
        RECT 1345.140 907.160 1345.400 907.420 ;
        RECT 1343.760 857.860 1344.020 858.120 ;
        RECT 1345.140 857.860 1345.400 858.120 ;
        RECT 1343.760 811.620 1344.020 811.880 ;
        RECT 1345.140 811.620 1345.400 811.880 ;
        RECT 1343.760 762.320 1344.020 762.580 ;
        RECT 1345.140 762.320 1345.400 762.580 ;
        RECT 1343.760 714.040 1344.020 714.300 ;
        RECT 1345.140 714.040 1345.400 714.300 ;
        RECT 1343.760 665.760 1344.020 666.020 ;
        RECT 1345.140 665.760 1345.400 666.020 ;
        RECT 1343.760 617.480 1344.020 617.740 ;
        RECT 1345.140 617.480 1345.400 617.740 ;
        RECT 1343.760 569.200 1344.020 569.460 ;
        RECT 1345.140 569.200 1345.400 569.460 ;
        RECT 1343.760 542.680 1344.020 542.940 ;
        RECT 1345.140 542.680 1345.400 542.940 ;
        RECT 1343.760 471.620 1344.020 471.880 ;
        RECT 1345.140 471.620 1345.400 471.880 ;
        RECT 1343.760 424.360 1344.020 424.620 ;
        RECT 1345.140 424.360 1345.400 424.620 ;
        RECT 1343.760 375.400 1344.020 375.660 ;
        RECT 1345.140 375.400 1345.400 375.660 ;
        RECT 1343.760 327.460 1344.020 327.720 ;
        RECT 1345.140 327.460 1345.400 327.720 ;
        RECT 1343.760 279.180 1344.020 279.440 ;
        RECT 1345.140 279.180 1345.400 279.440 ;
        RECT 1343.760 230.900 1344.020 231.160 ;
        RECT 1345.140 230.900 1345.400 231.160 ;
        RECT 1343.760 160.860 1344.020 161.120 ;
        RECT 1345.140 160.860 1345.400 161.120 ;
        RECT 1343.760 134.340 1344.020 134.600 ;
        RECT 1345.140 134.340 1345.400 134.600 ;
        RECT 1343.760 86.060 1344.020 86.320 ;
        RECT 1345.140 86.060 1345.400 86.320 ;
        RECT 1343.760 24.180 1344.020 24.440 ;
        RECT 2863.140 24.180 2863.400 24.440 ;
      LAYER met2 ;
        RECT 1342.240 1600.450 1342.520 1604.000 ;
        RECT 1342.240 1600.310 1343.960 1600.450 ;
        RECT 1342.240 1600.000 1342.520 1600.310 ;
        RECT 1343.820 1580.050 1343.960 1600.310 ;
        RECT 1343.820 1579.910 1345.340 1580.050 ;
        RECT 1345.200 1535.850 1345.340 1579.910 ;
        RECT 1344.280 1535.710 1345.340 1535.850 ;
        RECT 1344.280 1487.150 1344.420 1535.710 ;
        RECT 1344.220 1486.830 1344.480 1487.150 ;
        RECT 1345.140 1486.830 1345.400 1487.150 ;
        RECT 1345.200 1438.870 1345.340 1486.830 ;
        RECT 1344.220 1438.550 1344.480 1438.870 ;
        RECT 1345.140 1438.550 1345.400 1438.870 ;
        RECT 1344.280 1390.590 1344.420 1438.550 ;
        RECT 1344.220 1390.270 1344.480 1390.590 ;
        RECT 1345.140 1390.270 1345.400 1390.590 ;
        RECT 1345.200 1341.290 1345.340 1390.270 ;
        RECT 1343.760 1340.970 1344.020 1341.290 ;
        RECT 1345.140 1340.970 1345.400 1341.290 ;
        RECT 1343.820 1294.030 1343.960 1340.970 ;
        RECT 1343.760 1293.710 1344.020 1294.030 ;
        RECT 1345.140 1293.710 1345.400 1294.030 ;
        RECT 1345.200 1223.650 1345.340 1293.710 ;
        RECT 1343.760 1223.330 1344.020 1223.650 ;
        RECT 1345.140 1223.330 1345.400 1223.650 ;
        RECT 1343.820 1197.470 1343.960 1223.330 ;
        RECT 1343.760 1197.150 1344.020 1197.470 ;
        RECT 1345.140 1197.150 1345.400 1197.470 ;
        RECT 1345.200 1148.850 1345.340 1197.150 ;
        RECT 1343.760 1148.530 1344.020 1148.850 ;
        RECT 1345.140 1148.530 1345.400 1148.850 ;
        RECT 1343.820 1122.670 1343.960 1148.530 ;
        RECT 1343.760 1122.350 1344.020 1122.670 ;
        RECT 1345.140 1122.350 1345.400 1122.670 ;
        RECT 1345.200 1052.290 1345.340 1122.350 ;
        RECT 1343.760 1051.970 1344.020 1052.290 ;
        RECT 1345.140 1051.970 1345.400 1052.290 ;
        RECT 1343.820 1005.030 1343.960 1051.970 ;
        RECT 1343.760 1004.710 1344.020 1005.030 ;
        RECT 1345.140 1004.710 1345.400 1005.030 ;
        RECT 1345.200 955.730 1345.340 1004.710 ;
        RECT 1343.760 955.410 1344.020 955.730 ;
        RECT 1345.140 955.410 1345.400 955.730 ;
        RECT 1343.820 907.450 1343.960 955.410 ;
        RECT 1343.760 907.130 1344.020 907.450 ;
        RECT 1345.140 907.130 1345.400 907.450 ;
        RECT 1345.200 858.150 1345.340 907.130 ;
        RECT 1343.760 857.830 1344.020 858.150 ;
        RECT 1345.140 857.830 1345.400 858.150 ;
        RECT 1343.820 811.910 1343.960 857.830 ;
        RECT 1343.760 811.590 1344.020 811.910 ;
        RECT 1345.140 811.590 1345.400 811.910 ;
        RECT 1345.200 762.610 1345.340 811.590 ;
        RECT 1343.760 762.290 1344.020 762.610 ;
        RECT 1345.140 762.290 1345.400 762.610 ;
        RECT 1343.820 714.330 1343.960 762.290 ;
        RECT 1343.760 714.010 1344.020 714.330 ;
        RECT 1345.140 714.010 1345.400 714.330 ;
        RECT 1345.200 666.050 1345.340 714.010 ;
        RECT 1343.760 665.730 1344.020 666.050 ;
        RECT 1345.140 665.730 1345.400 666.050 ;
        RECT 1343.820 617.770 1343.960 665.730 ;
        RECT 1343.760 617.450 1344.020 617.770 ;
        RECT 1345.140 617.450 1345.400 617.770 ;
        RECT 1345.200 569.490 1345.340 617.450 ;
        RECT 1343.760 569.170 1344.020 569.490 ;
        RECT 1345.140 569.170 1345.400 569.490 ;
        RECT 1343.820 542.970 1343.960 569.170 ;
        RECT 1343.760 542.650 1344.020 542.970 ;
        RECT 1345.140 542.650 1345.400 542.970 ;
        RECT 1345.200 471.910 1345.340 542.650 ;
        RECT 1343.760 471.590 1344.020 471.910 ;
        RECT 1345.140 471.590 1345.400 471.910 ;
        RECT 1343.820 424.650 1343.960 471.590 ;
        RECT 1343.760 424.330 1344.020 424.650 ;
        RECT 1345.140 424.330 1345.400 424.650 ;
        RECT 1345.200 375.690 1345.340 424.330 ;
        RECT 1343.760 375.370 1344.020 375.690 ;
        RECT 1345.140 375.370 1345.400 375.690 ;
        RECT 1343.820 327.750 1343.960 375.370 ;
        RECT 1343.760 327.430 1344.020 327.750 ;
        RECT 1345.140 327.430 1345.400 327.750 ;
        RECT 1345.200 279.470 1345.340 327.430 ;
        RECT 1343.760 279.150 1344.020 279.470 ;
        RECT 1345.140 279.150 1345.400 279.470 ;
        RECT 1343.820 231.190 1343.960 279.150 ;
        RECT 1343.760 230.870 1344.020 231.190 ;
        RECT 1345.140 230.870 1345.400 231.190 ;
        RECT 1345.200 161.150 1345.340 230.870 ;
        RECT 1343.760 160.830 1344.020 161.150 ;
        RECT 1345.140 160.830 1345.400 161.150 ;
        RECT 1343.820 134.630 1343.960 160.830 ;
        RECT 1343.760 134.310 1344.020 134.630 ;
        RECT 1345.140 134.310 1345.400 134.630 ;
        RECT 1345.200 86.350 1345.340 134.310 ;
        RECT 1343.760 86.030 1344.020 86.350 ;
        RECT 1345.140 86.030 1345.400 86.350 ;
        RECT 1343.820 24.470 1343.960 86.030 ;
        RECT 1343.760 24.150 1344.020 24.470 ;
        RECT 2863.140 24.150 2863.400 24.470 ;
        RECT 2863.200 2.400 2863.340 24.150 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1348.680 1600.450 1348.960 1604.000 ;
        RECT 1348.680 1600.310 1349.940 1600.450 ;
        RECT 1348.680 1600.000 1348.960 1600.310 ;
        RECT 1349.800 1580.050 1349.940 1600.310 ;
        RECT 1349.800 1579.910 1352.240 1580.050 ;
        RECT 1352.100 24.325 1352.240 1579.910 ;
        RECT 1352.030 23.955 1352.310 24.325 ;
        RECT 2881.070 23.955 2881.350 24.325 ;
        RECT 2881.140 2.400 2881.280 23.955 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
      LAYER via2 ;
        RECT 1352.030 24.000 1352.310 24.280 ;
        RECT 2881.070 24.000 2881.350 24.280 ;
      LAYER met3 ;
        RECT 1352.005 24.290 1352.335 24.305 ;
        RECT 2881.045 24.290 2881.375 24.305 ;
        RECT 1352.005 23.990 2881.375 24.290 ;
        RECT 1352.005 23.975 1352.335 23.990 ;
        RECT 2881.045 23.975 2881.375 23.990 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1356.150 1579.880 1356.470 1579.940 ;
        RECT 1358.910 1579.880 1359.230 1579.940 ;
        RECT 1356.150 1579.740 1359.230 1579.880 ;
        RECT 1356.150 1579.680 1356.470 1579.740 ;
        RECT 1358.910 1579.680 1359.230 1579.740 ;
        RECT 1358.910 24.040 1359.230 24.100 ;
        RECT 2898.990 24.040 2899.310 24.100 ;
        RECT 1358.910 23.900 2899.310 24.040 ;
        RECT 1358.910 23.840 1359.230 23.900 ;
        RECT 2898.990 23.840 2899.310 23.900 ;
      LAYER via ;
        RECT 1356.180 1579.680 1356.440 1579.940 ;
        RECT 1358.940 1579.680 1359.200 1579.940 ;
        RECT 1358.940 23.840 1359.200 24.100 ;
        RECT 2899.020 23.840 2899.280 24.100 ;
      LAYER met2 ;
        RECT 1354.660 1600.450 1354.940 1604.000 ;
        RECT 1354.660 1600.310 1356.380 1600.450 ;
        RECT 1354.660 1600.000 1354.940 1600.310 ;
        RECT 1356.240 1579.970 1356.380 1600.310 ;
        RECT 1356.180 1579.650 1356.440 1579.970 ;
        RECT 1358.940 1579.650 1359.200 1579.970 ;
        RECT 1359.000 24.130 1359.140 1579.650 ;
        RECT 1358.940 23.810 1359.200 24.130 ;
        RECT 2899.020 23.810 2899.280 24.130 ;
        RECT 2899.080 2.400 2899.220 23.810 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 643.610 1589.740 643.930 1589.800 ;
        RECT 648.210 1589.740 648.530 1589.800 ;
        RECT 643.610 1589.600 648.530 1589.740 ;
        RECT 643.610 1589.540 643.930 1589.600 ;
        RECT 648.210 1589.540 648.530 1589.600 ;
        RECT 648.210 19.960 648.530 20.020 ;
        RECT 846.930 19.960 847.250 20.020 ;
        RECT 648.210 19.820 847.250 19.960 ;
        RECT 648.210 19.760 648.530 19.820 ;
        RECT 846.930 19.760 847.250 19.820 ;
      LAYER via ;
        RECT 643.640 1589.540 643.900 1589.800 ;
        RECT 648.240 1589.540 648.500 1589.800 ;
        RECT 648.240 19.760 648.500 20.020 ;
        RECT 846.960 19.760 847.220 20.020 ;
      LAYER met2 ;
        RECT 643.500 1600.380 643.780 1604.000 ;
        RECT 643.500 1600.000 643.840 1600.380 ;
        RECT 643.700 1589.830 643.840 1600.000 ;
        RECT 643.640 1589.510 643.900 1589.830 ;
        RECT 648.240 1589.510 648.500 1589.830 ;
        RECT 648.300 20.050 648.440 1589.510 ;
        RECT 648.240 19.730 648.500 20.050 ;
        RECT 846.960 19.730 847.220 20.050 ;
        RECT 847.020 2.400 847.160 19.730 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 649.590 1589.740 649.910 1589.800 ;
        RECT 655.110 1589.740 655.430 1589.800 ;
        RECT 649.590 1589.600 655.430 1589.740 ;
        RECT 649.590 1589.540 649.910 1589.600 ;
        RECT 655.110 1589.540 655.430 1589.600 ;
        RECT 655.110 18.940 655.430 19.000 ;
        RECT 864.870 18.940 865.190 19.000 ;
        RECT 655.110 18.800 865.190 18.940 ;
        RECT 655.110 18.740 655.430 18.800 ;
        RECT 864.870 18.740 865.190 18.800 ;
      LAYER via ;
        RECT 649.620 1589.540 649.880 1589.800 ;
        RECT 655.140 1589.540 655.400 1589.800 ;
        RECT 655.140 18.740 655.400 19.000 ;
        RECT 864.900 18.740 865.160 19.000 ;
      LAYER met2 ;
        RECT 649.480 1600.380 649.760 1604.000 ;
        RECT 649.480 1600.000 649.820 1600.380 ;
        RECT 649.680 1589.830 649.820 1600.000 ;
        RECT 649.620 1589.510 649.880 1589.830 ;
        RECT 655.140 1589.510 655.400 1589.830 ;
        RECT 655.200 19.030 655.340 1589.510 ;
        RECT 655.140 18.710 655.400 19.030 ;
        RECT 864.900 18.710 865.160 19.030 ;
        RECT 864.960 2.400 865.100 18.710 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 656.030 1589.400 656.350 1589.460 ;
        RECT 662.010 1589.400 662.330 1589.460 ;
        RECT 656.030 1589.260 662.330 1589.400 ;
        RECT 656.030 1589.200 656.350 1589.260 ;
        RECT 662.010 1589.200 662.330 1589.260 ;
        RECT 662.010 18.600 662.330 18.660 ;
        RECT 882.810 18.600 883.130 18.660 ;
        RECT 662.010 18.460 883.130 18.600 ;
        RECT 662.010 18.400 662.330 18.460 ;
        RECT 882.810 18.400 883.130 18.460 ;
      LAYER via ;
        RECT 656.060 1589.200 656.320 1589.460 ;
        RECT 662.040 1589.200 662.300 1589.460 ;
        RECT 662.040 18.400 662.300 18.660 ;
        RECT 882.840 18.400 883.100 18.660 ;
      LAYER met2 ;
        RECT 655.920 1600.380 656.200 1604.000 ;
        RECT 655.920 1600.000 656.260 1600.380 ;
        RECT 656.120 1589.490 656.260 1600.000 ;
        RECT 656.060 1589.170 656.320 1589.490 ;
        RECT 662.040 1589.170 662.300 1589.490 ;
        RECT 662.100 18.690 662.240 1589.170 ;
        RECT 662.040 18.370 662.300 18.690 ;
        RECT 882.840 18.370 883.100 18.690 ;
        RECT 882.900 2.400 883.040 18.370 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 696.585 1586.525 696.755 1588.055 ;
        RECT 703.945 1586.525 704.115 1588.055 ;
        RECT 714.525 1587.885 714.695 1588.735 ;
        RECT 759.145 14.365 759.315 15.555 ;
      LAYER mcon ;
        RECT 714.525 1588.565 714.695 1588.735 ;
        RECT 696.585 1587.885 696.755 1588.055 ;
        RECT 703.945 1587.885 704.115 1588.055 ;
        RECT 759.145 15.385 759.315 15.555 ;
      LAYER met1 ;
        RECT 660.630 1592.460 660.950 1592.520 ;
        RECT 662.010 1592.460 662.330 1592.520 ;
        RECT 660.630 1592.320 662.330 1592.460 ;
        RECT 660.630 1592.260 660.950 1592.320 ;
        RECT 662.010 1592.260 662.330 1592.320 ;
        RECT 714.465 1588.720 714.755 1588.765 ;
        RECT 727.790 1588.720 728.110 1588.780 ;
        RECT 714.465 1588.580 728.110 1588.720 ;
        RECT 714.465 1588.535 714.755 1588.580 ;
        RECT 727.790 1588.520 728.110 1588.580 ;
        RECT 660.630 1588.380 660.950 1588.440 ;
        RECT 660.630 1588.240 662.700 1588.380 ;
        RECT 660.630 1588.180 660.950 1588.240 ;
        RECT 662.560 1588.040 662.700 1588.240 ;
        RECT 696.525 1588.040 696.815 1588.085 ;
        RECT 662.560 1587.900 696.815 1588.040 ;
        RECT 696.525 1587.855 696.815 1587.900 ;
        RECT 703.885 1588.040 704.175 1588.085 ;
        RECT 714.465 1588.040 714.755 1588.085 ;
        RECT 703.885 1587.900 714.755 1588.040 ;
        RECT 703.885 1587.855 704.175 1587.900 ;
        RECT 714.465 1587.855 714.755 1587.900 ;
        RECT 696.525 1586.680 696.815 1586.725 ;
        RECT 703.885 1586.680 704.175 1586.725 ;
        RECT 696.525 1586.540 704.175 1586.680 ;
        RECT 696.525 1586.495 696.815 1586.540 ;
        RECT 703.885 1586.495 704.175 1586.540 ;
        RECT 727.330 15.540 727.650 15.600 ;
        RECT 759.085 15.540 759.375 15.585 ;
        RECT 727.330 15.400 759.375 15.540 ;
        RECT 727.330 15.340 727.650 15.400 ;
        RECT 759.085 15.355 759.375 15.400 ;
        RECT 759.085 14.520 759.375 14.565 ;
        RECT 900.750 14.520 901.070 14.580 ;
        RECT 759.085 14.380 901.070 14.520 ;
        RECT 759.085 14.335 759.375 14.380 ;
        RECT 900.750 14.320 901.070 14.380 ;
      LAYER via ;
        RECT 660.660 1592.260 660.920 1592.520 ;
        RECT 662.040 1592.260 662.300 1592.520 ;
        RECT 727.820 1588.520 728.080 1588.780 ;
        RECT 660.660 1588.180 660.920 1588.440 ;
        RECT 727.360 15.340 727.620 15.600 ;
        RECT 900.780 14.320 901.040 14.580 ;
      LAYER met2 ;
        RECT 661.900 1600.380 662.180 1604.000 ;
        RECT 661.900 1600.000 662.240 1600.380 ;
        RECT 662.100 1592.550 662.240 1600.000 ;
        RECT 660.660 1592.230 660.920 1592.550 ;
        RECT 662.040 1592.230 662.300 1592.550 ;
        RECT 660.720 1588.470 660.860 1592.230 ;
        RECT 727.820 1588.490 728.080 1588.810 ;
        RECT 660.660 1588.150 660.920 1588.470 ;
        RECT 727.880 24.210 728.020 1588.490 ;
        RECT 727.420 24.070 728.020 24.210 ;
        RECT 727.420 15.630 727.560 24.070 ;
        RECT 727.360 15.310 727.620 15.630 ;
        RECT 900.780 14.290 901.040 14.610 ;
        RECT 900.840 2.400 900.980 14.290 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 692.445 1587.205 692.615 1589.075 ;
        RECT 765.125 15.725 765.295 20.315 ;
        RECT 786.285 15.725 786.455 20.655 ;
      LAYER mcon ;
        RECT 692.445 1588.905 692.615 1589.075 ;
        RECT 786.285 20.485 786.455 20.655 ;
        RECT 765.125 20.145 765.295 20.315 ;
      LAYER met1 ;
        RECT 692.385 1589.060 692.675 1589.105 ;
        RECT 741.590 1589.060 741.910 1589.120 ;
        RECT 692.385 1588.920 741.910 1589.060 ;
        RECT 692.385 1588.875 692.675 1588.920 ;
        RECT 741.590 1588.860 741.910 1588.920 ;
        RECT 668.450 1587.360 668.770 1587.420 ;
        RECT 692.385 1587.360 692.675 1587.405 ;
        RECT 668.450 1587.220 692.675 1587.360 ;
        RECT 668.450 1587.160 668.770 1587.220 ;
        RECT 692.385 1587.175 692.675 1587.220 ;
        RECT 786.225 20.640 786.515 20.685 ;
        RECT 918.690 20.640 919.010 20.700 ;
        RECT 786.225 20.500 919.010 20.640 ;
        RECT 786.225 20.455 786.515 20.500 ;
        RECT 918.690 20.440 919.010 20.500 ;
        RECT 741.590 20.300 741.910 20.360 ;
        RECT 765.065 20.300 765.355 20.345 ;
        RECT 741.590 20.160 765.355 20.300 ;
        RECT 741.590 20.100 741.910 20.160 ;
        RECT 765.065 20.115 765.355 20.160 ;
        RECT 765.065 15.880 765.355 15.925 ;
        RECT 786.225 15.880 786.515 15.925 ;
        RECT 765.065 15.740 786.515 15.880 ;
        RECT 765.065 15.695 765.355 15.740 ;
        RECT 786.225 15.695 786.515 15.740 ;
      LAYER via ;
        RECT 741.620 1588.860 741.880 1589.120 ;
        RECT 668.480 1587.160 668.740 1587.420 ;
        RECT 918.720 20.440 918.980 20.700 ;
        RECT 741.620 20.100 741.880 20.360 ;
      LAYER met2 ;
        RECT 668.340 1600.380 668.620 1604.000 ;
        RECT 668.340 1600.000 668.680 1600.380 ;
        RECT 668.540 1587.450 668.680 1600.000 ;
        RECT 741.620 1588.830 741.880 1589.150 ;
        RECT 668.480 1587.130 668.740 1587.450 ;
        RECT 741.680 20.390 741.820 1588.830 ;
        RECT 918.720 20.410 918.980 20.730 ;
        RECT 741.620 20.070 741.880 20.390 ;
        RECT 918.780 2.400 918.920 20.410 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 714.065 1588.565 714.235 1589.415 ;
        RECT 736.605 1545.725 736.775 1589.415 ;
        RECT 755.465 1449.165 755.635 1497.275 ;
        RECT 755.465 1352.605 755.635 1400.715 ;
        RECT 755.465 1256.045 755.635 1304.155 ;
        RECT 755.465 772.905 755.635 821.015 ;
        RECT 755.465 676.345 755.635 724.455 ;
        RECT 755.465 579.785 755.635 627.895 ;
        RECT 755.465 483.225 755.635 531.335 ;
        RECT 755.465 386.325 755.635 434.775 ;
        RECT 755.465 289.765 755.635 337.875 ;
        RECT 755.465 193.205 755.635 241.315 ;
        RECT 755.465 96.645 755.635 144.755 ;
      LAYER mcon ;
        RECT 714.065 1589.245 714.235 1589.415 ;
        RECT 736.605 1589.245 736.775 1589.415 ;
        RECT 755.465 1497.105 755.635 1497.275 ;
        RECT 755.465 1400.545 755.635 1400.715 ;
        RECT 755.465 1303.985 755.635 1304.155 ;
        RECT 755.465 820.845 755.635 821.015 ;
        RECT 755.465 724.285 755.635 724.455 ;
        RECT 755.465 627.725 755.635 627.895 ;
        RECT 755.465 531.165 755.635 531.335 ;
        RECT 755.465 434.605 755.635 434.775 ;
        RECT 755.465 337.705 755.635 337.875 ;
        RECT 755.465 241.145 755.635 241.315 ;
        RECT 755.465 144.585 755.635 144.755 ;
      LAYER met1 ;
        RECT 714.005 1589.400 714.295 1589.445 ;
        RECT 736.545 1589.400 736.835 1589.445 ;
        RECT 714.005 1589.260 736.835 1589.400 ;
        RECT 714.005 1589.215 714.295 1589.260 ;
        RECT 736.545 1589.215 736.835 1589.260 ;
        RECT 674.430 1588.720 674.750 1588.780 ;
        RECT 714.005 1588.720 714.295 1588.765 ;
        RECT 674.430 1588.580 714.295 1588.720 ;
        RECT 674.430 1588.520 674.750 1588.580 ;
        RECT 714.005 1588.535 714.295 1588.580 ;
        RECT 736.545 1545.880 736.835 1545.925 ;
        RECT 755.390 1545.880 755.710 1545.940 ;
        RECT 736.545 1545.740 755.710 1545.880 ;
        RECT 736.545 1545.695 736.835 1545.740 ;
        RECT 755.390 1545.680 755.710 1545.740 ;
        RECT 755.390 1497.260 755.710 1497.320 ;
        RECT 755.195 1497.120 755.710 1497.260 ;
        RECT 755.390 1497.060 755.710 1497.120 ;
        RECT 755.390 1449.320 755.710 1449.380 ;
        RECT 755.195 1449.180 755.710 1449.320 ;
        RECT 755.390 1449.120 755.710 1449.180 ;
        RECT 755.390 1400.700 755.710 1400.760 ;
        RECT 755.195 1400.560 755.710 1400.700 ;
        RECT 755.390 1400.500 755.710 1400.560 ;
        RECT 755.390 1352.760 755.710 1352.820 ;
        RECT 755.195 1352.620 755.710 1352.760 ;
        RECT 755.390 1352.560 755.710 1352.620 ;
        RECT 755.390 1304.140 755.710 1304.200 ;
        RECT 755.195 1304.000 755.710 1304.140 ;
        RECT 755.390 1303.940 755.710 1304.000 ;
        RECT 755.390 1256.200 755.710 1256.260 ;
        RECT 755.195 1256.060 755.710 1256.200 ;
        RECT 755.390 1256.000 755.710 1256.060 ;
        RECT 754.930 1159.300 755.250 1159.360 ;
        RECT 755.390 1159.300 755.710 1159.360 ;
        RECT 754.930 1159.160 755.710 1159.300 ;
        RECT 754.930 1159.100 755.250 1159.160 ;
        RECT 755.390 1159.100 755.710 1159.160 ;
        RECT 754.930 1062.740 755.250 1062.800 ;
        RECT 755.390 1062.740 755.710 1062.800 ;
        RECT 754.930 1062.600 755.710 1062.740 ;
        RECT 754.930 1062.540 755.250 1062.600 ;
        RECT 755.390 1062.540 755.710 1062.600 ;
        RECT 754.930 966.180 755.250 966.240 ;
        RECT 755.390 966.180 755.710 966.240 ;
        RECT 754.930 966.040 755.710 966.180 ;
        RECT 754.930 965.980 755.250 966.040 ;
        RECT 755.390 965.980 755.710 966.040 ;
        RECT 754.930 869.620 755.250 869.680 ;
        RECT 755.390 869.620 755.710 869.680 ;
        RECT 754.930 869.480 755.710 869.620 ;
        RECT 754.930 869.420 755.250 869.480 ;
        RECT 755.390 869.420 755.710 869.480 ;
        RECT 755.390 821.000 755.710 821.060 ;
        RECT 755.195 820.860 755.710 821.000 ;
        RECT 755.390 820.800 755.710 820.860 ;
        RECT 755.390 773.060 755.710 773.120 ;
        RECT 755.195 772.920 755.710 773.060 ;
        RECT 755.390 772.860 755.710 772.920 ;
        RECT 755.390 724.440 755.710 724.500 ;
        RECT 755.195 724.300 755.710 724.440 ;
        RECT 755.390 724.240 755.710 724.300 ;
        RECT 755.390 676.500 755.710 676.560 ;
        RECT 755.195 676.360 755.710 676.500 ;
        RECT 755.390 676.300 755.710 676.360 ;
        RECT 755.390 627.880 755.710 627.940 ;
        RECT 755.195 627.740 755.710 627.880 ;
        RECT 755.390 627.680 755.710 627.740 ;
        RECT 755.390 579.940 755.710 580.000 ;
        RECT 755.195 579.800 755.710 579.940 ;
        RECT 755.390 579.740 755.710 579.800 ;
        RECT 755.390 531.320 755.710 531.380 ;
        RECT 755.195 531.180 755.710 531.320 ;
        RECT 755.390 531.120 755.710 531.180 ;
        RECT 755.390 483.380 755.710 483.440 ;
        RECT 755.195 483.240 755.710 483.380 ;
        RECT 755.390 483.180 755.710 483.240 ;
        RECT 755.390 434.760 755.710 434.820 ;
        RECT 755.195 434.620 755.710 434.760 ;
        RECT 755.390 434.560 755.710 434.620 ;
        RECT 755.390 386.480 755.710 386.540 ;
        RECT 755.195 386.340 755.710 386.480 ;
        RECT 755.390 386.280 755.710 386.340 ;
        RECT 755.390 337.860 755.710 337.920 ;
        RECT 755.195 337.720 755.710 337.860 ;
        RECT 755.390 337.660 755.710 337.720 ;
        RECT 755.390 289.920 755.710 289.980 ;
        RECT 755.195 289.780 755.710 289.920 ;
        RECT 755.390 289.720 755.710 289.780 ;
        RECT 755.390 241.300 755.710 241.360 ;
        RECT 755.195 241.160 755.710 241.300 ;
        RECT 755.390 241.100 755.710 241.160 ;
        RECT 755.390 193.360 755.710 193.420 ;
        RECT 755.195 193.220 755.710 193.360 ;
        RECT 755.390 193.160 755.710 193.220 ;
        RECT 755.390 144.740 755.710 144.800 ;
        RECT 755.195 144.600 755.710 144.740 ;
        RECT 755.390 144.540 755.710 144.600 ;
        RECT 755.390 96.800 755.710 96.860 ;
        RECT 755.195 96.660 755.710 96.800 ;
        RECT 755.390 96.600 755.710 96.660 ;
        RECT 765.970 15.200 766.290 15.260 ;
        RECT 936.170 15.200 936.490 15.260 ;
        RECT 765.970 15.060 936.490 15.200 ;
        RECT 765.970 15.000 766.290 15.060 ;
        RECT 936.170 15.000 936.490 15.060 ;
      LAYER via ;
        RECT 674.460 1588.520 674.720 1588.780 ;
        RECT 755.420 1545.680 755.680 1545.940 ;
        RECT 755.420 1497.060 755.680 1497.320 ;
        RECT 755.420 1449.120 755.680 1449.380 ;
        RECT 755.420 1400.500 755.680 1400.760 ;
        RECT 755.420 1352.560 755.680 1352.820 ;
        RECT 755.420 1303.940 755.680 1304.200 ;
        RECT 755.420 1256.000 755.680 1256.260 ;
        RECT 754.960 1159.100 755.220 1159.360 ;
        RECT 755.420 1159.100 755.680 1159.360 ;
        RECT 754.960 1062.540 755.220 1062.800 ;
        RECT 755.420 1062.540 755.680 1062.800 ;
        RECT 754.960 965.980 755.220 966.240 ;
        RECT 755.420 965.980 755.680 966.240 ;
        RECT 754.960 869.420 755.220 869.680 ;
        RECT 755.420 869.420 755.680 869.680 ;
        RECT 755.420 820.800 755.680 821.060 ;
        RECT 755.420 772.860 755.680 773.120 ;
        RECT 755.420 724.240 755.680 724.500 ;
        RECT 755.420 676.300 755.680 676.560 ;
        RECT 755.420 627.680 755.680 627.940 ;
        RECT 755.420 579.740 755.680 580.000 ;
        RECT 755.420 531.120 755.680 531.380 ;
        RECT 755.420 483.180 755.680 483.440 ;
        RECT 755.420 434.560 755.680 434.820 ;
        RECT 755.420 386.280 755.680 386.540 ;
        RECT 755.420 337.660 755.680 337.920 ;
        RECT 755.420 289.720 755.680 289.980 ;
        RECT 755.420 241.100 755.680 241.360 ;
        RECT 755.420 193.160 755.680 193.420 ;
        RECT 755.420 144.540 755.680 144.800 ;
        RECT 755.420 96.600 755.680 96.860 ;
        RECT 766.000 15.000 766.260 15.260 ;
        RECT 936.200 15.000 936.460 15.260 ;
      LAYER met2 ;
        RECT 674.320 1600.380 674.600 1604.000 ;
        RECT 674.320 1600.000 674.660 1600.380 ;
        RECT 674.520 1588.810 674.660 1600.000 ;
        RECT 674.460 1588.490 674.720 1588.810 ;
        RECT 755.420 1545.650 755.680 1545.970 ;
        RECT 755.480 1497.350 755.620 1545.650 ;
        RECT 755.420 1497.030 755.680 1497.350 ;
        RECT 755.420 1449.090 755.680 1449.410 ;
        RECT 755.480 1400.790 755.620 1449.090 ;
        RECT 755.420 1400.470 755.680 1400.790 ;
        RECT 755.420 1352.530 755.680 1352.850 ;
        RECT 755.480 1304.230 755.620 1352.530 ;
        RECT 755.420 1303.910 755.680 1304.230 ;
        RECT 755.420 1255.970 755.680 1256.290 ;
        RECT 755.480 1207.525 755.620 1255.970 ;
        RECT 755.410 1207.155 755.690 1207.525 ;
        RECT 754.950 1206.475 755.230 1206.845 ;
        RECT 755.020 1159.390 755.160 1206.475 ;
        RECT 754.960 1159.070 755.220 1159.390 ;
        RECT 755.420 1159.070 755.680 1159.390 ;
        RECT 755.480 1110.965 755.620 1159.070 ;
        RECT 755.410 1110.595 755.690 1110.965 ;
        RECT 754.950 1109.915 755.230 1110.285 ;
        RECT 755.020 1062.830 755.160 1109.915 ;
        RECT 754.960 1062.510 755.220 1062.830 ;
        RECT 755.420 1062.510 755.680 1062.830 ;
        RECT 755.480 1014.405 755.620 1062.510 ;
        RECT 755.410 1014.035 755.690 1014.405 ;
        RECT 754.950 1013.355 755.230 1013.725 ;
        RECT 755.020 966.270 755.160 1013.355 ;
        RECT 754.960 965.950 755.220 966.270 ;
        RECT 755.420 965.950 755.680 966.270 ;
        RECT 755.480 917.845 755.620 965.950 ;
        RECT 755.410 917.475 755.690 917.845 ;
        RECT 754.950 916.795 755.230 917.165 ;
        RECT 755.020 869.710 755.160 916.795 ;
        RECT 754.960 869.390 755.220 869.710 ;
        RECT 755.420 869.390 755.680 869.710 ;
        RECT 755.480 821.090 755.620 869.390 ;
        RECT 755.420 820.770 755.680 821.090 ;
        RECT 755.420 772.830 755.680 773.150 ;
        RECT 755.480 724.530 755.620 772.830 ;
        RECT 755.420 724.210 755.680 724.530 ;
        RECT 755.420 676.270 755.680 676.590 ;
        RECT 755.480 627.970 755.620 676.270 ;
        RECT 755.420 627.650 755.680 627.970 ;
        RECT 755.420 579.710 755.680 580.030 ;
        RECT 755.480 531.410 755.620 579.710 ;
        RECT 755.420 531.090 755.680 531.410 ;
        RECT 755.420 483.150 755.680 483.470 ;
        RECT 755.480 434.850 755.620 483.150 ;
        RECT 755.420 434.530 755.680 434.850 ;
        RECT 755.420 386.250 755.680 386.570 ;
        RECT 755.480 337.950 755.620 386.250 ;
        RECT 755.420 337.630 755.680 337.950 ;
        RECT 755.420 289.690 755.680 290.010 ;
        RECT 755.480 241.390 755.620 289.690 ;
        RECT 755.420 241.070 755.680 241.390 ;
        RECT 755.420 193.130 755.680 193.450 ;
        RECT 755.480 144.830 755.620 193.130 ;
        RECT 755.420 144.510 755.680 144.830 ;
        RECT 755.420 96.570 755.680 96.890 ;
        RECT 755.480 48.295 755.620 96.570 ;
        RECT 755.410 47.925 755.690 48.295 ;
        RECT 765.990 47.075 766.270 47.445 ;
        RECT 766.060 15.290 766.200 47.075 ;
        RECT 766.000 14.970 766.260 15.290 ;
        RECT 936.200 14.970 936.460 15.290 ;
        RECT 936.260 2.400 936.400 14.970 ;
        RECT 936.050 -4.800 936.610 2.400 ;
      LAYER via2 ;
        RECT 755.410 1207.200 755.690 1207.480 ;
        RECT 754.950 1206.520 755.230 1206.800 ;
        RECT 755.410 1110.640 755.690 1110.920 ;
        RECT 754.950 1109.960 755.230 1110.240 ;
        RECT 755.410 1014.080 755.690 1014.360 ;
        RECT 754.950 1013.400 755.230 1013.680 ;
        RECT 755.410 917.520 755.690 917.800 ;
        RECT 754.950 916.840 755.230 917.120 ;
        RECT 755.410 47.970 755.690 48.250 ;
        RECT 765.990 47.120 766.270 47.400 ;
      LAYER met3 ;
        RECT 755.385 1207.490 755.715 1207.505 ;
        RECT 755.385 1207.175 755.930 1207.490 ;
        RECT 754.925 1206.810 755.255 1206.825 ;
        RECT 755.630 1206.810 755.930 1207.175 ;
        RECT 754.925 1206.510 755.930 1206.810 ;
        RECT 754.925 1206.495 755.255 1206.510 ;
        RECT 755.385 1110.930 755.715 1110.945 ;
        RECT 755.385 1110.615 755.930 1110.930 ;
        RECT 754.925 1110.250 755.255 1110.265 ;
        RECT 755.630 1110.250 755.930 1110.615 ;
        RECT 754.925 1109.950 755.930 1110.250 ;
        RECT 754.925 1109.935 755.255 1109.950 ;
        RECT 755.385 1014.370 755.715 1014.385 ;
        RECT 755.385 1014.055 755.930 1014.370 ;
        RECT 754.925 1013.690 755.255 1013.705 ;
        RECT 755.630 1013.690 755.930 1014.055 ;
        RECT 754.925 1013.390 755.930 1013.690 ;
        RECT 754.925 1013.375 755.255 1013.390 ;
        RECT 755.385 917.810 755.715 917.825 ;
        RECT 755.385 917.495 755.930 917.810 ;
        RECT 754.925 917.130 755.255 917.145 ;
        RECT 755.630 917.130 755.930 917.495 ;
        RECT 754.925 916.830 755.930 917.130 ;
        RECT 754.925 916.815 755.255 916.830 ;
        RECT 755.385 48.260 755.715 48.275 ;
        RECT 754.710 47.960 755.715 48.260 ;
        RECT 754.710 47.410 755.010 47.960 ;
        RECT 755.385 47.945 755.715 47.960 ;
        RECT 765.965 47.410 766.295 47.425 ;
        RECT 754.710 47.110 766.295 47.410 ;
        RECT 765.965 47.095 766.295 47.110 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 709.925 1588.225 710.095 1589.415 ;
        RECT 776.165 16.745 776.335 19.635 ;
      LAYER mcon ;
        RECT 709.925 1589.245 710.095 1589.415 ;
        RECT 776.165 19.465 776.335 19.635 ;
      LAYER met1 ;
        RECT 680.870 1589.400 681.190 1589.460 ;
        RECT 709.865 1589.400 710.155 1589.445 ;
        RECT 680.870 1589.260 710.155 1589.400 ;
        RECT 680.870 1589.200 681.190 1589.260 ;
        RECT 709.865 1589.215 710.155 1589.260 ;
        RECT 709.865 1588.380 710.155 1588.425 ;
        RECT 709.865 1588.240 724.800 1588.380 ;
        RECT 709.865 1588.195 710.155 1588.240 ;
        RECT 724.660 1588.040 724.800 1588.240 ;
        RECT 755.390 1588.040 755.710 1588.100 ;
        RECT 724.660 1587.900 755.710 1588.040 ;
        RECT 755.390 1587.840 755.710 1587.900 ;
        RECT 776.105 19.620 776.395 19.665 ;
        RECT 954.110 19.620 954.430 19.680 ;
        RECT 776.105 19.480 954.430 19.620 ;
        RECT 776.105 19.435 776.395 19.480 ;
        RECT 954.110 19.420 954.430 19.480 ;
        RECT 756.310 16.900 756.630 16.960 ;
        RECT 776.105 16.900 776.395 16.945 ;
        RECT 756.310 16.760 776.395 16.900 ;
        RECT 756.310 16.700 756.630 16.760 ;
        RECT 776.105 16.715 776.395 16.760 ;
      LAYER via ;
        RECT 680.900 1589.200 681.160 1589.460 ;
        RECT 755.420 1587.840 755.680 1588.100 ;
        RECT 954.140 19.420 954.400 19.680 ;
        RECT 756.340 16.700 756.600 16.960 ;
      LAYER met2 ;
        RECT 680.760 1600.380 681.040 1604.000 ;
        RECT 680.760 1600.000 681.100 1600.380 ;
        RECT 680.960 1589.490 681.100 1600.000 ;
        RECT 680.900 1589.170 681.160 1589.490 ;
        RECT 755.420 1587.810 755.680 1588.130 ;
        RECT 755.480 1563.730 755.620 1587.810 ;
        RECT 755.480 1563.590 756.540 1563.730 ;
        RECT 756.400 16.990 756.540 1563.590 ;
        RECT 954.140 19.390 954.400 19.710 ;
        RECT 756.340 16.670 756.600 16.990 ;
        RECT 954.200 2.400 954.340 19.390 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 691.985 1588.905 692.155 1590.775 ;
      LAYER mcon ;
        RECT 691.985 1590.605 692.155 1590.775 ;
      LAYER met1 ;
        RECT 762.290 1591.440 762.610 1591.500 ;
        RECT 738.920 1591.300 762.610 1591.440 ;
        RECT 691.925 1590.760 692.215 1590.805 ;
        RECT 738.920 1590.760 739.060 1591.300 ;
        RECT 762.290 1591.240 762.610 1591.300 ;
        RECT 691.925 1590.620 739.060 1590.760 ;
        RECT 691.925 1590.575 692.215 1590.620 ;
        RECT 686.850 1589.060 687.170 1589.120 ;
        RECT 691.925 1589.060 692.215 1589.105 ;
        RECT 686.850 1588.920 692.215 1589.060 ;
        RECT 686.850 1588.860 687.170 1588.920 ;
        RECT 691.925 1588.875 692.215 1588.920 ;
        RECT 762.290 19.280 762.610 19.340 ;
        RECT 972.050 19.280 972.370 19.340 ;
        RECT 762.290 19.140 972.370 19.280 ;
        RECT 762.290 19.080 762.610 19.140 ;
        RECT 972.050 19.080 972.370 19.140 ;
      LAYER via ;
        RECT 762.320 1591.240 762.580 1591.500 ;
        RECT 686.880 1588.860 687.140 1589.120 ;
        RECT 762.320 19.080 762.580 19.340 ;
        RECT 972.080 19.080 972.340 19.340 ;
      LAYER met2 ;
        RECT 686.740 1600.380 687.020 1604.000 ;
        RECT 686.740 1600.000 687.080 1600.380 ;
        RECT 686.940 1589.150 687.080 1600.000 ;
        RECT 762.320 1591.210 762.580 1591.530 ;
        RECT 686.880 1588.830 687.140 1589.150 ;
        RECT 762.380 19.370 762.520 1591.210 ;
        RECT 762.320 19.050 762.580 19.370 ;
        RECT 972.080 19.050 972.340 19.370 ;
        RECT 972.140 2.400 972.280 19.050 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 575.530 1589.400 575.850 1589.460 ;
        RECT 579.210 1589.400 579.530 1589.460 ;
        RECT 575.530 1589.260 579.530 1589.400 ;
        RECT 575.530 1589.200 575.850 1589.260 ;
        RECT 579.210 1589.200 579.530 1589.260 ;
        RECT 579.210 18.940 579.530 19.000 ;
        RECT 650.970 18.940 651.290 19.000 ;
        RECT 579.210 18.800 651.290 18.940 ;
        RECT 579.210 18.740 579.530 18.800 ;
        RECT 650.970 18.740 651.290 18.800 ;
      LAYER via ;
        RECT 575.560 1589.200 575.820 1589.460 ;
        RECT 579.240 1589.200 579.500 1589.460 ;
        RECT 579.240 18.740 579.500 19.000 ;
        RECT 651.000 18.740 651.260 19.000 ;
      LAYER met2 ;
        RECT 575.420 1600.380 575.700 1604.000 ;
        RECT 575.420 1600.000 575.760 1600.380 ;
        RECT 575.620 1589.490 575.760 1600.000 ;
        RECT 575.560 1589.170 575.820 1589.490 ;
        RECT 579.240 1589.170 579.500 1589.490 ;
        RECT 579.300 19.030 579.440 1589.170 ;
        RECT 579.240 18.710 579.500 19.030 ;
        RECT 651.000 18.710 651.260 19.030 ;
        RECT 651.060 2.400 651.200 18.710 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 692.830 1587.360 693.150 1587.420 ;
        RECT 696.510 1587.360 696.830 1587.420 ;
        RECT 692.830 1587.220 696.830 1587.360 ;
        RECT 692.830 1587.160 693.150 1587.220 ;
        RECT 696.510 1587.160 696.830 1587.220 ;
        RECT 696.510 21.320 696.830 21.380 ;
        RECT 989.990 21.320 990.310 21.380 ;
        RECT 696.510 21.180 990.310 21.320 ;
        RECT 696.510 21.120 696.830 21.180 ;
        RECT 989.990 21.120 990.310 21.180 ;
      LAYER via ;
        RECT 692.860 1587.160 693.120 1587.420 ;
        RECT 696.540 1587.160 696.800 1587.420 ;
        RECT 696.540 21.120 696.800 21.380 ;
        RECT 990.020 21.120 990.280 21.380 ;
      LAYER met2 ;
        RECT 692.720 1600.380 693.000 1604.000 ;
        RECT 692.720 1600.000 693.060 1600.380 ;
        RECT 692.920 1587.450 693.060 1600.000 ;
        RECT 692.860 1587.130 693.120 1587.450 ;
        RECT 696.540 1587.130 696.800 1587.450 ;
        RECT 696.600 21.410 696.740 1587.130 ;
        RECT 696.540 21.090 696.800 21.410 ;
        RECT 990.020 21.090 990.280 21.410 ;
        RECT 990.080 2.400 990.220 21.090 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 699.270 1587.360 699.590 1587.420 ;
        RECT 702.950 1587.360 703.270 1587.420 ;
        RECT 699.270 1587.220 703.270 1587.360 ;
        RECT 699.270 1587.160 699.590 1587.220 ;
        RECT 702.950 1587.160 703.270 1587.220 ;
        RECT 702.950 21.660 703.270 21.720 ;
        RECT 1007.470 21.660 1007.790 21.720 ;
        RECT 702.950 21.520 1007.790 21.660 ;
        RECT 702.950 21.460 703.270 21.520 ;
        RECT 1007.470 21.460 1007.790 21.520 ;
      LAYER via ;
        RECT 699.300 1587.160 699.560 1587.420 ;
        RECT 702.980 1587.160 703.240 1587.420 ;
        RECT 702.980 21.460 703.240 21.720 ;
        RECT 1007.500 21.460 1007.760 21.720 ;
      LAYER met2 ;
        RECT 699.160 1600.380 699.440 1604.000 ;
        RECT 699.160 1600.000 699.500 1600.380 ;
        RECT 699.360 1587.450 699.500 1600.000 ;
        RECT 699.300 1587.130 699.560 1587.450 ;
        RECT 702.980 1587.130 703.240 1587.450 ;
        RECT 703.040 21.750 703.180 1587.130 ;
        RECT 702.980 21.430 703.240 21.750 ;
        RECT 1007.500 21.430 1007.760 21.750 ;
        RECT 1007.560 2.400 1007.700 21.430 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 705.250 1587.360 705.570 1587.420 ;
        RECT 710.310 1587.360 710.630 1587.420 ;
        RECT 705.250 1587.220 710.630 1587.360 ;
        RECT 705.250 1587.160 705.570 1587.220 ;
        RECT 710.310 1587.160 710.630 1587.220 ;
        RECT 710.310 22.000 710.630 22.060 ;
        RECT 1025.410 22.000 1025.730 22.060 ;
        RECT 710.310 21.860 1025.730 22.000 ;
        RECT 710.310 21.800 710.630 21.860 ;
        RECT 1025.410 21.800 1025.730 21.860 ;
      LAYER via ;
        RECT 705.280 1587.160 705.540 1587.420 ;
        RECT 710.340 1587.160 710.600 1587.420 ;
        RECT 710.340 21.800 710.600 22.060 ;
        RECT 1025.440 21.800 1025.700 22.060 ;
      LAYER met2 ;
        RECT 705.140 1600.380 705.420 1604.000 ;
        RECT 705.140 1600.000 705.480 1600.380 ;
        RECT 705.340 1587.450 705.480 1600.000 ;
        RECT 705.280 1587.130 705.540 1587.450 ;
        RECT 710.340 1587.130 710.600 1587.450 ;
        RECT 710.400 22.090 710.540 1587.130 ;
        RECT 710.340 21.770 710.600 22.090 ;
        RECT 1025.440 21.770 1025.700 22.090 ;
        RECT 1025.500 2.400 1025.640 21.770 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 711.690 1587.360 712.010 1587.420 ;
        RECT 717.210 1587.360 717.530 1587.420 ;
        RECT 711.690 1587.220 717.530 1587.360 ;
        RECT 711.690 1587.160 712.010 1587.220 ;
        RECT 717.210 1587.160 717.530 1587.220 ;
        RECT 717.210 22.340 717.530 22.400 ;
        RECT 1043.350 22.340 1043.670 22.400 ;
        RECT 717.210 22.200 1043.670 22.340 ;
        RECT 717.210 22.140 717.530 22.200 ;
        RECT 1043.350 22.140 1043.670 22.200 ;
      LAYER via ;
        RECT 711.720 1587.160 711.980 1587.420 ;
        RECT 717.240 1587.160 717.500 1587.420 ;
        RECT 717.240 22.140 717.500 22.400 ;
        RECT 1043.380 22.140 1043.640 22.400 ;
      LAYER met2 ;
        RECT 711.580 1600.380 711.860 1604.000 ;
        RECT 711.580 1600.000 711.920 1600.380 ;
        RECT 711.780 1587.450 711.920 1600.000 ;
        RECT 711.720 1587.130 711.980 1587.450 ;
        RECT 717.240 1587.130 717.500 1587.450 ;
        RECT 717.300 22.430 717.440 1587.130 ;
        RECT 717.240 22.110 717.500 22.430 ;
        RECT 1043.380 22.110 1043.640 22.430 ;
        RECT 1043.440 2.400 1043.580 22.110 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 717.670 1587.360 717.990 1587.420 ;
        RECT 723.190 1587.360 723.510 1587.420 ;
        RECT 717.670 1587.220 723.510 1587.360 ;
        RECT 717.670 1587.160 717.990 1587.220 ;
        RECT 723.190 1587.160 723.510 1587.220 ;
        RECT 723.190 22.680 723.510 22.740 ;
        RECT 1061.290 22.680 1061.610 22.740 ;
        RECT 723.190 22.540 1061.610 22.680 ;
        RECT 723.190 22.480 723.510 22.540 ;
        RECT 1061.290 22.480 1061.610 22.540 ;
      LAYER via ;
        RECT 717.700 1587.160 717.960 1587.420 ;
        RECT 723.220 1587.160 723.480 1587.420 ;
        RECT 723.220 22.480 723.480 22.740 ;
        RECT 1061.320 22.480 1061.580 22.740 ;
      LAYER met2 ;
        RECT 717.560 1600.380 717.840 1604.000 ;
        RECT 717.560 1600.000 717.900 1600.380 ;
        RECT 717.760 1587.450 717.900 1600.000 ;
        RECT 717.700 1587.130 717.960 1587.450 ;
        RECT 723.220 1587.130 723.480 1587.450 ;
        RECT 723.280 22.770 723.420 1587.130 ;
        RECT 723.220 22.450 723.480 22.770 ;
        RECT 1061.320 22.450 1061.580 22.770 ;
        RECT 1061.380 2.400 1061.520 22.450 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 723.650 23.020 723.970 23.080 ;
        RECT 1079.230 23.020 1079.550 23.080 ;
        RECT 723.650 22.880 1079.550 23.020 ;
        RECT 723.650 22.820 723.970 22.880 ;
        RECT 1079.230 22.820 1079.550 22.880 ;
      LAYER via ;
        RECT 723.680 22.820 723.940 23.080 ;
        RECT 1079.260 22.820 1079.520 23.080 ;
      LAYER met2 ;
        RECT 724.000 1600.380 724.280 1604.000 ;
        RECT 724.000 1600.000 724.340 1600.380 ;
        RECT 724.200 1588.720 724.340 1600.000 ;
        RECT 723.740 1588.580 724.340 1588.720 ;
        RECT 723.740 23.110 723.880 1588.580 ;
        RECT 723.680 22.790 723.940 23.110 ;
        RECT 1079.260 22.790 1079.520 23.110 ;
        RECT 1079.320 2.400 1079.460 22.790 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 731.010 23.360 731.330 23.420 ;
        RECT 1094.870 23.360 1095.190 23.420 ;
        RECT 731.010 23.220 1095.190 23.360 ;
        RECT 731.010 23.160 731.330 23.220 ;
        RECT 1094.870 23.160 1095.190 23.220 ;
      LAYER via ;
        RECT 731.040 23.160 731.300 23.420 ;
        RECT 1094.900 23.160 1095.160 23.420 ;
      LAYER met2 ;
        RECT 729.980 1600.450 730.260 1604.000 ;
        RECT 729.980 1600.310 731.240 1600.450 ;
        RECT 729.980 1600.000 730.260 1600.310 ;
        RECT 731.100 23.450 731.240 1600.310 ;
        RECT 731.040 23.130 731.300 23.450 ;
        RECT 1094.900 23.130 1095.160 23.450 ;
        RECT 1094.960 16.730 1095.100 23.130 ;
        RECT 1094.960 16.590 1096.940 16.730 ;
        RECT 1096.800 2.400 1096.940 16.590 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1076.545 23.545 1077.175 23.715 ;
        RECT 1077.005 22.525 1077.175 23.545 ;
      LAYER met1 ;
        RECT 737.910 23.700 738.230 23.760 ;
        RECT 1076.485 23.700 1076.775 23.745 ;
        RECT 737.910 23.560 1076.775 23.700 ;
        RECT 737.910 23.500 738.230 23.560 ;
        RECT 1076.485 23.515 1076.775 23.560 ;
        RECT 1114.650 23.020 1114.970 23.080 ;
        RECT 1079.780 22.880 1114.970 23.020 ;
        RECT 1076.945 22.680 1077.235 22.725 ;
        RECT 1079.780 22.680 1079.920 22.880 ;
        RECT 1114.650 22.820 1114.970 22.880 ;
        RECT 1076.945 22.540 1079.920 22.680 ;
        RECT 1076.945 22.495 1077.235 22.540 ;
      LAYER via ;
        RECT 737.940 23.500 738.200 23.760 ;
        RECT 1114.680 22.820 1114.940 23.080 ;
      LAYER met2 ;
        RECT 736.420 1600.450 736.700 1604.000 ;
        RECT 736.420 1600.310 737.680 1600.450 ;
        RECT 736.420 1600.000 736.700 1600.310 ;
        RECT 737.540 1580.050 737.680 1600.310 ;
        RECT 737.540 1579.910 738.140 1580.050 ;
        RECT 738.000 23.790 738.140 1579.910 ;
        RECT 737.940 23.470 738.200 23.790 ;
        RECT 1114.680 22.790 1114.940 23.110 ;
        RECT 1114.740 2.400 1114.880 22.790 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 742.510 1587.360 742.830 1587.420 ;
        RECT 744.810 1587.360 745.130 1587.420 ;
        RECT 742.510 1587.220 745.130 1587.360 ;
        RECT 742.510 1587.160 742.830 1587.220 ;
        RECT 744.810 1587.160 745.130 1587.220 ;
        RECT 744.810 27.440 745.130 27.500 ;
        RECT 1132.590 27.440 1132.910 27.500 ;
        RECT 744.810 27.300 1132.910 27.440 ;
        RECT 744.810 27.240 745.130 27.300 ;
        RECT 1132.590 27.240 1132.910 27.300 ;
      LAYER via ;
        RECT 742.540 1587.160 742.800 1587.420 ;
        RECT 744.840 1587.160 745.100 1587.420 ;
        RECT 744.840 27.240 745.100 27.500 ;
        RECT 1132.620 27.240 1132.880 27.500 ;
      LAYER met2 ;
        RECT 742.400 1600.380 742.680 1604.000 ;
        RECT 742.400 1600.000 742.740 1600.380 ;
        RECT 742.600 1587.450 742.740 1600.000 ;
        RECT 742.540 1587.130 742.800 1587.450 ;
        RECT 744.840 1587.130 745.100 1587.450 ;
        RECT 744.900 27.530 745.040 1587.130 ;
        RECT 744.840 27.210 745.100 27.530 ;
        RECT 1132.620 27.210 1132.880 27.530 ;
        RECT 1132.680 2.400 1132.820 27.210 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 748.950 1592.120 749.270 1592.180 ;
        RECT 751.250 1592.120 751.570 1592.180 ;
        RECT 748.950 1591.980 751.570 1592.120 ;
        RECT 748.950 1591.920 749.270 1591.980 ;
        RECT 751.250 1591.920 751.570 1591.980 ;
        RECT 751.250 26.760 751.570 26.820 ;
        RECT 1150.530 26.760 1150.850 26.820 ;
        RECT 751.250 26.620 1150.850 26.760 ;
        RECT 751.250 26.560 751.570 26.620 ;
        RECT 1150.530 26.560 1150.850 26.620 ;
      LAYER via ;
        RECT 748.980 1591.920 749.240 1592.180 ;
        RECT 751.280 1591.920 751.540 1592.180 ;
        RECT 751.280 26.560 751.540 26.820 ;
        RECT 1150.560 26.560 1150.820 26.820 ;
      LAYER met2 ;
        RECT 748.380 1600.450 748.660 1604.000 ;
        RECT 748.380 1600.310 749.180 1600.450 ;
        RECT 748.380 1600.000 748.660 1600.310 ;
        RECT 749.040 1592.210 749.180 1600.310 ;
        RECT 748.980 1591.890 749.240 1592.210 ;
        RECT 751.280 1591.890 751.540 1592.210 ;
        RECT 751.340 26.850 751.480 1591.890 ;
        RECT 751.280 26.530 751.540 26.850 ;
        RECT 1150.560 26.530 1150.820 26.850 ;
        RECT 1150.620 2.400 1150.760 26.530 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 581.510 1590.420 581.830 1590.480 ;
        RECT 586.110 1590.420 586.430 1590.480 ;
        RECT 581.510 1590.280 586.430 1590.420 ;
        RECT 581.510 1590.220 581.830 1590.280 ;
        RECT 586.110 1590.220 586.430 1590.280 ;
        RECT 584.730 25.400 585.050 25.460 ;
        RECT 586.110 25.400 586.430 25.460 ;
        RECT 584.730 25.260 586.430 25.400 ;
        RECT 584.730 25.200 585.050 25.260 ;
        RECT 586.110 25.200 586.430 25.260 ;
        RECT 584.730 14.180 585.050 14.240 ;
        RECT 668.910 14.180 669.230 14.240 ;
        RECT 584.730 14.040 669.230 14.180 ;
        RECT 584.730 13.980 585.050 14.040 ;
        RECT 668.910 13.980 669.230 14.040 ;
      LAYER via ;
        RECT 581.540 1590.220 581.800 1590.480 ;
        RECT 586.140 1590.220 586.400 1590.480 ;
        RECT 584.760 25.200 585.020 25.460 ;
        RECT 586.140 25.200 586.400 25.460 ;
        RECT 584.760 13.980 585.020 14.240 ;
        RECT 668.940 13.980 669.200 14.240 ;
      LAYER met2 ;
        RECT 581.400 1600.380 581.680 1604.000 ;
        RECT 581.400 1600.000 581.740 1600.380 ;
        RECT 581.600 1590.510 581.740 1600.000 ;
        RECT 581.540 1590.190 581.800 1590.510 ;
        RECT 586.140 1590.190 586.400 1590.510 ;
        RECT 586.200 25.490 586.340 1590.190 ;
        RECT 584.760 25.170 585.020 25.490 ;
        RECT 586.140 25.170 586.400 25.490 ;
        RECT 584.820 14.270 584.960 25.170 ;
        RECT 584.760 13.950 585.020 14.270 ;
        RECT 668.940 13.950 669.200 14.270 ;
        RECT 669.000 2.400 669.140 13.950 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 758.150 26.080 758.470 26.140 ;
        RECT 1168.470 26.080 1168.790 26.140 ;
        RECT 758.150 25.940 1168.790 26.080 ;
        RECT 758.150 25.880 758.470 25.940 ;
        RECT 1168.470 25.880 1168.790 25.940 ;
      LAYER via ;
        RECT 758.180 25.880 758.440 26.140 ;
        RECT 1168.500 25.880 1168.760 26.140 ;
      LAYER met2 ;
        RECT 754.820 1600.450 755.100 1604.000 ;
        RECT 754.820 1600.310 756.080 1600.450 ;
        RECT 754.820 1600.000 755.100 1600.310 ;
        RECT 755.940 1564.410 756.080 1600.310 ;
        RECT 755.940 1564.270 758.380 1564.410 ;
        RECT 758.240 26.170 758.380 1564.270 ;
        RECT 758.180 25.850 758.440 26.170 ;
        RECT 1168.500 25.850 1168.760 26.170 ;
        RECT 1168.560 2.400 1168.700 25.850 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 760.910 1587.700 761.230 1587.760 ;
        RECT 765.510 1587.700 765.830 1587.760 ;
        RECT 760.910 1587.560 765.830 1587.700 ;
        RECT 760.910 1587.500 761.230 1587.560 ;
        RECT 765.510 1587.500 765.830 1587.560 ;
        RECT 765.510 25.400 765.830 25.460 ;
        RECT 1185.950 25.400 1186.270 25.460 ;
        RECT 765.510 25.260 1186.270 25.400 ;
        RECT 765.510 25.200 765.830 25.260 ;
        RECT 1185.950 25.200 1186.270 25.260 ;
      LAYER via ;
        RECT 760.940 1587.500 761.200 1587.760 ;
        RECT 765.540 1587.500 765.800 1587.760 ;
        RECT 765.540 25.200 765.800 25.460 ;
        RECT 1185.980 25.200 1186.240 25.460 ;
      LAYER met2 ;
        RECT 760.800 1600.380 761.080 1604.000 ;
        RECT 760.800 1600.000 761.140 1600.380 ;
        RECT 761.000 1587.790 761.140 1600.000 ;
        RECT 760.940 1587.470 761.200 1587.790 ;
        RECT 765.540 1587.470 765.800 1587.790 ;
        RECT 765.600 25.490 765.740 1587.470 ;
        RECT 765.540 25.170 765.800 25.490 ;
        RECT 1185.980 25.170 1186.240 25.490 ;
        RECT 1186.040 2.400 1186.180 25.170 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 767.350 1587.360 767.670 1587.420 ;
        RECT 772.410 1587.360 772.730 1587.420 ;
        RECT 767.350 1587.220 772.730 1587.360 ;
        RECT 767.350 1587.160 767.670 1587.220 ;
        RECT 772.410 1587.160 772.730 1587.220 ;
        RECT 772.410 25.060 772.730 25.120 ;
        RECT 1203.890 25.060 1204.210 25.120 ;
        RECT 772.410 24.920 1204.210 25.060 ;
        RECT 772.410 24.860 772.730 24.920 ;
        RECT 1203.890 24.860 1204.210 24.920 ;
      LAYER via ;
        RECT 767.380 1587.160 767.640 1587.420 ;
        RECT 772.440 1587.160 772.700 1587.420 ;
        RECT 772.440 24.860 772.700 25.120 ;
        RECT 1203.920 24.860 1204.180 25.120 ;
      LAYER met2 ;
        RECT 767.240 1600.380 767.520 1604.000 ;
        RECT 767.240 1600.000 767.580 1600.380 ;
        RECT 767.440 1587.450 767.580 1600.000 ;
        RECT 767.380 1587.130 767.640 1587.450 ;
        RECT 772.440 1587.130 772.700 1587.450 ;
        RECT 772.500 25.150 772.640 1587.130 ;
        RECT 772.440 24.830 772.700 25.150 ;
        RECT 1203.920 24.830 1204.180 25.150 ;
        RECT 1203.980 2.400 1204.120 24.830 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 773.330 1587.700 773.650 1587.760 ;
        RECT 779.310 1587.700 779.630 1587.760 ;
        RECT 773.330 1587.560 779.630 1587.700 ;
        RECT 773.330 1587.500 773.650 1587.560 ;
        RECT 779.310 1587.500 779.630 1587.560 ;
        RECT 779.310 24.720 779.630 24.780 ;
        RECT 1221.830 24.720 1222.150 24.780 ;
        RECT 779.310 24.580 1222.150 24.720 ;
        RECT 779.310 24.520 779.630 24.580 ;
        RECT 1221.830 24.520 1222.150 24.580 ;
      LAYER via ;
        RECT 773.360 1587.500 773.620 1587.760 ;
        RECT 779.340 1587.500 779.600 1587.760 ;
        RECT 779.340 24.520 779.600 24.780 ;
        RECT 1221.860 24.520 1222.120 24.780 ;
      LAYER met2 ;
        RECT 773.220 1600.380 773.500 1604.000 ;
        RECT 773.220 1600.000 773.560 1600.380 ;
        RECT 773.420 1587.790 773.560 1600.000 ;
        RECT 773.360 1587.470 773.620 1587.790 ;
        RECT 779.340 1587.470 779.600 1587.790 ;
        RECT 779.400 24.810 779.540 1587.470 ;
        RECT 779.340 24.490 779.600 24.810 ;
        RECT 1221.860 24.490 1222.120 24.810 ;
        RECT 1221.920 2.400 1222.060 24.490 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.770 1587.700 780.090 1587.760 ;
        RECT 786.210 1587.700 786.530 1587.760 ;
        RECT 779.770 1587.560 786.530 1587.700 ;
        RECT 779.770 1587.500 780.090 1587.560 ;
        RECT 786.210 1587.500 786.530 1587.560 ;
        RECT 786.210 24.380 786.530 24.440 ;
        RECT 1239.770 24.380 1240.090 24.440 ;
        RECT 786.210 24.240 1240.090 24.380 ;
        RECT 786.210 24.180 786.530 24.240 ;
        RECT 1239.770 24.180 1240.090 24.240 ;
      LAYER via ;
        RECT 779.800 1587.500 780.060 1587.760 ;
        RECT 786.240 1587.500 786.500 1587.760 ;
        RECT 786.240 24.180 786.500 24.440 ;
        RECT 1239.800 24.180 1240.060 24.440 ;
      LAYER met2 ;
        RECT 779.660 1600.380 779.940 1604.000 ;
        RECT 779.660 1600.000 780.000 1600.380 ;
        RECT 779.860 1587.790 780.000 1600.000 ;
        RECT 779.800 1587.470 780.060 1587.790 ;
        RECT 786.240 1587.470 786.500 1587.790 ;
        RECT 786.300 24.470 786.440 1587.470 ;
        RECT 786.240 24.150 786.500 24.470 ;
        RECT 1239.800 24.150 1240.060 24.470 ;
        RECT 1239.860 2.400 1240.000 24.150 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 786.745 23.885 786.915 27.795 ;
        RECT 858.965 20.825 859.135 24.055 ;
        RECT 907.265 20.825 907.435 24.055 ;
        RECT 979.485 19.805 979.655 24.055 ;
        RECT 979.945 19.805 980.115 24.055 ;
        RECT 1147.845 22.185 1148.015 24.055 ;
        RECT 1172.225 22.525 1173.315 22.695 ;
        RECT 1195.685 22.525 1195.855 23.715 ;
        RECT 1239.385 23.545 1239.555 25.755 ;
        RECT 1172.225 22.185 1172.395 22.525 ;
      LAYER mcon ;
        RECT 786.745 27.625 786.915 27.795 ;
        RECT 1239.385 25.585 1239.555 25.755 ;
        RECT 858.965 23.885 859.135 24.055 ;
        RECT 907.265 23.885 907.435 24.055 ;
        RECT 979.485 23.885 979.655 24.055 ;
        RECT 979.945 23.885 980.115 24.055 ;
        RECT 1147.845 23.885 1148.015 24.055 ;
        RECT 1195.685 23.545 1195.855 23.715 ;
        RECT 1173.145 22.525 1173.315 22.695 ;
      LAYER met1 ;
        RECT 785.750 27.780 786.070 27.840 ;
        RECT 786.685 27.780 786.975 27.825 ;
        RECT 785.750 27.640 786.975 27.780 ;
        RECT 785.750 27.580 786.070 27.640 ;
        RECT 786.685 27.595 786.975 27.640 ;
        RECT 1239.325 25.740 1239.615 25.785 ;
        RECT 1257.250 25.740 1257.570 25.800 ;
        RECT 1239.325 25.600 1257.570 25.740 ;
        RECT 1239.325 25.555 1239.615 25.600 ;
        RECT 1257.250 25.540 1257.570 25.600 ;
        RECT 786.685 24.040 786.975 24.085 ;
        RECT 858.905 24.040 859.195 24.085 ;
        RECT 786.685 23.900 859.195 24.040 ;
        RECT 786.685 23.855 786.975 23.900 ;
        RECT 858.905 23.855 859.195 23.900 ;
        RECT 907.205 24.040 907.495 24.085 ;
        RECT 979.425 24.040 979.715 24.085 ;
        RECT 907.205 23.900 979.715 24.040 ;
        RECT 907.205 23.855 907.495 23.900 ;
        RECT 979.425 23.855 979.715 23.900 ;
        RECT 979.885 24.040 980.175 24.085 ;
        RECT 1075.550 24.040 1075.870 24.100 ;
        RECT 979.885 23.900 1075.870 24.040 ;
        RECT 979.885 23.855 980.175 23.900 ;
        RECT 1075.550 23.840 1075.870 23.900 ;
        RECT 1077.850 24.040 1078.170 24.100 ;
        RECT 1147.785 24.040 1148.075 24.085 ;
        RECT 1077.850 23.900 1148.075 24.040 ;
        RECT 1077.850 23.840 1078.170 23.900 ;
        RECT 1147.785 23.855 1148.075 23.900 ;
        RECT 1195.625 23.700 1195.915 23.745 ;
        RECT 1239.325 23.700 1239.615 23.745 ;
        RECT 1195.625 23.560 1239.615 23.700 ;
        RECT 1195.625 23.515 1195.915 23.560 ;
        RECT 1239.325 23.515 1239.615 23.560 ;
        RECT 1173.085 22.680 1173.375 22.725 ;
        RECT 1195.625 22.680 1195.915 22.725 ;
        RECT 1173.085 22.540 1195.915 22.680 ;
        RECT 1173.085 22.495 1173.375 22.540 ;
        RECT 1195.625 22.495 1195.915 22.540 ;
        RECT 1147.785 22.340 1148.075 22.385 ;
        RECT 1172.165 22.340 1172.455 22.385 ;
        RECT 1147.785 22.200 1172.455 22.340 ;
        RECT 1147.785 22.155 1148.075 22.200 ;
        RECT 1172.165 22.155 1172.455 22.200 ;
        RECT 858.905 20.980 859.195 21.025 ;
        RECT 907.205 20.980 907.495 21.025 ;
        RECT 858.905 20.840 907.495 20.980 ;
        RECT 858.905 20.795 859.195 20.840 ;
        RECT 907.205 20.795 907.495 20.840 ;
        RECT 979.425 19.960 979.715 20.005 ;
        RECT 979.885 19.960 980.175 20.005 ;
        RECT 979.425 19.820 980.175 19.960 ;
        RECT 979.425 19.775 979.715 19.820 ;
        RECT 979.885 19.775 980.175 19.820 ;
      LAYER via ;
        RECT 785.780 27.580 786.040 27.840 ;
        RECT 1257.280 25.540 1257.540 25.800 ;
        RECT 1075.580 23.840 1075.840 24.100 ;
        RECT 1077.880 23.840 1078.140 24.100 ;
      LAYER met2 ;
        RECT 785.640 1600.380 785.920 1604.000 ;
        RECT 785.640 1600.000 785.980 1600.380 ;
        RECT 785.840 27.870 785.980 1600.000 ;
        RECT 785.780 27.550 786.040 27.870 ;
        RECT 1257.280 25.510 1257.540 25.830 ;
        RECT 1075.580 23.810 1075.840 24.130 ;
        RECT 1077.880 23.810 1078.140 24.130 ;
        RECT 1075.640 23.645 1075.780 23.810 ;
        RECT 1077.940 23.645 1078.080 23.810 ;
        RECT 1075.570 23.275 1075.850 23.645 ;
        RECT 1077.870 23.275 1078.150 23.645 ;
        RECT 1257.340 2.400 1257.480 25.510 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
      LAYER via2 ;
        RECT 1075.570 23.320 1075.850 23.600 ;
        RECT 1077.870 23.320 1078.150 23.600 ;
      LAYER met3 ;
        RECT 1075.545 23.610 1075.875 23.625 ;
        RECT 1077.845 23.610 1078.175 23.625 ;
        RECT 1075.545 23.310 1078.175 23.610 ;
        RECT 1075.545 23.295 1075.875 23.310 ;
        RECT 1077.845 23.295 1078.175 23.310 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 792.080 1600.450 792.360 1604.000 ;
        RECT 792.080 1600.310 793.340 1600.450 ;
        RECT 792.080 1600.000 792.360 1600.310 ;
        RECT 793.200 27.045 793.340 1600.310 ;
        RECT 793.130 26.675 793.410 27.045 ;
        RECT 1275.210 26.675 1275.490 27.045 ;
        RECT 1275.280 2.400 1275.420 26.675 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
      LAYER via2 ;
        RECT 793.130 26.720 793.410 27.000 ;
        RECT 1275.210 26.720 1275.490 27.000 ;
      LAYER met3 ;
        RECT 793.105 27.010 793.435 27.025 ;
        RECT 1275.185 27.010 1275.515 27.025 ;
        RECT 793.105 26.710 1275.515 27.010 ;
        RECT 793.105 26.695 793.435 26.710 ;
        RECT 1275.185 26.695 1275.515 26.710 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 798.170 1587.360 798.490 1587.420 ;
        RECT 800.010 1587.360 800.330 1587.420 ;
        RECT 798.170 1587.220 800.330 1587.360 ;
        RECT 798.170 1587.160 798.490 1587.220 ;
        RECT 800.010 1587.160 800.330 1587.220 ;
      LAYER via ;
        RECT 798.200 1587.160 798.460 1587.420 ;
        RECT 800.040 1587.160 800.300 1587.420 ;
      LAYER met2 ;
        RECT 798.060 1600.380 798.340 1604.000 ;
        RECT 798.060 1600.000 798.400 1600.380 ;
        RECT 798.260 1587.450 798.400 1600.000 ;
        RECT 798.200 1587.130 798.460 1587.450 ;
        RECT 800.040 1587.130 800.300 1587.450 ;
        RECT 800.100 26.365 800.240 1587.130 ;
        RECT 800.030 25.995 800.310 26.365 ;
        RECT 1293.150 25.995 1293.430 26.365 ;
        RECT 1293.220 2.400 1293.360 25.995 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
      LAYER via2 ;
        RECT 800.030 26.040 800.310 26.320 ;
        RECT 1293.150 26.040 1293.430 26.320 ;
      LAYER met3 ;
        RECT 800.005 26.330 800.335 26.345 ;
        RECT 1293.125 26.330 1293.455 26.345 ;
        RECT 800.005 26.030 1293.455 26.330 ;
        RECT 800.005 26.015 800.335 26.030 ;
        RECT 1293.125 26.015 1293.455 26.030 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 804.150 1587.360 804.470 1587.420 ;
        RECT 806.910 1587.360 807.230 1587.420 ;
        RECT 804.150 1587.220 807.230 1587.360 ;
        RECT 804.150 1587.160 804.470 1587.220 ;
        RECT 806.910 1587.160 807.230 1587.220 ;
      LAYER via ;
        RECT 804.180 1587.160 804.440 1587.420 ;
        RECT 806.940 1587.160 807.200 1587.420 ;
      LAYER met2 ;
        RECT 804.040 1600.380 804.320 1604.000 ;
        RECT 804.040 1600.000 804.380 1600.380 ;
        RECT 804.240 1587.450 804.380 1600.000 ;
        RECT 804.180 1587.130 804.440 1587.450 ;
        RECT 806.940 1587.130 807.200 1587.450 ;
        RECT 807.000 25.685 807.140 1587.130 ;
        RECT 806.930 25.315 807.210 25.685 ;
        RECT 1311.090 25.315 1311.370 25.685 ;
        RECT 1311.160 2.400 1311.300 25.315 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
      LAYER via2 ;
        RECT 806.930 25.360 807.210 25.640 ;
        RECT 1311.090 25.360 1311.370 25.640 ;
      LAYER met3 ;
        RECT 806.905 25.650 807.235 25.665 ;
        RECT 1311.065 25.650 1311.395 25.665 ;
        RECT 806.905 25.350 1311.395 25.650 ;
        RECT 806.905 25.335 807.235 25.350 ;
        RECT 1311.065 25.335 1311.395 25.350 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 810.590 1587.360 810.910 1587.420 ;
        RECT 813.810 1587.360 814.130 1587.420 ;
        RECT 810.590 1587.220 814.130 1587.360 ;
        RECT 810.590 1587.160 810.910 1587.220 ;
        RECT 813.810 1587.160 814.130 1587.220 ;
      LAYER via ;
        RECT 810.620 1587.160 810.880 1587.420 ;
        RECT 813.840 1587.160 814.100 1587.420 ;
      LAYER met2 ;
        RECT 810.480 1600.380 810.760 1604.000 ;
        RECT 810.480 1600.000 810.820 1600.380 ;
        RECT 810.680 1587.450 810.820 1600.000 ;
        RECT 810.620 1587.130 810.880 1587.450 ;
        RECT 813.840 1587.130 814.100 1587.450 ;
        RECT 813.900 25.005 814.040 1587.130 ;
        RECT 813.830 24.635 814.110 25.005 ;
        RECT 1329.030 24.635 1329.310 25.005 ;
        RECT 1329.100 2.400 1329.240 24.635 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
      LAYER via2 ;
        RECT 813.830 24.680 814.110 24.960 ;
        RECT 1329.030 24.680 1329.310 24.960 ;
      LAYER met3 ;
        RECT 813.805 24.970 814.135 24.985 ;
        RECT 1329.005 24.970 1329.335 24.985 ;
        RECT 813.805 24.670 1329.335 24.970 ;
        RECT 813.805 24.655 814.135 24.670 ;
        RECT 1329.005 24.655 1329.335 24.670 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 638.165 16.405 638.335 17.595 ;
        RECT 664.845 13.685 665.015 17.595 ;
      LAYER mcon ;
        RECT 638.165 17.425 638.335 17.595 ;
        RECT 664.845 17.425 665.015 17.595 ;
      LAYER met1 ;
        RECT 587.950 1588.040 588.270 1588.100 ;
        RECT 592.550 1588.040 592.870 1588.100 ;
        RECT 587.950 1587.900 592.870 1588.040 ;
        RECT 587.950 1587.840 588.270 1587.900 ;
        RECT 592.550 1587.840 592.870 1587.900 ;
        RECT 638.105 17.580 638.395 17.625 ;
        RECT 664.785 17.580 665.075 17.625 ;
        RECT 638.105 17.440 665.075 17.580 ;
        RECT 638.105 17.395 638.395 17.440 ;
        RECT 664.785 17.395 665.075 17.440 ;
        RECT 592.550 16.900 592.870 16.960 ;
        RECT 592.550 16.760 609.800 16.900 ;
        RECT 592.550 16.700 592.870 16.760 ;
        RECT 609.660 16.560 609.800 16.760 ;
        RECT 638.105 16.560 638.395 16.605 ;
        RECT 609.660 16.420 638.395 16.560 ;
        RECT 638.105 16.375 638.395 16.420 ;
        RECT 686.390 14.180 686.710 14.240 ;
        RECT 669.460 14.040 686.710 14.180 ;
        RECT 664.785 13.840 665.075 13.885 ;
        RECT 669.460 13.840 669.600 14.040 ;
        RECT 686.390 13.980 686.710 14.040 ;
        RECT 664.785 13.700 669.600 13.840 ;
        RECT 664.785 13.655 665.075 13.700 ;
      LAYER via ;
        RECT 587.980 1587.840 588.240 1588.100 ;
        RECT 592.580 1587.840 592.840 1588.100 ;
        RECT 592.580 16.700 592.840 16.960 ;
        RECT 686.420 13.980 686.680 14.240 ;
      LAYER met2 ;
        RECT 587.840 1600.380 588.120 1604.000 ;
        RECT 587.840 1600.000 588.180 1600.380 ;
        RECT 588.040 1588.130 588.180 1600.000 ;
        RECT 587.980 1587.810 588.240 1588.130 ;
        RECT 592.580 1587.810 592.840 1588.130 ;
        RECT 592.640 16.990 592.780 1587.810 ;
        RECT 592.580 16.670 592.840 16.990 ;
        RECT 686.420 13.950 686.680 14.270 ;
        RECT 686.480 2.400 686.620 13.950 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 816.570 1587.360 816.890 1587.420 ;
        RECT 820.710 1587.360 821.030 1587.420 ;
        RECT 816.570 1587.220 821.030 1587.360 ;
        RECT 816.570 1587.160 816.890 1587.220 ;
        RECT 820.710 1587.160 821.030 1587.220 ;
      LAYER via ;
        RECT 816.600 1587.160 816.860 1587.420 ;
        RECT 820.740 1587.160 821.000 1587.420 ;
      LAYER met2 ;
        RECT 816.460 1600.380 816.740 1604.000 ;
        RECT 816.460 1600.000 816.800 1600.380 ;
        RECT 816.660 1587.450 816.800 1600.000 ;
        RECT 816.600 1587.130 816.860 1587.450 ;
        RECT 820.740 1587.130 821.000 1587.450 ;
        RECT 820.800 24.325 820.940 1587.130 ;
        RECT 820.730 23.955 821.010 24.325 ;
        RECT 1346.510 23.955 1346.790 24.325 ;
        RECT 1346.580 2.400 1346.720 23.955 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
      LAYER via2 ;
        RECT 820.730 24.000 821.010 24.280 ;
        RECT 1346.510 24.000 1346.790 24.280 ;
      LAYER met3 ;
        RECT 820.705 24.290 821.035 24.305 ;
        RECT 1346.485 24.290 1346.815 24.305 ;
        RECT 820.705 23.990 1346.815 24.290 ;
        RECT 820.705 23.975 821.035 23.990 ;
        RECT 1346.485 23.975 1346.815 23.990 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 823.010 1587.360 823.330 1587.420 ;
        RECT 826.690 1587.360 827.010 1587.420 ;
        RECT 823.010 1587.220 827.010 1587.360 ;
        RECT 823.010 1587.160 823.330 1587.220 ;
        RECT 826.690 1587.160 827.010 1587.220 ;
        RECT 826.690 62.460 827.010 62.520 ;
        RECT 1359.370 62.460 1359.690 62.520 ;
        RECT 826.690 62.320 1359.690 62.460 ;
        RECT 826.690 62.260 827.010 62.320 ;
        RECT 1359.370 62.260 1359.690 62.320 ;
        RECT 1359.370 2.960 1359.690 3.020 ;
        RECT 1364.430 2.960 1364.750 3.020 ;
        RECT 1359.370 2.820 1364.750 2.960 ;
        RECT 1359.370 2.760 1359.690 2.820 ;
        RECT 1364.430 2.760 1364.750 2.820 ;
      LAYER via ;
        RECT 823.040 1587.160 823.300 1587.420 ;
        RECT 826.720 1587.160 826.980 1587.420 ;
        RECT 826.720 62.260 826.980 62.520 ;
        RECT 1359.400 62.260 1359.660 62.520 ;
        RECT 1359.400 2.760 1359.660 3.020 ;
        RECT 1364.460 2.760 1364.720 3.020 ;
      LAYER met2 ;
        RECT 822.900 1600.380 823.180 1604.000 ;
        RECT 822.900 1600.000 823.240 1600.380 ;
        RECT 823.100 1587.450 823.240 1600.000 ;
        RECT 823.040 1587.130 823.300 1587.450 ;
        RECT 826.720 1587.130 826.980 1587.450 ;
        RECT 826.780 62.550 826.920 1587.130 ;
        RECT 826.720 62.230 826.980 62.550 ;
        RECT 1359.400 62.230 1359.660 62.550 ;
        RECT 1359.460 3.050 1359.600 62.230 ;
        RECT 1359.400 2.730 1359.660 3.050 ;
        RECT 1364.460 2.730 1364.720 3.050 ;
        RECT 1364.520 2.400 1364.660 2.730 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 828.990 1587.700 829.310 1587.760 ;
        RECT 834.510 1587.700 834.830 1587.760 ;
        RECT 828.990 1587.560 834.830 1587.700 ;
        RECT 828.990 1587.500 829.310 1587.560 ;
        RECT 834.510 1587.500 834.830 1587.560 ;
      LAYER via ;
        RECT 829.020 1587.500 829.280 1587.760 ;
        RECT 834.540 1587.500 834.800 1587.760 ;
      LAYER met2 ;
        RECT 828.880 1600.380 829.160 1604.000 ;
        RECT 828.880 1600.000 829.220 1600.380 ;
        RECT 829.080 1587.790 829.220 1600.000 ;
        RECT 829.020 1587.470 829.280 1587.790 ;
        RECT 834.540 1587.470 834.800 1587.790 ;
        RECT 834.600 27.725 834.740 1587.470 ;
        RECT 834.530 27.355 834.810 27.725 ;
        RECT 1382.390 27.355 1382.670 27.725 ;
        RECT 1382.460 2.400 1382.600 27.355 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
      LAYER via2 ;
        RECT 834.530 27.400 834.810 27.680 ;
        RECT 1382.390 27.400 1382.670 27.680 ;
      LAYER met3 ;
        RECT 834.505 27.690 834.835 27.705 ;
        RECT 1382.365 27.690 1382.695 27.705 ;
        RECT 834.505 27.390 1382.695 27.690 ;
        RECT 834.505 27.375 834.835 27.390 ;
        RECT 1382.365 27.375 1382.695 27.390 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 835.430 1587.360 835.750 1587.420 ;
        RECT 840.490 1587.360 840.810 1587.420 ;
        RECT 835.430 1587.220 840.810 1587.360 ;
        RECT 835.430 1587.160 835.750 1587.220 ;
        RECT 840.490 1587.160 840.810 1587.220 ;
        RECT 840.490 69.600 840.810 69.660 ;
        RECT 1393.870 69.600 1394.190 69.660 ;
        RECT 840.490 69.460 1394.190 69.600 ;
        RECT 840.490 69.400 840.810 69.460 ;
        RECT 1393.870 69.400 1394.190 69.460 ;
        RECT 1393.870 16.900 1394.190 16.960 ;
        RECT 1400.310 16.900 1400.630 16.960 ;
        RECT 1393.870 16.760 1400.630 16.900 ;
        RECT 1393.870 16.700 1394.190 16.760 ;
        RECT 1400.310 16.700 1400.630 16.760 ;
      LAYER via ;
        RECT 835.460 1587.160 835.720 1587.420 ;
        RECT 840.520 1587.160 840.780 1587.420 ;
        RECT 840.520 69.400 840.780 69.660 ;
        RECT 1393.900 69.400 1394.160 69.660 ;
        RECT 1393.900 16.700 1394.160 16.960 ;
        RECT 1400.340 16.700 1400.600 16.960 ;
      LAYER met2 ;
        RECT 835.320 1600.380 835.600 1604.000 ;
        RECT 835.320 1600.000 835.660 1600.380 ;
        RECT 835.520 1587.450 835.660 1600.000 ;
        RECT 835.460 1587.130 835.720 1587.450 ;
        RECT 840.520 1587.130 840.780 1587.450 ;
        RECT 840.580 69.690 840.720 1587.130 ;
        RECT 840.520 69.370 840.780 69.690 ;
        RECT 1393.900 69.370 1394.160 69.690 ;
        RECT 1393.960 16.990 1394.100 69.370 ;
        RECT 1393.900 16.670 1394.160 16.990 ;
        RECT 1400.340 16.670 1400.600 16.990 ;
        RECT 1400.400 2.400 1400.540 16.670 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.950 70.960 841.270 71.020 ;
        RECT 1414.570 70.960 1414.890 71.020 ;
        RECT 840.950 70.820 1414.890 70.960 ;
        RECT 840.950 70.760 841.270 70.820 ;
        RECT 1414.570 70.760 1414.890 70.820 ;
        RECT 1414.570 2.960 1414.890 3.020 ;
        RECT 1418.250 2.960 1418.570 3.020 ;
        RECT 1414.570 2.820 1418.570 2.960 ;
        RECT 1414.570 2.760 1414.890 2.820 ;
        RECT 1418.250 2.760 1418.570 2.820 ;
      LAYER via ;
        RECT 840.980 70.760 841.240 71.020 ;
        RECT 1414.600 70.760 1414.860 71.020 ;
        RECT 1414.600 2.760 1414.860 3.020 ;
        RECT 1418.280 2.760 1418.540 3.020 ;
      LAYER met2 ;
        RECT 841.300 1600.380 841.580 1604.000 ;
        RECT 841.300 1600.000 841.640 1600.380 ;
        RECT 841.500 1588.210 841.640 1600.000 ;
        RECT 841.040 1588.070 841.640 1588.210 ;
        RECT 841.040 71.050 841.180 1588.070 ;
        RECT 840.980 70.730 841.240 71.050 ;
        RECT 1414.600 70.730 1414.860 71.050 ;
        RECT 1414.660 3.050 1414.800 70.730 ;
        RECT 1414.600 2.730 1414.860 3.050 ;
        RECT 1418.280 2.730 1418.540 3.050 ;
        RECT 1418.340 2.400 1418.480 2.730 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 848.310 27.780 848.630 27.840 ;
        RECT 1434.810 27.780 1435.130 27.840 ;
        RECT 848.310 27.640 1435.130 27.780 ;
        RECT 848.310 27.580 848.630 27.640 ;
        RECT 1434.810 27.580 1435.130 27.640 ;
      LAYER via ;
        RECT 848.340 27.580 848.600 27.840 ;
        RECT 1434.840 27.580 1435.100 27.840 ;
      LAYER met2 ;
        RECT 847.740 1600.450 848.020 1604.000 ;
        RECT 847.740 1600.310 848.540 1600.450 ;
        RECT 847.740 1600.000 848.020 1600.310 ;
        RECT 848.400 27.870 848.540 1600.310 ;
        RECT 848.340 27.550 848.600 27.870 ;
        RECT 1434.840 27.550 1435.100 27.870 ;
        RECT 1434.900 26.930 1435.040 27.550 ;
        RECT 1434.900 26.790 1435.960 26.930 ;
        RECT 1435.820 2.400 1435.960 26.790 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 855.210 28.120 855.530 28.180 ;
        RECT 1453.670 28.120 1453.990 28.180 ;
        RECT 855.210 27.980 1453.990 28.120 ;
        RECT 855.210 27.920 855.530 27.980 ;
        RECT 1453.670 27.920 1453.990 27.980 ;
      LAYER via ;
        RECT 855.240 27.920 855.500 28.180 ;
        RECT 1453.700 27.920 1453.960 28.180 ;
      LAYER met2 ;
        RECT 853.720 1600.450 854.000 1604.000 ;
        RECT 853.720 1600.310 855.440 1600.450 ;
        RECT 853.720 1600.000 854.000 1600.310 ;
        RECT 855.300 28.210 855.440 1600.310 ;
        RECT 855.240 27.890 855.500 28.210 ;
        RECT 1453.700 27.890 1453.960 28.210 ;
        RECT 1453.760 2.400 1453.900 27.890 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 859.810 1587.700 860.130 1587.760 ;
        RECT 862.110 1587.700 862.430 1587.760 ;
        RECT 859.810 1587.560 862.430 1587.700 ;
        RECT 859.810 1587.500 860.130 1587.560 ;
        RECT 862.110 1587.500 862.430 1587.560 ;
        RECT 862.110 28.460 862.430 28.520 ;
        RECT 1471.610 28.460 1471.930 28.520 ;
        RECT 862.110 28.320 1471.930 28.460 ;
        RECT 862.110 28.260 862.430 28.320 ;
        RECT 1471.610 28.260 1471.930 28.320 ;
      LAYER via ;
        RECT 859.840 1587.500 860.100 1587.760 ;
        RECT 862.140 1587.500 862.400 1587.760 ;
        RECT 862.140 28.260 862.400 28.520 ;
        RECT 1471.640 28.260 1471.900 28.520 ;
      LAYER met2 ;
        RECT 859.700 1600.380 859.980 1604.000 ;
        RECT 859.700 1600.000 860.040 1600.380 ;
        RECT 859.900 1587.790 860.040 1600.000 ;
        RECT 859.840 1587.470 860.100 1587.790 ;
        RECT 862.140 1587.470 862.400 1587.790 ;
        RECT 862.200 28.550 862.340 1587.470 ;
        RECT 862.140 28.230 862.400 28.550 ;
        RECT 1471.640 28.230 1471.900 28.550 ;
        RECT 1471.700 2.400 1471.840 28.230 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 866.250 1587.700 866.570 1587.760 ;
        RECT 869.010 1587.700 869.330 1587.760 ;
        RECT 866.250 1587.560 869.330 1587.700 ;
        RECT 866.250 1587.500 866.570 1587.560 ;
        RECT 869.010 1587.500 869.330 1587.560 ;
        RECT 869.010 28.800 869.330 28.860 ;
        RECT 1489.550 28.800 1489.870 28.860 ;
        RECT 869.010 28.660 1489.870 28.800 ;
        RECT 869.010 28.600 869.330 28.660 ;
        RECT 1489.550 28.600 1489.870 28.660 ;
      LAYER via ;
        RECT 866.280 1587.500 866.540 1587.760 ;
        RECT 869.040 1587.500 869.300 1587.760 ;
        RECT 869.040 28.600 869.300 28.860 ;
        RECT 1489.580 28.600 1489.840 28.860 ;
      LAYER met2 ;
        RECT 866.140 1600.380 866.420 1604.000 ;
        RECT 866.140 1600.000 866.480 1600.380 ;
        RECT 866.340 1587.790 866.480 1600.000 ;
        RECT 866.280 1587.470 866.540 1587.790 ;
        RECT 869.040 1587.470 869.300 1587.790 ;
        RECT 869.100 28.890 869.240 1587.470 ;
        RECT 869.040 28.570 869.300 28.890 ;
        RECT 1489.580 28.570 1489.840 28.890 ;
        RECT 1489.640 2.400 1489.780 28.570 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 872.230 1587.360 872.550 1587.420 ;
        RECT 875.450 1587.360 875.770 1587.420 ;
        RECT 872.230 1587.220 875.770 1587.360 ;
        RECT 872.230 1587.160 872.550 1587.220 ;
        RECT 875.450 1587.160 875.770 1587.220 ;
        RECT 875.450 29.140 875.770 29.200 ;
        RECT 1507.030 29.140 1507.350 29.200 ;
        RECT 875.450 29.000 1507.350 29.140 ;
        RECT 875.450 28.940 875.770 29.000 ;
        RECT 1507.030 28.940 1507.350 29.000 ;
      LAYER via ;
        RECT 872.260 1587.160 872.520 1587.420 ;
        RECT 875.480 1587.160 875.740 1587.420 ;
        RECT 875.480 28.940 875.740 29.200 ;
        RECT 1507.060 28.940 1507.320 29.200 ;
      LAYER met2 ;
        RECT 872.120 1600.380 872.400 1604.000 ;
        RECT 872.120 1600.000 872.460 1600.380 ;
        RECT 872.320 1587.450 872.460 1600.000 ;
        RECT 872.260 1587.130 872.520 1587.450 ;
        RECT 875.480 1587.130 875.740 1587.450 ;
        RECT 875.540 29.230 875.680 1587.130 ;
        RECT 875.480 28.910 875.740 29.230 ;
        RECT 1507.060 28.910 1507.320 29.230 ;
        RECT 1507.120 2.400 1507.260 28.910 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 593.930 1590.080 594.250 1590.140 ;
        RECT 599.910 1590.080 600.230 1590.140 ;
        RECT 593.930 1589.940 600.230 1590.080 ;
        RECT 593.930 1589.880 594.250 1589.940 ;
        RECT 599.910 1589.880 600.230 1589.940 ;
        RECT 599.910 14.520 600.230 14.580 ;
        RECT 704.330 14.520 704.650 14.580 ;
        RECT 599.910 14.380 704.650 14.520 ;
        RECT 599.910 14.320 600.230 14.380 ;
        RECT 704.330 14.320 704.650 14.380 ;
      LAYER via ;
        RECT 593.960 1589.880 594.220 1590.140 ;
        RECT 599.940 1589.880 600.200 1590.140 ;
        RECT 599.940 14.320 600.200 14.580 ;
        RECT 704.360 14.320 704.620 14.580 ;
      LAYER met2 ;
        RECT 593.820 1600.380 594.100 1604.000 ;
        RECT 593.820 1600.000 594.160 1600.380 ;
        RECT 594.020 1590.170 594.160 1600.000 ;
        RECT 593.960 1589.850 594.220 1590.170 ;
        RECT 599.940 1589.850 600.200 1590.170 ;
        RECT 600.000 14.610 600.140 1589.850 ;
        RECT 599.940 14.290 600.200 14.610 ;
        RECT 704.360 14.290 704.620 14.610 ;
        RECT 704.420 2.400 704.560 14.290 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 878.670 1587.700 878.990 1587.760 ;
        RECT 882.810 1587.700 883.130 1587.760 ;
        RECT 878.670 1587.560 883.130 1587.700 ;
        RECT 878.670 1587.500 878.990 1587.560 ;
        RECT 882.810 1587.500 883.130 1587.560 ;
        RECT 882.810 29.480 883.130 29.540 ;
        RECT 1525.430 29.480 1525.750 29.540 ;
        RECT 882.810 29.340 1525.750 29.480 ;
        RECT 882.810 29.280 883.130 29.340 ;
        RECT 1525.430 29.280 1525.750 29.340 ;
      LAYER via ;
        RECT 878.700 1587.500 878.960 1587.760 ;
        RECT 882.840 1587.500 883.100 1587.760 ;
        RECT 882.840 29.280 883.100 29.540 ;
        RECT 1525.460 29.280 1525.720 29.540 ;
      LAYER met2 ;
        RECT 878.560 1600.380 878.840 1604.000 ;
        RECT 878.560 1600.000 878.900 1600.380 ;
        RECT 878.760 1587.790 878.900 1600.000 ;
        RECT 878.700 1587.470 878.960 1587.790 ;
        RECT 882.840 1587.470 883.100 1587.790 ;
        RECT 882.900 29.570 883.040 1587.470 ;
        RECT 882.840 29.250 883.100 29.570 ;
        RECT 1525.460 29.250 1525.720 29.570 ;
        RECT 1525.520 16.050 1525.660 29.250 ;
        RECT 1525.060 15.910 1525.660 16.050 ;
        RECT 1525.060 2.400 1525.200 15.910 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 884.650 1587.360 884.970 1587.420 ;
        RECT 889.710 1587.360 890.030 1587.420 ;
        RECT 884.650 1587.220 890.030 1587.360 ;
        RECT 884.650 1587.160 884.970 1587.220 ;
        RECT 889.710 1587.160 890.030 1587.220 ;
        RECT 889.710 29.820 890.030 29.880 ;
        RECT 1542.910 29.820 1543.230 29.880 ;
        RECT 889.710 29.680 1543.230 29.820 ;
        RECT 889.710 29.620 890.030 29.680 ;
        RECT 1542.910 29.620 1543.230 29.680 ;
      LAYER via ;
        RECT 884.680 1587.160 884.940 1587.420 ;
        RECT 889.740 1587.160 890.000 1587.420 ;
        RECT 889.740 29.620 890.000 29.880 ;
        RECT 1542.940 29.620 1543.200 29.880 ;
      LAYER met2 ;
        RECT 884.540 1600.380 884.820 1604.000 ;
        RECT 884.540 1600.000 884.880 1600.380 ;
        RECT 884.740 1587.450 884.880 1600.000 ;
        RECT 884.680 1587.130 884.940 1587.450 ;
        RECT 889.740 1587.130 890.000 1587.450 ;
        RECT 889.800 29.910 889.940 1587.130 ;
        RECT 889.740 29.590 890.000 29.910 ;
        RECT 1542.940 29.590 1543.200 29.910 ;
        RECT 1543.000 2.400 1543.140 29.590 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 891.090 1587.360 891.410 1587.420 ;
        RECT 895.690 1587.360 896.010 1587.420 ;
        RECT 891.090 1587.220 896.010 1587.360 ;
        RECT 891.090 1587.160 891.410 1587.220 ;
        RECT 895.690 1587.160 896.010 1587.220 ;
        RECT 896.150 30.160 896.470 30.220 ;
        RECT 1560.850 30.160 1561.170 30.220 ;
        RECT 896.150 30.020 1561.170 30.160 ;
        RECT 896.150 29.960 896.470 30.020 ;
        RECT 1560.850 29.960 1561.170 30.020 ;
      LAYER via ;
        RECT 891.120 1587.160 891.380 1587.420 ;
        RECT 895.720 1587.160 895.980 1587.420 ;
        RECT 896.180 29.960 896.440 30.220 ;
        RECT 1560.880 29.960 1561.140 30.220 ;
      LAYER met2 ;
        RECT 890.980 1600.380 891.260 1604.000 ;
        RECT 890.980 1600.000 891.320 1600.380 ;
        RECT 891.180 1587.450 891.320 1600.000 ;
        RECT 891.120 1587.130 891.380 1587.450 ;
        RECT 895.720 1587.130 895.980 1587.450 ;
        RECT 895.780 1579.370 895.920 1587.130 ;
        RECT 895.780 1579.230 896.380 1579.370 ;
        RECT 896.240 30.250 896.380 1579.230 ;
        RECT 896.180 29.930 896.440 30.250 ;
        RECT 1560.880 29.930 1561.140 30.250 ;
        RECT 1560.940 2.400 1561.080 29.930 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 897.070 1587.700 897.390 1587.760 ;
        RECT 903.510 1587.700 903.830 1587.760 ;
        RECT 897.070 1587.560 903.830 1587.700 ;
        RECT 897.070 1587.500 897.390 1587.560 ;
        RECT 903.510 1587.500 903.830 1587.560 ;
        RECT 903.510 30.500 903.830 30.560 ;
        RECT 1578.790 30.500 1579.110 30.560 ;
        RECT 903.510 30.360 1579.110 30.500 ;
        RECT 903.510 30.300 903.830 30.360 ;
        RECT 1578.790 30.300 1579.110 30.360 ;
      LAYER via ;
        RECT 897.100 1587.500 897.360 1587.760 ;
        RECT 903.540 1587.500 903.800 1587.760 ;
        RECT 903.540 30.300 903.800 30.560 ;
        RECT 1578.820 30.300 1579.080 30.560 ;
      LAYER met2 ;
        RECT 896.960 1600.380 897.240 1604.000 ;
        RECT 896.960 1600.000 897.300 1600.380 ;
        RECT 897.160 1587.790 897.300 1600.000 ;
        RECT 897.100 1587.470 897.360 1587.790 ;
        RECT 903.540 1587.470 903.800 1587.790 ;
        RECT 903.600 30.590 903.740 1587.470 ;
        RECT 903.540 30.270 903.800 30.590 ;
        RECT 1578.820 30.270 1579.080 30.590 ;
        RECT 1578.880 2.400 1579.020 30.270 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 903.050 34.240 903.370 34.300 ;
        RECT 1596.270 34.240 1596.590 34.300 ;
        RECT 903.050 34.100 1596.590 34.240 ;
        RECT 903.050 34.040 903.370 34.100 ;
        RECT 1596.270 34.040 1596.590 34.100 ;
      LAYER via ;
        RECT 903.080 34.040 903.340 34.300 ;
        RECT 1596.300 34.040 1596.560 34.300 ;
      LAYER met2 ;
        RECT 903.400 1600.380 903.680 1604.000 ;
        RECT 903.400 1600.000 903.740 1600.380 ;
        RECT 903.600 1588.210 903.740 1600.000 ;
        RECT 903.140 1588.070 903.740 1588.210 ;
        RECT 903.140 34.330 903.280 1588.070 ;
        RECT 903.080 34.010 903.340 34.330 ;
        RECT 1596.300 34.010 1596.560 34.330 ;
        RECT 1596.360 2.400 1596.500 34.010 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 910.410 33.900 910.730 33.960 ;
        RECT 1614.210 33.900 1614.530 33.960 ;
        RECT 910.410 33.760 1614.530 33.900 ;
        RECT 910.410 33.700 910.730 33.760 ;
        RECT 1614.210 33.700 1614.530 33.760 ;
      LAYER via ;
        RECT 910.440 33.700 910.700 33.960 ;
        RECT 1614.240 33.700 1614.500 33.960 ;
      LAYER met2 ;
        RECT 909.380 1600.450 909.660 1604.000 ;
        RECT 909.380 1600.310 910.640 1600.450 ;
        RECT 909.380 1600.000 909.660 1600.310 ;
        RECT 910.500 33.990 910.640 1600.310 ;
        RECT 910.440 33.670 910.700 33.990 ;
        RECT 1614.240 33.670 1614.500 33.990 ;
        RECT 1614.300 2.400 1614.440 33.670 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 917.310 33.560 917.630 33.620 ;
        RECT 1632.150 33.560 1632.470 33.620 ;
        RECT 917.310 33.420 1632.470 33.560 ;
        RECT 917.310 33.360 917.630 33.420 ;
        RECT 1632.150 33.360 1632.470 33.420 ;
      LAYER via ;
        RECT 917.340 33.360 917.600 33.620 ;
        RECT 1632.180 33.360 1632.440 33.620 ;
      LAYER met2 ;
        RECT 915.360 1600.450 915.640 1604.000 ;
        RECT 915.360 1600.310 917.080 1600.450 ;
        RECT 915.360 1600.000 915.640 1600.310 ;
        RECT 916.940 1580.050 917.080 1600.310 ;
        RECT 916.940 1579.910 917.540 1580.050 ;
        RECT 917.400 33.650 917.540 1579.910 ;
        RECT 917.340 33.330 917.600 33.650 ;
        RECT 1632.180 33.330 1632.440 33.650 ;
        RECT 1632.240 2.400 1632.380 33.330 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 921.910 1587.360 922.230 1587.420 ;
        RECT 923.750 1587.360 924.070 1587.420 ;
        RECT 921.910 1587.220 924.070 1587.360 ;
        RECT 921.910 1587.160 922.230 1587.220 ;
        RECT 923.750 1587.160 924.070 1587.220 ;
        RECT 923.750 33.220 924.070 33.280 ;
        RECT 1650.090 33.220 1650.410 33.280 ;
        RECT 923.750 33.080 1650.410 33.220 ;
        RECT 923.750 33.020 924.070 33.080 ;
        RECT 1650.090 33.020 1650.410 33.080 ;
      LAYER via ;
        RECT 921.940 1587.160 922.200 1587.420 ;
        RECT 923.780 1587.160 924.040 1587.420 ;
        RECT 923.780 33.020 924.040 33.280 ;
        RECT 1650.120 33.020 1650.380 33.280 ;
      LAYER met2 ;
        RECT 921.800 1600.380 922.080 1604.000 ;
        RECT 921.800 1600.000 922.140 1600.380 ;
        RECT 922.000 1587.450 922.140 1600.000 ;
        RECT 921.940 1587.130 922.200 1587.450 ;
        RECT 923.780 1587.130 924.040 1587.450 ;
        RECT 923.840 33.310 923.980 1587.130 ;
        RECT 923.780 32.990 924.040 33.310 ;
        RECT 1650.120 32.990 1650.380 33.310 ;
        RECT 1650.180 2.400 1650.320 32.990 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 927.890 1587.360 928.210 1587.420 ;
        RECT 931.110 1587.360 931.430 1587.420 ;
        RECT 927.890 1587.220 931.430 1587.360 ;
        RECT 927.890 1587.160 928.210 1587.220 ;
        RECT 931.110 1587.160 931.430 1587.220 ;
        RECT 931.110 32.880 931.430 32.940 ;
        RECT 1668.030 32.880 1668.350 32.940 ;
        RECT 931.110 32.740 1668.350 32.880 ;
        RECT 931.110 32.680 931.430 32.740 ;
        RECT 1668.030 32.680 1668.350 32.740 ;
      LAYER via ;
        RECT 927.920 1587.160 928.180 1587.420 ;
        RECT 931.140 1587.160 931.400 1587.420 ;
        RECT 931.140 32.680 931.400 32.940 ;
        RECT 1668.060 32.680 1668.320 32.940 ;
      LAYER met2 ;
        RECT 927.780 1600.380 928.060 1604.000 ;
        RECT 927.780 1600.000 928.120 1600.380 ;
        RECT 927.980 1587.450 928.120 1600.000 ;
        RECT 927.920 1587.130 928.180 1587.450 ;
        RECT 931.140 1587.130 931.400 1587.450 ;
        RECT 931.200 32.970 931.340 1587.130 ;
        RECT 931.140 32.650 931.400 32.970 ;
        RECT 1668.060 32.650 1668.320 32.970 ;
        RECT 1668.120 2.400 1668.260 32.650 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 934.330 1587.360 934.650 1587.420 ;
        RECT 937.550 1587.360 937.870 1587.420 ;
        RECT 934.330 1587.220 937.870 1587.360 ;
        RECT 934.330 1587.160 934.650 1587.220 ;
        RECT 937.550 1587.160 937.870 1587.220 ;
        RECT 937.550 32.540 937.870 32.600 ;
        RECT 1685.510 32.540 1685.830 32.600 ;
        RECT 937.550 32.400 1685.830 32.540 ;
        RECT 937.550 32.340 937.870 32.400 ;
        RECT 1685.510 32.340 1685.830 32.400 ;
      LAYER via ;
        RECT 934.360 1587.160 934.620 1587.420 ;
        RECT 937.580 1587.160 937.840 1587.420 ;
        RECT 937.580 32.340 937.840 32.600 ;
        RECT 1685.540 32.340 1685.800 32.600 ;
      LAYER met2 ;
        RECT 934.220 1600.380 934.500 1604.000 ;
        RECT 934.220 1600.000 934.560 1600.380 ;
        RECT 934.420 1587.450 934.560 1600.000 ;
        RECT 934.360 1587.130 934.620 1587.450 ;
        RECT 937.580 1587.130 937.840 1587.450 ;
        RECT 937.640 32.630 937.780 1587.130 ;
        RECT 937.580 32.310 937.840 32.630 ;
        RECT 1685.540 32.310 1685.800 32.630 ;
        RECT 1685.600 2.400 1685.740 32.310 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 684.625 1589.585 684.795 1591.455 ;
      LAYER mcon ;
        RECT 684.625 1591.285 684.795 1591.455 ;
      LAYER met1 ;
        RECT 600.370 1591.440 600.690 1591.500 ;
        RECT 684.565 1591.440 684.855 1591.485 ;
        RECT 600.370 1591.300 684.855 1591.440 ;
        RECT 600.370 1591.240 600.690 1591.300 ;
        RECT 684.565 1591.255 684.855 1591.300 ;
        RECT 684.565 1589.740 684.855 1589.785 ;
        RECT 707.090 1589.740 707.410 1589.800 ;
        RECT 684.565 1589.600 707.410 1589.740 ;
        RECT 684.565 1589.555 684.855 1589.600 ;
        RECT 707.090 1589.540 707.410 1589.600 ;
        RECT 707.090 17.580 707.410 17.640 ;
        RECT 722.270 17.580 722.590 17.640 ;
        RECT 707.090 17.440 722.590 17.580 ;
        RECT 707.090 17.380 707.410 17.440 ;
        RECT 722.270 17.380 722.590 17.440 ;
      LAYER via ;
        RECT 600.400 1591.240 600.660 1591.500 ;
        RECT 707.120 1589.540 707.380 1589.800 ;
        RECT 707.120 17.380 707.380 17.640 ;
        RECT 722.300 17.380 722.560 17.640 ;
      LAYER met2 ;
        RECT 600.260 1600.380 600.540 1604.000 ;
        RECT 600.260 1600.000 600.600 1600.380 ;
        RECT 600.460 1591.530 600.600 1600.000 ;
        RECT 600.400 1591.210 600.660 1591.530 ;
        RECT 707.120 1589.510 707.380 1589.830 ;
        RECT 707.180 17.670 707.320 1589.510 ;
        RECT 707.120 17.350 707.380 17.670 ;
        RECT 722.300 17.350 722.560 17.670 ;
        RECT 722.360 2.400 722.500 17.350 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 940.310 1587.360 940.630 1587.420 ;
        RECT 944.450 1587.360 944.770 1587.420 ;
        RECT 940.310 1587.220 944.770 1587.360 ;
        RECT 940.310 1587.160 940.630 1587.220 ;
        RECT 944.450 1587.160 944.770 1587.220 ;
        RECT 944.450 32.200 944.770 32.260 ;
        RECT 1703.450 32.200 1703.770 32.260 ;
        RECT 944.450 32.060 1703.770 32.200 ;
        RECT 944.450 32.000 944.770 32.060 ;
        RECT 1703.450 32.000 1703.770 32.060 ;
      LAYER via ;
        RECT 940.340 1587.160 940.600 1587.420 ;
        RECT 944.480 1587.160 944.740 1587.420 ;
        RECT 944.480 32.000 944.740 32.260 ;
        RECT 1703.480 32.000 1703.740 32.260 ;
      LAYER met2 ;
        RECT 940.200 1600.380 940.480 1604.000 ;
        RECT 940.200 1600.000 940.540 1600.380 ;
        RECT 940.400 1587.450 940.540 1600.000 ;
        RECT 940.340 1587.130 940.600 1587.450 ;
        RECT 944.480 1587.130 944.740 1587.450 ;
        RECT 944.540 32.290 944.680 1587.130 ;
        RECT 944.480 31.970 944.740 32.290 ;
        RECT 1703.480 31.970 1703.740 32.290 ;
        RECT 1703.540 2.400 1703.680 31.970 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 946.750 1587.360 947.070 1587.420 ;
        RECT 951.810 1587.360 952.130 1587.420 ;
        RECT 946.750 1587.220 952.130 1587.360 ;
        RECT 946.750 1587.160 947.070 1587.220 ;
        RECT 951.810 1587.160 952.130 1587.220 ;
        RECT 951.810 31.860 952.130 31.920 ;
        RECT 1721.390 31.860 1721.710 31.920 ;
        RECT 951.810 31.720 1721.710 31.860 ;
        RECT 951.810 31.660 952.130 31.720 ;
        RECT 1721.390 31.660 1721.710 31.720 ;
      LAYER via ;
        RECT 946.780 1587.160 947.040 1587.420 ;
        RECT 951.840 1587.160 952.100 1587.420 ;
        RECT 951.840 31.660 952.100 31.920 ;
        RECT 1721.420 31.660 1721.680 31.920 ;
      LAYER met2 ;
        RECT 946.640 1600.380 946.920 1604.000 ;
        RECT 946.640 1600.000 946.980 1600.380 ;
        RECT 946.840 1587.450 946.980 1600.000 ;
        RECT 946.780 1587.130 947.040 1587.450 ;
        RECT 951.840 1587.130 952.100 1587.450 ;
        RECT 951.900 31.950 952.040 1587.130 ;
        RECT 951.840 31.630 952.100 31.950 ;
        RECT 1721.420 31.630 1721.680 31.950 ;
        RECT 1721.480 2.400 1721.620 31.630 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 952.730 1587.360 953.050 1587.420 ;
        RECT 958.710 1587.360 959.030 1587.420 ;
        RECT 952.730 1587.220 959.030 1587.360 ;
        RECT 952.730 1587.160 953.050 1587.220 ;
        RECT 958.710 1587.160 959.030 1587.220 ;
        RECT 958.710 31.520 959.030 31.580 ;
        RECT 1739.330 31.520 1739.650 31.580 ;
        RECT 958.710 31.380 1739.650 31.520 ;
        RECT 958.710 31.320 959.030 31.380 ;
        RECT 1739.330 31.320 1739.650 31.380 ;
      LAYER via ;
        RECT 952.760 1587.160 953.020 1587.420 ;
        RECT 958.740 1587.160 959.000 1587.420 ;
        RECT 958.740 31.320 959.000 31.580 ;
        RECT 1739.360 31.320 1739.620 31.580 ;
      LAYER met2 ;
        RECT 952.620 1600.380 952.900 1604.000 ;
        RECT 952.620 1600.000 952.960 1600.380 ;
        RECT 952.820 1587.450 952.960 1600.000 ;
        RECT 952.760 1587.130 953.020 1587.450 ;
        RECT 958.740 1587.130 959.000 1587.450 ;
        RECT 958.800 31.610 958.940 1587.130 ;
        RECT 958.740 31.290 959.000 31.610 ;
        RECT 1739.360 31.290 1739.620 31.610 ;
        RECT 1739.420 2.400 1739.560 31.290 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 959.170 1588.380 959.490 1588.440 ;
        RECT 965.150 1588.380 965.470 1588.440 ;
        RECT 959.170 1588.240 965.470 1588.380 ;
        RECT 959.170 1588.180 959.490 1588.240 ;
        RECT 965.150 1588.180 965.470 1588.240 ;
        RECT 965.150 31.180 965.470 31.240 ;
        RECT 1756.810 31.180 1757.130 31.240 ;
        RECT 965.150 31.040 1757.130 31.180 ;
        RECT 965.150 30.980 965.470 31.040 ;
        RECT 1756.810 30.980 1757.130 31.040 ;
      LAYER via ;
        RECT 959.200 1588.180 959.460 1588.440 ;
        RECT 965.180 1588.180 965.440 1588.440 ;
        RECT 965.180 30.980 965.440 31.240 ;
        RECT 1756.840 30.980 1757.100 31.240 ;
      LAYER met2 ;
        RECT 959.060 1600.380 959.340 1604.000 ;
        RECT 959.060 1600.000 959.400 1600.380 ;
        RECT 959.260 1588.470 959.400 1600.000 ;
        RECT 959.200 1588.150 959.460 1588.470 ;
        RECT 965.180 1588.150 965.440 1588.470 ;
        RECT 965.240 31.270 965.380 1588.150 ;
        RECT 965.180 30.950 965.440 31.270 ;
        RECT 1756.840 30.950 1757.100 31.270 ;
        RECT 1756.900 2.400 1757.040 30.950 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 965.610 30.840 965.930 30.900 ;
        RECT 1774.750 30.840 1775.070 30.900 ;
        RECT 965.610 30.700 1775.070 30.840 ;
        RECT 965.610 30.640 965.930 30.700 ;
        RECT 1774.750 30.640 1775.070 30.700 ;
      LAYER via ;
        RECT 965.640 30.640 965.900 30.900 ;
        RECT 1774.780 30.640 1775.040 30.900 ;
      LAYER met2 ;
        RECT 965.040 1600.450 965.320 1604.000 ;
        RECT 965.040 1600.310 965.840 1600.450 ;
        RECT 965.040 1600.000 965.320 1600.310 ;
        RECT 965.700 30.930 965.840 1600.310 ;
        RECT 965.640 30.610 965.900 30.930 ;
        RECT 1774.780 30.610 1775.040 30.930 ;
        RECT 1774.840 2.400 1774.980 30.610 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.020 1600.450 971.300 1604.000 ;
        RECT 971.020 1600.310 972.280 1600.450 ;
        RECT 971.020 1600.000 971.300 1600.310 ;
        RECT 972.140 33.845 972.280 1600.310 ;
        RECT 972.070 33.475 972.350 33.845 ;
        RECT 1792.710 33.475 1792.990 33.845 ;
        RECT 1792.780 2.400 1792.920 33.475 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
      LAYER via2 ;
        RECT 972.070 33.520 972.350 33.800 ;
        RECT 1792.710 33.520 1792.990 33.800 ;
      LAYER met3 ;
        RECT 972.045 33.810 972.375 33.825 ;
        RECT 1792.685 33.810 1793.015 33.825 ;
        RECT 972.045 33.510 1793.015 33.810 ;
        RECT 972.045 33.495 972.375 33.510 ;
        RECT 1792.685 33.495 1793.015 33.510 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 977.570 1587.360 977.890 1587.420 ;
        RECT 979.410 1587.360 979.730 1587.420 ;
        RECT 977.570 1587.220 979.730 1587.360 ;
        RECT 977.570 1587.160 977.890 1587.220 ;
        RECT 979.410 1587.160 979.730 1587.220 ;
      LAYER via ;
        RECT 977.600 1587.160 977.860 1587.420 ;
        RECT 979.440 1587.160 979.700 1587.420 ;
      LAYER met2 ;
        RECT 977.460 1600.380 977.740 1604.000 ;
        RECT 977.460 1600.000 977.800 1600.380 ;
        RECT 977.660 1587.450 977.800 1600.000 ;
        RECT 977.600 1587.130 977.860 1587.450 ;
        RECT 979.440 1587.130 979.700 1587.450 ;
        RECT 979.500 33.165 979.640 1587.130 ;
        RECT 979.430 32.795 979.710 33.165 ;
        RECT 1810.650 32.795 1810.930 33.165 ;
        RECT 1810.720 2.400 1810.860 32.795 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
      LAYER via2 ;
        RECT 979.430 32.840 979.710 33.120 ;
        RECT 1810.650 32.840 1810.930 33.120 ;
      LAYER met3 ;
        RECT 979.405 33.130 979.735 33.145 ;
        RECT 1810.625 33.130 1810.955 33.145 ;
        RECT 979.405 32.830 1810.955 33.130 ;
        RECT 979.405 32.815 979.735 32.830 ;
        RECT 1810.625 32.815 1810.955 32.830 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 983.550 1587.360 983.870 1587.420 ;
        RECT 986.310 1587.360 986.630 1587.420 ;
        RECT 983.550 1587.220 986.630 1587.360 ;
        RECT 983.550 1587.160 983.870 1587.220 ;
        RECT 986.310 1587.160 986.630 1587.220 ;
      LAYER via ;
        RECT 983.580 1587.160 983.840 1587.420 ;
        RECT 986.340 1587.160 986.600 1587.420 ;
      LAYER met2 ;
        RECT 983.440 1600.380 983.720 1604.000 ;
        RECT 983.440 1600.000 983.780 1600.380 ;
        RECT 983.640 1587.450 983.780 1600.000 ;
        RECT 983.580 1587.130 983.840 1587.450 ;
        RECT 986.340 1587.130 986.600 1587.450 ;
        RECT 986.400 32.485 986.540 1587.130 ;
        RECT 986.330 32.115 986.610 32.485 ;
        RECT 1829.050 32.115 1829.330 32.485 ;
        RECT 1829.120 15.370 1829.260 32.115 ;
        RECT 1828.660 15.230 1829.260 15.370 ;
        RECT 1828.660 2.400 1828.800 15.230 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
      LAYER via2 ;
        RECT 986.330 32.160 986.610 32.440 ;
        RECT 1829.050 32.160 1829.330 32.440 ;
      LAYER met3 ;
        RECT 986.305 32.450 986.635 32.465 ;
        RECT 1829.025 32.450 1829.355 32.465 ;
        RECT 986.305 32.150 1829.355 32.450 ;
        RECT 986.305 32.135 986.635 32.150 ;
        RECT 1829.025 32.135 1829.355 32.150 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 989.990 1587.360 990.310 1587.420 ;
        RECT 993.210 1587.360 993.530 1587.420 ;
        RECT 989.990 1587.220 993.530 1587.360 ;
        RECT 989.990 1587.160 990.310 1587.220 ;
        RECT 993.210 1587.160 993.530 1587.220 ;
      LAYER via ;
        RECT 990.020 1587.160 990.280 1587.420 ;
        RECT 993.240 1587.160 993.500 1587.420 ;
      LAYER met2 ;
        RECT 989.880 1600.380 990.160 1604.000 ;
        RECT 989.880 1600.000 990.220 1600.380 ;
        RECT 990.080 1587.450 990.220 1600.000 ;
        RECT 990.020 1587.130 990.280 1587.450 ;
        RECT 993.240 1587.130 993.500 1587.450 ;
        RECT 993.300 31.805 993.440 1587.130 ;
        RECT 993.230 31.435 993.510 31.805 ;
        RECT 1846.070 31.435 1846.350 31.805 ;
        RECT 1846.140 2.400 1846.280 31.435 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
      LAYER via2 ;
        RECT 993.230 31.480 993.510 31.760 ;
        RECT 1846.070 31.480 1846.350 31.760 ;
      LAYER met3 ;
        RECT 993.205 31.770 993.535 31.785 ;
        RECT 1846.045 31.770 1846.375 31.785 ;
        RECT 993.205 31.470 1846.375 31.770 ;
        RECT 993.205 31.455 993.535 31.470 ;
        RECT 1846.045 31.455 1846.375 31.470 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 995.970 1587.360 996.290 1587.420 ;
        RECT 999.650 1587.360 999.970 1587.420 ;
        RECT 995.970 1587.220 999.970 1587.360 ;
        RECT 995.970 1587.160 996.290 1587.220 ;
        RECT 999.650 1587.160 999.970 1587.220 ;
      LAYER via ;
        RECT 996.000 1587.160 996.260 1587.420 ;
        RECT 999.680 1587.160 999.940 1587.420 ;
      LAYER met2 ;
        RECT 995.860 1600.380 996.140 1604.000 ;
        RECT 995.860 1600.000 996.200 1600.380 ;
        RECT 996.060 1587.450 996.200 1600.000 ;
        RECT 996.000 1587.130 996.260 1587.450 ;
        RECT 999.680 1587.130 999.940 1587.450 ;
        RECT 999.740 31.125 999.880 1587.130 ;
        RECT 999.670 30.755 999.950 31.125 ;
        RECT 1864.010 30.755 1864.290 31.125 ;
        RECT 1864.080 2.400 1864.220 30.755 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
      LAYER via2 ;
        RECT 999.670 30.800 999.950 31.080 ;
        RECT 1864.010 30.800 1864.290 31.080 ;
      LAYER met3 ;
        RECT 999.645 31.090 999.975 31.105 ;
        RECT 1863.985 31.090 1864.315 31.105 ;
        RECT 999.645 30.790 1864.315 31.090 ;
        RECT 999.645 30.775 999.975 30.790 ;
        RECT 1863.985 30.775 1864.315 30.790 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.350 1590.760 606.670 1590.820 ;
        RECT 606.350 1590.620 691.680 1590.760 ;
        RECT 606.350 1590.560 606.670 1590.620 ;
        RECT 691.540 1590.420 691.680 1590.620 ;
        RECT 728.250 1590.420 728.570 1590.480 ;
        RECT 691.540 1590.280 728.570 1590.420 ;
        RECT 728.250 1590.220 728.570 1590.280 ;
        RECT 728.250 17.580 728.570 17.640 ;
        RECT 740.210 17.580 740.530 17.640 ;
        RECT 728.250 17.440 740.530 17.580 ;
        RECT 728.250 17.380 728.570 17.440 ;
        RECT 740.210 17.380 740.530 17.440 ;
      LAYER via ;
        RECT 606.380 1590.560 606.640 1590.820 ;
        RECT 728.280 1590.220 728.540 1590.480 ;
        RECT 728.280 17.380 728.540 17.640 ;
        RECT 740.240 17.380 740.500 17.640 ;
      LAYER met2 ;
        RECT 606.240 1600.380 606.520 1604.000 ;
        RECT 606.240 1600.000 606.580 1600.380 ;
        RECT 606.440 1590.850 606.580 1600.000 ;
        RECT 606.380 1590.530 606.640 1590.850 ;
        RECT 728.280 1590.190 728.540 1590.510 ;
        RECT 728.340 17.670 728.480 1590.190 ;
        RECT 728.280 17.350 728.540 17.670 ;
        RECT 740.240 17.350 740.500 17.670 ;
        RECT 740.300 2.400 740.440 17.350 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1002.410 1587.360 1002.730 1587.420 ;
        RECT 1006.090 1587.360 1006.410 1587.420 ;
        RECT 1002.410 1587.220 1006.410 1587.360 ;
        RECT 1002.410 1587.160 1002.730 1587.220 ;
        RECT 1006.090 1587.160 1006.410 1587.220 ;
        RECT 1006.090 71.980 1006.410 72.040 ;
        RECT 1876.870 71.980 1877.190 72.040 ;
        RECT 1006.090 71.840 1877.190 71.980 ;
        RECT 1006.090 71.780 1006.410 71.840 ;
        RECT 1876.870 71.780 1877.190 71.840 ;
        RECT 1876.870 2.960 1877.190 3.020 ;
        RECT 1881.930 2.960 1882.250 3.020 ;
        RECT 1876.870 2.820 1882.250 2.960 ;
        RECT 1876.870 2.760 1877.190 2.820 ;
        RECT 1881.930 2.760 1882.250 2.820 ;
      LAYER via ;
        RECT 1002.440 1587.160 1002.700 1587.420 ;
        RECT 1006.120 1587.160 1006.380 1587.420 ;
        RECT 1006.120 71.780 1006.380 72.040 ;
        RECT 1876.900 71.780 1877.160 72.040 ;
        RECT 1876.900 2.760 1877.160 3.020 ;
        RECT 1881.960 2.760 1882.220 3.020 ;
      LAYER met2 ;
        RECT 1002.300 1600.380 1002.580 1604.000 ;
        RECT 1002.300 1600.000 1002.640 1600.380 ;
        RECT 1002.500 1587.450 1002.640 1600.000 ;
        RECT 1002.440 1587.130 1002.700 1587.450 ;
        RECT 1006.120 1587.130 1006.380 1587.450 ;
        RECT 1006.180 72.070 1006.320 1587.130 ;
        RECT 1006.120 71.750 1006.380 72.070 ;
        RECT 1876.900 71.750 1877.160 72.070 ;
        RECT 1876.960 3.050 1877.100 71.750 ;
        RECT 1876.900 2.730 1877.160 3.050 ;
        RECT 1881.960 2.730 1882.220 3.050 ;
        RECT 1882.020 2.400 1882.160 2.730 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1008.390 1587.360 1008.710 1587.420 ;
        RECT 1013.910 1587.360 1014.230 1587.420 ;
        RECT 1008.390 1587.220 1014.230 1587.360 ;
        RECT 1008.390 1587.160 1008.710 1587.220 ;
        RECT 1013.910 1587.160 1014.230 1587.220 ;
        RECT 1013.910 75.720 1014.230 75.780 ;
        RECT 1897.570 75.720 1897.890 75.780 ;
        RECT 1013.910 75.580 1897.890 75.720 ;
        RECT 1013.910 75.520 1014.230 75.580 ;
        RECT 1897.570 75.520 1897.890 75.580 ;
        RECT 1897.570 2.960 1897.890 3.020 ;
        RECT 1899.870 2.960 1900.190 3.020 ;
        RECT 1897.570 2.820 1900.190 2.960 ;
        RECT 1897.570 2.760 1897.890 2.820 ;
        RECT 1899.870 2.760 1900.190 2.820 ;
      LAYER via ;
        RECT 1008.420 1587.160 1008.680 1587.420 ;
        RECT 1013.940 1587.160 1014.200 1587.420 ;
        RECT 1013.940 75.520 1014.200 75.780 ;
        RECT 1897.600 75.520 1897.860 75.780 ;
        RECT 1897.600 2.760 1897.860 3.020 ;
        RECT 1899.900 2.760 1900.160 3.020 ;
      LAYER met2 ;
        RECT 1008.280 1600.380 1008.560 1604.000 ;
        RECT 1008.280 1600.000 1008.620 1600.380 ;
        RECT 1008.480 1587.450 1008.620 1600.000 ;
        RECT 1008.420 1587.130 1008.680 1587.450 ;
        RECT 1013.940 1587.130 1014.200 1587.450 ;
        RECT 1014.000 75.810 1014.140 1587.130 ;
        RECT 1013.940 75.490 1014.200 75.810 ;
        RECT 1897.600 75.490 1897.860 75.810 ;
        RECT 1897.660 3.050 1897.800 75.490 ;
        RECT 1897.600 2.730 1897.860 3.050 ;
        RECT 1899.900 2.730 1900.160 3.050 ;
        RECT 1899.960 2.400 1900.100 2.730 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1014.830 1588.720 1015.150 1588.780 ;
        RECT 1020.350 1588.720 1020.670 1588.780 ;
        RECT 1014.830 1588.580 1020.670 1588.720 ;
        RECT 1014.830 1588.520 1015.150 1588.580 ;
        RECT 1020.350 1588.520 1020.670 1588.580 ;
        RECT 1020.350 75.380 1020.670 75.440 ;
        RECT 1911.830 75.380 1912.150 75.440 ;
        RECT 1020.350 75.240 1912.150 75.380 ;
        RECT 1020.350 75.180 1020.670 75.240 ;
        RECT 1911.830 75.180 1912.150 75.240 ;
        RECT 1911.830 18.940 1912.150 19.000 ;
        RECT 1917.810 18.940 1918.130 19.000 ;
        RECT 1911.830 18.800 1918.130 18.940 ;
        RECT 1911.830 18.740 1912.150 18.800 ;
        RECT 1917.810 18.740 1918.130 18.800 ;
      LAYER via ;
        RECT 1014.860 1588.520 1015.120 1588.780 ;
        RECT 1020.380 1588.520 1020.640 1588.780 ;
        RECT 1020.380 75.180 1020.640 75.440 ;
        RECT 1911.860 75.180 1912.120 75.440 ;
        RECT 1911.860 18.740 1912.120 19.000 ;
        RECT 1917.840 18.740 1918.100 19.000 ;
      LAYER met2 ;
        RECT 1014.720 1600.380 1015.000 1604.000 ;
        RECT 1014.720 1600.000 1015.060 1600.380 ;
        RECT 1014.920 1588.810 1015.060 1600.000 ;
        RECT 1014.860 1588.490 1015.120 1588.810 ;
        RECT 1020.380 1588.490 1020.640 1588.810 ;
        RECT 1020.440 75.470 1020.580 1588.490 ;
        RECT 1020.380 75.150 1020.640 75.470 ;
        RECT 1911.860 75.150 1912.120 75.470 ;
        RECT 1911.920 19.030 1912.060 75.150 ;
        RECT 1911.860 18.710 1912.120 19.030 ;
        RECT 1917.840 18.710 1918.100 19.030 ;
        RECT 1917.900 2.400 1918.040 18.710 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1019.890 74.020 1020.210 74.080 ;
        RECT 1932.070 74.020 1932.390 74.080 ;
        RECT 1019.890 73.880 1932.390 74.020 ;
        RECT 1019.890 73.820 1020.210 73.880 ;
        RECT 1932.070 73.820 1932.390 73.880 ;
      LAYER via ;
        RECT 1019.920 73.820 1020.180 74.080 ;
        RECT 1932.100 73.820 1932.360 74.080 ;
      LAYER met2 ;
        RECT 1020.700 1600.450 1020.980 1604.000 ;
        RECT 1019.980 1600.310 1020.980 1600.450 ;
        RECT 1019.980 74.110 1020.120 1600.310 ;
        RECT 1020.700 1600.000 1020.980 1600.310 ;
        RECT 1019.920 73.790 1020.180 74.110 ;
        RECT 1932.100 73.790 1932.360 74.110 ;
        RECT 1932.160 16.730 1932.300 73.790 ;
        RECT 1932.160 16.590 1935.520 16.730 ;
        RECT 1935.380 2.400 1935.520 16.590 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1027.710 35.260 1028.030 35.320 ;
        RECT 1953.230 35.260 1953.550 35.320 ;
        RECT 1027.710 35.120 1953.550 35.260 ;
        RECT 1027.710 35.060 1028.030 35.120 ;
        RECT 1953.230 35.060 1953.550 35.120 ;
      LAYER via ;
        RECT 1027.740 35.060 1028.000 35.320 ;
        RECT 1953.260 35.060 1953.520 35.320 ;
      LAYER met2 ;
        RECT 1026.680 1600.450 1026.960 1604.000 ;
        RECT 1026.680 1600.310 1027.940 1600.450 ;
        RECT 1026.680 1600.000 1026.960 1600.310 ;
        RECT 1027.800 35.350 1027.940 1600.310 ;
        RECT 1027.740 35.030 1028.000 35.350 ;
        RECT 1953.260 35.030 1953.520 35.350 ;
        RECT 1953.320 2.400 1953.460 35.030 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1034.610 35.600 1034.930 35.660 ;
        RECT 1971.170 35.600 1971.490 35.660 ;
        RECT 1034.610 35.460 1971.490 35.600 ;
        RECT 1034.610 35.400 1034.930 35.460 ;
        RECT 1971.170 35.400 1971.490 35.460 ;
      LAYER via ;
        RECT 1034.640 35.400 1034.900 35.660 ;
        RECT 1971.200 35.400 1971.460 35.660 ;
      LAYER met2 ;
        RECT 1033.120 1600.450 1033.400 1604.000 ;
        RECT 1033.120 1600.310 1034.380 1600.450 ;
        RECT 1033.120 1600.000 1033.400 1600.310 ;
        RECT 1034.240 1580.050 1034.380 1600.310 ;
        RECT 1034.240 1579.910 1034.840 1580.050 ;
        RECT 1034.700 35.690 1034.840 1579.910 ;
        RECT 1034.640 35.370 1034.900 35.690 ;
        RECT 1971.200 35.370 1971.460 35.690 ;
        RECT 1971.260 2.400 1971.400 35.370 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.050 35.940 1041.370 36.000 ;
        RECT 1989.110 35.940 1989.430 36.000 ;
        RECT 1041.050 35.800 1989.430 35.940 ;
        RECT 1041.050 35.740 1041.370 35.800 ;
        RECT 1989.110 35.740 1989.430 35.800 ;
      LAYER via ;
        RECT 1041.080 35.740 1041.340 36.000 ;
        RECT 1989.140 35.740 1989.400 36.000 ;
      LAYER met2 ;
        RECT 1039.100 1600.450 1039.380 1604.000 ;
        RECT 1039.100 1600.310 1040.820 1600.450 ;
        RECT 1039.100 1600.000 1039.380 1600.310 ;
        RECT 1040.680 1580.050 1040.820 1600.310 ;
        RECT 1040.680 1579.910 1041.280 1580.050 ;
        RECT 1041.140 36.030 1041.280 1579.910 ;
        RECT 1041.080 35.710 1041.340 36.030 ;
        RECT 1989.140 35.710 1989.400 36.030 ;
        RECT 1989.200 2.400 1989.340 35.710 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1045.650 1587.360 1045.970 1587.420 ;
        RECT 1048.410 1587.360 1048.730 1587.420 ;
        RECT 1045.650 1587.220 1048.730 1587.360 ;
        RECT 1045.650 1587.160 1045.970 1587.220 ;
        RECT 1048.410 1587.160 1048.730 1587.220 ;
        RECT 1048.410 36.280 1048.730 36.340 ;
        RECT 2006.590 36.280 2006.910 36.340 ;
        RECT 1048.410 36.140 2006.910 36.280 ;
        RECT 1048.410 36.080 1048.730 36.140 ;
        RECT 2006.590 36.080 2006.910 36.140 ;
      LAYER via ;
        RECT 1045.680 1587.160 1045.940 1587.420 ;
        RECT 1048.440 1587.160 1048.700 1587.420 ;
        RECT 1048.440 36.080 1048.700 36.340 ;
        RECT 2006.620 36.080 2006.880 36.340 ;
      LAYER met2 ;
        RECT 1045.540 1600.380 1045.820 1604.000 ;
        RECT 1045.540 1600.000 1045.880 1600.380 ;
        RECT 1045.740 1587.450 1045.880 1600.000 ;
        RECT 1045.680 1587.130 1045.940 1587.450 ;
        RECT 1048.440 1587.130 1048.700 1587.450 ;
        RECT 1048.500 36.370 1048.640 1587.130 ;
        RECT 1048.440 36.050 1048.700 36.370 ;
        RECT 2006.620 36.050 2006.880 36.370 ;
        RECT 2006.680 2.400 2006.820 36.050 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1051.630 1587.360 1051.950 1587.420 ;
        RECT 1055.310 1587.360 1055.630 1587.420 ;
        RECT 1051.630 1587.220 1055.630 1587.360 ;
        RECT 1051.630 1587.160 1051.950 1587.220 ;
        RECT 1055.310 1587.160 1055.630 1587.220 ;
        RECT 1055.310 36.620 1055.630 36.680 ;
        RECT 2024.530 36.620 2024.850 36.680 ;
        RECT 1055.310 36.480 2024.850 36.620 ;
        RECT 1055.310 36.420 1055.630 36.480 ;
        RECT 2024.530 36.420 2024.850 36.480 ;
      LAYER via ;
        RECT 1051.660 1587.160 1051.920 1587.420 ;
        RECT 1055.340 1587.160 1055.600 1587.420 ;
        RECT 1055.340 36.420 1055.600 36.680 ;
        RECT 2024.560 36.420 2024.820 36.680 ;
      LAYER met2 ;
        RECT 1051.520 1600.380 1051.800 1604.000 ;
        RECT 1051.520 1600.000 1051.860 1600.380 ;
        RECT 1051.720 1587.450 1051.860 1600.000 ;
        RECT 1051.660 1587.130 1051.920 1587.450 ;
        RECT 1055.340 1587.130 1055.600 1587.450 ;
        RECT 1055.400 36.710 1055.540 1587.130 ;
        RECT 1055.340 36.390 1055.600 36.710 ;
        RECT 2024.560 36.390 2024.820 36.710 ;
        RECT 2024.620 2.400 2024.760 36.390 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1058.070 1590.080 1058.390 1590.140 ;
        RECT 1062.210 1590.080 1062.530 1590.140 ;
        RECT 1058.070 1589.940 1062.530 1590.080 ;
        RECT 1058.070 1589.880 1058.390 1589.940 ;
        RECT 1062.210 1589.880 1062.530 1589.940 ;
        RECT 1062.210 36.960 1062.530 37.020 ;
        RECT 2042.930 36.960 2043.250 37.020 ;
        RECT 1062.210 36.820 2043.250 36.960 ;
        RECT 1062.210 36.760 1062.530 36.820 ;
        RECT 2042.930 36.760 2043.250 36.820 ;
      LAYER via ;
        RECT 1058.100 1589.880 1058.360 1590.140 ;
        RECT 1062.240 1589.880 1062.500 1590.140 ;
        RECT 1062.240 36.760 1062.500 37.020 ;
        RECT 2042.960 36.760 2043.220 37.020 ;
      LAYER met2 ;
        RECT 1057.960 1600.380 1058.240 1604.000 ;
        RECT 1057.960 1600.000 1058.300 1600.380 ;
        RECT 1058.160 1590.170 1058.300 1600.000 ;
        RECT 1058.100 1589.850 1058.360 1590.170 ;
        RECT 1062.240 1589.850 1062.500 1590.170 ;
        RECT 1062.300 37.050 1062.440 1589.850 ;
        RECT 1062.240 36.730 1062.500 37.050 ;
        RECT 2042.960 36.730 2043.220 37.050 ;
        RECT 2043.020 17.410 2043.160 36.730 ;
        RECT 2042.560 17.270 2043.160 17.410 ;
        RECT 2042.560 2.400 2042.700 17.270 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 613.250 19.280 613.570 19.340 ;
        RECT 757.690 19.280 758.010 19.340 ;
        RECT 613.250 19.140 758.010 19.280 ;
        RECT 613.250 19.080 613.570 19.140 ;
        RECT 757.690 19.080 758.010 19.140 ;
      LAYER via ;
        RECT 613.280 19.080 613.540 19.340 ;
        RECT 757.720 19.080 757.980 19.340 ;
      LAYER met2 ;
        RECT 612.680 1600.450 612.960 1604.000 ;
        RECT 612.680 1600.310 613.480 1600.450 ;
        RECT 612.680 1600.000 612.960 1600.310 ;
        RECT 613.340 19.370 613.480 1600.310 ;
        RECT 613.280 19.050 613.540 19.370 ;
        RECT 757.720 19.050 757.980 19.370 ;
        RECT 757.780 2.400 757.920 19.050 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1064.050 1587.360 1064.370 1587.420 ;
        RECT 1068.650 1587.360 1068.970 1587.420 ;
        RECT 1064.050 1587.220 1068.970 1587.360 ;
        RECT 1064.050 1587.160 1064.370 1587.220 ;
        RECT 1068.650 1587.160 1068.970 1587.220 ;
        RECT 1068.650 37.300 1068.970 37.360 ;
        RECT 2060.410 37.300 2060.730 37.360 ;
        RECT 1068.650 37.160 2060.730 37.300 ;
        RECT 1068.650 37.100 1068.970 37.160 ;
        RECT 2060.410 37.100 2060.730 37.160 ;
      LAYER via ;
        RECT 1064.080 1587.160 1064.340 1587.420 ;
        RECT 1068.680 1587.160 1068.940 1587.420 ;
        RECT 1068.680 37.100 1068.940 37.360 ;
        RECT 2060.440 37.100 2060.700 37.360 ;
      LAYER met2 ;
        RECT 1063.940 1600.380 1064.220 1604.000 ;
        RECT 1063.940 1600.000 1064.280 1600.380 ;
        RECT 1064.140 1587.450 1064.280 1600.000 ;
        RECT 1064.080 1587.130 1064.340 1587.450 ;
        RECT 1068.680 1587.130 1068.940 1587.450 ;
        RECT 1068.740 37.390 1068.880 1587.130 ;
        RECT 1068.680 37.070 1068.940 37.390 ;
        RECT 2060.440 37.070 2060.700 37.390 ;
        RECT 2060.500 2.400 2060.640 37.070 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1070.490 1590.080 1070.810 1590.140 ;
        RECT 1076.010 1590.080 1076.330 1590.140 ;
        RECT 1070.490 1589.940 1076.330 1590.080 ;
        RECT 1070.490 1589.880 1070.810 1589.940 ;
        RECT 1076.010 1589.880 1076.330 1589.940 ;
        RECT 1076.010 37.640 1076.330 37.700 ;
        RECT 2078.350 37.640 2078.670 37.700 ;
        RECT 1076.010 37.500 2078.670 37.640 ;
        RECT 1076.010 37.440 1076.330 37.500 ;
        RECT 2078.350 37.440 2078.670 37.500 ;
      LAYER via ;
        RECT 1070.520 1589.880 1070.780 1590.140 ;
        RECT 1076.040 1589.880 1076.300 1590.140 ;
        RECT 1076.040 37.440 1076.300 37.700 ;
        RECT 2078.380 37.440 2078.640 37.700 ;
      LAYER met2 ;
        RECT 1070.380 1600.380 1070.660 1604.000 ;
        RECT 1070.380 1600.000 1070.720 1600.380 ;
        RECT 1070.580 1590.170 1070.720 1600.000 ;
        RECT 1070.520 1589.850 1070.780 1590.170 ;
        RECT 1076.040 1589.850 1076.300 1590.170 ;
        RECT 1076.100 37.730 1076.240 1589.850 ;
        RECT 1076.040 37.410 1076.300 37.730 ;
        RECT 2078.380 37.410 2078.640 37.730 ;
        RECT 2078.440 2.400 2078.580 37.410 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.470 1590.760 1076.790 1590.820 ;
        RECT 1082.450 1590.760 1082.770 1590.820 ;
        RECT 1076.470 1590.620 1082.770 1590.760 ;
        RECT 1076.470 1590.560 1076.790 1590.620 ;
        RECT 1082.450 1590.560 1082.770 1590.620 ;
        RECT 1082.450 41.380 1082.770 41.440 ;
        RECT 2095.830 41.380 2096.150 41.440 ;
        RECT 1082.450 41.240 2096.150 41.380 ;
        RECT 1082.450 41.180 1082.770 41.240 ;
        RECT 2095.830 41.180 2096.150 41.240 ;
      LAYER via ;
        RECT 1076.500 1590.560 1076.760 1590.820 ;
        RECT 1082.480 1590.560 1082.740 1590.820 ;
        RECT 1082.480 41.180 1082.740 41.440 ;
        RECT 2095.860 41.180 2096.120 41.440 ;
      LAYER met2 ;
        RECT 1076.360 1600.380 1076.640 1604.000 ;
        RECT 1076.360 1600.000 1076.700 1600.380 ;
        RECT 1076.560 1590.850 1076.700 1600.000 ;
        RECT 1076.500 1590.530 1076.760 1590.850 ;
        RECT 1082.480 1590.530 1082.740 1590.850 ;
        RECT 1082.540 41.470 1082.680 1590.530 ;
        RECT 1082.480 41.150 1082.740 41.470 ;
        RECT 2095.860 41.150 2096.120 41.470 ;
        RECT 2095.920 2.400 2096.060 41.150 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1082.910 41.040 1083.230 41.100 ;
        RECT 2113.770 41.040 2114.090 41.100 ;
        RECT 1082.910 40.900 2114.090 41.040 ;
        RECT 1082.910 40.840 1083.230 40.900 ;
        RECT 2113.770 40.840 2114.090 40.900 ;
      LAYER via ;
        RECT 1082.940 40.840 1083.200 41.100 ;
        RECT 2113.800 40.840 2114.060 41.100 ;
      LAYER met2 ;
        RECT 1082.340 1600.450 1082.620 1604.000 ;
        RECT 1082.340 1600.310 1083.140 1600.450 ;
        RECT 1082.340 1600.000 1082.620 1600.310 ;
        RECT 1083.000 41.130 1083.140 1600.310 ;
        RECT 1082.940 40.810 1083.200 41.130 ;
        RECT 2113.800 40.810 2114.060 41.130 ;
        RECT 2113.860 2.400 2114.000 40.810 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1089.810 40.700 1090.130 40.760 ;
        RECT 2131.710 40.700 2132.030 40.760 ;
        RECT 1089.810 40.560 2132.030 40.700 ;
        RECT 1089.810 40.500 1090.130 40.560 ;
        RECT 2131.710 40.500 2132.030 40.560 ;
      LAYER via ;
        RECT 1089.840 40.500 1090.100 40.760 ;
        RECT 2131.740 40.500 2132.000 40.760 ;
      LAYER met2 ;
        RECT 1088.780 1600.450 1089.060 1604.000 ;
        RECT 1088.780 1600.310 1090.040 1600.450 ;
        RECT 1088.780 1600.000 1089.060 1600.310 ;
        RECT 1089.900 40.790 1090.040 1600.310 ;
        RECT 1089.840 40.470 1090.100 40.790 ;
        RECT 2131.740 40.470 2132.000 40.790 ;
        RECT 2131.800 2.400 2131.940 40.470 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.250 40.360 1096.570 40.420 ;
        RECT 2149.650 40.360 2149.970 40.420 ;
        RECT 1096.250 40.220 2149.970 40.360 ;
        RECT 1096.250 40.160 1096.570 40.220 ;
        RECT 2149.650 40.160 2149.970 40.220 ;
      LAYER via ;
        RECT 1096.280 40.160 1096.540 40.420 ;
        RECT 2149.680 40.160 2149.940 40.420 ;
      LAYER met2 ;
        RECT 1094.760 1600.450 1095.040 1604.000 ;
        RECT 1094.760 1600.310 1096.480 1600.450 ;
        RECT 1094.760 1600.000 1095.040 1600.310 ;
        RECT 1096.340 40.450 1096.480 1600.310 ;
        RECT 1096.280 40.130 1096.540 40.450 ;
        RECT 2149.680 40.130 2149.940 40.450 ;
        RECT 2149.740 2.400 2149.880 40.130 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1101.310 1590.760 1101.630 1590.820 ;
        RECT 1103.610 1590.760 1103.930 1590.820 ;
        RECT 1101.310 1590.620 1103.930 1590.760 ;
        RECT 1101.310 1590.560 1101.630 1590.620 ;
        RECT 1103.610 1590.560 1103.930 1590.620 ;
        RECT 1103.610 40.020 1103.930 40.080 ;
        RECT 2167.590 40.020 2167.910 40.080 ;
        RECT 1103.610 39.880 2167.910 40.020 ;
        RECT 1103.610 39.820 1103.930 39.880 ;
        RECT 2167.590 39.820 2167.910 39.880 ;
      LAYER via ;
        RECT 1101.340 1590.560 1101.600 1590.820 ;
        RECT 1103.640 1590.560 1103.900 1590.820 ;
        RECT 1103.640 39.820 1103.900 40.080 ;
        RECT 2167.620 39.820 2167.880 40.080 ;
      LAYER met2 ;
        RECT 1101.200 1600.380 1101.480 1604.000 ;
        RECT 1101.200 1600.000 1101.540 1600.380 ;
        RECT 1101.400 1590.850 1101.540 1600.000 ;
        RECT 1101.340 1590.530 1101.600 1590.850 ;
        RECT 1103.640 1590.530 1103.900 1590.850 ;
        RECT 1103.700 40.110 1103.840 1590.530 ;
        RECT 1103.640 39.790 1103.900 40.110 ;
        RECT 2167.620 39.790 2167.880 40.110 ;
        RECT 2167.680 2.400 2167.820 39.790 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1107.290 1590.080 1107.610 1590.140 ;
        RECT 1110.050 1590.080 1110.370 1590.140 ;
        RECT 1107.290 1589.940 1110.370 1590.080 ;
        RECT 1107.290 1589.880 1107.610 1589.940 ;
        RECT 1110.050 1589.880 1110.370 1589.940 ;
        RECT 1110.050 39.680 1110.370 39.740 ;
        RECT 2185.070 39.680 2185.390 39.740 ;
        RECT 1110.050 39.540 2185.390 39.680 ;
        RECT 1110.050 39.480 1110.370 39.540 ;
        RECT 2185.070 39.480 2185.390 39.540 ;
      LAYER via ;
        RECT 1107.320 1589.880 1107.580 1590.140 ;
        RECT 1110.080 1589.880 1110.340 1590.140 ;
        RECT 1110.080 39.480 1110.340 39.740 ;
        RECT 2185.100 39.480 2185.360 39.740 ;
      LAYER met2 ;
        RECT 1107.180 1600.380 1107.460 1604.000 ;
        RECT 1107.180 1600.000 1107.520 1600.380 ;
        RECT 1107.380 1590.170 1107.520 1600.000 ;
        RECT 1107.320 1589.850 1107.580 1590.170 ;
        RECT 1110.080 1589.850 1110.340 1590.170 ;
        RECT 1110.140 39.770 1110.280 1589.850 ;
        RECT 1110.080 39.450 1110.340 39.770 ;
        RECT 2185.100 39.450 2185.360 39.770 ;
        RECT 2185.160 2.400 2185.300 39.450 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1113.730 1590.080 1114.050 1590.140 ;
        RECT 1117.410 1590.080 1117.730 1590.140 ;
        RECT 1113.730 1589.940 1117.730 1590.080 ;
        RECT 1113.730 1589.880 1114.050 1589.940 ;
        RECT 1117.410 1589.880 1117.730 1589.940 ;
        RECT 1117.410 39.340 1117.730 39.400 ;
        RECT 2203.010 39.340 2203.330 39.400 ;
        RECT 1117.410 39.200 2203.330 39.340 ;
        RECT 1117.410 39.140 1117.730 39.200 ;
        RECT 2203.010 39.140 2203.330 39.200 ;
      LAYER via ;
        RECT 1113.760 1589.880 1114.020 1590.140 ;
        RECT 1117.440 1589.880 1117.700 1590.140 ;
        RECT 1117.440 39.140 1117.700 39.400 ;
        RECT 2203.040 39.140 2203.300 39.400 ;
      LAYER met2 ;
        RECT 1113.620 1600.380 1113.900 1604.000 ;
        RECT 1113.620 1600.000 1113.960 1600.380 ;
        RECT 1113.820 1590.170 1113.960 1600.000 ;
        RECT 1113.760 1589.850 1114.020 1590.170 ;
        RECT 1117.440 1589.850 1117.700 1590.170 ;
        RECT 1117.500 39.430 1117.640 1589.850 ;
        RECT 1117.440 39.110 1117.700 39.430 ;
        RECT 2203.040 39.110 2203.300 39.430 ;
        RECT 2203.100 2.400 2203.240 39.110 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1119.710 1590.080 1120.030 1590.140 ;
        RECT 1123.850 1590.080 1124.170 1590.140 ;
        RECT 1119.710 1589.940 1124.170 1590.080 ;
        RECT 1119.710 1589.880 1120.030 1589.940 ;
        RECT 1123.850 1589.880 1124.170 1589.940 ;
        RECT 1123.850 39.000 1124.170 39.060 ;
        RECT 2220.950 39.000 2221.270 39.060 ;
        RECT 1123.850 38.860 2221.270 39.000 ;
        RECT 1123.850 38.800 1124.170 38.860 ;
        RECT 2220.950 38.800 2221.270 38.860 ;
      LAYER via ;
        RECT 1119.740 1589.880 1120.000 1590.140 ;
        RECT 1123.880 1589.880 1124.140 1590.140 ;
        RECT 1123.880 38.800 1124.140 39.060 ;
        RECT 2220.980 38.800 2221.240 39.060 ;
      LAYER met2 ;
        RECT 1119.600 1600.380 1119.880 1604.000 ;
        RECT 1119.600 1600.000 1119.940 1600.380 ;
        RECT 1119.800 1590.170 1119.940 1600.000 ;
        RECT 1119.740 1589.850 1120.000 1590.170 ;
        RECT 1123.880 1589.850 1124.140 1590.170 ;
        RECT 1123.940 39.090 1124.080 1589.850 ;
        RECT 1123.880 38.770 1124.140 39.090 ;
        RECT 2220.980 38.770 2221.240 39.090 ;
        RECT 2221.040 2.400 2221.180 38.770 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 618.770 1592.120 619.090 1592.180 ;
        RECT 736.990 1592.120 737.310 1592.180 ;
        RECT 618.770 1591.980 737.310 1592.120 ;
        RECT 618.770 1591.920 619.090 1591.980 ;
        RECT 736.990 1591.920 737.310 1591.980 ;
        RECT 739.290 1590.760 739.610 1590.820 ;
        RECT 754.470 1590.760 754.790 1590.820 ;
        RECT 739.290 1590.620 754.790 1590.760 ;
        RECT 739.290 1590.560 739.610 1590.620 ;
        RECT 754.470 1590.560 754.790 1590.620 ;
        RECT 754.470 1563.220 754.790 1563.280 ;
        RECT 755.850 1563.220 756.170 1563.280 ;
        RECT 754.470 1563.080 756.170 1563.220 ;
        RECT 754.470 1563.020 754.790 1563.080 ;
        RECT 755.850 1563.020 756.170 1563.080 ;
        RECT 755.850 19.620 756.170 19.680 ;
        RECT 775.630 19.620 775.950 19.680 ;
        RECT 755.850 19.480 775.950 19.620 ;
        RECT 755.850 19.420 756.170 19.480 ;
        RECT 775.630 19.420 775.950 19.480 ;
      LAYER via ;
        RECT 618.800 1591.920 619.060 1592.180 ;
        RECT 737.020 1591.920 737.280 1592.180 ;
        RECT 739.320 1590.560 739.580 1590.820 ;
        RECT 754.500 1590.560 754.760 1590.820 ;
        RECT 754.500 1563.020 754.760 1563.280 ;
        RECT 755.880 1563.020 756.140 1563.280 ;
        RECT 755.880 19.420 756.140 19.680 ;
        RECT 775.660 19.420 775.920 19.680 ;
      LAYER met2 ;
        RECT 618.660 1600.380 618.940 1604.000 ;
        RECT 618.660 1600.000 619.000 1600.380 ;
        RECT 618.860 1592.210 619.000 1600.000 ;
        RECT 618.800 1591.890 619.060 1592.210 ;
        RECT 737.020 1591.890 737.280 1592.210 ;
        RECT 737.080 1591.045 737.220 1591.890 ;
        RECT 737.010 1590.675 737.290 1591.045 ;
        RECT 739.310 1590.675 739.590 1591.045 ;
        RECT 739.320 1590.530 739.580 1590.675 ;
        RECT 754.500 1590.530 754.760 1590.850 ;
        RECT 754.560 1563.310 754.700 1590.530 ;
        RECT 754.500 1562.990 754.760 1563.310 ;
        RECT 755.880 1562.990 756.140 1563.310 ;
        RECT 755.940 19.710 756.080 1562.990 ;
        RECT 755.880 19.390 756.140 19.710 ;
        RECT 775.660 19.390 775.920 19.710 ;
        RECT 775.720 2.400 775.860 19.390 ;
        RECT 775.510 -4.800 776.070 2.400 ;
      LAYER via2 ;
        RECT 737.010 1590.720 737.290 1591.000 ;
        RECT 739.310 1590.720 739.590 1591.000 ;
      LAYER met3 ;
        RECT 736.985 1591.010 737.315 1591.025 ;
        RECT 739.285 1591.010 739.615 1591.025 ;
        RECT 736.985 1590.710 739.615 1591.010 ;
        RECT 736.985 1590.695 737.315 1590.710 ;
        RECT 739.285 1590.695 739.615 1590.710 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1124.770 1535.340 1125.090 1535.400 ;
        RECT 1130.750 1535.340 1131.070 1535.400 ;
        RECT 1124.770 1535.200 1131.070 1535.340 ;
        RECT 1124.770 1535.140 1125.090 1535.200 ;
        RECT 1130.750 1535.140 1131.070 1535.200 ;
        RECT 1130.750 38.660 1131.070 38.720 ;
        RECT 2238.890 38.660 2239.210 38.720 ;
        RECT 1130.750 38.520 2239.210 38.660 ;
        RECT 1130.750 38.460 1131.070 38.520 ;
        RECT 2238.890 38.460 2239.210 38.520 ;
      LAYER via ;
        RECT 1124.800 1535.140 1125.060 1535.400 ;
        RECT 1130.780 1535.140 1131.040 1535.400 ;
        RECT 1130.780 38.460 1131.040 38.720 ;
        RECT 2238.920 38.460 2239.180 38.720 ;
      LAYER met2 ;
        RECT 1126.040 1600.450 1126.320 1604.000 ;
        RECT 1124.860 1600.310 1126.320 1600.450 ;
        RECT 1124.860 1535.430 1125.000 1600.310 ;
        RECT 1126.040 1600.000 1126.320 1600.310 ;
        RECT 1124.800 1535.110 1125.060 1535.430 ;
        RECT 1130.780 1535.110 1131.040 1535.430 ;
        RECT 1130.840 38.750 1130.980 1535.110 ;
        RECT 1130.780 38.430 1131.040 38.750 ;
        RECT 2238.920 38.430 2239.180 38.750 ;
        RECT 2238.980 2.400 2239.120 38.430 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1132.130 1590.080 1132.450 1590.140 ;
        RECT 1138.110 1590.080 1138.430 1590.140 ;
        RECT 1132.130 1589.940 1138.430 1590.080 ;
        RECT 1132.130 1589.880 1132.450 1589.940 ;
        RECT 1138.110 1589.880 1138.430 1589.940 ;
        RECT 1138.110 38.320 1138.430 38.380 ;
        RECT 2256.830 38.320 2257.150 38.380 ;
        RECT 1138.110 38.180 2257.150 38.320 ;
        RECT 1138.110 38.120 1138.430 38.180 ;
        RECT 2256.830 38.120 2257.150 38.180 ;
      LAYER via ;
        RECT 1132.160 1589.880 1132.420 1590.140 ;
        RECT 1138.140 1589.880 1138.400 1590.140 ;
        RECT 1138.140 38.120 1138.400 38.380 ;
        RECT 2256.860 38.120 2257.120 38.380 ;
      LAYER met2 ;
        RECT 1132.020 1600.380 1132.300 1604.000 ;
        RECT 1132.020 1600.000 1132.360 1600.380 ;
        RECT 1132.220 1590.170 1132.360 1600.000 ;
        RECT 1132.160 1589.850 1132.420 1590.170 ;
        RECT 1138.140 1589.850 1138.400 1590.170 ;
        RECT 1138.200 38.410 1138.340 1589.850 ;
        RECT 1138.140 38.090 1138.400 38.410 ;
        RECT 2256.860 38.090 2257.120 38.410 ;
        RECT 2256.920 7.210 2257.060 38.090 ;
        RECT 2256.460 7.070 2257.060 7.210 ;
        RECT 2256.460 2.400 2256.600 7.070 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1137.650 37.980 1137.970 38.040 ;
        RECT 2274.310 37.980 2274.630 38.040 ;
        RECT 1137.650 37.840 2274.630 37.980 ;
        RECT 1137.650 37.780 1137.970 37.840 ;
        RECT 2274.310 37.780 2274.630 37.840 ;
      LAYER via ;
        RECT 1137.680 37.780 1137.940 38.040 ;
        RECT 2274.340 37.780 2274.600 38.040 ;
      LAYER met2 ;
        RECT 1138.000 1600.380 1138.280 1604.000 ;
        RECT 1138.000 1600.000 1138.340 1600.380 ;
        RECT 1138.200 1590.930 1138.340 1600.000 ;
        RECT 1137.740 1590.790 1138.340 1590.930 ;
        RECT 1137.740 38.070 1137.880 1590.790 ;
        RECT 1137.680 37.750 1137.940 38.070 ;
        RECT 2274.340 37.750 2274.600 38.070 ;
        RECT 2274.400 2.400 2274.540 37.750 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.440 1600.380 1144.720 1604.000 ;
        RECT 1144.440 1600.000 1144.780 1600.380 ;
        RECT 1144.640 41.325 1144.780 1600.000 ;
        RECT 1144.570 40.955 1144.850 41.325 ;
        RECT 2292.270 40.955 2292.550 41.325 ;
        RECT 2292.340 2.400 2292.480 40.955 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
      LAYER via2 ;
        RECT 1144.570 41.000 1144.850 41.280 ;
        RECT 2292.270 41.000 2292.550 41.280 ;
      LAYER met3 ;
        RECT 1144.545 41.290 1144.875 41.305 ;
        RECT 2292.245 41.290 2292.575 41.305 ;
        RECT 1144.545 40.990 2292.575 41.290 ;
        RECT 1144.545 40.975 1144.875 40.990 ;
        RECT 2292.245 40.975 2292.575 40.990 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.420 1600.450 1150.700 1604.000 ;
        RECT 1150.420 1600.310 1152.140 1600.450 ;
        RECT 1150.420 1600.000 1150.700 1600.310 ;
        RECT 1152.000 40.645 1152.140 1600.310 ;
        RECT 1151.930 40.275 1152.210 40.645 ;
        RECT 2310.210 40.275 2310.490 40.645 ;
        RECT 2310.280 2.400 2310.420 40.275 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
      LAYER via2 ;
        RECT 1151.930 40.320 1152.210 40.600 ;
        RECT 2310.210 40.320 2310.490 40.600 ;
      LAYER met3 ;
        RECT 1151.905 40.610 1152.235 40.625 ;
        RECT 2310.185 40.610 2310.515 40.625 ;
        RECT 1151.905 40.310 2310.515 40.610 ;
        RECT 1151.905 40.295 1152.235 40.310 ;
        RECT 2310.185 40.295 2310.515 40.310 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.860 1600.450 1157.140 1604.000 ;
        RECT 1156.860 1600.310 1157.660 1600.450 ;
        RECT 1156.860 1600.000 1157.140 1600.310 ;
        RECT 1157.520 1590.930 1157.660 1600.310 ;
        RECT 1157.520 1590.790 1158.120 1590.930 ;
        RECT 1157.980 1579.370 1158.120 1590.790 ;
        RECT 1157.980 1579.230 1158.580 1579.370 ;
        RECT 1158.440 39.965 1158.580 1579.230 ;
        RECT 1158.370 39.595 1158.650 39.965 ;
        RECT 2328.150 39.595 2328.430 39.965 ;
        RECT 2328.220 2.400 2328.360 39.595 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
      LAYER via2 ;
        RECT 1158.370 39.640 1158.650 39.920 ;
        RECT 2328.150 39.640 2328.430 39.920 ;
      LAYER met3 ;
        RECT 1158.345 39.930 1158.675 39.945 ;
        RECT 2328.125 39.930 2328.455 39.945 ;
        RECT 1158.345 39.630 2328.455 39.930 ;
        RECT 1158.345 39.615 1158.675 39.630 ;
        RECT 2328.125 39.615 2328.455 39.630 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1160.190 1511.200 1160.510 1511.260 ;
        RECT 1165.710 1511.200 1166.030 1511.260 ;
        RECT 1160.190 1511.060 1166.030 1511.200 ;
        RECT 1160.190 1511.000 1160.510 1511.060 ;
        RECT 1165.710 1511.000 1166.030 1511.060 ;
      LAYER via ;
        RECT 1160.220 1511.000 1160.480 1511.260 ;
        RECT 1165.740 1511.000 1166.000 1511.260 ;
      LAYER met2 ;
        RECT 1162.840 1600.450 1163.120 1604.000 ;
        RECT 1162.120 1600.310 1163.120 1600.450 ;
        RECT 1162.120 1580.050 1162.260 1600.310 ;
        RECT 1162.840 1600.000 1163.120 1600.310 ;
        RECT 1160.280 1579.910 1162.260 1580.050 ;
        RECT 1160.280 1511.290 1160.420 1579.910 ;
        RECT 1160.220 1510.970 1160.480 1511.290 ;
        RECT 1165.740 1510.970 1166.000 1511.290 ;
        RECT 1165.800 39.285 1165.940 1510.970 ;
        RECT 1165.730 38.915 1166.010 39.285 ;
        RECT 2345.630 38.915 2345.910 39.285 ;
        RECT 2345.700 2.400 2345.840 38.915 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
      LAYER via2 ;
        RECT 1165.730 38.960 1166.010 39.240 ;
        RECT 2345.630 38.960 2345.910 39.240 ;
      LAYER met3 ;
        RECT 1165.705 39.250 1166.035 39.265 ;
        RECT 2345.605 39.250 2345.935 39.265 ;
        RECT 1165.705 38.950 2345.935 39.250 ;
        RECT 1165.705 38.935 1166.035 38.950 ;
        RECT 2345.605 38.935 2345.935 38.950 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1167.090 1511.340 1167.410 1511.600 ;
        RECT 1167.180 1511.200 1167.320 1511.340 ;
        RECT 1172.150 1511.200 1172.470 1511.260 ;
        RECT 1167.180 1511.060 1172.470 1511.200 ;
        RECT 1172.150 1511.000 1172.470 1511.060 ;
      LAYER via ;
        RECT 1167.120 1511.340 1167.380 1511.600 ;
        RECT 1172.180 1511.000 1172.440 1511.260 ;
      LAYER met2 ;
        RECT 1169.280 1600.450 1169.560 1604.000 ;
        RECT 1168.100 1600.310 1169.560 1600.450 ;
        RECT 1168.100 1580.050 1168.240 1600.310 ;
        RECT 1169.280 1600.000 1169.560 1600.310 ;
        RECT 1167.180 1579.910 1168.240 1580.050 ;
        RECT 1167.180 1511.630 1167.320 1579.910 ;
        RECT 1167.120 1511.310 1167.380 1511.630 ;
        RECT 1172.180 1510.970 1172.440 1511.290 ;
        RECT 1172.240 50.050 1172.380 1510.970 ;
        RECT 1171.780 49.910 1172.380 50.050 ;
        RECT 1171.780 38.605 1171.920 49.910 ;
        RECT 1171.710 38.235 1171.990 38.605 ;
        RECT 2363.570 38.235 2363.850 38.605 ;
        RECT 2363.640 2.400 2363.780 38.235 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
      LAYER via2 ;
        RECT 1171.710 38.280 1171.990 38.560 ;
        RECT 2363.570 38.280 2363.850 38.560 ;
      LAYER met3 ;
        RECT 1171.685 38.570 1172.015 38.585 ;
        RECT 2363.545 38.570 2363.875 38.585 ;
        RECT 1171.685 38.270 2363.875 38.570 ;
        RECT 1171.685 38.255 1172.015 38.270 ;
        RECT 2363.545 38.255 2363.875 38.270 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.260 1600.450 1175.540 1604.000 ;
        RECT 1175.260 1600.310 1176.980 1600.450 ;
        RECT 1175.260 1600.000 1175.540 1600.310 ;
        RECT 1176.840 1579.370 1176.980 1600.310 ;
        RECT 1176.840 1579.230 1179.740 1579.370 ;
        RECT 1179.600 37.925 1179.740 1579.230 ;
        RECT 1179.530 37.555 1179.810 37.925 ;
        RECT 2381.510 37.555 2381.790 37.925 ;
        RECT 2381.580 2.400 2381.720 37.555 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
      LAYER via2 ;
        RECT 1179.530 37.600 1179.810 37.880 ;
        RECT 2381.510 37.600 2381.790 37.880 ;
      LAYER met3 ;
        RECT 1179.505 37.890 1179.835 37.905 ;
        RECT 2381.485 37.890 2381.815 37.905 ;
        RECT 1179.505 37.590 2381.815 37.890 ;
        RECT 1179.505 37.575 1179.835 37.590 ;
        RECT 2381.485 37.575 2381.815 37.590 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1180.965 1538.925 1181.135 1587.035 ;
      LAYER mcon ;
        RECT 1180.965 1586.865 1181.135 1587.035 ;
      LAYER met1 ;
        RECT 1180.890 1587.020 1181.210 1587.080 ;
        RECT 1180.695 1586.880 1181.210 1587.020 ;
        RECT 1180.890 1586.820 1181.210 1586.880 ;
        RECT 1180.890 1539.080 1181.210 1539.140 ;
        RECT 1180.695 1538.940 1181.210 1539.080 ;
        RECT 1180.890 1538.880 1181.210 1538.940 ;
        RECT 1180.890 1533.640 1181.210 1533.700 ;
        RECT 1185.490 1533.640 1185.810 1533.700 ;
        RECT 1180.890 1533.500 1185.810 1533.640 ;
        RECT 1180.890 1533.440 1181.210 1533.500 ;
        RECT 1185.490 1533.440 1185.810 1533.500 ;
        RECT 1185.490 73.340 1185.810 73.400 ;
        RECT 2394.370 73.340 2394.690 73.400 ;
        RECT 1185.490 73.200 2394.690 73.340 ;
        RECT 1185.490 73.140 1185.810 73.200 ;
        RECT 2394.370 73.140 2394.690 73.200 ;
        RECT 2394.370 2.960 2394.690 3.020 ;
        RECT 2399.430 2.960 2399.750 3.020 ;
        RECT 2394.370 2.820 2399.750 2.960 ;
        RECT 2394.370 2.760 2394.690 2.820 ;
        RECT 2399.430 2.760 2399.750 2.820 ;
      LAYER via ;
        RECT 1180.920 1586.820 1181.180 1587.080 ;
        RECT 1180.920 1538.880 1181.180 1539.140 ;
        RECT 1180.920 1533.440 1181.180 1533.700 ;
        RECT 1185.520 1533.440 1185.780 1533.700 ;
        RECT 1185.520 73.140 1185.780 73.400 ;
        RECT 2394.400 73.140 2394.660 73.400 ;
        RECT 2394.400 2.760 2394.660 3.020 ;
        RECT 2399.460 2.760 2399.720 3.020 ;
      LAYER met2 ;
        RECT 1181.700 1600.450 1181.980 1604.000 ;
        RECT 1180.980 1600.310 1181.980 1600.450 ;
        RECT 1180.980 1587.110 1181.120 1600.310 ;
        RECT 1181.700 1600.000 1181.980 1600.310 ;
        RECT 1180.920 1586.790 1181.180 1587.110 ;
        RECT 1180.920 1538.850 1181.180 1539.170 ;
        RECT 1180.980 1533.730 1181.120 1538.850 ;
        RECT 1180.920 1533.410 1181.180 1533.730 ;
        RECT 1185.520 1533.410 1185.780 1533.730 ;
        RECT 1185.580 1448.810 1185.720 1533.410 ;
        RECT 1185.580 1448.670 1186.180 1448.810 ;
        RECT 1186.040 134.370 1186.180 1448.670 ;
        RECT 1185.580 134.230 1186.180 134.370 ;
        RECT 1185.580 73.430 1185.720 134.230 ;
        RECT 1185.520 73.110 1185.780 73.430 ;
        RECT 2394.400 73.110 2394.660 73.430 ;
        RECT 2394.460 3.050 2394.600 73.110 ;
        RECT 2394.400 2.730 2394.660 3.050 ;
        RECT 2399.460 2.730 2399.720 3.050 ;
        RECT 2399.520 2.400 2399.660 2.730 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 639.545 16.745 639.715 20.995 ;
        RECT 745.345 16.065 745.515 16.915 ;
      LAYER mcon ;
        RECT 639.545 20.825 639.715 20.995 ;
        RECT 745.345 16.745 745.515 16.915 ;
      LAYER met1 ;
        RECT 639.485 20.980 639.775 21.025 ;
        RECT 637.720 20.840 639.775 20.980 ;
        RECT 626.590 20.640 626.910 20.700 ;
        RECT 637.720 20.640 637.860 20.840 ;
        RECT 639.485 20.795 639.775 20.840 ;
        RECT 626.590 20.500 637.860 20.640 ;
        RECT 626.590 20.440 626.910 20.500 ;
        RECT 639.485 16.900 639.775 16.945 ;
        RECT 745.285 16.900 745.575 16.945 ;
        RECT 639.485 16.760 745.575 16.900 ;
        RECT 639.485 16.715 639.775 16.760 ;
        RECT 745.285 16.715 745.575 16.760 ;
        RECT 745.285 16.220 745.575 16.265 ;
        RECT 793.570 16.220 793.890 16.280 ;
        RECT 745.285 16.080 793.890 16.220 ;
        RECT 745.285 16.035 745.575 16.080 ;
        RECT 793.570 16.020 793.890 16.080 ;
      LAYER via ;
        RECT 626.620 20.440 626.880 20.700 ;
        RECT 793.600 16.020 793.860 16.280 ;
      LAYER met2 ;
        RECT 625.100 1600.450 625.380 1604.000 ;
        RECT 625.100 1600.310 625.900 1600.450 ;
        RECT 625.100 1600.000 625.380 1600.310 ;
        RECT 625.760 1590.250 625.900 1600.310 ;
        RECT 625.760 1590.110 626.820 1590.250 ;
        RECT 626.680 20.730 626.820 1590.110 ;
        RECT 626.620 20.410 626.880 20.730 ;
        RECT 793.600 15.990 793.860 16.310 ;
        RECT 793.660 2.400 793.800 15.990 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 571.390 20.300 571.710 20.360 ;
        RECT 637.630 20.300 637.950 20.360 ;
        RECT 571.390 20.160 637.950 20.300 ;
        RECT 571.390 20.100 571.710 20.160 ;
        RECT 637.630 20.100 637.950 20.160 ;
      LAYER via ;
        RECT 571.420 20.100 571.680 20.360 ;
        RECT 637.660 20.100 637.920 20.360 ;
      LAYER met2 ;
        RECT 571.280 1600.380 571.560 1604.000 ;
        RECT 571.280 1600.000 571.620 1600.380 ;
        RECT 571.480 20.390 571.620 1600.000 ;
        RECT 571.420 20.070 571.680 20.390 ;
        RECT 637.660 20.130 637.920 20.390 ;
        RECT 637.660 20.070 639.240 20.130 ;
        RECT 637.720 19.990 639.240 20.070 ;
        RECT 639.100 2.400 639.240 19.990 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1188.250 1594.160 1188.570 1594.220 ;
        RECT 1190.090 1594.160 1190.410 1594.220 ;
        RECT 1188.250 1594.020 1190.410 1594.160 ;
        RECT 1188.250 1593.960 1188.570 1594.020 ;
        RECT 1190.090 1593.960 1190.410 1594.020 ;
        RECT 1188.250 1587.020 1188.570 1587.080 ;
        RECT 1192.850 1587.020 1193.170 1587.080 ;
        RECT 1188.250 1586.880 1193.170 1587.020 ;
        RECT 1188.250 1586.820 1188.570 1586.880 ;
        RECT 1192.850 1586.820 1193.170 1586.880 ;
        RECT 1192.850 73.000 1193.170 73.060 ;
        RECT 2421.970 73.000 2422.290 73.060 ;
        RECT 1192.850 72.860 2422.290 73.000 ;
        RECT 1192.850 72.800 1193.170 72.860 ;
        RECT 2421.970 72.800 2422.290 72.860 ;
      LAYER via ;
        RECT 1188.280 1593.960 1188.540 1594.220 ;
        RECT 1190.120 1593.960 1190.380 1594.220 ;
        RECT 1188.280 1586.820 1188.540 1587.080 ;
        RECT 1192.880 1586.820 1193.140 1587.080 ;
        RECT 1192.880 72.800 1193.140 73.060 ;
        RECT 2422.000 72.800 2422.260 73.060 ;
      LAYER met2 ;
        RECT 1189.980 1600.380 1190.260 1604.000 ;
        RECT 1189.980 1600.000 1190.320 1600.380 ;
        RECT 1190.180 1594.250 1190.320 1600.000 ;
        RECT 1188.280 1593.930 1188.540 1594.250 ;
        RECT 1190.120 1593.930 1190.380 1594.250 ;
        RECT 1188.340 1587.110 1188.480 1593.930 ;
        RECT 1188.280 1586.790 1188.540 1587.110 ;
        RECT 1192.880 1586.790 1193.140 1587.110 ;
        RECT 1192.940 73.090 1193.080 1586.790 ;
        RECT 1192.880 72.770 1193.140 73.090 ;
        RECT 2422.000 72.770 2422.260 73.090 ;
        RECT 2422.060 17.410 2422.200 72.770 ;
        RECT 2422.060 17.270 2423.120 17.410 ;
        RECT 2422.980 2.400 2423.120 17.270 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1194.765 1538.925 1194.935 1587.035 ;
      LAYER mcon ;
        RECT 1194.765 1586.865 1194.935 1587.035 ;
      LAYER met1 ;
        RECT 1194.690 1587.020 1195.010 1587.080 ;
        RECT 1194.495 1586.880 1195.010 1587.020 ;
        RECT 1194.690 1586.820 1195.010 1586.880 ;
        RECT 1194.690 1539.080 1195.010 1539.140 ;
        RECT 1194.495 1538.940 1195.010 1539.080 ;
        RECT 1194.690 1538.880 1195.010 1538.940 ;
        RECT 1194.690 1511.000 1195.010 1511.260 ;
        RECT 1194.780 1510.860 1194.920 1511.000 ;
        RECT 1198.830 1510.860 1199.150 1510.920 ;
        RECT 1194.780 1510.720 1199.150 1510.860 ;
        RECT 1198.830 1510.660 1199.150 1510.720 ;
        RECT 1198.370 72.320 1198.690 72.380 ;
        RECT 2435.770 72.320 2436.090 72.380 ;
        RECT 1198.370 72.180 2436.090 72.320 ;
        RECT 1198.370 72.120 1198.690 72.180 ;
        RECT 2435.770 72.120 2436.090 72.180 ;
      LAYER via ;
        RECT 1194.720 1586.820 1194.980 1587.080 ;
        RECT 1194.720 1538.880 1194.980 1539.140 ;
        RECT 1194.720 1511.000 1194.980 1511.260 ;
        RECT 1198.860 1510.660 1199.120 1510.920 ;
        RECT 1198.400 72.120 1198.660 72.380 ;
        RECT 2435.800 72.120 2436.060 72.380 ;
      LAYER met2 ;
        RECT 1195.960 1600.450 1196.240 1604.000 ;
        RECT 1195.240 1600.310 1196.240 1600.450 ;
        RECT 1195.240 1594.330 1195.380 1600.310 ;
        RECT 1195.960 1600.000 1196.240 1600.310 ;
        RECT 1194.780 1594.190 1195.380 1594.330 ;
        RECT 1194.780 1587.110 1194.920 1594.190 ;
        RECT 1194.720 1586.790 1194.980 1587.110 ;
        RECT 1194.720 1538.850 1194.980 1539.170 ;
        RECT 1194.780 1511.290 1194.920 1538.850 ;
        RECT 1194.720 1510.970 1194.980 1511.290 ;
        RECT 1198.860 1510.630 1199.120 1510.950 ;
        RECT 1198.920 1390.330 1199.060 1510.630 ;
        RECT 1198.460 1390.190 1199.060 1390.330 ;
        RECT 1198.460 72.410 1198.600 1390.190 ;
        RECT 1198.400 72.090 1198.660 72.410 ;
        RECT 2435.800 72.090 2436.060 72.410 ;
        RECT 2435.860 17.410 2436.000 72.090 ;
        RECT 2435.860 17.270 2441.060 17.410 ;
        RECT 2440.920 2.400 2441.060 17.270 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1203.430 1600.960 1203.750 1601.020 ;
        RECT 1206.650 1600.960 1206.970 1601.020 ;
        RECT 1203.430 1600.820 1206.970 1600.960 ;
        RECT 1203.430 1600.760 1203.750 1600.820 ;
        RECT 1206.650 1600.760 1206.970 1600.820 ;
        RECT 1206.650 42.060 1206.970 42.120 ;
        RECT 2458.770 42.060 2459.090 42.120 ;
        RECT 1206.650 41.920 2459.090 42.060 ;
        RECT 1206.650 41.860 1206.970 41.920 ;
        RECT 2458.770 41.860 2459.090 41.920 ;
      LAYER via ;
        RECT 1203.460 1600.760 1203.720 1601.020 ;
        RECT 1206.680 1600.760 1206.940 1601.020 ;
        RECT 1206.680 41.860 1206.940 42.120 ;
        RECT 2458.800 41.860 2459.060 42.120 ;
      LAYER met2 ;
        RECT 1201.940 1601.130 1202.220 1604.000 ;
        RECT 1201.940 1601.050 1203.660 1601.130 ;
        RECT 1201.940 1600.990 1203.720 1601.050 ;
        RECT 1201.940 1600.000 1202.220 1600.990 ;
        RECT 1203.460 1600.730 1203.720 1600.990 ;
        RECT 1206.680 1600.730 1206.940 1601.050 ;
        RECT 1206.740 42.150 1206.880 1600.730 ;
        RECT 1206.680 41.830 1206.940 42.150 ;
        RECT 2458.800 41.830 2459.060 42.150 ;
        RECT 2458.860 2.400 2459.000 41.830 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1245.365 42.245 1245.535 44.115 ;
      LAYER mcon ;
        RECT 1245.365 43.945 1245.535 44.115 ;
      LAYER met1 ;
        RECT 1209.410 1600.960 1209.730 1601.020 ;
        RECT 1213.550 1600.960 1213.870 1601.020 ;
        RECT 1209.410 1600.820 1213.870 1600.960 ;
        RECT 1209.410 1600.760 1209.730 1600.820 ;
        RECT 1213.550 1600.760 1213.870 1600.820 ;
        RECT 1213.550 44.100 1213.870 44.160 ;
        RECT 1245.305 44.100 1245.595 44.145 ;
        RECT 1213.550 43.960 1245.595 44.100 ;
        RECT 1213.550 43.900 1213.870 43.960 ;
        RECT 1245.305 43.915 1245.595 43.960 ;
        RECT 1245.305 42.400 1245.595 42.445 ;
        RECT 2476.710 42.400 2477.030 42.460 ;
        RECT 1245.305 42.260 2477.030 42.400 ;
        RECT 1245.305 42.215 1245.595 42.260 ;
        RECT 2476.710 42.200 2477.030 42.260 ;
      LAYER via ;
        RECT 1209.440 1600.760 1209.700 1601.020 ;
        RECT 1213.580 1600.760 1213.840 1601.020 ;
        RECT 1213.580 43.900 1213.840 44.160 ;
        RECT 2476.740 42.200 2477.000 42.460 ;
      LAYER met2 ;
        RECT 1208.380 1601.130 1208.660 1604.000 ;
        RECT 1208.380 1601.050 1209.640 1601.130 ;
        RECT 1208.380 1600.990 1209.700 1601.050 ;
        RECT 1208.380 1600.000 1208.660 1600.990 ;
        RECT 1209.440 1600.730 1209.700 1600.990 ;
        RECT 1213.580 1600.730 1213.840 1601.050 ;
        RECT 1213.640 44.190 1213.780 1600.730 ;
        RECT 1213.580 43.870 1213.840 44.190 ;
        RECT 2476.740 42.170 2477.000 42.490 ;
        RECT 2476.800 2.400 2476.940 42.170 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1245.825 42.585 1245.995 46.835 ;
      LAYER mcon ;
        RECT 1245.825 46.665 1245.995 46.835 ;
      LAYER met1 ;
        RECT 1219.990 46.820 1220.310 46.880 ;
        RECT 1245.765 46.820 1246.055 46.865 ;
        RECT 1219.990 46.680 1246.055 46.820 ;
        RECT 1219.990 46.620 1220.310 46.680 ;
        RECT 1245.765 46.635 1246.055 46.680 ;
        RECT 1245.765 42.740 1246.055 42.785 ;
        RECT 2494.650 42.740 2494.970 42.800 ;
        RECT 1245.765 42.600 2494.970 42.740 ;
        RECT 1245.765 42.555 1246.055 42.600 ;
        RECT 2494.650 42.540 2494.970 42.600 ;
      LAYER via ;
        RECT 1220.020 46.620 1220.280 46.880 ;
        RECT 2494.680 42.540 2494.940 42.800 ;
      LAYER met2 ;
        RECT 1214.360 1600.450 1214.640 1604.000 ;
        RECT 1214.360 1600.310 1215.160 1600.450 ;
        RECT 1214.360 1600.000 1214.640 1600.310 ;
        RECT 1215.020 1535.340 1215.160 1600.310 ;
        RECT 1215.020 1535.200 1220.220 1535.340 ;
        RECT 1220.080 46.910 1220.220 1535.200 ;
        RECT 1220.020 46.590 1220.280 46.910 ;
        RECT 2494.680 42.510 2494.940 42.830 ;
        RECT 2494.740 2.400 2494.880 42.510 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1220.450 1580.360 1220.770 1580.620 ;
        RECT 1220.540 1579.600 1220.680 1580.360 ;
        RECT 1220.450 1579.340 1220.770 1579.600 ;
        RECT 1246.670 43.080 1246.990 43.140 ;
        RECT 2512.130 43.080 2512.450 43.140 ;
        RECT 1246.670 42.940 2512.450 43.080 ;
        RECT 1246.670 42.880 1246.990 42.940 ;
        RECT 2512.130 42.880 2512.450 42.940 ;
      LAYER via ;
        RECT 1220.480 1580.360 1220.740 1580.620 ;
        RECT 1220.480 1579.340 1220.740 1579.600 ;
        RECT 1246.700 42.880 1246.960 43.140 ;
        RECT 2512.160 42.880 2512.420 43.140 ;
      LAYER met2 ;
        RECT 1220.800 1600.380 1221.080 1604.000 ;
        RECT 1220.800 1600.000 1221.140 1600.380 ;
        RECT 1221.000 1597.220 1221.140 1600.000 ;
        RECT 1220.540 1597.080 1221.140 1597.220 ;
        RECT 1220.540 1580.650 1220.680 1597.080 ;
        RECT 1220.480 1580.330 1220.740 1580.650 ;
        RECT 1220.480 1579.310 1220.740 1579.630 ;
        RECT 1220.540 46.085 1220.680 1579.310 ;
        RECT 1220.470 45.715 1220.750 46.085 ;
        RECT 1246.690 45.715 1246.970 46.085 ;
        RECT 1246.760 43.170 1246.900 45.715 ;
        RECT 1246.700 42.850 1246.960 43.170 ;
        RECT 2512.160 42.850 2512.420 43.170 ;
        RECT 2512.220 2.400 2512.360 42.850 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
      LAYER via2 ;
        RECT 1220.470 45.760 1220.750 46.040 ;
        RECT 1246.690 45.760 1246.970 46.040 ;
      LAYER met3 ;
        RECT 1220.445 46.050 1220.775 46.065 ;
        RECT 1246.665 46.050 1246.995 46.065 ;
        RECT 1220.445 45.750 1246.995 46.050 ;
        RECT 1220.445 45.735 1220.775 45.750 ;
        RECT 1246.665 45.735 1246.995 45.750 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1247.205 43.265 1247.375 47.175 ;
      LAYER mcon ;
        RECT 1247.205 47.005 1247.375 47.175 ;
      LAYER met1 ;
        RECT 1221.370 1600.960 1221.690 1601.020 ;
        RECT 1225.510 1600.960 1225.830 1601.020 ;
        RECT 1221.370 1600.820 1225.830 1600.960 ;
        RECT 1221.370 1600.760 1221.690 1600.820 ;
        RECT 1225.510 1600.760 1225.830 1600.820 ;
        RECT 1221.370 1535.340 1221.690 1535.400 ;
        RECT 1227.350 1535.340 1227.670 1535.400 ;
        RECT 1221.370 1535.200 1227.670 1535.340 ;
        RECT 1221.370 1535.140 1221.690 1535.200 ;
        RECT 1227.350 1535.140 1227.670 1535.200 ;
        RECT 1227.350 47.160 1227.670 47.220 ;
        RECT 1247.145 47.160 1247.435 47.205 ;
        RECT 1227.350 47.020 1247.435 47.160 ;
        RECT 1227.350 46.960 1227.670 47.020 ;
        RECT 1247.145 46.975 1247.435 47.020 ;
        RECT 1247.145 43.420 1247.435 43.465 ;
        RECT 2530.070 43.420 2530.390 43.480 ;
        RECT 1247.145 43.280 2530.390 43.420 ;
        RECT 1247.145 43.235 1247.435 43.280 ;
        RECT 2530.070 43.220 2530.390 43.280 ;
      LAYER via ;
        RECT 1221.400 1600.760 1221.660 1601.020 ;
        RECT 1225.540 1600.760 1225.800 1601.020 ;
        RECT 1221.400 1535.140 1221.660 1535.400 ;
        RECT 1227.380 1535.140 1227.640 1535.400 ;
        RECT 1227.380 46.960 1227.640 47.220 ;
        RECT 2530.100 43.220 2530.360 43.480 ;
      LAYER met2 ;
        RECT 1226.780 1601.130 1227.060 1604.000 ;
        RECT 1225.600 1601.050 1227.060 1601.130 ;
        RECT 1221.400 1600.730 1221.660 1601.050 ;
        RECT 1225.540 1600.990 1227.060 1601.050 ;
        RECT 1225.540 1600.730 1225.800 1600.990 ;
        RECT 1221.460 1535.430 1221.600 1600.730 ;
        RECT 1226.780 1600.000 1227.060 1600.990 ;
        RECT 1221.400 1535.110 1221.660 1535.430 ;
        RECT 1227.380 1535.110 1227.640 1535.430 ;
        RECT 1227.440 47.250 1227.580 1535.110 ;
        RECT 1227.380 46.930 1227.640 47.250 ;
        RECT 2530.100 43.190 2530.360 43.510 ;
        RECT 2530.160 2.400 2530.300 43.190 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1246.745 43.605 1246.915 46.495 ;
      LAYER mcon ;
        RECT 1246.745 46.325 1246.915 46.495 ;
      LAYER met1 ;
        RECT 1228.270 1600.960 1228.590 1601.020 ;
        RECT 1231.950 1600.960 1232.270 1601.020 ;
        RECT 1228.270 1600.820 1232.270 1600.960 ;
        RECT 1228.270 1600.760 1228.590 1600.820 ;
        RECT 1231.950 1600.760 1232.270 1600.820 ;
        RECT 1228.270 1535.340 1228.590 1535.400 ;
        RECT 1234.250 1535.340 1234.570 1535.400 ;
        RECT 1228.270 1535.200 1234.570 1535.340 ;
        RECT 1228.270 1535.140 1228.590 1535.200 ;
        RECT 1234.250 1535.140 1234.570 1535.200 ;
        RECT 1234.250 46.480 1234.570 46.540 ;
        RECT 1246.685 46.480 1246.975 46.525 ;
        RECT 1234.250 46.340 1246.975 46.480 ;
        RECT 1234.250 46.280 1234.570 46.340 ;
        RECT 1246.685 46.295 1246.975 46.340 ;
        RECT 1246.685 43.760 1246.975 43.805 ;
        RECT 2548.010 43.760 2548.330 43.820 ;
        RECT 1246.685 43.620 2548.330 43.760 ;
        RECT 1246.685 43.575 1246.975 43.620 ;
        RECT 2548.010 43.560 2548.330 43.620 ;
      LAYER via ;
        RECT 1228.300 1600.760 1228.560 1601.020 ;
        RECT 1231.980 1600.760 1232.240 1601.020 ;
        RECT 1228.300 1535.140 1228.560 1535.400 ;
        RECT 1234.280 1535.140 1234.540 1535.400 ;
        RECT 1234.280 46.280 1234.540 46.540 ;
        RECT 2548.040 43.560 2548.300 43.820 ;
      LAYER met2 ;
        RECT 1233.220 1601.130 1233.500 1604.000 ;
        RECT 1232.040 1601.050 1233.500 1601.130 ;
        RECT 1228.300 1600.730 1228.560 1601.050 ;
        RECT 1231.980 1600.990 1233.500 1601.050 ;
        RECT 1231.980 1600.730 1232.240 1600.990 ;
        RECT 1228.360 1535.430 1228.500 1600.730 ;
        RECT 1233.220 1600.000 1233.500 1600.990 ;
        RECT 1228.300 1535.110 1228.560 1535.430 ;
        RECT 1234.280 1535.110 1234.540 1535.430 ;
        RECT 1234.340 46.570 1234.480 1535.110 ;
        RECT 1234.280 46.250 1234.540 46.570 ;
        RECT 2548.040 43.530 2548.300 43.850 ;
        RECT 2548.100 2.400 2548.240 43.530 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1241.225 1442.025 1241.395 1490.475 ;
        RECT 1241.225 89.845 1241.395 137.955 ;
      LAYER mcon ;
        RECT 1241.225 1490.305 1241.395 1490.475 ;
        RECT 1241.225 137.785 1241.395 137.955 ;
      LAYER met1 ;
        RECT 1240.690 1587.020 1241.010 1587.080 ;
        RECT 1241.610 1587.020 1241.930 1587.080 ;
        RECT 1240.690 1586.880 1241.930 1587.020 ;
        RECT 1240.690 1586.820 1241.010 1586.880 ;
        RECT 1241.610 1586.820 1241.930 1586.880 ;
        RECT 1241.150 1490.460 1241.470 1490.520 ;
        RECT 1240.955 1490.320 1241.470 1490.460 ;
        RECT 1241.150 1490.260 1241.470 1490.320 ;
        RECT 1241.150 1442.180 1241.470 1442.240 ;
        RECT 1240.955 1442.040 1241.470 1442.180 ;
        RECT 1241.150 1441.980 1241.470 1442.040 ;
        RECT 1241.150 717.640 1241.470 717.700 ;
        RECT 1242.070 717.640 1242.390 717.700 ;
        RECT 1241.150 717.500 1242.390 717.640 ;
        RECT 1241.150 717.440 1241.470 717.500 ;
        RECT 1242.070 717.440 1242.390 717.500 ;
        RECT 1241.150 137.940 1241.470 138.000 ;
        RECT 1240.955 137.800 1241.470 137.940 ;
        RECT 1241.150 137.740 1241.470 137.800 ;
        RECT 1241.150 90.000 1241.470 90.060 ;
        RECT 1240.955 89.860 1241.470 90.000 ;
        RECT 1241.150 89.800 1241.470 89.860 ;
        RECT 1241.150 85.580 1241.470 85.640 ;
        RECT 1242.070 85.580 1242.390 85.640 ;
        RECT 1241.150 85.440 1242.390 85.580 ;
        RECT 1241.150 85.380 1241.470 85.440 ;
        RECT 1242.070 85.380 1242.390 85.440 ;
        RECT 2565.950 44.100 2566.270 44.160 ;
        RECT 1245.840 43.960 2566.270 44.100 ;
        RECT 1242.070 43.760 1242.390 43.820 ;
        RECT 1245.840 43.760 1245.980 43.960 ;
        RECT 2565.950 43.900 2566.270 43.960 ;
        RECT 1242.070 43.620 1245.980 43.760 ;
        RECT 1242.070 43.560 1242.390 43.620 ;
      LAYER via ;
        RECT 1240.720 1586.820 1240.980 1587.080 ;
        RECT 1241.640 1586.820 1241.900 1587.080 ;
        RECT 1241.180 1490.260 1241.440 1490.520 ;
        RECT 1241.180 1441.980 1241.440 1442.240 ;
        RECT 1241.180 717.440 1241.440 717.700 ;
        RECT 1242.100 717.440 1242.360 717.700 ;
        RECT 1241.180 137.740 1241.440 138.000 ;
        RECT 1241.180 89.800 1241.440 90.060 ;
        RECT 1241.180 85.380 1241.440 85.640 ;
        RECT 1242.100 85.380 1242.360 85.640 ;
        RECT 1242.100 43.560 1242.360 43.820 ;
        RECT 2565.980 43.900 2566.240 44.160 ;
      LAYER met2 ;
        RECT 1239.200 1600.450 1239.480 1604.000 ;
        RECT 1239.200 1600.310 1240.920 1600.450 ;
        RECT 1239.200 1600.000 1239.480 1600.310 ;
        RECT 1240.780 1587.110 1240.920 1600.310 ;
        RECT 1240.720 1586.790 1240.980 1587.110 ;
        RECT 1241.640 1586.790 1241.900 1587.110 ;
        RECT 1241.700 1558.290 1241.840 1586.790 ;
        RECT 1241.240 1558.150 1241.840 1558.290 ;
        RECT 1241.240 1490.550 1241.380 1558.150 ;
        RECT 1241.180 1490.230 1241.440 1490.550 ;
        RECT 1241.180 1441.950 1241.440 1442.270 ;
        RECT 1241.240 717.730 1241.380 1441.950 ;
        RECT 1241.180 717.410 1241.440 717.730 ;
        RECT 1242.100 717.410 1242.360 717.730 ;
        RECT 1242.160 669.645 1242.300 717.410 ;
        RECT 1241.170 669.275 1241.450 669.645 ;
        RECT 1242.090 669.275 1242.370 669.645 ;
        RECT 1241.240 138.030 1241.380 669.275 ;
        RECT 1241.180 137.710 1241.440 138.030 ;
        RECT 1241.180 89.770 1241.440 90.090 ;
        RECT 1241.240 85.670 1241.380 89.770 ;
        RECT 1241.180 85.350 1241.440 85.670 ;
        RECT 1242.100 85.350 1242.360 85.670 ;
        RECT 1242.160 43.850 1242.300 85.350 ;
        RECT 2565.980 43.870 2566.240 44.190 ;
        RECT 1242.100 43.530 1242.360 43.850 ;
        RECT 2566.040 2.400 2566.180 43.870 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
      LAYER via2 ;
        RECT 1241.170 669.320 1241.450 669.600 ;
        RECT 1242.090 669.320 1242.370 669.600 ;
      LAYER met3 ;
        RECT 1241.145 669.610 1241.475 669.625 ;
        RECT 1242.065 669.610 1242.395 669.625 ;
        RECT 1241.145 669.310 1242.395 669.610 ;
        RECT 1241.145 669.295 1241.475 669.310 ;
        RECT 1242.065 669.295 1242.395 669.310 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1248.125 1304.325 1248.295 1352.435 ;
        RECT 1248.125 89.845 1248.295 137.955 ;
        RECT 1293.665 44.285 1293.835 46.835 ;
      LAYER mcon ;
        RECT 1248.125 1352.265 1248.295 1352.435 ;
        RECT 1248.125 137.785 1248.295 137.955 ;
        RECT 1293.665 46.665 1293.835 46.835 ;
      LAYER met1 ;
        RECT 1247.130 1449.320 1247.450 1449.380 ;
        RECT 1248.050 1449.320 1248.370 1449.380 ;
        RECT 1247.130 1449.180 1248.370 1449.320 ;
        RECT 1247.130 1449.120 1247.450 1449.180 ;
        RECT 1248.050 1449.120 1248.370 1449.180 ;
        RECT 1248.050 1352.420 1248.370 1352.480 ;
        RECT 1247.855 1352.280 1248.370 1352.420 ;
        RECT 1248.050 1352.220 1248.370 1352.280 ;
        RECT 1248.050 1304.480 1248.370 1304.540 ;
        RECT 1247.855 1304.340 1248.370 1304.480 ;
        RECT 1248.050 1304.280 1248.370 1304.340 ;
        RECT 1247.130 717.640 1247.450 717.700 ;
        RECT 1248.050 717.640 1248.370 717.700 ;
        RECT 1247.130 717.500 1248.370 717.640 ;
        RECT 1247.130 717.440 1247.450 717.500 ;
        RECT 1248.050 717.440 1248.370 717.500 ;
        RECT 1248.050 137.940 1248.370 138.000 ;
        RECT 1247.855 137.800 1248.370 137.940 ;
        RECT 1248.050 137.740 1248.370 137.800 ;
        RECT 1248.050 90.000 1248.370 90.060 ;
        RECT 1247.855 89.860 1248.370 90.000 ;
        RECT 1248.050 89.800 1248.370 89.860 ;
        RECT 1247.590 46.820 1247.910 46.880 ;
        RECT 1293.605 46.820 1293.895 46.865 ;
        RECT 1247.590 46.680 1293.895 46.820 ;
        RECT 1247.590 46.620 1247.910 46.680 ;
        RECT 1293.605 46.635 1293.895 46.680 ;
        RECT 1293.605 44.440 1293.895 44.485 ;
        RECT 2583.890 44.440 2584.210 44.500 ;
        RECT 1293.605 44.300 2584.210 44.440 ;
        RECT 1293.605 44.255 1293.895 44.300 ;
        RECT 2583.890 44.240 2584.210 44.300 ;
      LAYER via ;
        RECT 1247.160 1449.120 1247.420 1449.380 ;
        RECT 1248.080 1449.120 1248.340 1449.380 ;
        RECT 1248.080 1352.220 1248.340 1352.480 ;
        RECT 1248.080 1304.280 1248.340 1304.540 ;
        RECT 1247.160 717.440 1247.420 717.700 ;
        RECT 1248.080 717.440 1248.340 717.700 ;
        RECT 1248.080 137.740 1248.340 138.000 ;
        RECT 1248.080 89.800 1248.340 90.060 ;
        RECT 1247.620 46.620 1247.880 46.880 ;
        RECT 2583.920 44.240 2584.180 44.500 ;
      LAYER met2 ;
        RECT 1245.640 1600.450 1245.920 1604.000 ;
        RECT 1245.640 1600.310 1246.440 1600.450 ;
        RECT 1245.640 1600.000 1245.920 1600.310 ;
        RECT 1246.300 1594.330 1246.440 1600.310 ;
        RECT 1246.300 1594.190 1246.900 1594.330 ;
        RECT 1246.760 1557.610 1246.900 1594.190 ;
        RECT 1246.760 1557.470 1247.360 1557.610 ;
        RECT 1247.220 1449.410 1247.360 1557.470 ;
        RECT 1247.160 1449.090 1247.420 1449.410 ;
        RECT 1248.080 1449.090 1248.340 1449.410 ;
        RECT 1248.140 1352.510 1248.280 1449.090 ;
        RECT 1248.080 1352.190 1248.340 1352.510 ;
        RECT 1248.080 1304.250 1248.340 1304.570 ;
        RECT 1248.140 717.730 1248.280 1304.250 ;
        RECT 1247.160 717.410 1247.420 717.730 ;
        RECT 1248.080 717.410 1248.340 717.730 ;
        RECT 1247.220 669.645 1247.360 717.410 ;
        RECT 1247.150 669.275 1247.430 669.645 ;
        RECT 1248.070 669.275 1248.350 669.645 ;
        RECT 1248.140 138.030 1248.280 669.275 ;
        RECT 1248.080 137.710 1248.340 138.030 ;
        RECT 1248.080 89.770 1248.340 90.090 ;
        RECT 1248.140 67.730 1248.280 89.770 ;
        RECT 1247.220 67.590 1248.280 67.730 ;
        RECT 1247.220 61.610 1247.360 67.590 ;
        RECT 1247.220 61.470 1247.820 61.610 ;
        RECT 1247.680 46.910 1247.820 61.470 ;
        RECT 1247.620 46.590 1247.880 46.910 ;
        RECT 2583.920 44.210 2584.180 44.530 ;
        RECT 2583.980 2.400 2584.120 44.210 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
      LAYER via2 ;
        RECT 1247.150 669.320 1247.430 669.600 ;
        RECT 1248.070 669.320 1248.350 669.600 ;
      LAYER met3 ;
        RECT 1247.125 669.610 1247.455 669.625 ;
        RECT 1248.045 669.610 1248.375 669.625 ;
        RECT 1247.125 669.310 1248.375 669.610 ;
        RECT 1247.125 669.295 1247.455 669.310 ;
        RECT 1248.045 669.295 1248.375 669.310 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 714.065 1591.285 714.235 1593.495 ;
        RECT 737.525 1591.285 737.695 1592.135 ;
        RECT 769.725 14.025 770.355 14.195 ;
        RECT 770.185 13.685 770.355 14.025 ;
        RECT 794.105 13.685 794.275 14.875 ;
      LAYER mcon ;
        RECT 714.065 1593.325 714.235 1593.495 ;
        RECT 737.525 1591.965 737.695 1592.135 ;
        RECT 794.105 14.705 794.275 14.875 ;
      LAYER met1 ;
        RECT 633.030 1593.480 633.350 1593.540 ;
        RECT 714.005 1593.480 714.295 1593.525 ;
        RECT 633.030 1593.340 714.295 1593.480 ;
        RECT 633.030 1593.280 633.350 1593.340 ;
        RECT 714.005 1593.295 714.295 1593.340 ;
        RECT 737.465 1592.120 737.755 1592.165 ;
        RECT 748.490 1592.120 748.810 1592.180 ;
        RECT 737.465 1591.980 748.810 1592.120 ;
        RECT 737.465 1591.935 737.755 1591.980 ;
        RECT 748.490 1591.920 748.810 1591.980 ;
        RECT 714.005 1591.440 714.295 1591.485 ;
        RECT 737.465 1591.440 737.755 1591.485 ;
        RECT 714.005 1591.300 737.755 1591.440 ;
        RECT 714.005 1591.255 714.295 1591.300 ;
        RECT 737.465 1591.255 737.755 1591.300 ;
        RECT 794.045 14.860 794.335 14.905 ;
        RECT 817.490 14.860 817.810 14.920 ;
        RECT 794.045 14.720 817.810 14.860 ;
        RECT 794.045 14.675 794.335 14.720 ;
        RECT 817.490 14.660 817.810 14.720 ;
        RECT 748.490 14.180 748.810 14.240 ;
        RECT 769.665 14.180 769.955 14.225 ;
        RECT 748.490 14.040 769.955 14.180 ;
        RECT 748.490 13.980 748.810 14.040 ;
        RECT 769.665 13.995 769.955 14.040 ;
        RECT 776.180 14.040 782.760 14.180 ;
        RECT 770.125 13.840 770.415 13.885 ;
        RECT 776.180 13.840 776.320 14.040 ;
        RECT 770.125 13.700 776.320 13.840 ;
        RECT 782.620 13.840 782.760 14.040 ;
        RECT 794.045 13.840 794.335 13.885 ;
        RECT 782.620 13.700 794.335 13.840 ;
        RECT 770.125 13.655 770.415 13.700 ;
        RECT 794.045 13.655 794.335 13.700 ;
      LAYER via ;
        RECT 633.060 1593.280 633.320 1593.540 ;
        RECT 748.520 1591.920 748.780 1592.180 ;
        RECT 817.520 14.660 817.780 14.920 ;
        RECT 748.520 13.980 748.780 14.240 ;
      LAYER met2 ;
        RECT 632.920 1600.380 633.200 1604.000 ;
        RECT 632.920 1600.000 633.260 1600.380 ;
        RECT 633.120 1593.570 633.260 1600.000 ;
        RECT 633.060 1593.250 633.320 1593.570 ;
        RECT 748.520 1591.890 748.780 1592.210 ;
        RECT 748.580 14.270 748.720 1591.890 ;
        RECT 817.520 14.630 817.780 14.950 ;
        RECT 748.520 13.950 748.780 14.270 ;
        RECT 817.580 2.400 817.720 14.630 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1255.025 1304.325 1255.195 1352.435 ;
        RECT 1255.025 186.405 1255.195 234.515 ;
      LAYER mcon ;
        RECT 1255.025 1352.265 1255.195 1352.435 ;
        RECT 1255.025 234.345 1255.195 234.515 ;
      LAYER met1 ;
        RECT 1252.650 1569.680 1252.970 1569.740 ;
        RECT 1254.950 1569.680 1255.270 1569.740 ;
        RECT 1252.650 1569.540 1255.270 1569.680 ;
        RECT 1252.650 1569.480 1252.970 1569.540 ;
        RECT 1254.950 1569.480 1255.270 1569.540 ;
        RECT 1254.030 1497.600 1254.350 1497.660 ;
        RECT 1254.950 1497.600 1255.270 1497.660 ;
        RECT 1254.030 1497.460 1255.270 1497.600 ;
        RECT 1254.030 1497.400 1254.350 1497.460 ;
        RECT 1254.950 1497.400 1255.270 1497.460 ;
        RECT 1254.030 1449.320 1254.350 1449.380 ;
        RECT 1254.950 1449.320 1255.270 1449.380 ;
        RECT 1254.030 1449.180 1255.270 1449.320 ;
        RECT 1254.030 1449.120 1254.350 1449.180 ;
        RECT 1254.950 1449.120 1255.270 1449.180 ;
        RECT 1254.950 1352.420 1255.270 1352.480 ;
        RECT 1254.755 1352.280 1255.270 1352.420 ;
        RECT 1254.950 1352.220 1255.270 1352.280 ;
        RECT 1254.950 1304.480 1255.270 1304.540 ;
        RECT 1254.755 1304.340 1255.270 1304.480 ;
        RECT 1254.950 1304.280 1255.270 1304.340 ;
        RECT 1254.030 1152.500 1254.350 1152.560 ;
        RECT 1254.950 1152.500 1255.270 1152.560 ;
        RECT 1254.030 1152.360 1255.270 1152.500 ;
        RECT 1254.030 1152.300 1254.350 1152.360 ;
        RECT 1254.950 1152.300 1255.270 1152.360 ;
        RECT 1254.030 910.760 1254.350 910.820 ;
        RECT 1254.950 910.760 1255.270 910.820 ;
        RECT 1254.030 910.620 1255.270 910.760 ;
        RECT 1254.030 910.560 1254.350 910.620 ;
        RECT 1254.950 910.560 1255.270 910.620 ;
        RECT 1254.030 814.200 1254.350 814.260 ;
        RECT 1254.950 814.200 1255.270 814.260 ;
        RECT 1254.030 814.060 1255.270 814.200 ;
        RECT 1254.030 814.000 1254.350 814.060 ;
        RECT 1254.950 814.000 1255.270 814.060 ;
        RECT 1254.950 717.640 1255.270 717.700 ;
        RECT 1255.870 717.640 1256.190 717.700 ;
        RECT 1254.950 717.500 1256.190 717.640 ;
        RECT 1254.950 717.440 1255.270 717.500 ;
        RECT 1255.870 717.440 1256.190 717.500 ;
        RECT 1254.950 234.500 1255.270 234.560 ;
        RECT 1254.755 234.360 1255.270 234.500 ;
        RECT 1254.950 234.300 1255.270 234.360 ;
        RECT 1254.950 186.560 1255.270 186.620 ;
        RECT 1254.755 186.420 1255.270 186.560 ;
        RECT 1254.950 186.360 1255.270 186.420 ;
        RECT 1254.030 99.520 1254.350 99.580 ;
        RECT 1254.950 99.520 1255.270 99.580 ;
        RECT 1254.030 99.380 1255.270 99.520 ;
        RECT 1254.030 99.320 1254.350 99.380 ;
        RECT 1254.950 99.320 1255.270 99.380 ;
        RECT 1254.490 48.180 1254.810 48.240 ;
        RECT 2601.830 48.180 2602.150 48.240 ;
        RECT 1254.490 48.040 2602.150 48.180 ;
        RECT 1254.490 47.980 1254.810 48.040 ;
        RECT 2601.830 47.980 2602.150 48.040 ;
      LAYER via ;
        RECT 1252.680 1569.480 1252.940 1569.740 ;
        RECT 1254.980 1569.480 1255.240 1569.740 ;
        RECT 1254.060 1497.400 1254.320 1497.660 ;
        RECT 1254.980 1497.400 1255.240 1497.660 ;
        RECT 1254.060 1449.120 1254.320 1449.380 ;
        RECT 1254.980 1449.120 1255.240 1449.380 ;
        RECT 1254.980 1352.220 1255.240 1352.480 ;
        RECT 1254.980 1304.280 1255.240 1304.540 ;
        RECT 1254.060 1152.300 1254.320 1152.560 ;
        RECT 1254.980 1152.300 1255.240 1152.560 ;
        RECT 1254.060 910.560 1254.320 910.820 ;
        RECT 1254.980 910.560 1255.240 910.820 ;
        RECT 1254.060 814.000 1254.320 814.260 ;
        RECT 1254.980 814.000 1255.240 814.260 ;
        RECT 1254.980 717.440 1255.240 717.700 ;
        RECT 1255.900 717.440 1256.160 717.700 ;
        RECT 1254.980 234.300 1255.240 234.560 ;
        RECT 1254.980 186.360 1255.240 186.620 ;
        RECT 1254.060 99.320 1254.320 99.580 ;
        RECT 1254.980 99.320 1255.240 99.580 ;
        RECT 1254.520 47.980 1254.780 48.240 ;
        RECT 2601.860 47.980 2602.120 48.240 ;
      LAYER met2 ;
        RECT 1251.620 1600.450 1251.900 1604.000 ;
        RECT 1251.620 1600.310 1252.880 1600.450 ;
        RECT 1251.620 1600.000 1251.900 1600.310 ;
        RECT 1252.740 1569.770 1252.880 1600.310 ;
        RECT 1252.680 1569.450 1252.940 1569.770 ;
        RECT 1254.980 1569.450 1255.240 1569.770 ;
        RECT 1255.040 1497.690 1255.180 1569.450 ;
        RECT 1254.060 1497.370 1254.320 1497.690 ;
        RECT 1254.980 1497.370 1255.240 1497.690 ;
        RECT 1254.120 1449.410 1254.260 1497.370 ;
        RECT 1254.060 1449.090 1254.320 1449.410 ;
        RECT 1254.980 1449.090 1255.240 1449.410 ;
        RECT 1255.040 1352.510 1255.180 1449.090 ;
        RECT 1254.980 1352.190 1255.240 1352.510 ;
        RECT 1254.980 1304.250 1255.240 1304.570 ;
        RECT 1255.040 1200.725 1255.180 1304.250 ;
        RECT 1254.050 1200.355 1254.330 1200.725 ;
        RECT 1254.970 1200.355 1255.250 1200.725 ;
        RECT 1254.120 1152.590 1254.260 1200.355 ;
        RECT 1254.060 1152.270 1254.320 1152.590 ;
        RECT 1254.980 1152.270 1255.240 1152.590 ;
        RECT 1255.040 1104.165 1255.180 1152.270 ;
        RECT 1254.050 1103.795 1254.330 1104.165 ;
        RECT 1254.970 1103.795 1255.250 1104.165 ;
        RECT 1254.120 1055.885 1254.260 1103.795 ;
        RECT 1254.050 1055.515 1254.330 1055.885 ;
        RECT 1254.970 1055.515 1255.250 1055.885 ;
        RECT 1255.040 910.850 1255.180 1055.515 ;
        RECT 1254.060 910.530 1254.320 910.850 ;
        RECT 1254.980 910.530 1255.240 910.850 ;
        RECT 1254.120 862.765 1254.260 910.530 ;
        RECT 1254.050 862.395 1254.330 862.765 ;
        RECT 1254.970 862.395 1255.250 862.765 ;
        RECT 1255.040 814.290 1255.180 862.395 ;
        RECT 1254.060 813.970 1254.320 814.290 ;
        RECT 1254.980 813.970 1255.240 814.290 ;
        RECT 1254.120 766.205 1254.260 813.970 ;
        RECT 1254.050 765.835 1254.330 766.205 ;
        RECT 1254.970 765.835 1255.250 766.205 ;
        RECT 1255.040 717.730 1255.180 765.835 ;
        RECT 1254.980 717.410 1255.240 717.730 ;
        RECT 1255.900 717.410 1256.160 717.730 ;
        RECT 1255.960 669.645 1256.100 717.410 ;
        RECT 1254.970 669.275 1255.250 669.645 ;
        RECT 1255.890 669.275 1256.170 669.645 ;
        RECT 1255.040 234.590 1255.180 669.275 ;
        RECT 1254.980 234.270 1255.240 234.590 ;
        RECT 1254.980 186.330 1255.240 186.650 ;
        RECT 1255.040 99.610 1255.180 186.330 ;
        RECT 1254.060 99.290 1254.320 99.610 ;
        RECT 1254.980 99.290 1255.240 99.610 ;
        RECT 1254.120 61.610 1254.260 99.290 ;
        RECT 1254.120 61.470 1254.720 61.610 ;
        RECT 1254.580 48.270 1254.720 61.470 ;
        RECT 1254.520 47.950 1254.780 48.270 ;
        RECT 2601.860 47.950 2602.120 48.270 ;
        RECT 2601.920 7.210 2602.060 47.950 ;
        RECT 2601.460 7.070 2602.060 7.210 ;
        RECT 2601.460 2.400 2601.600 7.070 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
      LAYER via2 ;
        RECT 1254.050 1200.400 1254.330 1200.680 ;
        RECT 1254.970 1200.400 1255.250 1200.680 ;
        RECT 1254.050 1103.840 1254.330 1104.120 ;
        RECT 1254.970 1103.840 1255.250 1104.120 ;
        RECT 1254.050 1055.560 1254.330 1055.840 ;
        RECT 1254.970 1055.560 1255.250 1055.840 ;
        RECT 1254.050 862.440 1254.330 862.720 ;
        RECT 1254.970 862.440 1255.250 862.720 ;
        RECT 1254.050 765.880 1254.330 766.160 ;
        RECT 1254.970 765.880 1255.250 766.160 ;
        RECT 1254.970 669.320 1255.250 669.600 ;
        RECT 1255.890 669.320 1256.170 669.600 ;
      LAYER met3 ;
        RECT 1254.025 1200.690 1254.355 1200.705 ;
        RECT 1254.945 1200.690 1255.275 1200.705 ;
        RECT 1254.025 1200.390 1255.275 1200.690 ;
        RECT 1254.025 1200.375 1254.355 1200.390 ;
        RECT 1254.945 1200.375 1255.275 1200.390 ;
        RECT 1254.025 1104.130 1254.355 1104.145 ;
        RECT 1254.945 1104.130 1255.275 1104.145 ;
        RECT 1254.025 1103.830 1255.275 1104.130 ;
        RECT 1254.025 1103.815 1254.355 1103.830 ;
        RECT 1254.945 1103.815 1255.275 1103.830 ;
        RECT 1254.025 1055.850 1254.355 1055.865 ;
        RECT 1254.945 1055.850 1255.275 1055.865 ;
        RECT 1254.025 1055.550 1255.275 1055.850 ;
        RECT 1254.025 1055.535 1254.355 1055.550 ;
        RECT 1254.945 1055.535 1255.275 1055.550 ;
        RECT 1254.025 862.730 1254.355 862.745 ;
        RECT 1254.945 862.730 1255.275 862.745 ;
        RECT 1254.025 862.430 1255.275 862.730 ;
        RECT 1254.025 862.415 1254.355 862.430 ;
        RECT 1254.945 862.415 1255.275 862.430 ;
        RECT 1254.025 766.170 1254.355 766.185 ;
        RECT 1254.945 766.170 1255.275 766.185 ;
        RECT 1254.025 765.870 1255.275 766.170 ;
        RECT 1254.025 765.855 1254.355 765.870 ;
        RECT 1254.945 765.855 1255.275 765.870 ;
        RECT 1254.945 669.610 1255.275 669.625 ;
        RECT 1255.865 669.610 1256.195 669.625 ;
        RECT 1254.945 669.310 1256.195 669.610 ;
        RECT 1254.945 669.295 1255.275 669.310 ;
        RECT 1255.865 669.295 1256.195 669.310 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1261.465 1304.325 1261.635 1352.435 ;
        RECT 1261.465 1207.425 1261.635 1255.875 ;
        RECT 1261.465 959.225 1261.635 1007.335 ;
        RECT 1261.465 572.645 1261.635 620.755 ;
        RECT 1260.545 476.085 1260.715 524.195 ;
        RECT 1261.465 379.525 1261.635 427.635 ;
        RECT 1261.465 282.965 1261.635 331.075 ;
        RECT 1261.465 186.405 1261.635 234.515 ;
      LAYER mcon ;
        RECT 1261.465 1352.265 1261.635 1352.435 ;
        RECT 1261.465 1255.705 1261.635 1255.875 ;
        RECT 1261.465 1007.165 1261.635 1007.335 ;
        RECT 1261.465 620.585 1261.635 620.755 ;
        RECT 1260.545 524.025 1260.715 524.195 ;
        RECT 1261.465 427.465 1261.635 427.635 ;
        RECT 1261.465 330.905 1261.635 331.075 ;
        RECT 1261.465 234.345 1261.635 234.515 ;
      LAYER met1 ;
        RECT 1257.250 1597.220 1257.570 1597.280 ;
        RECT 1258.170 1597.220 1258.490 1597.280 ;
        RECT 1257.250 1597.080 1258.490 1597.220 ;
        RECT 1257.250 1597.020 1257.570 1597.080 ;
        RECT 1258.170 1597.020 1258.490 1597.080 ;
        RECT 1256.330 1545.880 1256.650 1545.940 ;
        RECT 1257.250 1545.880 1257.570 1545.940 ;
        RECT 1256.330 1545.740 1257.570 1545.880 ;
        RECT 1256.330 1545.680 1256.650 1545.740 ;
        RECT 1257.250 1545.680 1257.570 1545.740 ;
        RECT 1261.390 1352.420 1261.710 1352.480 ;
        RECT 1261.195 1352.280 1261.710 1352.420 ;
        RECT 1261.390 1352.220 1261.710 1352.280 ;
        RECT 1261.390 1304.480 1261.710 1304.540 ;
        RECT 1261.195 1304.340 1261.710 1304.480 ;
        RECT 1261.390 1304.280 1261.710 1304.340 ;
        RECT 1261.390 1255.860 1261.710 1255.920 ;
        RECT 1261.195 1255.720 1261.710 1255.860 ;
        RECT 1261.390 1255.660 1261.710 1255.720 ;
        RECT 1261.390 1207.580 1261.710 1207.640 ;
        RECT 1261.195 1207.440 1261.710 1207.580 ;
        RECT 1261.390 1207.380 1261.710 1207.440 ;
        RECT 1260.470 1152.500 1260.790 1152.560 ;
        RECT 1261.390 1152.500 1261.710 1152.560 ;
        RECT 1260.470 1152.360 1261.710 1152.500 ;
        RECT 1260.470 1152.300 1260.790 1152.360 ;
        RECT 1261.390 1152.300 1261.710 1152.360 ;
        RECT 1261.390 1007.320 1261.710 1007.380 ;
        RECT 1261.195 1007.180 1261.710 1007.320 ;
        RECT 1261.390 1007.120 1261.710 1007.180 ;
        RECT 1261.390 959.380 1261.710 959.440 ;
        RECT 1261.195 959.240 1261.710 959.380 ;
        RECT 1261.390 959.180 1261.710 959.240 ;
        RECT 1260.470 910.760 1260.790 910.820 ;
        RECT 1261.390 910.760 1261.710 910.820 ;
        RECT 1260.470 910.620 1261.710 910.760 ;
        RECT 1260.470 910.560 1260.790 910.620 ;
        RECT 1261.390 910.560 1261.710 910.620 ;
        RECT 1260.470 814.200 1260.790 814.260 ;
        RECT 1261.390 814.200 1261.710 814.260 ;
        RECT 1260.470 814.060 1261.710 814.200 ;
        RECT 1260.470 814.000 1260.790 814.060 ;
        RECT 1261.390 814.000 1261.710 814.060 ;
        RECT 1260.470 717.640 1260.790 717.700 ;
        RECT 1261.390 717.640 1261.710 717.700 ;
        RECT 1260.470 717.500 1261.710 717.640 ;
        RECT 1260.470 717.440 1260.790 717.500 ;
        RECT 1261.390 717.440 1261.710 717.500 ;
        RECT 1261.390 620.740 1261.710 620.800 ;
        RECT 1261.195 620.600 1261.710 620.740 ;
        RECT 1261.390 620.540 1261.710 620.600 ;
        RECT 1261.390 572.800 1261.710 572.860 ;
        RECT 1261.195 572.660 1261.710 572.800 ;
        RECT 1261.390 572.600 1261.710 572.660 ;
        RECT 1260.485 524.180 1260.775 524.225 ;
        RECT 1261.390 524.180 1261.710 524.240 ;
        RECT 1260.485 524.040 1261.710 524.180 ;
        RECT 1260.485 523.995 1260.775 524.040 ;
        RECT 1261.390 523.980 1261.710 524.040 ;
        RECT 1260.470 476.240 1260.790 476.300 ;
        RECT 1260.275 476.100 1260.790 476.240 ;
        RECT 1260.470 476.040 1260.790 476.100 ;
        RECT 1261.390 427.620 1261.710 427.680 ;
        RECT 1261.195 427.480 1261.710 427.620 ;
        RECT 1261.390 427.420 1261.710 427.480 ;
        RECT 1261.390 379.680 1261.710 379.740 ;
        RECT 1261.195 379.540 1261.710 379.680 ;
        RECT 1261.390 379.480 1261.710 379.540 ;
        RECT 1261.390 331.060 1261.710 331.120 ;
        RECT 1261.195 330.920 1261.710 331.060 ;
        RECT 1261.390 330.860 1261.710 330.920 ;
        RECT 1261.390 283.120 1261.710 283.180 ;
        RECT 1261.195 282.980 1261.710 283.120 ;
        RECT 1261.390 282.920 1261.710 282.980 ;
        RECT 1261.390 234.500 1261.710 234.560 ;
        RECT 1261.195 234.360 1261.710 234.500 ;
        RECT 1261.390 234.300 1261.710 234.360 ;
        RECT 1261.390 186.560 1261.710 186.620 ;
        RECT 1261.195 186.420 1261.710 186.560 ;
        RECT 1261.390 186.360 1261.710 186.420 ;
        RECT 1260.930 47.840 1261.250 47.900 ;
        RECT 2619.310 47.840 2619.630 47.900 ;
        RECT 1260.930 47.700 2619.630 47.840 ;
        RECT 1260.930 47.640 1261.250 47.700 ;
        RECT 2619.310 47.640 2619.630 47.700 ;
      LAYER via ;
        RECT 1257.280 1597.020 1257.540 1597.280 ;
        RECT 1258.200 1597.020 1258.460 1597.280 ;
        RECT 1256.360 1545.680 1256.620 1545.940 ;
        RECT 1257.280 1545.680 1257.540 1545.940 ;
        RECT 1261.420 1352.220 1261.680 1352.480 ;
        RECT 1261.420 1304.280 1261.680 1304.540 ;
        RECT 1261.420 1255.660 1261.680 1255.920 ;
        RECT 1261.420 1207.380 1261.680 1207.640 ;
        RECT 1260.500 1152.300 1260.760 1152.560 ;
        RECT 1261.420 1152.300 1261.680 1152.560 ;
        RECT 1261.420 1007.120 1261.680 1007.380 ;
        RECT 1261.420 959.180 1261.680 959.440 ;
        RECT 1260.500 910.560 1260.760 910.820 ;
        RECT 1261.420 910.560 1261.680 910.820 ;
        RECT 1260.500 814.000 1260.760 814.260 ;
        RECT 1261.420 814.000 1261.680 814.260 ;
        RECT 1260.500 717.440 1260.760 717.700 ;
        RECT 1261.420 717.440 1261.680 717.700 ;
        RECT 1261.420 620.540 1261.680 620.800 ;
        RECT 1261.420 572.600 1261.680 572.860 ;
        RECT 1261.420 523.980 1261.680 524.240 ;
        RECT 1260.500 476.040 1260.760 476.300 ;
        RECT 1261.420 427.420 1261.680 427.680 ;
        RECT 1261.420 379.480 1261.680 379.740 ;
        RECT 1261.420 330.860 1261.680 331.120 ;
        RECT 1261.420 282.920 1261.680 283.180 ;
        RECT 1261.420 234.300 1261.680 234.560 ;
        RECT 1261.420 186.360 1261.680 186.620 ;
        RECT 1260.960 47.640 1261.220 47.900 ;
        RECT 2619.340 47.640 2619.600 47.900 ;
      LAYER met2 ;
        RECT 1257.600 1600.450 1257.880 1604.000 ;
        RECT 1257.600 1600.310 1258.400 1600.450 ;
        RECT 1257.600 1600.000 1257.880 1600.310 ;
        RECT 1258.260 1597.310 1258.400 1600.310 ;
        RECT 1257.280 1596.990 1257.540 1597.310 ;
        RECT 1258.200 1596.990 1258.460 1597.310 ;
        RECT 1257.340 1545.970 1257.480 1596.990 ;
        RECT 1256.360 1545.650 1256.620 1545.970 ;
        RECT 1257.280 1545.650 1257.540 1545.970 ;
        RECT 1256.420 1535.170 1256.560 1545.650 ;
        RECT 1256.420 1535.030 1257.020 1535.170 ;
        RECT 1256.880 1486.890 1257.020 1535.030 ;
        RECT 1256.880 1486.750 1261.620 1486.890 ;
        RECT 1261.480 1352.510 1261.620 1486.750 ;
        RECT 1261.420 1352.190 1261.680 1352.510 ;
        RECT 1261.420 1304.250 1261.680 1304.570 ;
        RECT 1261.480 1255.950 1261.620 1304.250 ;
        RECT 1261.420 1255.630 1261.680 1255.950 ;
        RECT 1261.420 1207.350 1261.680 1207.670 ;
        RECT 1261.480 1200.725 1261.620 1207.350 ;
        RECT 1260.490 1200.355 1260.770 1200.725 ;
        RECT 1261.410 1200.355 1261.690 1200.725 ;
        RECT 1260.560 1152.590 1260.700 1200.355 ;
        RECT 1260.500 1152.270 1260.760 1152.590 ;
        RECT 1261.420 1152.270 1261.680 1152.590 ;
        RECT 1261.480 1104.165 1261.620 1152.270 ;
        RECT 1260.490 1103.795 1260.770 1104.165 ;
        RECT 1261.410 1103.795 1261.690 1104.165 ;
        RECT 1260.560 1055.885 1260.700 1103.795 ;
        RECT 1260.490 1055.515 1260.770 1055.885 ;
        RECT 1261.410 1055.515 1261.690 1055.885 ;
        RECT 1261.480 1007.410 1261.620 1055.515 ;
        RECT 1261.420 1007.090 1261.680 1007.410 ;
        RECT 1261.420 959.150 1261.680 959.470 ;
        RECT 1261.480 910.850 1261.620 959.150 ;
        RECT 1260.500 910.530 1260.760 910.850 ;
        RECT 1261.420 910.530 1261.680 910.850 ;
        RECT 1260.560 862.765 1260.700 910.530 ;
        RECT 1260.490 862.395 1260.770 862.765 ;
        RECT 1261.410 862.395 1261.690 862.765 ;
        RECT 1261.480 814.290 1261.620 862.395 ;
        RECT 1260.500 813.970 1260.760 814.290 ;
        RECT 1261.420 813.970 1261.680 814.290 ;
        RECT 1260.560 766.205 1260.700 813.970 ;
        RECT 1260.490 765.835 1260.770 766.205 ;
        RECT 1261.410 765.835 1261.690 766.205 ;
        RECT 1261.480 717.730 1261.620 765.835 ;
        RECT 1260.500 717.410 1260.760 717.730 ;
        RECT 1261.420 717.410 1261.680 717.730 ;
        RECT 1260.560 669.645 1260.700 717.410 ;
        RECT 1260.490 669.275 1260.770 669.645 ;
        RECT 1261.410 669.275 1261.690 669.645 ;
        RECT 1261.480 620.830 1261.620 669.275 ;
        RECT 1261.420 620.510 1261.680 620.830 ;
        RECT 1261.420 572.570 1261.680 572.890 ;
        RECT 1261.480 524.270 1261.620 572.570 ;
        RECT 1261.420 523.950 1261.680 524.270 ;
        RECT 1260.500 476.010 1260.760 476.330 ;
        RECT 1260.560 435.045 1260.700 476.010 ;
        RECT 1260.490 434.675 1260.770 435.045 ;
        RECT 1261.410 434.675 1261.690 435.045 ;
        RECT 1261.480 427.710 1261.620 434.675 ;
        RECT 1261.420 427.390 1261.680 427.710 ;
        RECT 1261.420 379.450 1261.680 379.770 ;
        RECT 1261.480 331.150 1261.620 379.450 ;
        RECT 1261.420 330.830 1261.680 331.150 ;
        RECT 1261.420 282.890 1261.680 283.210 ;
        RECT 1261.480 234.590 1261.620 282.890 ;
        RECT 1261.420 234.270 1261.680 234.590 ;
        RECT 1261.420 186.330 1261.680 186.650 ;
        RECT 1261.480 62.290 1261.620 186.330 ;
        RECT 1260.560 62.150 1261.620 62.290 ;
        RECT 1260.560 61.610 1260.700 62.150 ;
        RECT 1260.560 61.470 1261.160 61.610 ;
        RECT 1261.020 47.930 1261.160 61.470 ;
        RECT 1260.960 47.610 1261.220 47.930 ;
        RECT 2619.340 47.610 2619.600 47.930 ;
        RECT 2619.400 2.400 2619.540 47.610 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
      LAYER via2 ;
        RECT 1260.490 1200.400 1260.770 1200.680 ;
        RECT 1261.410 1200.400 1261.690 1200.680 ;
        RECT 1260.490 1103.840 1260.770 1104.120 ;
        RECT 1261.410 1103.840 1261.690 1104.120 ;
        RECT 1260.490 1055.560 1260.770 1055.840 ;
        RECT 1261.410 1055.560 1261.690 1055.840 ;
        RECT 1260.490 862.440 1260.770 862.720 ;
        RECT 1261.410 862.440 1261.690 862.720 ;
        RECT 1260.490 765.880 1260.770 766.160 ;
        RECT 1261.410 765.880 1261.690 766.160 ;
        RECT 1260.490 669.320 1260.770 669.600 ;
        RECT 1261.410 669.320 1261.690 669.600 ;
        RECT 1260.490 434.720 1260.770 435.000 ;
        RECT 1261.410 434.720 1261.690 435.000 ;
      LAYER met3 ;
        RECT 1260.465 1200.690 1260.795 1200.705 ;
        RECT 1261.385 1200.690 1261.715 1200.705 ;
        RECT 1260.465 1200.390 1261.715 1200.690 ;
        RECT 1260.465 1200.375 1260.795 1200.390 ;
        RECT 1261.385 1200.375 1261.715 1200.390 ;
        RECT 1260.465 1104.130 1260.795 1104.145 ;
        RECT 1261.385 1104.130 1261.715 1104.145 ;
        RECT 1260.465 1103.830 1261.715 1104.130 ;
        RECT 1260.465 1103.815 1260.795 1103.830 ;
        RECT 1261.385 1103.815 1261.715 1103.830 ;
        RECT 1260.465 1055.850 1260.795 1055.865 ;
        RECT 1261.385 1055.850 1261.715 1055.865 ;
        RECT 1260.465 1055.550 1261.715 1055.850 ;
        RECT 1260.465 1055.535 1260.795 1055.550 ;
        RECT 1261.385 1055.535 1261.715 1055.550 ;
        RECT 1260.465 862.730 1260.795 862.745 ;
        RECT 1261.385 862.730 1261.715 862.745 ;
        RECT 1260.465 862.430 1261.715 862.730 ;
        RECT 1260.465 862.415 1260.795 862.430 ;
        RECT 1261.385 862.415 1261.715 862.430 ;
        RECT 1260.465 766.170 1260.795 766.185 ;
        RECT 1261.385 766.170 1261.715 766.185 ;
        RECT 1260.465 765.870 1261.715 766.170 ;
        RECT 1260.465 765.855 1260.795 765.870 ;
        RECT 1261.385 765.855 1261.715 765.870 ;
        RECT 1260.465 669.610 1260.795 669.625 ;
        RECT 1261.385 669.610 1261.715 669.625 ;
        RECT 1260.465 669.310 1261.715 669.610 ;
        RECT 1260.465 669.295 1260.795 669.310 ;
        RECT 1261.385 669.295 1261.715 669.310 ;
        RECT 1260.465 435.010 1260.795 435.025 ;
        RECT 1261.385 435.010 1261.715 435.025 ;
        RECT 1260.465 434.710 1261.715 435.010 ;
        RECT 1260.465 434.695 1260.795 434.710 ;
        RECT 1261.385 434.695 1261.715 434.710 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1265.070 1600.960 1265.390 1601.020 ;
        RECT 1268.750 1600.960 1269.070 1601.020 ;
        RECT 1265.070 1600.820 1269.070 1600.960 ;
        RECT 1265.070 1600.760 1265.390 1600.820 ;
        RECT 1268.750 1600.760 1269.070 1600.820 ;
        RECT 1268.750 47.500 1269.070 47.560 ;
        RECT 2637.250 47.500 2637.570 47.560 ;
        RECT 1268.750 47.360 2637.570 47.500 ;
        RECT 1268.750 47.300 1269.070 47.360 ;
        RECT 2637.250 47.300 2637.570 47.360 ;
      LAYER via ;
        RECT 1265.100 1600.760 1265.360 1601.020 ;
        RECT 1268.780 1600.760 1269.040 1601.020 ;
        RECT 1268.780 47.300 1269.040 47.560 ;
        RECT 2637.280 47.300 2637.540 47.560 ;
      LAYER met2 ;
        RECT 1264.040 1601.130 1264.320 1604.000 ;
        RECT 1264.040 1601.050 1265.300 1601.130 ;
        RECT 1264.040 1600.990 1265.360 1601.050 ;
        RECT 1264.040 1600.000 1264.320 1600.990 ;
        RECT 1265.100 1600.730 1265.360 1600.990 ;
        RECT 1268.780 1600.730 1269.040 1601.050 ;
        RECT 1268.840 47.590 1268.980 1600.730 ;
        RECT 1268.780 47.270 1269.040 47.590 ;
        RECT 2637.280 47.270 2637.540 47.590 ;
        RECT 2637.340 2.400 2637.480 47.270 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1275.725 55.165 1275.895 65.535 ;
        RECT 1295.045 45.645 1295.215 47.175 ;
      LAYER mcon ;
        RECT 1275.725 65.365 1275.895 65.535 ;
        RECT 1295.045 47.005 1295.215 47.175 ;
      LAYER met1 ;
        RECT 1269.670 1535.340 1269.990 1535.400 ;
        RECT 1275.650 1535.340 1275.970 1535.400 ;
        RECT 1269.670 1535.200 1275.970 1535.340 ;
        RECT 1269.670 1535.140 1269.990 1535.200 ;
        RECT 1275.650 1535.140 1275.970 1535.200 ;
        RECT 1275.650 65.520 1275.970 65.580 ;
        RECT 1275.455 65.380 1275.970 65.520 ;
        RECT 1275.650 65.320 1275.970 65.380 ;
        RECT 1275.650 55.320 1275.970 55.380 ;
        RECT 1275.455 55.180 1275.970 55.320 ;
        RECT 1275.650 55.120 1275.970 55.180 ;
        RECT 1294.985 47.160 1295.275 47.205 ;
        RECT 2655.190 47.160 2655.510 47.220 ;
        RECT 1294.985 47.020 2655.510 47.160 ;
        RECT 1294.985 46.975 1295.275 47.020 ;
        RECT 2655.190 46.960 2655.510 47.020 ;
        RECT 1275.650 45.800 1275.970 45.860 ;
        RECT 1294.985 45.800 1295.275 45.845 ;
        RECT 1275.650 45.660 1295.275 45.800 ;
        RECT 1275.650 45.600 1275.970 45.660 ;
        RECT 1294.985 45.615 1295.275 45.660 ;
      LAYER via ;
        RECT 1269.700 1535.140 1269.960 1535.400 ;
        RECT 1275.680 1535.140 1275.940 1535.400 ;
        RECT 1275.680 65.320 1275.940 65.580 ;
        RECT 1275.680 55.120 1275.940 55.380 ;
        RECT 2655.220 46.960 2655.480 47.220 ;
        RECT 1275.680 45.600 1275.940 45.860 ;
      LAYER met2 ;
        RECT 1270.020 1601.130 1270.300 1604.000 ;
        RECT 1269.300 1600.990 1270.300 1601.130 ;
        RECT 1269.300 1597.050 1269.440 1600.990 ;
        RECT 1270.020 1600.000 1270.300 1600.990 ;
        RECT 1269.300 1596.910 1269.900 1597.050 ;
        RECT 1269.760 1535.430 1269.900 1596.910 ;
        RECT 1269.700 1535.110 1269.960 1535.430 ;
        RECT 1275.680 1535.110 1275.940 1535.430 ;
        RECT 1275.740 65.610 1275.880 1535.110 ;
        RECT 1275.680 65.290 1275.940 65.610 ;
        RECT 1275.680 55.090 1275.940 55.410 ;
        RECT 1275.740 45.890 1275.880 55.090 ;
        RECT 2655.220 46.930 2655.480 47.250 ;
        RECT 1275.680 45.570 1275.940 45.890 ;
        RECT 2655.280 2.400 2655.420 46.930 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1277.030 1535.340 1277.350 1535.400 ;
        RECT 1282.090 1535.340 1282.410 1535.400 ;
        RECT 1277.030 1535.200 1282.410 1535.340 ;
        RECT 1277.030 1535.140 1277.350 1535.200 ;
        RECT 1282.090 1535.140 1282.410 1535.200 ;
        RECT 1282.090 47.160 1282.410 47.220 ;
        RECT 1282.090 47.020 1294.740 47.160 ;
        RECT 1282.090 46.960 1282.410 47.020 ;
        RECT 1294.600 46.820 1294.740 47.020 ;
        RECT 2672.670 46.820 2672.990 46.880 ;
        RECT 1294.600 46.680 2672.990 46.820 ;
        RECT 2672.670 46.620 2672.990 46.680 ;
      LAYER via ;
        RECT 1277.060 1535.140 1277.320 1535.400 ;
        RECT 1282.120 1535.140 1282.380 1535.400 ;
        RECT 1282.120 46.960 1282.380 47.220 ;
        RECT 2672.700 46.620 2672.960 46.880 ;
      LAYER met2 ;
        RECT 1276.460 1600.450 1276.740 1604.000 ;
        RECT 1276.460 1600.310 1277.260 1600.450 ;
        RECT 1276.460 1600.000 1276.740 1600.310 ;
        RECT 1277.120 1535.430 1277.260 1600.310 ;
        RECT 1277.060 1535.110 1277.320 1535.430 ;
        RECT 1282.120 1535.110 1282.380 1535.430 ;
        RECT 1282.180 47.250 1282.320 1535.110 ;
        RECT 1282.120 46.930 1282.380 47.250 ;
        RECT 2672.700 46.590 2672.960 46.910 ;
        RECT 2672.760 2.400 2672.900 46.590 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1282.090 1594.160 1282.410 1594.220 ;
        RECT 1283.010 1594.160 1283.330 1594.220 ;
        RECT 1282.090 1594.020 1283.330 1594.160 ;
        RECT 1282.090 1593.960 1282.410 1594.020 ;
        RECT 1283.010 1593.960 1283.330 1594.020 ;
        RECT 1276.570 1575.120 1276.890 1575.180 ;
        RECT 1282.090 1575.120 1282.410 1575.180 ;
        RECT 1276.570 1574.980 1282.410 1575.120 ;
        RECT 1276.570 1574.920 1276.890 1574.980 ;
        RECT 1282.090 1574.920 1282.410 1574.980 ;
        RECT 1276.570 1535.680 1276.890 1535.740 ;
        RECT 1282.550 1535.680 1282.870 1535.740 ;
        RECT 1276.570 1535.540 1282.870 1535.680 ;
        RECT 1276.570 1535.480 1276.890 1535.540 ;
        RECT 1282.550 1535.480 1282.870 1535.540 ;
        RECT 1282.550 46.480 1282.870 46.540 ;
        RECT 2690.610 46.480 2690.930 46.540 ;
        RECT 1282.550 46.340 2690.930 46.480 ;
        RECT 1282.550 46.280 1282.870 46.340 ;
        RECT 2690.610 46.280 2690.930 46.340 ;
      LAYER via ;
        RECT 1282.120 1593.960 1282.380 1594.220 ;
        RECT 1283.040 1593.960 1283.300 1594.220 ;
        RECT 1276.600 1574.920 1276.860 1575.180 ;
        RECT 1282.120 1574.920 1282.380 1575.180 ;
        RECT 1276.600 1535.480 1276.860 1535.740 ;
        RECT 1282.580 1535.480 1282.840 1535.740 ;
        RECT 1282.580 46.280 1282.840 46.540 ;
        RECT 2690.640 46.280 2690.900 46.540 ;
      LAYER met2 ;
        RECT 1282.440 1600.450 1282.720 1604.000 ;
        RECT 1282.440 1600.310 1283.240 1600.450 ;
        RECT 1282.440 1600.000 1282.720 1600.310 ;
        RECT 1283.100 1594.250 1283.240 1600.310 ;
        RECT 1282.120 1593.930 1282.380 1594.250 ;
        RECT 1283.040 1593.930 1283.300 1594.250 ;
        RECT 1282.180 1575.210 1282.320 1593.930 ;
        RECT 1276.600 1574.890 1276.860 1575.210 ;
        RECT 1282.120 1574.890 1282.380 1575.210 ;
        RECT 1276.660 1535.770 1276.800 1574.890 ;
        RECT 1276.600 1535.450 1276.860 1535.770 ;
        RECT 1282.580 1535.450 1282.840 1535.770 ;
        RECT 1282.640 46.570 1282.780 1535.450 ;
        RECT 1282.580 46.250 1282.840 46.570 ;
        RECT 2690.640 46.250 2690.900 46.570 ;
        RECT 2690.700 2.400 2690.840 46.250 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1287.150 1575.120 1287.470 1575.180 ;
        RECT 1289.450 1575.120 1289.770 1575.180 ;
        RECT 1287.150 1574.980 1289.770 1575.120 ;
        RECT 1287.150 1574.920 1287.470 1574.980 ;
        RECT 1289.450 1574.920 1289.770 1574.980 ;
        RECT 1289.450 46.140 1289.770 46.200 ;
        RECT 2708.550 46.140 2708.870 46.200 ;
        RECT 1289.450 46.000 2708.870 46.140 ;
        RECT 1289.450 45.940 1289.770 46.000 ;
        RECT 2708.550 45.940 2708.870 46.000 ;
      LAYER via ;
        RECT 1287.180 1574.920 1287.440 1575.180 ;
        RECT 1289.480 1574.920 1289.740 1575.180 ;
        RECT 1289.480 45.940 1289.740 46.200 ;
        RECT 2708.580 45.940 2708.840 46.200 ;
      LAYER met2 ;
        RECT 1288.880 1600.450 1289.160 1604.000 ;
        RECT 1287.240 1600.310 1289.160 1600.450 ;
        RECT 1287.240 1575.210 1287.380 1600.310 ;
        RECT 1288.880 1600.000 1289.160 1600.310 ;
        RECT 1287.180 1574.890 1287.440 1575.210 ;
        RECT 1289.480 1574.890 1289.740 1575.210 ;
        RECT 1289.540 46.230 1289.680 1574.890 ;
        RECT 1289.480 45.910 1289.740 46.230 ;
        RECT 2708.580 45.910 2708.840 46.230 ;
        RECT 2708.640 2.400 2708.780 45.910 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1296.425 1449.165 1296.595 1487.415 ;
        RECT 1296.425 1304.325 1296.595 1352.435 ;
        RECT 1296.425 476.085 1296.595 524.195 ;
        RECT 1296.425 379.525 1296.595 427.635 ;
        RECT 1296.425 282.965 1296.595 331.075 ;
        RECT 1296.425 186.405 1296.595 234.515 ;
      LAYER mcon ;
        RECT 1296.425 1487.245 1296.595 1487.415 ;
        RECT 1296.425 1352.265 1296.595 1352.435 ;
        RECT 1296.425 524.025 1296.595 524.195 ;
        RECT 1296.425 427.465 1296.595 427.635 ;
        RECT 1296.425 330.905 1296.595 331.075 ;
        RECT 1296.425 234.345 1296.595 234.515 ;
      LAYER met1 ;
        RECT 1295.890 1545.880 1296.210 1545.940 ;
        RECT 1296.350 1545.880 1296.670 1545.940 ;
        RECT 1295.890 1545.740 1296.670 1545.880 ;
        RECT 1295.890 1545.680 1296.210 1545.740 ;
        RECT 1296.350 1545.680 1296.670 1545.740 ;
        RECT 1295.890 1511.340 1296.210 1511.600 ;
        RECT 1295.980 1510.920 1296.120 1511.340 ;
        RECT 1295.890 1510.660 1296.210 1510.920 ;
        RECT 1295.890 1487.400 1296.210 1487.460 ;
        RECT 1296.365 1487.400 1296.655 1487.445 ;
        RECT 1295.890 1487.260 1296.655 1487.400 ;
        RECT 1295.890 1487.200 1296.210 1487.260 ;
        RECT 1296.365 1487.215 1296.655 1487.260 ;
        RECT 1296.350 1449.320 1296.670 1449.380 ;
        RECT 1296.155 1449.180 1296.670 1449.320 ;
        RECT 1296.350 1449.120 1296.670 1449.180 ;
        RECT 1296.350 1352.420 1296.670 1352.480 ;
        RECT 1296.155 1352.280 1296.670 1352.420 ;
        RECT 1296.350 1352.220 1296.670 1352.280 ;
        RECT 1296.350 1304.480 1296.670 1304.540 ;
        RECT 1296.155 1304.340 1296.670 1304.480 ;
        RECT 1296.350 1304.280 1296.670 1304.340 ;
        RECT 1295.430 1152.500 1295.750 1152.560 ;
        RECT 1296.350 1152.500 1296.670 1152.560 ;
        RECT 1295.430 1152.360 1296.670 1152.500 ;
        RECT 1295.430 1152.300 1295.750 1152.360 ;
        RECT 1296.350 1152.300 1296.670 1152.360 ;
        RECT 1295.430 910.760 1295.750 910.820 ;
        RECT 1296.350 910.760 1296.670 910.820 ;
        RECT 1295.430 910.620 1296.670 910.760 ;
        RECT 1295.430 910.560 1295.750 910.620 ;
        RECT 1296.350 910.560 1296.670 910.620 ;
        RECT 1295.430 814.200 1295.750 814.260 ;
        RECT 1296.350 814.200 1296.670 814.260 ;
        RECT 1295.430 814.060 1296.670 814.200 ;
        RECT 1295.430 814.000 1295.750 814.060 ;
        RECT 1296.350 814.000 1296.670 814.060 ;
        RECT 1295.430 717.640 1295.750 717.700 ;
        RECT 1296.350 717.640 1296.670 717.700 ;
        RECT 1295.430 717.500 1296.670 717.640 ;
        RECT 1295.430 717.440 1295.750 717.500 ;
        RECT 1296.350 717.440 1296.670 717.500 ;
        RECT 1295.430 572.800 1295.750 572.860 ;
        RECT 1296.350 572.800 1296.670 572.860 ;
        RECT 1295.430 572.660 1296.670 572.800 ;
        RECT 1295.430 572.600 1295.750 572.660 ;
        RECT 1296.350 572.600 1296.670 572.660 ;
        RECT 1296.350 524.180 1296.670 524.240 ;
        RECT 1296.155 524.040 1296.670 524.180 ;
        RECT 1296.350 523.980 1296.670 524.040 ;
        RECT 1296.350 476.240 1296.670 476.300 ;
        RECT 1296.155 476.100 1296.670 476.240 ;
        RECT 1296.350 476.040 1296.670 476.100 ;
        RECT 1296.350 427.620 1296.670 427.680 ;
        RECT 1296.155 427.480 1296.670 427.620 ;
        RECT 1296.350 427.420 1296.670 427.480 ;
        RECT 1296.350 379.680 1296.670 379.740 ;
        RECT 1296.155 379.540 1296.670 379.680 ;
        RECT 1296.350 379.480 1296.670 379.540 ;
        RECT 1296.350 331.060 1296.670 331.120 ;
        RECT 1296.155 330.920 1296.670 331.060 ;
        RECT 1296.350 330.860 1296.670 330.920 ;
        RECT 1296.350 283.120 1296.670 283.180 ;
        RECT 1296.155 282.980 1296.670 283.120 ;
        RECT 1296.350 282.920 1296.670 282.980 ;
        RECT 1296.350 234.500 1296.670 234.560 ;
        RECT 1296.155 234.360 1296.670 234.500 ;
        RECT 1296.350 234.300 1296.670 234.360 ;
        RECT 1296.350 186.560 1296.670 186.620 ;
        RECT 1296.155 186.420 1296.670 186.560 ;
        RECT 1296.350 186.360 1296.670 186.420 ;
      LAYER via ;
        RECT 1295.920 1545.680 1296.180 1545.940 ;
        RECT 1296.380 1545.680 1296.640 1545.940 ;
        RECT 1295.920 1511.340 1296.180 1511.600 ;
        RECT 1295.920 1510.660 1296.180 1510.920 ;
        RECT 1295.920 1487.200 1296.180 1487.460 ;
        RECT 1296.380 1449.120 1296.640 1449.380 ;
        RECT 1296.380 1352.220 1296.640 1352.480 ;
        RECT 1296.380 1304.280 1296.640 1304.540 ;
        RECT 1295.460 1152.300 1295.720 1152.560 ;
        RECT 1296.380 1152.300 1296.640 1152.560 ;
        RECT 1295.460 910.560 1295.720 910.820 ;
        RECT 1296.380 910.560 1296.640 910.820 ;
        RECT 1295.460 814.000 1295.720 814.260 ;
        RECT 1296.380 814.000 1296.640 814.260 ;
        RECT 1295.460 717.440 1295.720 717.700 ;
        RECT 1296.380 717.440 1296.640 717.700 ;
        RECT 1295.460 572.600 1295.720 572.860 ;
        RECT 1296.380 572.600 1296.640 572.860 ;
        RECT 1296.380 523.980 1296.640 524.240 ;
        RECT 1296.380 476.040 1296.640 476.300 ;
        RECT 1296.380 427.420 1296.640 427.680 ;
        RECT 1296.380 379.480 1296.640 379.740 ;
        RECT 1296.380 330.860 1296.640 331.120 ;
        RECT 1296.380 282.920 1296.640 283.180 ;
        RECT 1296.380 234.300 1296.640 234.560 ;
        RECT 1296.380 186.360 1296.640 186.620 ;
      LAYER met2 ;
        RECT 1294.860 1600.450 1295.140 1604.000 ;
        RECT 1294.860 1600.310 1296.120 1600.450 ;
        RECT 1294.860 1600.000 1295.140 1600.310 ;
        RECT 1295.980 1593.650 1296.120 1600.310 ;
        RECT 1295.980 1593.510 1296.580 1593.650 ;
        RECT 1296.440 1545.970 1296.580 1593.510 ;
        RECT 1295.920 1545.650 1296.180 1545.970 ;
        RECT 1296.380 1545.650 1296.640 1545.970 ;
        RECT 1295.980 1511.630 1296.120 1545.650 ;
        RECT 1295.920 1511.310 1296.180 1511.630 ;
        RECT 1295.920 1510.630 1296.180 1510.950 ;
        RECT 1295.980 1487.490 1296.120 1510.630 ;
        RECT 1295.920 1487.170 1296.180 1487.490 ;
        RECT 1296.380 1449.090 1296.640 1449.410 ;
        RECT 1296.440 1352.510 1296.580 1449.090 ;
        RECT 1296.380 1352.190 1296.640 1352.510 ;
        RECT 1296.380 1304.250 1296.640 1304.570 ;
        RECT 1296.440 1200.725 1296.580 1304.250 ;
        RECT 1295.450 1200.355 1295.730 1200.725 ;
        RECT 1296.370 1200.355 1296.650 1200.725 ;
        RECT 1295.520 1152.590 1295.660 1200.355 ;
        RECT 1295.460 1152.270 1295.720 1152.590 ;
        RECT 1296.380 1152.270 1296.640 1152.590 ;
        RECT 1296.440 1104.165 1296.580 1152.270 ;
        RECT 1295.450 1103.795 1295.730 1104.165 ;
        RECT 1296.370 1103.795 1296.650 1104.165 ;
        RECT 1295.520 1055.885 1295.660 1103.795 ;
        RECT 1295.450 1055.515 1295.730 1055.885 ;
        RECT 1296.370 1055.515 1296.650 1055.885 ;
        RECT 1296.440 910.850 1296.580 1055.515 ;
        RECT 1295.460 910.530 1295.720 910.850 ;
        RECT 1296.380 910.530 1296.640 910.850 ;
        RECT 1295.520 862.765 1295.660 910.530 ;
        RECT 1295.450 862.395 1295.730 862.765 ;
        RECT 1296.370 862.395 1296.650 862.765 ;
        RECT 1296.440 814.290 1296.580 862.395 ;
        RECT 1295.460 813.970 1295.720 814.290 ;
        RECT 1296.380 813.970 1296.640 814.290 ;
        RECT 1295.520 766.205 1295.660 813.970 ;
        RECT 1295.450 765.835 1295.730 766.205 ;
        RECT 1296.370 765.835 1296.650 766.205 ;
        RECT 1296.440 717.730 1296.580 765.835 ;
        RECT 1295.460 717.410 1295.720 717.730 ;
        RECT 1296.380 717.410 1296.640 717.730 ;
        RECT 1295.520 628.165 1295.660 717.410 ;
        RECT 1295.450 627.795 1295.730 628.165 ;
        RECT 1296.370 627.795 1296.650 628.165 ;
        RECT 1296.440 572.890 1296.580 627.795 ;
        RECT 1295.460 572.570 1295.720 572.890 ;
        RECT 1296.380 572.570 1296.640 572.890 ;
        RECT 1295.520 531.605 1295.660 572.570 ;
        RECT 1295.450 531.235 1295.730 531.605 ;
        RECT 1296.370 531.235 1296.650 531.605 ;
        RECT 1296.440 524.270 1296.580 531.235 ;
        RECT 1296.380 523.950 1296.640 524.270 ;
        RECT 1296.380 476.010 1296.640 476.330 ;
        RECT 1296.440 427.710 1296.580 476.010 ;
        RECT 1296.380 427.390 1296.640 427.710 ;
        RECT 1296.380 379.450 1296.640 379.770 ;
        RECT 1296.440 331.150 1296.580 379.450 ;
        RECT 1296.380 330.830 1296.640 331.150 ;
        RECT 1296.380 282.890 1296.640 283.210 ;
        RECT 1296.440 234.590 1296.580 282.890 ;
        RECT 1296.380 234.270 1296.640 234.590 ;
        RECT 1296.380 186.330 1296.640 186.650 ;
        RECT 1296.440 65.010 1296.580 186.330 ;
        RECT 1295.980 64.870 1296.580 65.010 ;
        RECT 1295.980 48.125 1296.120 64.870 ;
        RECT 1295.910 47.755 1296.190 48.125 ;
        RECT 2726.510 47.755 2726.790 48.125 ;
        RECT 2726.580 2.400 2726.720 47.755 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
      LAYER via2 ;
        RECT 1295.450 1200.400 1295.730 1200.680 ;
        RECT 1296.370 1200.400 1296.650 1200.680 ;
        RECT 1295.450 1103.840 1295.730 1104.120 ;
        RECT 1296.370 1103.840 1296.650 1104.120 ;
        RECT 1295.450 1055.560 1295.730 1055.840 ;
        RECT 1296.370 1055.560 1296.650 1055.840 ;
        RECT 1295.450 862.440 1295.730 862.720 ;
        RECT 1296.370 862.440 1296.650 862.720 ;
        RECT 1295.450 765.880 1295.730 766.160 ;
        RECT 1296.370 765.880 1296.650 766.160 ;
        RECT 1295.450 627.840 1295.730 628.120 ;
        RECT 1296.370 627.840 1296.650 628.120 ;
        RECT 1295.450 531.280 1295.730 531.560 ;
        RECT 1296.370 531.280 1296.650 531.560 ;
        RECT 1295.910 47.800 1296.190 48.080 ;
        RECT 2726.510 47.800 2726.790 48.080 ;
      LAYER met3 ;
        RECT 1295.425 1200.690 1295.755 1200.705 ;
        RECT 1296.345 1200.690 1296.675 1200.705 ;
        RECT 1295.425 1200.390 1296.675 1200.690 ;
        RECT 1295.425 1200.375 1295.755 1200.390 ;
        RECT 1296.345 1200.375 1296.675 1200.390 ;
        RECT 1295.425 1104.130 1295.755 1104.145 ;
        RECT 1296.345 1104.130 1296.675 1104.145 ;
        RECT 1295.425 1103.830 1296.675 1104.130 ;
        RECT 1295.425 1103.815 1295.755 1103.830 ;
        RECT 1296.345 1103.815 1296.675 1103.830 ;
        RECT 1295.425 1055.850 1295.755 1055.865 ;
        RECT 1296.345 1055.850 1296.675 1055.865 ;
        RECT 1295.425 1055.550 1296.675 1055.850 ;
        RECT 1295.425 1055.535 1295.755 1055.550 ;
        RECT 1296.345 1055.535 1296.675 1055.550 ;
        RECT 1295.425 862.730 1295.755 862.745 ;
        RECT 1296.345 862.730 1296.675 862.745 ;
        RECT 1295.425 862.430 1296.675 862.730 ;
        RECT 1295.425 862.415 1295.755 862.430 ;
        RECT 1296.345 862.415 1296.675 862.430 ;
        RECT 1295.425 766.170 1295.755 766.185 ;
        RECT 1296.345 766.170 1296.675 766.185 ;
        RECT 1295.425 765.870 1296.675 766.170 ;
        RECT 1295.425 765.855 1295.755 765.870 ;
        RECT 1296.345 765.855 1296.675 765.870 ;
        RECT 1295.425 628.130 1295.755 628.145 ;
        RECT 1296.345 628.130 1296.675 628.145 ;
        RECT 1295.425 627.830 1296.675 628.130 ;
        RECT 1295.425 627.815 1295.755 627.830 ;
        RECT 1296.345 627.815 1296.675 627.830 ;
        RECT 1295.425 531.570 1295.755 531.585 ;
        RECT 1296.345 531.570 1296.675 531.585 ;
        RECT 1295.425 531.270 1296.675 531.570 ;
        RECT 1295.425 531.255 1295.755 531.270 ;
        RECT 1296.345 531.255 1296.675 531.270 ;
        RECT 1295.885 48.090 1296.215 48.105 ;
        RECT 2726.485 48.090 2726.815 48.105 ;
        RECT 1295.885 47.790 2726.815 48.090 ;
        RECT 1295.885 47.775 1296.215 47.790 ;
        RECT 2726.485 47.775 2726.815 47.790 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1297.270 1579.880 1297.590 1579.940 ;
        RECT 1300.030 1579.880 1300.350 1579.940 ;
        RECT 1297.270 1579.740 1300.350 1579.880 ;
        RECT 1297.270 1579.680 1297.590 1579.740 ;
        RECT 1300.030 1579.680 1300.350 1579.740 ;
        RECT 1297.270 1535.000 1297.590 1535.060 ;
        RECT 1303.250 1535.000 1303.570 1535.060 ;
        RECT 1297.270 1534.860 1303.570 1535.000 ;
        RECT 1297.270 1534.800 1297.590 1534.860 ;
        RECT 1303.250 1534.800 1303.570 1534.860 ;
        RECT 1303.250 45.800 1303.570 45.860 ;
        RECT 2744.430 45.800 2744.750 45.860 ;
        RECT 1303.250 45.660 2744.750 45.800 ;
        RECT 1303.250 45.600 1303.570 45.660 ;
        RECT 2744.430 45.600 2744.750 45.660 ;
      LAYER via ;
        RECT 1297.300 1579.680 1297.560 1579.940 ;
        RECT 1300.060 1579.680 1300.320 1579.940 ;
        RECT 1297.300 1534.800 1297.560 1535.060 ;
        RECT 1303.280 1534.800 1303.540 1535.060 ;
        RECT 1303.280 45.600 1303.540 45.860 ;
        RECT 2744.460 45.600 2744.720 45.860 ;
      LAYER met2 ;
        RECT 1301.300 1600.450 1301.580 1604.000 ;
        RECT 1300.120 1600.310 1301.580 1600.450 ;
        RECT 1300.120 1579.970 1300.260 1600.310 ;
        RECT 1301.300 1600.000 1301.580 1600.310 ;
        RECT 1297.300 1579.650 1297.560 1579.970 ;
        RECT 1300.060 1579.650 1300.320 1579.970 ;
        RECT 1297.360 1535.090 1297.500 1579.650 ;
        RECT 1297.300 1534.770 1297.560 1535.090 ;
        RECT 1303.280 1534.770 1303.540 1535.090 ;
        RECT 1303.340 45.890 1303.480 1534.770 ;
        RECT 1303.280 45.570 1303.540 45.890 ;
        RECT 2744.460 45.570 2744.720 45.890 ;
        RECT 2744.520 2.400 2744.660 45.570 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1309.765 148.325 1309.935 165.835 ;
      LAYER mcon ;
        RECT 1309.765 165.665 1309.935 165.835 ;
      LAYER met1 ;
        RECT 1307.850 1594.160 1308.170 1594.220 ;
        RECT 1308.310 1594.160 1308.630 1594.220 ;
        RECT 1307.850 1594.020 1308.630 1594.160 ;
        RECT 1307.850 1593.960 1308.170 1594.020 ;
        RECT 1308.310 1593.960 1308.630 1594.020 ;
        RECT 1310.150 331.060 1310.470 331.120 ;
        RECT 1311.070 331.060 1311.390 331.120 ;
        RECT 1310.150 330.920 1311.390 331.060 ;
        RECT 1310.150 330.860 1310.470 330.920 ;
        RECT 1311.070 330.860 1311.390 330.920 ;
        RECT 1310.150 247.080 1310.470 247.140 ;
        RECT 1311.070 247.080 1311.390 247.140 ;
        RECT 1310.150 246.940 1311.390 247.080 ;
        RECT 1310.150 246.880 1310.470 246.940 ;
        RECT 1311.070 246.880 1311.390 246.940 ;
        RECT 1310.150 166.160 1310.470 166.220 ;
        RECT 1309.320 166.020 1310.470 166.160 ;
        RECT 1309.320 165.820 1309.460 166.020 ;
        RECT 1310.150 165.960 1310.470 166.020 ;
        RECT 1309.705 165.820 1309.995 165.865 ;
        RECT 1309.320 165.680 1309.995 165.820 ;
        RECT 1309.705 165.635 1309.995 165.680 ;
        RECT 1309.705 148.480 1309.995 148.525 ;
        RECT 1310.150 148.480 1310.470 148.540 ;
        RECT 1309.705 148.340 1310.470 148.480 ;
        RECT 1309.705 148.295 1309.995 148.340 ;
        RECT 1310.150 148.280 1310.470 148.340 ;
        RECT 1310.150 116.860 1310.470 116.920 ;
        RECT 1311.070 116.860 1311.390 116.920 ;
        RECT 1310.150 116.720 1311.390 116.860 ;
        RECT 1310.150 116.660 1310.470 116.720 ;
        RECT 1311.070 116.660 1311.390 116.720 ;
      LAYER via ;
        RECT 1307.880 1593.960 1308.140 1594.220 ;
        RECT 1308.340 1593.960 1308.600 1594.220 ;
        RECT 1310.180 330.860 1310.440 331.120 ;
        RECT 1311.100 330.860 1311.360 331.120 ;
        RECT 1310.180 246.880 1310.440 247.140 ;
        RECT 1311.100 246.880 1311.360 247.140 ;
        RECT 1310.180 165.960 1310.440 166.220 ;
        RECT 1310.180 148.280 1310.440 148.540 ;
        RECT 1310.180 116.660 1310.440 116.920 ;
        RECT 1311.100 116.660 1311.360 116.920 ;
      LAYER met2 ;
        RECT 1307.280 1600.450 1307.560 1604.000 ;
        RECT 1307.280 1600.310 1308.080 1600.450 ;
        RECT 1307.280 1600.000 1307.560 1600.310 ;
        RECT 1307.940 1594.250 1308.080 1600.310 ;
        RECT 1307.880 1593.930 1308.140 1594.250 ;
        RECT 1308.340 1593.930 1308.600 1594.250 ;
        RECT 1308.400 1569.680 1308.540 1593.930 ;
        RECT 1308.400 1569.540 1309.000 1569.680 ;
        RECT 1308.860 1545.370 1309.000 1569.540 ;
        RECT 1308.860 1545.230 1310.380 1545.370 ;
        RECT 1310.240 331.150 1310.380 1545.230 ;
        RECT 1310.180 330.830 1310.440 331.150 ;
        RECT 1311.100 330.830 1311.360 331.150 ;
        RECT 1311.160 247.170 1311.300 330.830 ;
        RECT 1310.180 246.850 1310.440 247.170 ;
        RECT 1311.100 246.850 1311.360 247.170 ;
        RECT 1310.240 166.250 1310.380 246.850 ;
        RECT 1310.180 165.930 1310.440 166.250 ;
        RECT 1310.180 148.250 1310.440 148.570 ;
        RECT 1310.240 116.950 1310.380 148.250 ;
        RECT 1310.180 116.630 1310.440 116.950 ;
        RECT 1311.100 116.630 1311.360 116.950 ;
        RECT 1311.160 69.205 1311.300 116.630 ;
        RECT 1311.090 68.835 1311.370 69.205 ;
        RECT 1312.010 68.835 1312.290 69.205 ;
        RECT 1312.080 47.445 1312.220 68.835 ;
        RECT 1312.010 47.075 1312.290 47.445 ;
        RECT 2761.930 47.075 2762.210 47.445 ;
        RECT 2762.000 2.400 2762.140 47.075 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
      LAYER via2 ;
        RECT 1311.090 68.880 1311.370 69.160 ;
        RECT 1312.010 68.880 1312.290 69.160 ;
        RECT 1312.010 47.120 1312.290 47.400 ;
        RECT 2761.930 47.120 2762.210 47.400 ;
      LAYER met3 ;
        RECT 1311.065 69.170 1311.395 69.185 ;
        RECT 1311.985 69.170 1312.315 69.185 ;
        RECT 1311.065 68.870 1312.315 69.170 ;
        RECT 1311.065 68.855 1311.395 68.870 ;
        RECT 1311.985 68.855 1312.315 68.870 ;
        RECT 1311.985 47.410 1312.315 47.425 ;
        RECT 2761.905 47.410 2762.235 47.425 ;
        RECT 1311.985 47.110 2762.235 47.410 ;
        RECT 1311.985 47.095 1312.315 47.110 ;
        RECT 2761.905 47.095 2762.235 47.110 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 639.470 1592.800 639.790 1592.860 ;
        RECT 824.390 1592.800 824.710 1592.860 ;
        RECT 639.470 1592.660 824.710 1592.800 ;
        RECT 639.470 1592.600 639.790 1592.660 ;
        RECT 824.390 1592.600 824.710 1592.660 ;
        RECT 824.390 17.920 824.710 17.980 ;
        RECT 835.430 17.920 835.750 17.980 ;
        RECT 824.390 17.780 835.750 17.920 ;
        RECT 824.390 17.720 824.710 17.780 ;
        RECT 835.430 17.720 835.750 17.780 ;
      LAYER via ;
        RECT 639.500 1592.600 639.760 1592.860 ;
        RECT 824.420 1592.600 824.680 1592.860 ;
        RECT 824.420 17.720 824.680 17.980 ;
        RECT 835.460 17.720 835.720 17.980 ;
      LAYER met2 ;
        RECT 639.360 1600.380 639.640 1604.000 ;
        RECT 639.360 1600.000 639.700 1600.380 ;
        RECT 639.560 1592.890 639.700 1600.000 ;
        RECT 639.500 1592.570 639.760 1592.890 ;
        RECT 824.420 1592.570 824.680 1592.890 ;
        RECT 824.480 18.010 824.620 1592.570 ;
        RECT 824.420 17.690 824.680 18.010 ;
        RECT 835.460 17.690 835.720 18.010 ;
        RECT 835.520 2.400 835.660 17.690 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1311.070 1563.560 1311.390 1563.620 ;
        RECT 1312.450 1563.560 1312.770 1563.620 ;
        RECT 1311.070 1563.420 1312.770 1563.560 ;
        RECT 1311.070 1563.360 1311.390 1563.420 ;
        RECT 1312.450 1563.360 1312.770 1563.420 ;
        RECT 1311.070 1535.340 1311.390 1535.400 ;
        RECT 1316.590 1535.340 1316.910 1535.400 ;
        RECT 1311.070 1535.200 1316.910 1535.340 ;
        RECT 1311.070 1535.140 1311.390 1535.200 ;
        RECT 1316.590 1535.140 1316.910 1535.200 ;
      LAYER via ;
        RECT 1311.100 1563.360 1311.360 1563.620 ;
        RECT 1312.480 1563.360 1312.740 1563.620 ;
        RECT 1311.100 1535.140 1311.360 1535.400 ;
        RECT 1316.620 1535.140 1316.880 1535.400 ;
      LAYER met2 ;
        RECT 1313.260 1600.450 1313.540 1604.000 ;
        RECT 1312.540 1600.310 1313.540 1600.450 ;
        RECT 1312.540 1563.650 1312.680 1600.310 ;
        RECT 1313.260 1600.000 1313.540 1600.310 ;
        RECT 1311.100 1563.330 1311.360 1563.650 ;
        RECT 1312.480 1563.330 1312.740 1563.650 ;
        RECT 1311.160 1535.430 1311.300 1563.330 ;
        RECT 1311.100 1535.110 1311.360 1535.430 ;
        RECT 1316.620 1535.110 1316.880 1535.430 ;
        RECT 1316.680 66.370 1316.820 1535.110 ;
        RECT 1316.220 66.230 1316.820 66.370 ;
        RECT 1316.220 46.765 1316.360 66.230 ;
        RECT 1316.150 46.395 1316.430 46.765 ;
        RECT 2779.870 46.395 2780.150 46.765 ;
        RECT 2779.940 2.400 2780.080 46.395 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
      LAYER via2 ;
        RECT 1316.150 46.440 1316.430 46.720 ;
        RECT 2779.870 46.440 2780.150 46.720 ;
      LAYER met3 ;
        RECT 1316.125 46.730 1316.455 46.745 ;
        RECT 2779.845 46.730 2780.175 46.745 ;
        RECT 1316.125 46.430 2780.175 46.730 ;
        RECT 1316.125 46.415 1316.455 46.430 ;
        RECT 2779.845 46.415 2780.175 46.430 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1320.730 1569.680 1321.050 1569.740 ;
        RECT 1323.490 1569.680 1323.810 1569.740 ;
        RECT 1320.730 1569.540 1323.810 1569.680 ;
        RECT 1320.730 1569.480 1321.050 1569.540 ;
        RECT 1323.490 1569.480 1323.810 1569.540 ;
        RECT 1323.490 1545.340 1323.810 1545.600 ;
        RECT 1323.580 1545.200 1323.720 1545.340 ;
        RECT 1323.950 1545.200 1324.270 1545.260 ;
        RECT 1323.580 1545.060 1324.270 1545.200 ;
        RECT 1323.950 1545.000 1324.270 1545.060 ;
        RECT 1323.950 717.640 1324.270 717.700 ;
        RECT 1324.870 717.640 1325.190 717.700 ;
        RECT 1323.950 717.500 1325.190 717.640 ;
        RECT 1323.950 717.440 1324.270 717.500 ;
        RECT 1324.870 717.440 1325.190 717.500 ;
      LAYER via ;
        RECT 1320.760 1569.480 1321.020 1569.740 ;
        RECT 1323.520 1569.480 1323.780 1569.740 ;
        RECT 1323.520 1545.340 1323.780 1545.600 ;
        RECT 1323.980 1545.000 1324.240 1545.260 ;
        RECT 1323.980 717.440 1324.240 717.700 ;
        RECT 1324.900 717.440 1325.160 717.700 ;
      LAYER met2 ;
        RECT 1319.700 1600.450 1319.980 1604.000 ;
        RECT 1319.700 1600.310 1320.960 1600.450 ;
        RECT 1319.700 1600.000 1319.980 1600.310 ;
        RECT 1320.820 1569.770 1320.960 1600.310 ;
        RECT 1320.760 1569.450 1321.020 1569.770 ;
        RECT 1323.520 1569.450 1323.780 1569.770 ;
        RECT 1323.580 1545.630 1323.720 1569.450 ;
        RECT 1323.520 1545.310 1323.780 1545.630 ;
        RECT 1323.980 1544.970 1324.240 1545.290 ;
        RECT 1324.040 717.730 1324.180 1544.970 ;
        RECT 1323.980 717.410 1324.240 717.730 ;
        RECT 1324.900 717.410 1325.160 717.730 ;
        RECT 1324.960 669.645 1325.100 717.410 ;
        RECT 1323.970 669.275 1324.250 669.645 ;
        RECT 1324.890 669.275 1325.170 669.645 ;
        RECT 1324.040 46.085 1324.180 669.275 ;
        RECT 1323.970 45.715 1324.250 46.085 ;
        RECT 2797.810 45.715 2798.090 46.085 ;
        RECT 2797.880 2.400 2798.020 45.715 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
      LAYER via2 ;
        RECT 1323.970 669.320 1324.250 669.600 ;
        RECT 1324.890 669.320 1325.170 669.600 ;
        RECT 1323.970 45.760 1324.250 46.040 ;
        RECT 2797.810 45.760 2798.090 46.040 ;
      LAYER met3 ;
        RECT 1323.945 669.610 1324.275 669.625 ;
        RECT 1324.865 669.610 1325.195 669.625 ;
        RECT 1323.945 669.310 1325.195 669.610 ;
        RECT 1323.945 669.295 1324.275 669.310 ;
        RECT 1324.865 669.295 1325.195 669.310 ;
        RECT 1323.945 46.050 1324.275 46.065 ;
        RECT 2797.785 46.050 2798.115 46.065 ;
        RECT 1323.945 45.750 2798.115 46.050 ;
        RECT 1323.945 45.735 1324.275 45.750 ;
        RECT 2797.785 45.735 2798.115 45.750 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1326.250 1579.880 1326.570 1579.940 ;
        RECT 1330.390 1579.880 1330.710 1579.940 ;
        RECT 1326.250 1579.740 1330.710 1579.880 ;
        RECT 1326.250 1579.680 1326.570 1579.740 ;
        RECT 1330.390 1579.680 1330.710 1579.740 ;
        RECT 1330.390 1497.600 1330.710 1497.660 ;
        RECT 1330.850 1497.600 1331.170 1497.660 ;
        RECT 1330.390 1497.460 1331.170 1497.600 ;
        RECT 1330.390 1497.400 1330.710 1497.460 ;
        RECT 1330.850 1497.400 1331.170 1497.460 ;
      LAYER via ;
        RECT 1326.280 1579.680 1326.540 1579.940 ;
        RECT 1330.420 1579.680 1330.680 1579.940 ;
        RECT 1330.420 1497.400 1330.680 1497.660 ;
        RECT 1330.880 1497.400 1331.140 1497.660 ;
      LAYER met2 ;
        RECT 1325.680 1600.450 1325.960 1604.000 ;
        RECT 1325.680 1600.310 1326.480 1600.450 ;
        RECT 1325.680 1600.000 1325.960 1600.310 ;
        RECT 1326.340 1579.970 1326.480 1600.310 ;
        RECT 1326.280 1579.650 1326.540 1579.970 ;
        RECT 1330.420 1579.650 1330.680 1579.970 ;
        RECT 1330.480 1497.690 1330.620 1579.650 ;
        RECT 1330.420 1497.370 1330.680 1497.690 ;
        RECT 1330.880 1497.370 1331.140 1497.690 ;
        RECT 1330.940 65.010 1331.080 1497.370 ;
        RECT 1330.480 64.870 1331.080 65.010 ;
        RECT 1330.480 48.010 1330.620 64.870 ;
        RECT 1330.480 47.870 1331.080 48.010 ;
        RECT 1330.940 45.405 1331.080 47.870 ;
        RECT 1330.870 45.035 1331.150 45.405 ;
        RECT 2815.750 45.035 2816.030 45.405 ;
        RECT 2815.820 2.400 2815.960 45.035 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
      LAYER via2 ;
        RECT 1330.870 45.080 1331.150 45.360 ;
        RECT 2815.750 45.080 2816.030 45.360 ;
      LAYER met3 ;
        RECT 1330.845 45.370 1331.175 45.385 ;
        RECT 2815.725 45.370 2816.055 45.385 ;
        RECT 1330.845 45.070 2816.055 45.370 ;
        RECT 1330.845 45.055 1331.175 45.070 ;
        RECT 2815.725 45.055 2816.055 45.070 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1333.150 1600.960 1333.470 1601.020 ;
        RECT 1337.290 1600.960 1337.610 1601.020 ;
        RECT 1333.150 1600.820 1337.610 1600.960 ;
        RECT 1333.150 1600.760 1333.470 1600.820 ;
        RECT 1337.290 1600.760 1337.610 1600.820 ;
        RECT 1337.290 45.460 1337.610 45.520 ;
        RECT 2833.670 45.460 2833.990 45.520 ;
        RECT 1337.290 45.320 2833.990 45.460 ;
        RECT 1337.290 45.260 1337.610 45.320 ;
        RECT 2833.670 45.260 2833.990 45.320 ;
      LAYER via ;
        RECT 1333.180 1600.760 1333.440 1601.020 ;
        RECT 1337.320 1600.760 1337.580 1601.020 ;
        RECT 1337.320 45.260 1337.580 45.520 ;
        RECT 2833.700 45.260 2833.960 45.520 ;
      LAYER met2 ;
        RECT 1332.120 1601.130 1332.400 1604.000 ;
        RECT 1332.120 1601.050 1333.380 1601.130 ;
        RECT 1332.120 1600.990 1333.440 1601.050 ;
        RECT 1332.120 1600.000 1332.400 1600.990 ;
        RECT 1333.180 1600.730 1333.440 1600.990 ;
        RECT 1337.320 1600.730 1337.580 1601.050 ;
        RECT 1337.380 45.550 1337.520 1600.730 ;
        RECT 1337.320 45.230 1337.580 45.550 ;
        RECT 2833.700 45.230 2833.960 45.550 ;
        RECT 2833.760 2.400 2833.900 45.230 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1336.830 1597.220 1337.150 1597.280 ;
        RECT 1337.750 1597.220 1338.070 1597.280 ;
        RECT 1336.830 1597.080 1338.070 1597.220 ;
        RECT 1336.830 1597.020 1337.150 1597.080 ;
        RECT 1337.750 1597.020 1338.070 1597.080 ;
        RECT 1332.230 1579.540 1332.550 1579.600 ;
        RECT 1337.750 1579.540 1338.070 1579.600 ;
        RECT 1332.230 1579.400 1338.070 1579.540 ;
        RECT 1332.230 1579.340 1332.550 1579.400 ;
        RECT 1337.750 1579.340 1338.070 1579.400 ;
        RECT 1332.230 1535.000 1332.550 1535.060 ;
        RECT 1337.750 1535.000 1338.070 1535.060 ;
        RECT 1332.230 1534.860 1338.070 1535.000 ;
        RECT 1332.230 1534.800 1332.550 1534.860 ;
        RECT 1337.750 1534.800 1338.070 1534.860 ;
        RECT 1337.750 45.120 1338.070 45.180 ;
        RECT 2851.150 45.120 2851.470 45.180 ;
        RECT 1337.750 44.980 2851.470 45.120 ;
        RECT 1337.750 44.920 1338.070 44.980 ;
        RECT 2851.150 44.920 2851.470 44.980 ;
      LAYER via ;
        RECT 1336.860 1597.020 1337.120 1597.280 ;
        RECT 1337.780 1597.020 1338.040 1597.280 ;
        RECT 1332.260 1579.340 1332.520 1579.600 ;
        RECT 1337.780 1579.340 1338.040 1579.600 ;
        RECT 1332.260 1534.800 1332.520 1535.060 ;
        RECT 1337.780 1534.800 1338.040 1535.060 ;
        RECT 1337.780 44.920 1338.040 45.180 ;
        RECT 2851.180 44.920 2851.440 45.180 ;
      LAYER met2 ;
        RECT 1338.100 1601.810 1338.380 1604.000 ;
        RECT 1336.920 1601.670 1338.380 1601.810 ;
        RECT 1336.920 1597.310 1337.060 1601.670 ;
        RECT 1338.100 1600.000 1338.380 1601.670 ;
        RECT 1336.860 1596.990 1337.120 1597.310 ;
        RECT 1337.780 1596.990 1338.040 1597.310 ;
        RECT 1337.840 1579.630 1337.980 1596.990 ;
        RECT 1332.260 1579.310 1332.520 1579.630 ;
        RECT 1337.780 1579.310 1338.040 1579.630 ;
        RECT 1332.320 1535.090 1332.460 1579.310 ;
        RECT 1332.260 1534.770 1332.520 1535.090 ;
        RECT 1337.780 1534.770 1338.040 1535.090 ;
        RECT 1337.840 45.210 1337.980 1534.770 ;
        RECT 1337.780 44.890 1338.040 45.210 ;
        RECT 2851.180 44.890 2851.440 45.210 ;
        RECT 2851.240 2.400 2851.380 44.890 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.670 1587.020 1338.990 1587.080 ;
        RECT 1344.650 1587.020 1344.970 1587.080 ;
        RECT 1338.670 1586.880 1344.970 1587.020 ;
        RECT 1338.670 1586.820 1338.990 1586.880 ;
        RECT 1344.650 1586.820 1344.970 1586.880 ;
        RECT 1338.670 1535.340 1338.990 1535.400 ;
        RECT 1344.650 1535.340 1344.970 1535.400 ;
        RECT 1338.670 1535.200 1344.970 1535.340 ;
        RECT 1338.670 1535.140 1338.990 1535.200 ;
        RECT 1344.650 1535.140 1344.970 1535.200 ;
      LAYER via ;
        RECT 1338.700 1586.820 1338.960 1587.080 ;
        RECT 1344.680 1586.820 1344.940 1587.080 ;
        RECT 1338.700 1535.140 1338.960 1535.400 ;
        RECT 1344.680 1535.140 1344.940 1535.400 ;
      LAYER met2 ;
        RECT 1344.540 1600.380 1344.820 1604.000 ;
        RECT 1344.540 1600.000 1344.880 1600.380 ;
        RECT 1344.740 1587.110 1344.880 1600.000 ;
        RECT 1338.700 1586.790 1338.960 1587.110 ;
        RECT 1344.680 1586.790 1344.940 1587.110 ;
        RECT 1338.760 1535.430 1338.900 1586.790 ;
        RECT 1338.700 1535.110 1338.960 1535.430 ;
        RECT 1344.680 1535.110 1344.940 1535.430 ;
        RECT 1344.740 44.725 1344.880 1535.110 ;
        RECT 1344.670 44.355 1344.950 44.725 ;
        RECT 2869.110 44.355 2869.390 44.725 ;
        RECT 2869.180 2.400 2869.320 44.355 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
      LAYER via2 ;
        RECT 1344.670 44.400 1344.950 44.680 ;
        RECT 2869.110 44.400 2869.390 44.680 ;
      LAYER met3 ;
        RECT 1344.645 44.690 1344.975 44.705 ;
        RECT 2869.085 44.690 2869.415 44.705 ;
        RECT 1344.645 44.390 2869.415 44.690 ;
        RECT 1344.645 44.375 1344.975 44.390 ;
        RECT 2869.085 44.375 2869.415 44.390 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1345.570 1600.960 1345.890 1601.020 ;
        RECT 1349.250 1600.960 1349.570 1601.020 ;
        RECT 1345.570 1600.820 1349.570 1600.960 ;
        RECT 1345.570 1600.760 1345.890 1600.820 ;
        RECT 1349.250 1600.760 1349.570 1600.820 ;
        RECT 1345.570 1528.880 1345.890 1528.940 ;
        RECT 1351.090 1528.880 1351.410 1528.940 ;
        RECT 1345.570 1528.740 1351.410 1528.880 ;
        RECT 1345.570 1528.680 1345.890 1528.740 ;
        RECT 1351.090 1528.680 1351.410 1528.740 ;
        RECT 2884.270 2.960 2884.590 3.020 ;
        RECT 2887.030 2.960 2887.350 3.020 ;
        RECT 2884.270 2.820 2887.350 2.960 ;
        RECT 2884.270 2.760 2884.590 2.820 ;
        RECT 2887.030 2.760 2887.350 2.820 ;
      LAYER via ;
        RECT 1345.600 1600.760 1345.860 1601.020 ;
        RECT 1349.280 1600.760 1349.540 1601.020 ;
        RECT 1345.600 1528.680 1345.860 1528.940 ;
        RECT 1351.120 1528.680 1351.380 1528.940 ;
        RECT 2884.300 2.760 2884.560 3.020 ;
        RECT 2887.060 2.760 2887.320 3.020 ;
      LAYER met2 ;
        RECT 1350.520 1601.130 1350.800 1604.000 ;
        RECT 1349.340 1601.050 1350.800 1601.130 ;
        RECT 1345.600 1600.730 1345.860 1601.050 ;
        RECT 1349.280 1600.990 1350.800 1601.050 ;
        RECT 1349.280 1600.730 1349.540 1600.990 ;
        RECT 1345.660 1528.970 1345.800 1600.730 ;
        RECT 1350.520 1600.000 1350.800 1600.990 ;
        RECT 1345.600 1528.650 1345.860 1528.970 ;
        RECT 1351.120 1528.650 1351.380 1528.970 ;
        RECT 1351.180 73.965 1351.320 1528.650 ;
        RECT 1351.110 73.595 1351.390 73.965 ;
        RECT 2884.290 73.595 2884.570 73.965 ;
        RECT 2884.360 3.050 2884.500 73.595 ;
        RECT 2884.300 2.730 2884.560 3.050 ;
        RECT 2887.060 2.730 2887.320 3.050 ;
        RECT 2887.120 2.400 2887.260 2.730 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
      LAYER via2 ;
        RECT 1351.110 73.640 1351.390 73.920 ;
        RECT 2884.290 73.640 2884.570 73.920 ;
      LAYER met3 ;
        RECT 1351.085 73.930 1351.415 73.945 ;
        RECT 2884.265 73.930 2884.595 73.945 ;
        RECT 1351.085 73.630 2884.595 73.930 ;
        RECT 1351.085 73.615 1351.415 73.630 ;
        RECT 2884.265 73.615 2884.595 73.630 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1358.450 44.780 1358.770 44.840 ;
        RECT 2905.430 44.780 2905.750 44.840 ;
        RECT 1358.450 44.640 2905.750 44.780 ;
        RECT 1358.450 44.580 1358.770 44.640 ;
        RECT 2905.430 44.580 2905.750 44.640 ;
      LAYER via ;
        RECT 1358.480 44.580 1358.740 44.840 ;
        RECT 2905.460 44.580 2905.720 44.840 ;
      LAYER met2 ;
        RECT 1356.960 1600.450 1357.240 1604.000 ;
        RECT 1356.960 1600.310 1358.220 1600.450 ;
        RECT 1356.960 1600.000 1357.240 1600.310 ;
        RECT 1358.080 1579.370 1358.220 1600.310 ;
        RECT 1358.080 1579.230 1358.680 1579.370 ;
        RECT 1358.540 44.870 1358.680 1579.230 ;
        RECT 1358.480 44.550 1358.740 44.870 ;
        RECT 2905.460 44.550 2905.720 44.870 ;
        RECT 2905.520 7.210 2905.660 44.550 ;
        RECT 2905.060 7.070 2905.660 7.210 ;
        RECT 2905.060 2.400 2905.200 7.070 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 645.450 1589.060 645.770 1589.120 ;
        RECT 647.290 1589.060 647.610 1589.120 ;
        RECT 645.450 1588.920 647.610 1589.060 ;
        RECT 645.450 1588.860 645.770 1588.920 ;
        RECT 647.290 1588.860 647.610 1588.920 ;
        RECT 647.290 32.880 647.610 32.940 ;
        RECT 852.910 32.880 853.230 32.940 ;
        RECT 647.290 32.740 853.230 32.880 ;
        RECT 647.290 32.680 647.610 32.740 ;
        RECT 852.910 32.680 853.230 32.740 ;
      LAYER via ;
        RECT 645.480 1588.860 645.740 1589.120 ;
        RECT 647.320 1588.860 647.580 1589.120 ;
        RECT 647.320 32.680 647.580 32.940 ;
        RECT 852.940 32.680 853.200 32.940 ;
      LAYER met2 ;
        RECT 645.340 1600.380 645.620 1604.000 ;
        RECT 645.340 1600.000 645.680 1600.380 ;
        RECT 645.540 1589.150 645.680 1600.000 ;
        RECT 645.480 1588.830 645.740 1589.150 ;
        RECT 647.320 1588.830 647.580 1589.150 ;
        RECT 647.380 32.970 647.520 1588.830 ;
        RECT 647.320 32.650 647.580 32.970 ;
        RECT 852.940 32.650 853.200 32.970 ;
        RECT 853.000 2.400 853.140 32.650 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 651.890 1589.060 652.210 1589.120 ;
        RECT 654.190 1589.060 654.510 1589.120 ;
        RECT 651.890 1588.920 654.510 1589.060 ;
        RECT 651.890 1588.860 652.210 1588.920 ;
        RECT 654.190 1588.860 654.510 1588.920 ;
        RECT 654.190 32.540 654.510 32.600 ;
        RECT 870.850 32.540 871.170 32.600 ;
        RECT 654.190 32.400 871.170 32.540 ;
        RECT 654.190 32.340 654.510 32.400 ;
        RECT 870.850 32.340 871.170 32.400 ;
      LAYER via ;
        RECT 651.920 1588.860 652.180 1589.120 ;
        RECT 654.220 1588.860 654.480 1589.120 ;
        RECT 654.220 32.340 654.480 32.600 ;
        RECT 870.880 32.340 871.140 32.600 ;
      LAYER met2 ;
        RECT 651.780 1600.380 652.060 1604.000 ;
        RECT 651.780 1600.000 652.120 1600.380 ;
        RECT 651.980 1589.150 652.120 1600.000 ;
        RECT 651.920 1588.830 652.180 1589.150 ;
        RECT 654.220 1588.830 654.480 1589.150 ;
        RECT 654.280 32.630 654.420 1588.830 ;
        RECT 654.220 32.310 654.480 32.630 ;
        RECT 870.880 32.310 871.140 32.630 ;
        RECT 870.940 2.400 871.080 32.310 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 657.870 1589.060 658.190 1589.120 ;
        RECT 661.090 1589.060 661.410 1589.120 ;
        RECT 657.870 1588.920 661.410 1589.060 ;
        RECT 657.870 1588.860 658.190 1588.920 ;
        RECT 661.090 1588.860 661.410 1588.920 ;
        RECT 661.090 32.200 661.410 32.260 ;
        RECT 888.790 32.200 889.110 32.260 ;
        RECT 661.090 32.060 889.110 32.200 ;
        RECT 661.090 32.000 661.410 32.060 ;
        RECT 888.790 32.000 889.110 32.060 ;
      LAYER via ;
        RECT 657.900 1588.860 658.160 1589.120 ;
        RECT 661.120 1588.860 661.380 1589.120 ;
        RECT 661.120 32.000 661.380 32.260 ;
        RECT 888.820 32.000 889.080 32.260 ;
      LAYER met2 ;
        RECT 657.760 1600.380 658.040 1604.000 ;
        RECT 657.760 1600.000 658.100 1600.380 ;
        RECT 657.960 1589.150 658.100 1600.000 ;
        RECT 657.900 1588.830 658.160 1589.150 ;
        RECT 661.120 1588.830 661.380 1589.150 ;
        RECT 661.180 32.290 661.320 1588.830 ;
        RECT 661.120 31.970 661.380 32.290 ;
        RECT 888.820 31.970 889.080 32.290 ;
        RECT 888.880 2.400 889.020 31.970 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 664.310 1590.080 664.630 1590.140 ;
        RECT 668.910 1590.080 669.230 1590.140 ;
        RECT 664.310 1589.940 669.230 1590.080 ;
        RECT 664.310 1589.880 664.630 1589.940 ;
        RECT 668.910 1589.880 669.230 1589.940 ;
        RECT 668.910 31.860 669.230 31.920 ;
        RECT 906.730 31.860 907.050 31.920 ;
        RECT 668.910 31.720 907.050 31.860 ;
        RECT 668.910 31.660 669.230 31.720 ;
        RECT 906.730 31.660 907.050 31.720 ;
      LAYER via ;
        RECT 664.340 1589.880 664.600 1590.140 ;
        RECT 668.940 1589.880 669.200 1590.140 ;
        RECT 668.940 31.660 669.200 31.920 ;
        RECT 906.760 31.660 907.020 31.920 ;
      LAYER met2 ;
        RECT 664.200 1600.380 664.480 1604.000 ;
        RECT 664.200 1600.000 664.540 1600.380 ;
        RECT 664.400 1590.170 664.540 1600.000 ;
        RECT 664.340 1589.850 664.600 1590.170 ;
        RECT 668.940 1589.850 669.200 1590.170 ;
        RECT 669.000 31.950 669.140 1589.850 ;
        RECT 668.940 31.630 669.200 31.950 ;
        RECT 906.760 31.630 907.020 31.950 ;
        RECT 906.820 2.400 906.960 31.630 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 670.290 1589.060 670.610 1589.120 ;
        RECT 675.810 1589.060 676.130 1589.120 ;
        RECT 670.290 1588.920 676.130 1589.060 ;
        RECT 670.290 1588.860 670.610 1588.920 ;
        RECT 675.810 1588.860 676.130 1588.920 ;
        RECT 675.810 31.520 676.130 31.580 ;
        RECT 924.210 31.520 924.530 31.580 ;
        RECT 675.810 31.380 924.530 31.520 ;
        RECT 675.810 31.320 676.130 31.380 ;
        RECT 924.210 31.320 924.530 31.380 ;
      LAYER via ;
        RECT 670.320 1588.860 670.580 1589.120 ;
        RECT 675.840 1588.860 676.100 1589.120 ;
        RECT 675.840 31.320 676.100 31.580 ;
        RECT 924.240 31.320 924.500 31.580 ;
      LAYER met2 ;
        RECT 670.180 1600.380 670.460 1604.000 ;
        RECT 670.180 1600.000 670.520 1600.380 ;
        RECT 670.380 1589.150 670.520 1600.000 ;
        RECT 670.320 1588.830 670.580 1589.150 ;
        RECT 675.840 1588.830 676.100 1589.150 ;
        RECT 675.900 31.610 676.040 1588.830 ;
        RECT 675.840 31.290 676.100 31.610 ;
        RECT 924.240 31.290 924.500 31.610 ;
        RECT 924.300 2.400 924.440 31.290 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 676.730 1590.080 677.050 1590.140 ;
        RECT 682.710 1590.080 683.030 1590.140 ;
        RECT 676.730 1589.940 683.030 1590.080 ;
        RECT 676.730 1589.880 677.050 1589.940 ;
        RECT 682.710 1589.880 683.030 1589.940 ;
        RECT 682.710 31.180 683.030 31.240 ;
        RECT 942.150 31.180 942.470 31.240 ;
        RECT 682.710 31.040 942.470 31.180 ;
        RECT 682.710 30.980 683.030 31.040 ;
        RECT 942.150 30.980 942.470 31.040 ;
      LAYER via ;
        RECT 676.760 1589.880 677.020 1590.140 ;
        RECT 682.740 1589.880 683.000 1590.140 ;
        RECT 682.740 30.980 683.000 31.240 ;
        RECT 942.180 30.980 942.440 31.240 ;
      LAYER met2 ;
        RECT 676.620 1600.380 676.900 1604.000 ;
        RECT 676.620 1600.000 676.960 1600.380 ;
        RECT 676.820 1590.170 676.960 1600.000 ;
        RECT 676.760 1589.850 677.020 1590.170 ;
        RECT 682.740 1589.850 683.000 1590.170 ;
        RECT 682.800 31.270 682.940 1589.850 ;
        RECT 682.740 30.950 683.000 31.270 ;
        RECT 942.180 30.950 942.440 31.270 ;
        RECT 942.240 2.400 942.380 30.950 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 682.250 30.840 682.570 30.900 ;
        RECT 960.090 30.840 960.410 30.900 ;
        RECT 682.250 30.700 960.410 30.840 ;
        RECT 682.250 30.640 682.570 30.700 ;
        RECT 960.090 30.640 960.410 30.700 ;
      LAYER via ;
        RECT 682.280 30.640 682.540 30.900 ;
        RECT 960.120 30.640 960.380 30.900 ;
      LAYER met2 ;
        RECT 682.600 1600.380 682.880 1604.000 ;
        RECT 682.600 1600.000 682.940 1600.380 ;
        RECT 682.800 1590.930 682.940 1600.000 ;
        RECT 682.340 1590.790 682.940 1590.930 ;
        RECT 682.340 30.930 682.480 1590.790 ;
        RECT 682.280 30.610 682.540 30.930 ;
        RECT 960.120 30.610 960.380 30.930 ;
        RECT 960.180 2.400 960.320 30.610 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 769.650 1588.040 769.970 1588.100 ;
        RECT 755.940 1587.900 769.970 1588.040 ;
        RECT 688.690 1587.700 689.010 1587.760 ;
        RECT 755.940 1587.700 756.080 1587.900 ;
        RECT 769.650 1587.840 769.970 1587.900 ;
        RECT 688.690 1587.560 756.080 1587.700 ;
        RECT 688.690 1587.500 689.010 1587.560 ;
        RECT 769.190 15.540 769.510 15.600 ;
        RECT 978.030 15.540 978.350 15.600 ;
        RECT 769.190 15.400 978.350 15.540 ;
        RECT 769.190 15.340 769.510 15.400 ;
        RECT 978.030 15.340 978.350 15.400 ;
      LAYER via ;
        RECT 688.720 1587.500 688.980 1587.760 ;
        RECT 769.680 1587.840 769.940 1588.100 ;
        RECT 769.220 15.340 769.480 15.600 ;
        RECT 978.060 15.340 978.320 15.600 ;
      LAYER met2 ;
        RECT 688.580 1600.380 688.860 1604.000 ;
        RECT 688.580 1600.000 688.920 1600.380 ;
        RECT 688.780 1587.790 688.920 1600.000 ;
        RECT 769.680 1587.810 769.940 1588.130 ;
        RECT 688.720 1587.470 688.980 1587.790 ;
        RECT 769.740 19.450 769.880 1587.810 ;
        RECT 769.280 19.310 769.880 19.450 ;
        RECT 769.280 15.630 769.420 19.310 ;
        RECT 769.220 15.310 769.480 15.630 ;
        RECT 978.060 15.310 978.320 15.630 ;
        RECT 978.120 2.400 978.260 15.310 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 578.750 18.600 579.070 18.660 ;
        RECT 656.950 18.600 657.270 18.660 ;
        RECT 578.750 18.460 657.270 18.600 ;
        RECT 578.750 18.400 579.070 18.460 ;
        RECT 656.950 18.400 657.270 18.460 ;
      LAYER via ;
        RECT 578.780 18.400 579.040 18.660 ;
        RECT 656.980 18.400 657.240 18.660 ;
      LAYER met2 ;
        RECT 577.260 1600.450 577.540 1604.000 ;
        RECT 577.260 1600.310 578.980 1600.450 ;
        RECT 577.260 1600.000 577.540 1600.310 ;
        RECT 578.840 18.690 578.980 1600.310 ;
        RECT 578.780 18.370 579.040 18.690 ;
        RECT 656.980 18.370 657.240 18.690 ;
        RECT 657.040 2.400 657.180 18.370 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 742.125 1587.205 742.295 1589.075 ;
      LAYER mcon ;
        RECT 742.125 1588.905 742.295 1589.075 ;
      LAYER met1 ;
        RECT 742.065 1589.060 742.355 1589.105 ;
        RECT 742.065 1588.920 744.580 1589.060 ;
        RECT 742.065 1588.875 742.355 1588.920 ;
        RECT 744.440 1588.720 744.580 1588.920 ;
        RECT 776.090 1588.720 776.410 1588.780 ;
        RECT 744.440 1588.580 776.410 1588.720 ;
        RECT 776.090 1588.520 776.410 1588.580 ;
        RECT 742.065 1587.360 742.355 1587.405 ;
        RECT 737.540 1587.220 742.355 1587.360 ;
        RECT 696.050 1587.020 696.370 1587.080 ;
        RECT 737.540 1587.020 737.680 1587.220 ;
        RECT 742.065 1587.175 742.355 1587.220 ;
        RECT 696.050 1586.880 737.680 1587.020 ;
        RECT 696.050 1586.820 696.370 1586.880 ;
        RECT 776.090 18.260 776.410 18.320 ;
        RECT 995.970 18.260 996.290 18.320 ;
        RECT 776.090 18.120 996.290 18.260 ;
        RECT 776.090 18.060 776.410 18.120 ;
        RECT 995.970 18.060 996.290 18.120 ;
      LAYER via ;
        RECT 776.120 1588.520 776.380 1588.780 ;
        RECT 696.080 1586.820 696.340 1587.080 ;
        RECT 776.120 18.060 776.380 18.320 ;
        RECT 996.000 18.060 996.260 18.320 ;
      LAYER met2 ;
        RECT 695.020 1600.450 695.300 1604.000 ;
        RECT 695.020 1600.310 696.280 1600.450 ;
        RECT 695.020 1600.000 695.300 1600.310 ;
        RECT 696.140 1587.110 696.280 1600.310 ;
        RECT 776.120 1588.490 776.380 1588.810 ;
        RECT 696.080 1586.790 696.340 1587.110 ;
        RECT 776.180 18.350 776.320 1588.490 ;
        RECT 776.120 18.030 776.380 18.350 ;
        RECT 996.000 18.030 996.260 18.350 ;
        RECT 996.060 2.400 996.200 18.030 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 702.490 40.020 702.810 40.080 ;
        RECT 1013.450 40.020 1013.770 40.080 ;
        RECT 702.490 39.880 1013.770 40.020 ;
        RECT 702.490 39.820 702.810 39.880 ;
        RECT 1013.450 39.820 1013.770 39.880 ;
      LAYER via ;
        RECT 702.520 39.820 702.780 40.080 ;
        RECT 1013.480 39.820 1013.740 40.080 ;
      LAYER met2 ;
        RECT 701.000 1600.450 701.280 1604.000 ;
        RECT 701.000 1600.310 702.720 1600.450 ;
        RECT 701.000 1600.000 701.280 1600.310 ;
        RECT 702.580 40.110 702.720 1600.310 ;
        RECT 702.520 39.790 702.780 40.110 ;
        RECT 1013.480 39.790 1013.740 40.110 ;
        RECT 1013.540 2.400 1013.680 39.790 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 709.850 39.680 710.170 39.740 ;
        RECT 1031.390 39.680 1031.710 39.740 ;
        RECT 709.850 39.540 1031.710 39.680 ;
        RECT 709.850 39.480 710.170 39.540 ;
        RECT 1031.390 39.480 1031.710 39.540 ;
      LAYER via ;
        RECT 709.880 39.480 710.140 39.740 ;
        RECT 1031.420 39.480 1031.680 39.740 ;
      LAYER met2 ;
        RECT 707.440 1600.450 707.720 1604.000 ;
        RECT 707.440 1600.310 708.240 1600.450 ;
        RECT 707.440 1600.000 707.720 1600.310 ;
        RECT 708.100 1580.050 708.240 1600.310 ;
        RECT 708.100 1579.910 710.080 1580.050 ;
        RECT 709.940 39.770 710.080 1579.910 ;
        RECT 709.880 39.450 710.140 39.770 ;
        RECT 1031.420 39.450 1031.680 39.770 ;
        RECT 1031.480 2.400 1031.620 39.450 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 716.750 39.340 717.070 39.400 ;
        RECT 1049.330 39.340 1049.650 39.400 ;
        RECT 716.750 39.200 1049.650 39.340 ;
        RECT 716.750 39.140 717.070 39.200 ;
        RECT 1049.330 39.140 1049.650 39.200 ;
      LAYER via ;
        RECT 716.780 39.140 717.040 39.400 ;
        RECT 1049.360 39.140 1049.620 39.400 ;
      LAYER met2 ;
        RECT 713.420 1600.450 713.700 1604.000 ;
        RECT 713.420 1600.310 714.680 1600.450 ;
        RECT 713.420 1600.000 713.700 1600.310 ;
        RECT 714.540 1580.050 714.680 1600.310 ;
        RECT 714.540 1579.910 716.980 1580.050 ;
        RECT 716.840 39.430 716.980 1579.910 ;
        RECT 716.780 39.110 717.040 39.430 ;
        RECT 1049.360 39.110 1049.620 39.430 ;
        RECT 1049.420 2.400 1049.560 39.110 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 722.730 39.000 723.050 39.060 ;
        RECT 1067.270 39.000 1067.590 39.060 ;
        RECT 722.730 38.860 1067.590 39.000 ;
        RECT 722.730 38.800 723.050 38.860 ;
        RECT 1067.270 38.800 1067.590 38.860 ;
      LAYER via ;
        RECT 722.760 38.800 723.020 39.060 ;
        RECT 1067.300 38.800 1067.560 39.060 ;
      LAYER met2 ;
        RECT 719.860 1600.450 720.140 1604.000 ;
        RECT 719.860 1600.310 720.660 1600.450 ;
        RECT 719.860 1600.000 720.140 1600.310 ;
        RECT 720.520 1580.050 720.660 1600.310 ;
        RECT 720.520 1579.910 722.960 1580.050 ;
        RECT 722.820 39.090 722.960 1579.910 ;
        RECT 722.760 38.770 723.020 39.090 ;
        RECT 1067.300 38.770 1067.560 39.090 ;
        RECT 1067.360 2.400 1067.500 38.770 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 725.950 1587.360 726.270 1587.420 ;
        RECT 730.550 1587.360 730.870 1587.420 ;
        RECT 725.950 1587.220 730.870 1587.360 ;
        RECT 725.950 1587.160 726.270 1587.220 ;
        RECT 730.550 1587.160 730.870 1587.220 ;
        RECT 730.550 38.660 730.870 38.720 ;
        RECT 1085.210 38.660 1085.530 38.720 ;
        RECT 730.550 38.520 1085.530 38.660 ;
        RECT 730.550 38.460 730.870 38.520 ;
        RECT 1085.210 38.460 1085.530 38.520 ;
      LAYER via ;
        RECT 725.980 1587.160 726.240 1587.420 ;
        RECT 730.580 1587.160 730.840 1587.420 ;
        RECT 730.580 38.460 730.840 38.720 ;
        RECT 1085.240 38.460 1085.500 38.720 ;
      LAYER met2 ;
        RECT 725.840 1600.380 726.120 1604.000 ;
        RECT 725.840 1600.000 726.180 1600.380 ;
        RECT 726.040 1587.450 726.180 1600.000 ;
        RECT 725.980 1587.130 726.240 1587.450 ;
        RECT 730.580 1587.130 730.840 1587.450 ;
        RECT 730.640 38.750 730.780 1587.130 ;
        RECT 730.580 38.430 730.840 38.750 ;
        RECT 1085.240 38.430 1085.500 38.750 ;
        RECT 1085.300 2.400 1085.440 38.430 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 732.390 1587.360 732.710 1587.420 ;
        RECT 736.990 1587.360 737.310 1587.420 ;
        RECT 732.390 1587.220 737.310 1587.360 ;
        RECT 732.390 1587.160 732.710 1587.220 ;
        RECT 736.990 1587.160 737.310 1587.220 ;
        RECT 737.450 38.320 737.770 38.380 ;
        RECT 1102.690 38.320 1103.010 38.380 ;
        RECT 737.450 38.180 1103.010 38.320 ;
        RECT 737.450 38.120 737.770 38.180 ;
        RECT 1102.690 38.120 1103.010 38.180 ;
      LAYER via ;
        RECT 732.420 1587.160 732.680 1587.420 ;
        RECT 737.020 1587.160 737.280 1587.420 ;
        RECT 737.480 38.120 737.740 38.380 ;
        RECT 1102.720 38.120 1102.980 38.380 ;
      LAYER met2 ;
        RECT 732.280 1600.380 732.560 1604.000 ;
        RECT 732.280 1600.000 732.620 1600.380 ;
        RECT 732.480 1587.450 732.620 1600.000 ;
        RECT 732.420 1587.130 732.680 1587.450 ;
        RECT 737.020 1587.130 737.280 1587.450 ;
        RECT 737.080 1579.370 737.220 1587.130 ;
        RECT 737.080 1579.230 737.680 1579.370 ;
        RECT 737.540 38.410 737.680 1579.230 ;
        RECT 737.480 38.090 737.740 38.410 ;
        RECT 1102.720 38.090 1102.980 38.410 ;
        RECT 1102.780 2.400 1102.920 38.090 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 738.370 1588.720 738.690 1588.780 ;
        RECT 743.890 1588.720 744.210 1588.780 ;
        RECT 738.370 1588.580 744.210 1588.720 ;
        RECT 738.370 1588.520 738.690 1588.580 ;
        RECT 743.890 1588.520 744.210 1588.580 ;
        RECT 743.890 37.980 744.210 38.040 ;
        RECT 1120.630 37.980 1120.950 38.040 ;
        RECT 743.890 37.840 1120.950 37.980 ;
        RECT 743.890 37.780 744.210 37.840 ;
        RECT 1120.630 37.780 1120.950 37.840 ;
      LAYER via ;
        RECT 738.400 1588.520 738.660 1588.780 ;
        RECT 743.920 1588.520 744.180 1588.780 ;
        RECT 743.920 37.780 744.180 38.040 ;
        RECT 1120.660 37.780 1120.920 38.040 ;
      LAYER met2 ;
        RECT 738.260 1600.380 738.540 1604.000 ;
        RECT 738.260 1600.000 738.600 1600.380 ;
        RECT 738.460 1588.810 738.600 1600.000 ;
        RECT 738.400 1588.490 738.660 1588.810 ;
        RECT 743.920 1588.490 744.180 1588.810 ;
        RECT 743.980 38.070 744.120 1588.490 ;
        RECT 743.920 37.750 744.180 38.070 ;
        RECT 1120.660 37.750 1120.920 38.070 ;
        RECT 1120.720 2.400 1120.860 37.750 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 744.350 27.100 744.670 27.160 ;
        RECT 1138.570 27.100 1138.890 27.160 ;
        RECT 744.350 26.960 1138.890 27.100 ;
        RECT 744.350 26.900 744.670 26.960 ;
        RECT 1138.570 26.900 1138.890 26.960 ;
      LAYER via ;
        RECT 744.380 26.900 744.640 27.160 ;
        RECT 1138.600 26.900 1138.860 27.160 ;
      LAYER met2 ;
        RECT 744.240 1600.380 744.520 1604.000 ;
        RECT 744.240 1600.000 744.580 1600.380 ;
        RECT 744.440 27.190 744.580 1600.000 ;
        RECT 744.380 26.870 744.640 27.190 ;
        RECT 1138.600 26.870 1138.860 27.190 ;
        RECT 1138.660 2.400 1138.800 26.870 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 751.710 26.420 752.030 26.480 ;
        RECT 1156.510 26.420 1156.830 26.480 ;
        RECT 751.710 26.280 1156.830 26.420 ;
        RECT 751.710 26.220 752.030 26.280 ;
        RECT 1156.510 26.220 1156.830 26.280 ;
      LAYER via ;
        RECT 751.740 26.220 752.000 26.480 ;
        RECT 1156.540 26.220 1156.800 26.480 ;
      LAYER met2 ;
        RECT 750.680 1600.450 750.960 1604.000 ;
        RECT 750.680 1600.310 751.940 1600.450 ;
        RECT 750.680 1600.000 750.960 1600.310 ;
        RECT 751.800 26.510 751.940 1600.310 ;
        RECT 751.740 26.190 752.000 26.510 ;
        RECT 1156.540 26.190 1156.800 26.510 ;
        RECT 1156.600 2.400 1156.740 26.190 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 585.190 15.200 585.510 15.260 ;
        RECT 674.430 15.200 674.750 15.260 ;
        RECT 585.190 15.060 674.750 15.200 ;
        RECT 585.190 15.000 585.510 15.060 ;
        RECT 674.430 15.000 674.750 15.060 ;
      LAYER via ;
        RECT 585.220 15.000 585.480 15.260 ;
        RECT 674.460 15.000 674.720 15.260 ;
      LAYER met2 ;
        RECT 583.700 1600.450 583.980 1604.000 ;
        RECT 583.700 1600.310 584.500 1600.450 ;
        RECT 583.700 1600.000 583.980 1600.310 ;
        RECT 584.360 1590.250 584.500 1600.310 ;
        RECT 584.360 1590.110 585.420 1590.250 ;
        RECT 585.280 15.290 585.420 1590.110 ;
        RECT 585.220 14.970 585.480 15.290 ;
        RECT 674.460 14.970 674.720 15.290 ;
        RECT 674.520 2.400 674.660 14.970 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 758.610 25.740 758.930 25.800 ;
        RECT 1173.990 25.740 1174.310 25.800 ;
        RECT 758.610 25.600 1174.310 25.740 ;
        RECT 758.610 25.540 758.930 25.600 ;
        RECT 1173.990 25.540 1174.310 25.600 ;
      LAYER via ;
        RECT 758.640 25.540 758.900 25.800 ;
        RECT 1174.020 25.540 1174.280 25.800 ;
      LAYER met2 ;
        RECT 756.660 1600.450 756.940 1604.000 ;
        RECT 756.660 1600.310 758.380 1600.450 ;
        RECT 756.660 1600.000 756.940 1600.310 ;
        RECT 758.240 1580.050 758.380 1600.310 ;
        RECT 758.240 1579.910 758.840 1580.050 ;
        RECT 758.700 25.830 758.840 1579.910 ;
        RECT 758.640 25.510 758.900 25.830 ;
        RECT 1174.020 25.510 1174.280 25.830 ;
        RECT 1174.080 2.400 1174.220 25.510 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 764.590 43.760 764.910 43.820 ;
        RECT 1191.930 43.760 1192.250 43.820 ;
        RECT 764.590 43.620 1192.250 43.760 ;
        RECT 764.590 43.560 764.910 43.620 ;
        RECT 1191.930 43.560 1192.250 43.620 ;
      LAYER via ;
        RECT 764.620 43.560 764.880 43.820 ;
        RECT 1191.960 43.560 1192.220 43.820 ;
      LAYER met2 ;
        RECT 763.100 1600.450 763.380 1604.000 ;
        RECT 763.100 1600.310 764.360 1600.450 ;
        RECT 763.100 1600.000 763.380 1600.310 ;
        RECT 764.220 1580.050 764.360 1600.310 ;
        RECT 764.220 1579.910 764.820 1580.050 ;
        RECT 764.680 43.850 764.820 1579.910 ;
        RECT 764.620 43.530 764.880 43.850 ;
        RECT 1191.960 43.530 1192.220 43.850 ;
        RECT 1192.020 2.400 1192.160 43.530 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 769.190 1591.780 769.510 1591.840 ;
        RECT 771.490 1591.780 771.810 1591.840 ;
        RECT 769.190 1591.640 771.810 1591.780 ;
        RECT 769.190 1591.580 769.510 1591.640 ;
        RECT 771.490 1591.580 771.810 1591.640 ;
        RECT 771.490 44.440 771.810 44.500 ;
        RECT 771.490 44.300 1193.080 44.440 ;
        RECT 771.490 44.240 771.810 44.300 ;
        RECT 1192.940 43.760 1193.080 44.300 ;
        RECT 1209.870 43.760 1210.190 43.820 ;
        RECT 1192.940 43.620 1210.190 43.760 ;
        RECT 1209.870 43.560 1210.190 43.620 ;
      LAYER via ;
        RECT 769.220 1591.580 769.480 1591.840 ;
        RECT 771.520 1591.580 771.780 1591.840 ;
        RECT 771.520 44.240 771.780 44.500 ;
        RECT 1209.900 43.560 1210.160 43.820 ;
      LAYER met2 ;
        RECT 769.080 1600.380 769.360 1604.000 ;
        RECT 769.080 1600.000 769.420 1600.380 ;
        RECT 769.280 1591.870 769.420 1600.000 ;
        RECT 769.220 1591.550 769.480 1591.870 ;
        RECT 771.520 1591.550 771.780 1591.870 ;
        RECT 771.580 44.530 771.720 1591.550 ;
        RECT 771.520 44.210 771.780 44.530 ;
        RECT 1209.900 43.530 1210.160 43.850 ;
        RECT 1209.960 2.400 1210.100 43.530 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1196.605 47.005 1196.775 47.855 ;
      LAYER mcon ;
        RECT 1196.605 47.685 1196.775 47.855 ;
      LAYER met1 ;
        RECT 775.630 1587.360 775.950 1587.420 ;
        RECT 778.850 1587.360 779.170 1587.420 ;
        RECT 775.630 1587.220 779.170 1587.360 ;
        RECT 775.630 1587.160 775.950 1587.220 ;
        RECT 778.850 1587.160 779.170 1587.220 ;
        RECT 778.850 47.840 779.170 47.900 ;
        RECT 1196.545 47.840 1196.835 47.885 ;
        RECT 778.850 47.700 1196.835 47.840 ;
        RECT 778.850 47.640 779.170 47.700 ;
        RECT 1196.545 47.655 1196.835 47.700 ;
        RECT 1227.810 47.500 1228.130 47.560 ;
        RECT 1224.680 47.360 1228.130 47.500 ;
        RECT 1196.545 47.160 1196.835 47.205 ;
        RECT 1224.680 47.160 1224.820 47.360 ;
        RECT 1227.810 47.300 1228.130 47.360 ;
        RECT 1196.545 47.020 1224.820 47.160 ;
        RECT 1196.545 46.975 1196.835 47.020 ;
      LAYER via ;
        RECT 775.660 1587.160 775.920 1587.420 ;
        RECT 778.880 1587.160 779.140 1587.420 ;
        RECT 778.880 47.640 779.140 47.900 ;
        RECT 1227.840 47.300 1228.100 47.560 ;
      LAYER met2 ;
        RECT 775.520 1600.380 775.800 1604.000 ;
        RECT 775.520 1600.000 775.860 1600.380 ;
        RECT 775.720 1587.450 775.860 1600.000 ;
        RECT 775.660 1587.130 775.920 1587.450 ;
        RECT 778.880 1587.130 779.140 1587.450 ;
        RECT 778.940 47.930 779.080 1587.130 ;
        RECT 778.880 47.610 779.140 47.930 ;
        RECT 1227.840 47.270 1228.100 47.590 ;
        RECT 1227.900 2.400 1228.040 47.270 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1196.145 44.285 1196.315 47.175 ;
      LAYER mcon ;
        RECT 1196.145 47.005 1196.315 47.175 ;
      LAYER met1 ;
        RECT 781.610 1587.360 781.930 1587.420 ;
        RECT 785.290 1587.360 785.610 1587.420 ;
        RECT 781.610 1587.220 785.610 1587.360 ;
        RECT 781.610 1587.160 781.930 1587.220 ;
        RECT 785.290 1587.160 785.610 1587.220 ;
        RECT 785.290 47.160 785.610 47.220 ;
        RECT 1196.085 47.160 1196.375 47.205 ;
        RECT 785.290 47.020 1196.375 47.160 ;
        RECT 785.290 46.960 785.610 47.020 ;
        RECT 1196.085 46.975 1196.375 47.020 ;
        RECT 1196.085 44.440 1196.375 44.485 ;
        RECT 1243.910 44.440 1244.230 44.500 ;
        RECT 1196.085 44.300 1244.230 44.440 ;
        RECT 1196.085 44.255 1196.375 44.300 ;
        RECT 1243.910 44.240 1244.230 44.300 ;
      LAYER via ;
        RECT 781.640 1587.160 781.900 1587.420 ;
        RECT 785.320 1587.160 785.580 1587.420 ;
        RECT 785.320 46.960 785.580 47.220 ;
        RECT 1243.940 44.240 1244.200 44.500 ;
      LAYER met2 ;
        RECT 781.500 1600.380 781.780 1604.000 ;
        RECT 781.500 1600.000 781.840 1600.380 ;
        RECT 781.700 1587.450 781.840 1600.000 ;
        RECT 781.640 1587.130 781.900 1587.450 ;
        RECT 785.320 1587.130 785.580 1587.450 ;
        RECT 785.380 47.250 785.520 1587.130 ;
        RECT 785.320 46.930 785.580 47.250 ;
        RECT 1244.000 44.530 1245.060 44.610 ;
        RECT 1243.940 44.470 1245.060 44.530 ;
        RECT 1243.940 44.210 1244.200 44.470 ;
        RECT 1244.920 42.570 1245.060 44.470 ;
        RECT 1244.920 42.430 1245.980 42.570 ;
        RECT 1245.840 2.400 1245.980 42.430 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1244.905 47.005 1246.455 47.175 ;
        RECT 1244.905 45.985 1245.075 47.005 ;
        RECT 1246.285 46.665 1246.455 47.005 ;
      LAYER met1 ;
        RECT 788.970 1579.540 789.290 1579.600 ;
        RECT 792.190 1579.540 792.510 1579.600 ;
        RECT 788.970 1579.400 792.510 1579.540 ;
        RECT 788.970 1579.340 789.290 1579.400 ;
        RECT 792.190 1579.340 792.510 1579.400 ;
        RECT 1246.225 46.820 1246.515 46.865 ;
        RECT 1246.225 46.680 1247.360 46.820 ;
        RECT 1246.225 46.635 1246.515 46.680 ;
        RECT 1247.220 46.480 1247.360 46.680 ;
        RECT 1263.230 46.480 1263.550 46.540 ;
        RECT 1247.220 46.340 1263.550 46.480 ;
        RECT 1263.230 46.280 1263.550 46.340 ;
        RECT 792.190 46.140 792.510 46.200 ;
        RECT 1244.845 46.140 1245.135 46.185 ;
        RECT 792.190 46.000 1245.135 46.140 ;
        RECT 792.190 45.940 792.510 46.000 ;
        RECT 1244.845 45.955 1245.135 46.000 ;
      LAYER via ;
        RECT 789.000 1579.340 789.260 1579.600 ;
        RECT 792.220 1579.340 792.480 1579.600 ;
        RECT 1263.260 46.280 1263.520 46.540 ;
        RECT 792.220 45.940 792.480 46.200 ;
      LAYER met2 ;
        RECT 787.940 1600.450 788.220 1604.000 ;
        RECT 787.940 1600.310 789.200 1600.450 ;
        RECT 787.940 1600.000 788.220 1600.310 ;
        RECT 789.060 1579.630 789.200 1600.310 ;
        RECT 789.000 1579.310 789.260 1579.630 ;
        RECT 792.220 1579.310 792.480 1579.630 ;
        RECT 792.280 46.230 792.420 1579.310 ;
        RECT 1263.260 46.250 1263.520 46.570 ;
        RECT 792.220 45.910 792.480 46.230 ;
        RECT 1263.320 2.400 1263.460 46.250 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 794.030 1587.700 794.350 1587.760 ;
        RECT 799.550 1587.700 799.870 1587.760 ;
        RECT 794.030 1587.560 799.870 1587.700 ;
        RECT 794.030 1587.500 794.350 1587.560 ;
        RECT 799.550 1587.500 799.870 1587.560 ;
        RECT 1281.170 46.140 1281.490 46.200 ;
        RECT 1245.380 46.000 1281.490 46.140 ;
        RECT 799.550 45.800 799.870 45.860 ;
        RECT 1245.380 45.800 1245.520 46.000 ;
        RECT 1281.170 45.940 1281.490 46.000 ;
        RECT 799.550 45.660 1245.520 45.800 ;
        RECT 799.550 45.600 799.870 45.660 ;
      LAYER via ;
        RECT 794.060 1587.500 794.320 1587.760 ;
        RECT 799.580 1587.500 799.840 1587.760 ;
        RECT 799.580 45.600 799.840 45.860 ;
        RECT 1281.200 45.940 1281.460 46.200 ;
      LAYER met2 ;
        RECT 793.920 1600.380 794.200 1604.000 ;
        RECT 793.920 1600.000 794.260 1600.380 ;
        RECT 794.120 1587.790 794.260 1600.000 ;
        RECT 794.060 1587.470 794.320 1587.790 ;
        RECT 799.580 1587.470 799.840 1587.790 ;
        RECT 799.640 45.890 799.780 1587.470 ;
        RECT 1281.200 45.910 1281.460 46.230 ;
        RECT 799.580 45.570 799.840 45.890 ;
        RECT 1281.260 2.400 1281.400 45.910 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1275.265 44.285 1275.435 45.815 ;
        RECT 1295.505 45.475 1295.675 45.815 ;
        RECT 1294.125 45.305 1295.675 45.475 ;
        RECT 1293.205 44.115 1293.375 44.455 ;
        RECT 1294.125 44.115 1294.295 45.305 ;
        RECT 1293.205 43.945 1294.295 44.115 ;
      LAYER mcon ;
        RECT 1275.265 45.645 1275.435 45.815 ;
        RECT 1295.505 45.645 1295.675 45.815 ;
        RECT 1293.205 44.285 1293.375 44.455 ;
      LAYER met1 ;
        RECT 1275.205 45.800 1275.495 45.845 ;
        RECT 1245.840 45.660 1275.495 45.800 ;
        RECT 799.090 45.460 799.410 45.520 ;
        RECT 1245.840 45.460 1245.980 45.660 ;
        RECT 1275.205 45.615 1275.495 45.660 ;
        RECT 1295.445 45.800 1295.735 45.845 ;
        RECT 1299.110 45.800 1299.430 45.860 ;
        RECT 1295.445 45.660 1299.430 45.800 ;
        RECT 1295.445 45.615 1295.735 45.660 ;
        RECT 1299.110 45.600 1299.430 45.660 ;
        RECT 799.090 45.320 1245.980 45.460 ;
        RECT 799.090 45.260 799.410 45.320 ;
        RECT 1275.205 44.440 1275.495 44.485 ;
        RECT 1293.145 44.440 1293.435 44.485 ;
        RECT 1275.205 44.300 1293.435 44.440 ;
        RECT 1275.205 44.255 1275.495 44.300 ;
        RECT 1293.145 44.255 1293.435 44.300 ;
      LAYER via ;
        RECT 799.120 45.260 799.380 45.520 ;
        RECT 1299.140 45.600 1299.400 45.860 ;
      LAYER met2 ;
        RECT 799.900 1600.450 800.180 1604.000 ;
        RECT 799.180 1600.310 800.180 1600.450 ;
        RECT 799.180 45.550 799.320 1600.310 ;
        RECT 799.900 1600.000 800.180 1600.310 ;
        RECT 1299.140 45.570 1299.400 45.890 ;
        RECT 799.120 45.230 799.380 45.550 ;
        RECT 1299.200 2.400 1299.340 45.570 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 806.450 34.920 806.770 34.980 ;
        RECT 1317.050 34.920 1317.370 34.980 ;
        RECT 806.450 34.780 1317.370 34.920 ;
        RECT 806.450 34.720 806.770 34.780 ;
        RECT 1317.050 34.720 1317.370 34.780 ;
      LAYER via ;
        RECT 806.480 34.720 806.740 34.980 ;
        RECT 1317.080 34.720 1317.340 34.980 ;
      LAYER met2 ;
        RECT 806.340 1600.380 806.620 1604.000 ;
        RECT 806.340 1600.000 806.680 1600.380 ;
        RECT 806.540 35.010 806.680 1600.000 ;
        RECT 806.480 34.690 806.740 35.010 ;
        RECT 1317.080 34.690 1317.340 35.010 ;
        RECT 1317.140 2.400 1317.280 34.690 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 813.350 45.120 813.670 45.180 ;
        RECT 1334.990 45.120 1335.310 45.180 ;
        RECT 813.350 44.980 1335.310 45.120 ;
        RECT 813.350 44.920 813.670 44.980 ;
        RECT 1334.990 44.920 1335.310 44.980 ;
      LAYER via ;
        RECT 813.380 44.920 813.640 45.180 ;
        RECT 1335.020 44.920 1335.280 45.180 ;
      LAYER met2 ;
        RECT 812.320 1600.450 812.600 1604.000 ;
        RECT 812.320 1600.310 813.580 1600.450 ;
        RECT 812.320 1600.000 812.600 1600.310 ;
        RECT 813.440 45.210 813.580 1600.310 ;
        RECT 813.380 44.890 813.640 45.210 ;
        RECT 1335.020 44.890 1335.280 45.210 ;
        RECT 1335.080 2.400 1335.220 44.890 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 665.305 14.705 665.475 17.255 ;
      LAYER mcon ;
        RECT 665.305 17.085 665.475 17.255 ;
      LAYER met1 ;
        RECT 593.010 17.240 593.330 17.300 ;
        RECT 665.245 17.240 665.535 17.285 ;
        RECT 593.010 17.100 665.535 17.240 ;
        RECT 593.010 17.040 593.330 17.100 ;
        RECT 665.245 17.055 665.535 17.100 ;
        RECT 665.245 14.860 665.535 14.905 ;
        RECT 692.370 14.860 692.690 14.920 ;
        RECT 665.245 14.720 692.690 14.860 ;
        RECT 665.245 14.675 665.535 14.720 ;
        RECT 692.370 14.660 692.690 14.720 ;
      LAYER via ;
        RECT 593.040 17.040 593.300 17.300 ;
        RECT 692.400 14.660 692.660 14.920 ;
      LAYER met2 ;
        RECT 589.680 1600.450 589.960 1604.000 ;
        RECT 589.680 1600.310 591.400 1600.450 ;
        RECT 589.680 1600.000 589.960 1600.310 ;
        RECT 591.260 1590.250 591.400 1600.310 ;
        RECT 591.260 1590.110 593.240 1590.250 ;
        RECT 593.100 17.330 593.240 1590.110 ;
        RECT 593.040 17.010 593.300 17.330 ;
        RECT 692.400 14.630 692.660 14.950 ;
        RECT 692.460 2.400 692.600 14.630 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 818.870 1587.700 819.190 1587.760 ;
        RECT 820.250 1587.700 820.570 1587.760 ;
        RECT 818.870 1587.560 820.570 1587.700 ;
        RECT 818.870 1587.500 819.190 1587.560 ;
        RECT 820.250 1587.500 820.570 1587.560 ;
        RECT 820.250 44.780 820.570 44.840 ;
        RECT 1352.470 44.780 1352.790 44.840 ;
        RECT 820.250 44.640 1352.790 44.780 ;
        RECT 820.250 44.580 820.570 44.640 ;
        RECT 1352.470 44.580 1352.790 44.640 ;
      LAYER via ;
        RECT 818.900 1587.500 819.160 1587.760 ;
        RECT 820.280 1587.500 820.540 1587.760 ;
        RECT 820.280 44.580 820.540 44.840 ;
        RECT 1352.500 44.580 1352.760 44.840 ;
      LAYER met2 ;
        RECT 818.760 1600.380 819.040 1604.000 ;
        RECT 818.760 1600.000 819.100 1600.380 ;
        RECT 818.960 1587.790 819.100 1600.000 ;
        RECT 818.900 1587.470 819.160 1587.790 ;
        RECT 820.280 1587.470 820.540 1587.790 ;
        RECT 820.340 44.870 820.480 1587.470 ;
        RECT 820.280 44.550 820.540 44.870 ;
        RECT 1352.500 44.550 1352.760 44.870 ;
        RECT 1352.560 2.400 1352.700 44.550 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1027.325 41.565 1028.875 41.735 ;
      LAYER mcon ;
        RECT 1028.705 41.565 1028.875 41.735 ;
      LAYER met1 ;
        RECT 824.850 1587.700 825.170 1587.760 ;
        RECT 827.610 1587.700 827.930 1587.760 ;
        RECT 824.850 1587.560 827.930 1587.700 ;
        RECT 824.850 1587.500 825.170 1587.560 ;
        RECT 827.610 1587.500 827.930 1587.560 ;
        RECT 827.610 41.720 827.930 41.780 ;
        RECT 1027.265 41.720 1027.555 41.765 ;
        RECT 827.610 41.580 1027.555 41.720 ;
        RECT 827.610 41.520 827.930 41.580 ;
        RECT 1027.265 41.535 1027.555 41.580 ;
        RECT 1028.645 41.720 1028.935 41.765 ;
        RECT 1370.410 41.720 1370.730 41.780 ;
        RECT 1028.645 41.580 1370.730 41.720 ;
        RECT 1028.645 41.535 1028.935 41.580 ;
        RECT 1370.410 41.520 1370.730 41.580 ;
      LAYER via ;
        RECT 824.880 1587.500 825.140 1587.760 ;
        RECT 827.640 1587.500 827.900 1587.760 ;
        RECT 827.640 41.520 827.900 41.780 ;
        RECT 1370.440 41.520 1370.700 41.780 ;
      LAYER met2 ;
        RECT 824.740 1600.380 825.020 1604.000 ;
        RECT 824.740 1600.000 825.080 1600.380 ;
        RECT 824.940 1587.790 825.080 1600.000 ;
        RECT 824.880 1587.470 825.140 1587.790 ;
        RECT 827.640 1587.470 827.900 1587.790 ;
        RECT 827.700 41.810 827.840 1587.470 ;
        RECT 827.640 41.490 827.900 41.810 ;
        RECT 1370.440 41.490 1370.700 41.810 ;
        RECT 1370.500 2.400 1370.640 41.490 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 831.290 1587.360 831.610 1587.420 ;
        RECT 834.050 1587.360 834.370 1587.420 ;
        RECT 831.290 1587.220 834.370 1587.360 ;
        RECT 831.290 1587.160 831.610 1587.220 ;
        RECT 834.050 1587.160 834.370 1587.220 ;
        RECT 834.050 69.260 834.370 69.320 ;
        RECT 1386.970 69.260 1387.290 69.320 ;
        RECT 834.050 69.120 1387.290 69.260 ;
        RECT 834.050 69.060 834.370 69.120 ;
        RECT 1386.970 69.060 1387.290 69.120 ;
        RECT 1386.970 2.960 1387.290 3.020 ;
        RECT 1388.350 2.960 1388.670 3.020 ;
        RECT 1386.970 2.820 1388.670 2.960 ;
        RECT 1386.970 2.760 1387.290 2.820 ;
        RECT 1388.350 2.760 1388.670 2.820 ;
      LAYER via ;
        RECT 831.320 1587.160 831.580 1587.420 ;
        RECT 834.080 1587.160 834.340 1587.420 ;
        RECT 834.080 69.060 834.340 69.320 ;
        RECT 1387.000 69.060 1387.260 69.320 ;
        RECT 1387.000 2.760 1387.260 3.020 ;
        RECT 1388.380 2.760 1388.640 3.020 ;
      LAYER met2 ;
        RECT 831.180 1600.380 831.460 1604.000 ;
        RECT 831.180 1600.000 831.520 1600.380 ;
        RECT 831.380 1587.450 831.520 1600.000 ;
        RECT 831.320 1587.130 831.580 1587.450 ;
        RECT 834.080 1587.130 834.340 1587.450 ;
        RECT 834.140 69.350 834.280 1587.130 ;
        RECT 834.080 69.030 834.340 69.350 ;
        RECT 1387.000 69.030 1387.260 69.350 ;
        RECT 1387.060 3.050 1387.200 69.030 ;
        RECT 1387.000 2.730 1387.260 3.050 ;
        RECT 1388.380 2.730 1388.640 3.050 ;
        RECT 1388.440 2.400 1388.580 2.730 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 837.270 1587.700 837.590 1587.760 ;
        RECT 841.410 1587.700 841.730 1587.760 ;
        RECT 837.270 1587.560 841.730 1587.700 ;
        RECT 837.270 1587.500 837.590 1587.560 ;
        RECT 841.410 1587.500 841.730 1587.560 ;
        RECT 841.410 69.940 841.730 70.000 ;
        RECT 1400.770 69.940 1401.090 70.000 ;
        RECT 841.410 69.800 1401.090 69.940 ;
        RECT 841.410 69.740 841.730 69.800 ;
        RECT 1400.770 69.740 1401.090 69.800 ;
        RECT 1400.770 2.960 1401.090 3.020 ;
        RECT 1406.290 2.960 1406.610 3.020 ;
        RECT 1400.770 2.820 1406.610 2.960 ;
        RECT 1400.770 2.760 1401.090 2.820 ;
        RECT 1406.290 2.760 1406.610 2.820 ;
      LAYER via ;
        RECT 837.300 1587.500 837.560 1587.760 ;
        RECT 841.440 1587.500 841.700 1587.760 ;
        RECT 841.440 69.740 841.700 70.000 ;
        RECT 1400.800 69.740 1401.060 70.000 ;
        RECT 1400.800 2.760 1401.060 3.020 ;
        RECT 1406.320 2.760 1406.580 3.020 ;
      LAYER met2 ;
        RECT 837.160 1600.380 837.440 1604.000 ;
        RECT 837.160 1600.000 837.500 1600.380 ;
        RECT 837.360 1587.790 837.500 1600.000 ;
        RECT 837.300 1587.470 837.560 1587.790 ;
        RECT 841.440 1587.470 841.700 1587.790 ;
        RECT 841.500 70.030 841.640 1587.470 ;
        RECT 841.440 69.710 841.700 70.030 ;
        RECT 1400.800 69.710 1401.060 70.030 ;
        RECT 1400.860 3.050 1401.000 69.710 ;
        RECT 1400.800 2.730 1401.060 3.050 ;
        RECT 1406.320 2.730 1406.580 3.050 ;
        RECT 1406.380 2.400 1406.520 2.730 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 843.710 1587.360 844.030 1587.420 ;
        RECT 847.850 1587.360 848.170 1587.420 ;
        RECT 843.710 1587.220 848.170 1587.360 ;
        RECT 843.710 1587.160 844.030 1587.220 ;
        RECT 847.850 1587.160 848.170 1587.220 ;
        RECT 847.850 71.300 848.170 71.360 ;
        RECT 1421.470 71.300 1421.790 71.360 ;
        RECT 847.850 71.160 1421.790 71.300 ;
        RECT 847.850 71.100 848.170 71.160 ;
        RECT 1421.470 71.100 1421.790 71.160 ;
      LAYER via ;
        RECT 843.740 1587.160 844.000 1587.420 ;
        RECT 847.880 1587.160 848.140 1587.420 ;
        RECT 847.880 71.100 848.140 71.360 ;
        RECT 1421.500 71.100 1421.760 71.360 ;
      LAYER met2 ;
        RECT 843.600 1600.380 843.880 1604.000 ;
        RECT 843.600 1600.000 843.940 1600.380 ;
        RECT 843.800 1587.450 843.940 1600.000 ;
        RECT 843.740 1587.130 844.000 1587.450 ;
        RECT 847.880 1587.130 848.140 1587.450 ;
        RECT 847.940 71.390 848.080 1587.130 ;
        RECT 847.880 71.070 848.140 71.390 ;
        RECT 1421.500 71.070 1421.760 71.390 ;
        RECT 1421.560 3.130 1421.700 71.070 ;
        RECT 1421.560 2.990 1424.000 3.130 ;
        RECT 1423.860 2.400 1424.000 2.990 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 849.690 1587.360 850.010 1587.420 ;
        RECT 854.750 1587.360 855.070 1587.420 ;
        RECT 849.690 1587.220 855.070 1587.360 ;
        RECT 849.690 1587.160 850.010 1587.220 ;
        RECT 854.750 1587.160 855.070 1587.220 ;
        RECT 854.750 71.640 855.070 71.700 ;
        RECT 1435.270 71.640 1435.590 71.700 ;
        RECT 854.750 71.500 1435.590 71.640 ;
        RECT 854.750 71.440 855.070 71.500 ;
        RECT 1435.270 71.440 1435.590 71.500 ;
        RECT 1435.270 27.780 1435.590 27.840 ;
        RECT 1441.710 27.780 1442.030 27.840 ;
        RECT 1435.270 27.640 1442.030 27.780 ;
        RECT 1435.270 27.580 1435.590 27.640 ;
        RECT 1441.710 27.580 1442.030 27.640 ;
      LAYER via ;
        RECT 849.720 1587.160 849.980 1587.420 ;
        RECT 854.780 1587.160 855.040 1587.420 ;
        RECT 854.780 71.440 855.040 71.700 ;
        RECT 1435.300 71.440 1435.560 71.700 ;
        RECT 1435.300 27.580 1435.560 27.840 ;
        RECT 1441.740 27.580 1442.000 27.840 ;
      LAYER met2 ;
        RECT 849.580 1600.380 849.860 1604.000 ;
        RECT 849.580 1600.000 849.920 1600.380 ;
        RECT 849.780 1587.450 849.920 1600.000 ;
        RECT 849.720 1587.130 849.980 1587.450 ;
        RECT 854.780 1587.130 855.040 1587.450 ;
        RECT 854.840 71.730 854.980 1587.130 ;
        RECT 854.780 71.410 855.040 71.730 ;
        RECT 1435.300 71.410 1435.560 71.730 ;
        RECT 1435.360 27.870 1435.500 71.410 ;
        RECT 1435.300 27.550 1435.560 27.870 ;
        RECT 1441.740 27.550 1442.000 27.870 ;
        RECT 1441.800 2.400 1441.940 27.550 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 856.130 1587.360 856.450 1587.420 ;
        RECT 861.190 1587.360 861.510 1587.420 ;
        RECT 856.130 1587.220 861.510 1587.360 ;
        RECT 856.130 1587.160 856.450 1587.220 ;
        RECT 861.190 1587.160 861.510 1587.220 ;
        RECT 861.190 48.520 861.510 48.580 ;
        RECT 1455.970 48.520 1456.290 48.580 ;
        RECT 861.190 48.380 1456.290 48.520 ;
        RECT 861.190 48.320 861.510 48.380 ;
        RECT 1455.970 48.320 1456.290 48.380 ;
        RECT 1455.970 2.960 1456.290 3.020 ;
        RECT 1459.650 2.960 1459.970 3.020 ;
        RECT 1455.970 2.820 1459.970 2.960 ;
        RECT 1455.970 2.760 1456.290 2.820 ;
        RECT 1459.650 2.760 1459.970 2.820 ;
      LAYER via ;
        RECT 856.160 1587.160 856.420 1587.420 ;
        RECT 861.220 1587.160 861.480 1587.420 ;
        RECT 861.220 48.320 861.480 48.580 ;
        RECT 1456.000 48.320 1456.260 48.580 ;
        RECT 1456.000 2.760 1456.260 3.020 ;
        RECT 1459.680 2.760 1459.940 3.020 ;
      LAYER met2 ;
        RECT 856.020 1600.380 856.300 1604.000 ;
        RECT 856.020 1600.000 856.360 1600.380 ;
        RECT 856.220 1587.450 856.360 1600.000 ;
        RECT 856.160 1587.130 856.420 1587.450 ;
        RECT 861.220 1587.130 861.480 1587.450 ;
        RECT 861.280 48.610 861.420 1587.130 ;
        RECT 861.220 48.290 861.480 48.610 ;
        RECT 1456.000 48.290 1456.260 48.610 ;
        RECT 1456.060 3.050 1456.200 48.290 ;
        RECT 1456.000 2.730 1456.260 3.050 ;
        RECT 1459.680 2.730 1459.940 3.050 ;
        RECT 1459.740 2.400 1459.880 2.730 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 861.650 48.860 861.970 48.920 ;
        RECT 1476.670 48.860 1476.990 48.920 ;
        RECT 861.650 48.720 1476.990 48.860 ;
        RECT 861.650 48.660 861.970 48.720 ;
        RECT 1476.670 48.660 1476.990 48.720 ;
        RECT 1476.670 2.960 1476.990 3.020 ;
        RECT 1477.590 2.960 1477.910 3.020 ;
        RECT 1476.670 2.820 1477.910 2.960 ;
        RECT 1476.670 2.760 1476.990 2.820 ;
        RECT 1477.590 2.760 1477.910 2.820 ;
      LAYER via ;
        RECT 861.680 48.660 861.940 48.920 ;
        RECT 1476.700 48.660 1476.960 48.920 ;
        RECT 1476.700 2.760 1476.960 3.020 ;
        RECT 1477.620 2.760 1477.880 3.020 ;
      LAYER met2 ;
        RECT 862.000 1600.380 862.280 1604.000 ;
        RECT 862.000 1600.000 862.340 1600.380 ;
        RECT 862.200 1588.210 862.340 1600.000 ;
        RECT 861.740 1588.070 862.340 1588.210 ;
        RECT 861.740 48.950 861.880 1588.070 ;
        RECT 861.680 48.630 861.940 48.950 ;
        RECT 1476.700 48.630 1476.960 48.950 ;
        RECT 1476.760 3.050 1476.900 48.630 ;
        RECT 1476.700 2.730 1476.960 3.050 ;
        RECT 1477.620 2.730 1477.880 3.050 ;
        RECT 1477.680 2.400 1477.820 2.730 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 868.550 49.200 868.870 49.260 ;
        RECT 1490.470 49.200 1490.790 49.260 ;
        RECT 868.550 49.060 1490.790 49.200 ;
        RECT 868.550 49.000 868.870 49.060 ;
        RECT 1490.470 49.000 1490.790 49.060 ;
        RECT 1490.470 2.960 1490.790 3.020 ;
        RECT 1495.530 2.960 1495.850 3.020 ;
        RECT 1490.470 2.820 1495.850 2.960 ;
        RECT 1490.470 2.760 1490.790 2.820 ;
        RECT 1495.530 2.760 1495.850 2.820 ;
      LAYER via ;
        RECT 868.580 49.000 868.840 49.260 ;
        RECT 1490.500 49.000 1490.760 49.260 ;
        RECT 1490.500 2.760 1490.760 3.020 ;
        RECT 1495.560 2.760 1495.820 3.020 ;
      LAYER met2 ;
        RECT 867.980 1600.450 868.260 1604.000 ;
        RECT 867.980 1600.310 868.780 1600.450 ;
        RECT 867.980 1600.000 868.260 1600.310 ;
        RECT 868.640 49.290 868.780 1600.310 ;
        RECT 868.580 48.970 868.840 49.290 ;
        RECT 1490.500 48.970 1490.760 49.290 ;
        RECT 1490.560 3.050 1490.700 48.970 ;
        RECT 1490.500 2.730 1490.760 3.050 ;
        RECT 1495.560 2.730 1495.820 3.050 ;
        RECT 1495.620 2.400 1495.760 2.730 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 874.990 49.540 875.310 49.600 ;
        RECT 1511.170 49.540 1511.490 49.600 ;
        RECT 874.990 49.400 1511.490 49.540 ;
        RECT 874.990 49.340 875.310 49.400 ;
        RECT 1511.170 49.340 1511.490 49.400 ;
      LAYER via ;
        RECT 875.020 49.340 875.280 49.600 ;
        RECT 1511.200 49.340 1511.460 49.600 ;
      LAYER met2 ;
        RECT 874.420 1600.450 874.700 1604.000 ;
        RECT 874.420 1600.310 875.220 1600.450 ;
        RECT 874.420 1600.000 874.700 1600.310 ;
        RECT 875.080 49.630 875.220 1600.310 ;
        RECT 875.020 49.310 875.280 49.630 ;
        RECT 1511.200 49.310 1511.460 49.630 ;
        RECT 1511.260 3.130 1511.400 49.310 ;
        RECT 1511.260 2.990 1513.240 3.130 ;
        RECT 1513.100 2.400 1513.240 2.990 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 596.230 1590.420 596.550 1590.480 ;
        RECT 599.450 1590.420 599.770 1590.480 ;
        RECT 596.230 1590.280 599.770 1590.420 ;
        RECT 596.230 1590.220 596.550 1590.280 ;
        RECT 599.450 1590.220 599.770 1590.280 ;
        RECT 599.450 15.540 599.770 15.600 ;
        RECT 710.310 15.540 710.630 15.600 ;
        RECT 599.450 15.400 710.630 15.540 ;
        RECT 599.450 15.340 599.770 15.400 ;
        RECT 710.310 15.340 710.630 15.400 ;
      LAYER via ;
        RECT 596.260 1590.220 596.520 1590.480 ;
        RECT 599.480 1590.220 599.740 1590.480 ;
        RECT 599.480 15.340 599.740 15.600 ;
        RECT 710.340 15.340 710.600 15.600 ;
      LAYER met2 ;
        RECT 596.120 1600.380 596.400 1604.000 ;
        RECT 596.120 1600.000 596.460 1600.380 ;
        RECT 596.320 1590.510 596.460 1600.000 ;
        RECT 596.260 1590.190 596.520 1590.510 ;
        RECT 599.480 1590.190 599.740 1590.510 ;
        RECT 599.540 15.630 599.680 1590.190 ;
        RECT 599.480 15.310 599.740 15.630 ;
        RECT 710.340 15.310 710.600 15.630 ;
        RECT 710.400 2.400 710.540 15.310 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 881.890 49.880 882.210 49.940 ;
        RECT 1524.970 49.880 1525.290 49.940 ;
        RECT 881.890 49.740 1525.290 49.880 ;
        RECT 881.890 49.680 882.210 49.740 ;
        RECT 1524.970 49.680 1525.290 49.740 ;
        RECT 1524.970 16.900 1525.290 16.960 ;
        RECT 1530.950 16.900 1531.270 16.960 ;
        RECT 1524.970 16.760 1531.270 16.900 ;
        RECT 1524.970 16.700 1525.290 16.760 ;
        RECT 1530.950 16.700 1531.270 16.760 ;
      LAYER via ;
        RECT 881.920 49.680 882.180 49.940 ;
        RECT 1525.000 49.680 1525.260 49.940 ;
        RECT 1525.000 16.700 1525.260 16.960 ;
        RECT 1530.980 16.700 1531.240 16.960 ;
      LAYER met2 ;
        RECT 880.400 1600.450 880.680 1604.000 ;
        RECT 880.400 1600.310 882.120 1600.450 ;
        RECT 880.400 1600.000 880.680 1600.310 ;
        RECT 881.980 49.970 882.120 1600.310 ;
        RECT 881.920 49.650 882.180 49.970 ;
        RECT 1525.000 49.650 1525.260 49.970 ;
        RECT 1525.060 16.990 1525.200 49.650 ;
        RECT 1525.000 16.670 1525.260 16.990 ;
        RECT 1530.980 16.670 1531.240 16.990 ;
        RECT 1531.040 2.400 1531.180 16.670 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 886.950 1587.700 887.270 1587.760 ;
        RECT 889.250 1587.700 889.570 1587.760 ;
        RECT 886.950 1587.560 889.570 1587.700 ;
        RECT 886.950 1587.500 887.270 1587.560 ;
        RECT 889.250 1587.500 889.570 1587.560 ;
        RECT 889.250 50.220 889.570 50.280 ;
        RECT 1545.670 50.220 1545.990 50.280 ;
        RECT 889.250 50.080 1545.990 50.220 ;
        RECT 889.250 50.020 889.570 50.080 ;
        RECT 1545.670 50.020 1545.990 50.080 ;
        RECT 1545.670 2.960 1545.990 3.020 ;
        RECT 1548.890 2.960 1549.210 3.020 ;
        RECT 1545.670 2.820 1549.210 2.960 ;
        RECT 1545.670 2.760 1545.990 2.820 ;
        RECT 1548.890 2.760 1549.210 2.820 ;
      LAYER via ;
        RECT 886.980 1587.500 887.240 1587.760 ;
        RECT 889.280 1587.500 889.540 1587.760 ;
        RECT 889.280 50.020 889.540 50.280 ;
        RECT 1545.700 50.020 1545.960 50.280 ;
        RECT 1545.700 2.760 1545.960 3.020 ;
        RECT 1548.920 2.760 1549.180 3.020 ;
      LAYER met2 ;
        RECT 886.840 1600.380 887.120 1604.000 ;
        RECT 886.840 1600.000 887.180 1600.380 ;
        RECT 887.040 1587.790 887.180 1600.000 ;
        RECT 886.980 1587.470 887.240 1587.790 ;
        RECT 889.280 1587.470 889.540 1587.790 ;
        RECT 889.340 50.310 889.480 1587.470 ;
        RECT 889.280 49.990 889.540 50.310 ;
        RECT 1545.700 49.990 1545.960 50.310 ;
        RECT 1545.760 3.050 1545.900 49.990 ;
        RECT 1545.700 2.730 1545.960 3.050 ;
        RECT 1548.920 2.730 1549.180 3.050 ;
        RECT 1548.980 2.400 1549.120 2.730 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 892.930 1587.700 893.250 1587.760 ;
        RECT 895.230 1587.700 895.550 1587.760 ;
        RECT 892.930 1587.560 895.550 1587.700 ;
        RECT 892.930 1587.500 893.250 1587.560 ;
        RECT 895.230 1587.500 895.550 1587.560 ;
        RECT 895.690 50.560 896.010 50.620 ;
        RECT 1566.830 50.560 1567.150 50.620 ;
        RECT 895.690 50.420 1567.150 50.560 ;
        RECT 895.690 50.360 896.010 50.420 ;
        RECT 1566.830 50.360 1567.150 50.420 ;
      LAYER via ;
        RECT 892.960 1587.500 893.220 1587.760 ;
        RECT 895.260 1587.500 895.520 1587.760 ;
        RECT 895.720 50.360 895.980 50.620 ;
        RECT 1566.860 50.360 1567.120 50.620 ;
      LAYER met2 ;
        RECT 892.820 1600.380 893.100 1604.000 ;
        RECT 892.820 1600.000 893.160 1600.380 ;
        RECT 893.020 1587.790 893.160 1600.000 ;
        RECT 892.960 1587.470 893.220 1587.790 ;
        RECT 895.260 1587.470 895.520 1587.790 ;
        RECT 895.320 1578.690 895.460 1587.470 ;
        RECT 895.320 1578.550 895.920 1578.690 ;
        RECT 895.780 50.650 895.920 1578.550 ;
        RECT 895.720 50.330 895.980 50.650 ;
        RECT 1566.860 50.330 1567.120 50.650 ;
        RECT 1566.920 2.400 1567.060 50.330 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 899.370 1587.360 899.690 1587.420 ;
        RECT 902.590 1587.360 902.910 1587.420 ;
        RECT 899.370 1587.220 902.910 1587.360 ;
        RECT 899.370 1587.160 899.690 1587.220 ;
        RECT 902.590 1587.160 902.910 1587.220 ;
        RECT 902.590 50.900 902.910 50.960 ;
        RECT 1580.170 50.900 1580.490 50.960 ;
        RECT 902.590 50.760 1580.490 50.900 ;
        RECT 902.590 50.700 902.910 50.760 ;
        RECT 1580.170 50.700 1580.490 50.760 ;
        RECT 1580.170 2.960 1580.490 3.020 ;
        RECT 1584.770 2.960 1585.090 3.020 ;
        RECT 1580.170 2.820 1585.090 2.960 ;
        RECT 1580.170 2.760 1580.490 2.820 ;
        RECT 1584.770 2.760 1585.090 2.820 ;
      LAYER via ;
        RECT 899.400 1587.160 899.660 1587.420 ;
        RECT 902.620 1587.160 902.880 1587.420 ;
        RECT 902.620 50.700 902.880 50.960 ;
        RECT 1580.200 50.700 1580.460 50.960 ;
        RECT 1580.200 2.760 1580.460 3.020 ;
        RECT 1584.800 2.760 1585.060 3.020 ;
      LAYER met2 ;
        RECT 899.260 1600.380 899.540 1604.000 ;
        RECT 899.260 1600.000 899.600 1600.380 ;
        RECT 899.460 1587.450 899.600 1600.000 ;
        RECT 899.400 1587.130 899.660 1587.450 ;
        RECT 902.620 1587.130 902.880 1587.450 ;
        RECT 902.680 50.990 902.820 1587.130 ;
        RECT 902.620 50.670 902.880 50.990 ;
        RECT 1580.200 50.670 1580.460 50.990 ;
        RECT 1580.260 3.050 1580.400 50.670 ;
        RECT 1580.200 2.730 1580.460 3.050 ;
        RECT 1584.800 2.730 1585.060 3.050 ;
        RECT 1584.860 2.400 1585.000 2.730 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 905.350 1587.360 905.670 1587.420 ;
        RECT 908.110 1587.360 908.430 1587.420 ;
        RECT 905.350 1587.220 908.430 1587.360 ;
        RECT 905.350 1587.160 905.670 1587.220 ;
        RECT 908.110 1587.160 908.430 1587.220 ;
        RECT 909.490 51.240 909.810 51.300 ;
        RECT 1600.870 51.240 1601.190 51.300 ;
        RECT 909.490 51.100 1601.190 51.240 ;
        RECT 909.490 51.040 909.810 51.100 ;
        RECT 1600.870 51.040 1601.190 51.100 ;
      LAYER via ;
        RECT 905.380 1587.160 905.640 1587.420 ;
        RECT 908.140 1587.160 908.400 1587.420 ;
        RECT 909.520 51.040 909.780 51.300 ;
        RECT 1600.900 51.040 1601.160 51.300 ;
      LAYER met2 ;
        RECT 905.240 1600.380 905.520 1604.000 ;
        RECT 905.240 1600.000 905.580 1600.380 ;
        RECT 905.440 1587.450 905.580 1600.000 ;
        RECT 905.380 1587.130 905.640 1587.450 ;
        RECT 908.140 1587.130 908.400 1587.450 ;
        RECT 908.200 1579.370 908.340 1587.130 ;
        RECT 908.200 1579.230 909.720 1579.370 ;
        RECT 909.580 51.330 909.720 1579.230 ;
        RECT 909.520 51.010 909.780 51.330 ;
        RECT 1600.900 51.010 1601.160 51.330 ;
        RECT 1600.960 3.130 1601.100 51.010 ;
        RECT 1600.960 2.990 1602.480 3.130 ;
        RECT 1602.340 2.400 1602.480 2.990 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 911.790 1587.360 912.110 1587.420 ;
        RECT 915.930 1587.360 916.250 1587.420 ;
        RECT 911.790 1587.220 916.250 1587.360 ;
        RECT 911.790 1587.160 912.110 1587.220 ;
        RECT 915.930 1587.160 916.250 1587.220 ;
        RECT 916.850 54.980 917.170 55.040 ;
        RECT 1614.670 54.980 1614.990 55.040 ;
        RECT 916.850 54.840 1614.990 54.980 ;
        RECT 916.850 54.780 917.170 54.840 ;
        RECT 1614.670 54.780 1614.990 54.840 ;
        RECT 1614.670 2.960 1614.990 3.020 ;
        RECT 1620.190 2.960 1620.510 3.020 ;
        RECT 1614.670 2.820 1620.510 2.960 ;
        RECT 1614.670 2.760 1614.990 2.820 ;
        RECT 1620.190 2.760 1620.510 2.820 ;
      LAYER via ;
        RECT 911.820 1587.160 912.080 1587.420 ;
        RECT 915.960 1587.160 916.220 1587.420 ;
        RECT 916.880 54.780 917.140 55.040 ;
        RECT 1614.700 54.780 1614.960 55.040 ;
        RECT 1614.700 2.760 1614.960 3.020 ;
        RECT 1620.220 2.760 1620.480 3.020 ;
      LAYER met2 ;
        RECT 911.680 1600.380 911.960 1604.000 ;
        RECT 911.680 1600.000 912.020 1600.380 ;
        RECT 911.880 1587.450 912.020 1600.000 ;
        RECT 911.820 1587.130 912.080 1587.450 ;
        RECT 915.960 1587.130 916.220 1587.450 ;
        RECT 916.020 1579.370 916.160 1587.130 ;
        RECT 916.020 1579.230 917.080 1579.370 ;
        RECT 916.940 55.070 917.080 1579.230 ;
        RECT 916.880 54.750 917.140 55.070 ;
        RECT 1614.700 54.750 1614.960 55.070 ;
        RECT 1614.760 3.050 1614.900 54.750 ;
        RECT 1614.700 2.730 1614.960 3.050 ;
        RECT 1620.220 2.730 1620.480 3.050 ;
        RECT 1620.280 2.400 1620.420 2.730 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 917.770 1587.700 918.090 1587.760 ;
        RECT 923.290 1587.700 923.610 1587.760 ;
        RECT 917.770 1587.560 923.610 1587.700 ;
        RECT 917.770 1587.500 918.090 1587.560 ;
        RECT 923.290 1587.500 923.610 1587.560 ;
        RECT 923.290 54.640 923.610 54.700 ;
        RECT 1635.370 54.640 1635.690 54.700 ;
        RECT 923.290 54.500 1635.690 54.640 ;
        RECT 923.290 54.440 923.610 54.500 ;
        RECT 1635.370 54.440 1635.690 54.500 ;
        RECT 1635.370 2.960 1635.690 3.020 ;
        RECT 1638.130 2.960 1638.450 3.020 ;
        RECT 1635.370 2.820 1638.450 2.960 ;
        RECT 1635.370 2.760 1635.690 2.820 ;
        RECT 1638.130 2.760 1638.450 2.820 ;
      LAYER via ;
        RECT 917.800 1587.500 918.060 1587.760 ;
        RECT 923.320 1587.500 923.580 1587.760 ;
        RECT 923.320 54.440 923.580 54.700 ;
        RECT 1635.400 54.440 1635.660 54.700 ;
        RECT 1635.400 2.760 1635.660 3.020 ;
        RECT 1638.160 2.760 1638.420 3.020 ;
      LAYER met2 ;
        RECT 917.660 1600.380 917.940 1604.000 ;
        RECT 917.660 1600.000 918.000 1600.380 ;
        RECT 917.860 1587.790 918.000 1600.000 ;
        RECT 917.800 1587.470 918.060 1587.790 ;
        RECT 923.320 1587.470 923.580 1587.790 ;
        RECT 923.380 54.730 923.520 1587.470 ;
        RECT 923.320 54.410 923.580 54.730 ;
        RECT 1635.400 54.410 1635.660 54.730 ;
        RECT 1635.460 3.050 1635.600 54.410 ;
        RECT 1635.400 2.730 1635.660 3.050 ;
        RECT 1638.160 2.730 1638.420 3.050 ;
        RECT 1638.220 2.400 1638.360 2.730 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 922.830 54.300 923.150 54.360 ;
        RECT 1656.530 54.300 1656.850 54.360 ;
        RECT 922.830 54.160 1656.850 54.300 ;
        RECT 922.830 54.100 923.150 54.160 ;
        RECT 1656.530 54.100 1656.850 54.160 ;
      LAYER via ;
        RECT 922.860 54.100 923.120 54.360 ;
        RECT 1656.560 54.100 1656.820 54.360 ;
      LAYER met2 ;
        RECT 923.640 1600.450 923.920 1604.000 ;
        RECT 922.920 1600.310 923.920 1600.450 ;
        RECT 922.920 54.390 923.060 1600.310 ;
        RECT 923.640 1600.000 923.920 1600.310 ;
        RECT 922.860 54.070 923.120 54.390 ;
        RECT 1656.560 54.070 1656.820 54.390 ;
        RECT 1656.620 3.130 1656.760 54.070 ;
        RECT 1656.160 2.990 1656.760 3.130 ;
        RECT 1656.160 2.400 1656.300 2.990 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 930.650 53.960 930.970 54.020 ;
        RECT 1669.870 53.960 1670.190 54.020 ;
        RECT 930.650 53.820 1670.190 53.960 ;
        RECT 930.650 53.760 930.970 53.820 ;
        RECT 1669.870 53.760 1670.190 53.820 ;
        RECT 1669.870 2.960 1670.190 3.020 ;
        RECT 1673.550 2.960 1673.870 3.020 ;
        RECT 1669.870 2.820 1673.870 2.960 ;
        RECT 1669.870 2.760 1670.190 2.820 ;
        RECT 1673.550 2.760 1673.870 2.820 ;
      LAYER via ;
        RECT 930.680 53.760 930.940 54.020 ;
        RECT 1669.900 53.760 1670.160 54.020 ;
        RECT 1669.900 2.760 1670.160 3.020 ;
        RECT 1673.580 2.760 1673.840 3.020 ;
      LAYER met2 ;
        RECT 930.080 1600.450 930.360 1604.000 ;
        RECT 930.080 1600.310 930.880 1600.450 ;
        RECT 930.080 1600.000 930.360 1600.310 ;
        RECT 930.740 54.050 930.880 1600.310 ;
        RECT 930.680 53.730 930.940 54.050 ;
        RECT 1669.900 53.730 1670.160 54.050 ;
        RECT 1669.960 3.050 1670.100 53.730 ;
        RECT 1669.900 2.730 1670.160 3.050 ;
        RECT 1673.580 2.730 1673.840 3.050 ;
        RECT 1673.640 2.400 1673.780 2.730 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 937.090 53.620 937.410 53.680 ;
        RECT 1690.570 53.620 1690.890 53.680 ;
        RECT 937.090 53.480 1690.890 53.620 ;
        RECT 937.090 53.420 937.410 53.480 ;
        RECT 1690.570 53.420 1690.890 53.480 ;
      LAYER via ;
        RECT 937.120 53.420 937.380 53.680 ;
        RECT 1690.600 53.420 1690.860 53.680 ;
      LAYER met2 ;
        RECT 936.060 1600.450 936.340 1604.000 ;
        RECT 936.060 1600.310 937.320 1600.450 ;
        RECT 936.060 1600.000 936.340 1600.310 ;
        RECT 937.180 53.710 937.320 1600.310 ;
        RECT 937.120 53.390 937.380 53.710 ;
        RECT 1690.600 53.390 1690.860 53.710 ;
        RECT 1690.660 3.130 1690.800 53.390 ;
        RECT 1690.660 2.990 1691.720 3.130 ;
        RECT 1691.580 2.400 1691.720 2.990 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 602.210 1588.040 602.530 1588.100 ;
        RECT 606.810 1588.040 607.130 1588.100 ;
        RECT 602.210 1587.900 607.130 1588.040 ;
        RECT 602.210 1587.840 602.530 1587.900 ;
        RECT 606.810 1587.840 607.130 1587.900 ;
        RECT 727.790 20.640 728.110 20.700 ;
        RECT 638.180 20.500 728.110 20.640 ;
        RECT 606.810 19.620 607.130 19.680 ;
        RECT 638.180 19.620 638.320 20.500 ;
        RECT 727.790 20.440 728.110 20.500 ;
        RECT 606.810 19.480 638.320 19.620 ;
        RECT 606.810 19.420 607.130 19.480 ;
      LAYER via ;
        RECT 602.240 1587.840 602.500 1588.100 ;
        RECT 606.840 1587.840 607.100 1588.100 ;
        RECT 606.840 19.420 607.100 19.680 ;
        RECT 727.820 20.440 728.080 20.700 ;
      LAYER met2 ;
        RECT 602.100 1600.380 602.380 1604.000 ;
        RECT 602.100 1600.000 602.440 1600.380 ;
        RECT 602.300 1588.130 602.440 1600.000 ;
        RECT 602.240 1587.810 602.500 1588.130 ;
        RECT 606.840 1587.810 607.100 1588.130 ;
        RECT 606.900 19.710 607.040 1587.810 ;
        RECT 727.820 20.410 728.080 20.730 ;
        RECT 606.840 19.390 607.100 19.710 ;
        RECT 727.880 16.730 728.020 20.410 ;
        RECT 727.880 16.590 728.480 16.730 ;
        RECT 728.340 2.400 728.480 16.590 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 943.990 53.280 944.310 53.340 ;
        RECT 1704.370 53.280 1704.690 53.340 ;
        RECT 943.990 53.140 1704.690 53.280 ;
        RECT 943.990 53.080 944.310 53.140 ;
        RECT 1704.370 53.080 1704.690 53.140 ;
        RECT 1704.370 2.960 1704.690 3.020 ;
        RECT 1709.430 2.960 1709.750 3.020 ;
        RECT 1704.370 2.820 1709.750 2.960 ;
        RECT 1704.370 2.760 1704.690 2.820 ;
        RECT 1709.430 2.760 1709.750 2.820 ;
      LAYER via ;
        RECT 944.020 53.080 944.280 53.340 ;
        RECT 1704.400 53.080 1704.660 53.340 ;
        RECT 1704.400 2.760 1704.660 3.020 ;
        RECT 1709.460 2.760 1709.720 3.020 ;
      LAYER met2 ;
        RECT 942.500 1600.450 942.780 1604.000 ;
        RECT 942.500 1600.310 943.300 1600.450 ;
        RECT 942.500 1600.000 942.780 1600.310 ;
        RECT 943.160 1580.050 943.300 1600.310 ;
        RECT 943.160 1579.910 944.220 1580.050 ;
        RECT 944.080 53.370 944.220 1579.910 ;
        RECT 944.020 53.050 944.280 53.370 ;
        RECT 1704.400 53.050 1704.660 53.370 ;
        RECT 1704.460 3.050 1704.600 53.050 ;
        RECT 1704.400 2.730 1704.660 3.050 ;
        RECT 1709.460 2.730 1709.720 3.050 ;
        RECT 1709.520 2.400 1709.660 2.730 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 948.590 1588.380 948.910 1588.440 ;
        RECT 951.350 1588.380 951.670 1588.440 ;
        RECT 948.590 1588.240 951.670 1588.380 ;
        RECT 948.590 1588.180 948.910 1588.240 ;
        RECT 951.350 1588.180 951.670 1588.240 ;
        RECT 951.350 52.940 951.670 53.000 ;
        RECT 1725.070 52.940 1725.390 53.000 ;
        RECT 951.350 52.800 1725.390 52.940 ;
        RECT 951.350 52.740 951.670 52.800 ;
        RECT 1725.070 52.740 1725.390 52.800 ;
      LAYER via ;
        RECT 948.620 1588.180 948.880 1588.440 ;
        RECT 951.380 1588.180 951.640 1588.440 ;
        RECT 951.380 52.740 951.640 53.000 ;
        RECT 1725.100 52.740 1725.360 53.000 ;
      LAYER met2 ;
        RECT 948.480 1600.380 948.760 1604.000 ;
        RECT 948.480 1600.000 948.820 1600.380 ;
        RECT 948.680 1588.470 948.820 1600.000 ;
        RECT 948.620 1588.150 948.880 1588.470 ;
        RECT 951.380 1588.150 951.640 1588.470 ;
        RECT 951.440 53.030 951.580 1588.150 ;
        RECT 951.380 52.710 951.640 53.030 ;
        RECT 1725.100 52.710 1725.360 53.030 ;
        RECT 1725.160 21.490 1725.300 52.710 ;
        RECT 1725.160 21.350 1727.140 21.490 ;
        RECT 1727.000 3.130 1727.140 21.350 ;
        RECT 1727.000 2.990 1727.600 3.130 ;
        RECT 1727.460 2.400 1727.600 2.990 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 955.030 1588.380 955.350 1588.440 ;
        RECT 957.790 1588.380 958.110 1588.440 ;
        RECT 955.030 1588.240 958.110 1588.380 ;
        RECT 955.030 1588.180 955.350 1588.240 ;
        RECT 957.790 1588.180 958.110 1588.240 ;
        RECT 957.790 52.600 958.110 52.660 ;
        RECT 1738.870 52.600 1739.190 52.660 ;
        RECT 957.790 52.460 1739.190 52.600 ;
        RECT 957.790 52.400 958.110 52.460 ;
        RECT 1738.870 52.400 1739.190 52.460 ;
        RECT 1738.870 16.560 1739.190 16.620 ;
        RECT 1745.310 16.560 1745.630 16.620 ;
        RECT 1738.870 16.420 1745.630 16.560 ;
        RECT 1738.870 16.360 1739.190 16.420 ;
        RECT 1745.310 16.360 1745.630 16.420 ;
      LAYER via ;
        RECT 955.060 1588.180 955.320 1588.440 ;
        RECT 957.820 1588.180 958.080 1588.440 ;
        RECT 957.820 52.400 958.080 52.660 ;
        RECT 1738.900 52.400 1739.160 52.660 ;
        RECT 1738.900 16.360 1739.160 16.620 ;
        RECT 1745.340 16.360 1745.600 16.620 ;
      LAYER met2 ;
        RECT 954.920 1600.380 955.200 1604.000 ;
        RECT 954.920 1600.000 955.260 1600.380 ;
        RECT 955.120 1588.470 955.260 1600.000 ;
        RECT 955.060 1588.150 955.320 1588.470 ;
        RECT 957.820 1588.150 958.080 1588.470 ;
        RECT 957.880 52.690 958.020 1588.150 ;
        RECT 957.820 52.370 958.080 52.690 ;
        RECT 1738.900 52.370 1739.160 52.690 ;
        RECT 1738.960 16.650 1739.100 52.370 ;
        RECT 1738.900 16.330 1739.160 16.650 ;
        RECT 1745.340 16.330 1745.600 16.650 ;
        RECT 1745.400 2.400 1745.540 16.330 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 961.010 1587.360 961.330 1587.420 ;
        RECT 964.690 1587.360 965.010 1587.420 ;
        RECT 961.010 1587.220 965.010 1587.360 ;
        RECT 961.010 1587.160 961.330 1587.220 ;
        RECT 964.690 1587.160 965.010 1587.220 ;
        RECT 964.690 52.260 965.010 52.320 ;
        RECT 1759.570 52.260 1759.890 52.320 ;
        RECT 964.690 52.120 1759.890 52.260 ;
        RECT 964.690 52.060 965.010 52.120 ;
        RECT 1759.570 52.060 1759.890 52.120 ;
        RECT 1759.570 2.960 1759.890 3.020 ;
        RECT 1762.790 2.960 1763.110 3.020 ;
        RECT 1759.570 2.820 1763.110 2.960 ;
        RECT 1759.570 2.760 1759.890 2.820 ;
        RECT 1762.790 2.760 1763.110 2.820 ;
      LAYER via ;
        RECT 961.040 1587.160 961.300 1587.420 ;
        RECT 964.720 1587.160 964.980 1587.420 ;
        RECT 964.720 52.060 964.980 52.320 ;
        RECT 1759.600 52.060 1759.860 52.320 ;
        RECT 1759.600 2.760 1759.860 3.020 ;
        RECT 1762.820 2.760 1763.080 3.020 ;
      LAYER met2 ;
        RECT 960.900 1600.380 961.180 1604.000 ;
        RECT 960.900 1600.000 961.240 1600.380 ;
        RECT 961.100 1587.450 961.240 1600.000 ;
        RECT 961.040 1587.130 961.300 1587.450 ;
        RECT 964.720 1587.130 964.980 1587.450 ;
        RECT 964.780 52.350 964.920 1587.130 ;
        RECT 964.720 52.030 964.980 52.350 ;
        RECT 1759.600 52.030 1759.860 52.350 ;
        RECT 1759.660 3.050 1759.800 52.030 ;
        RECT 1759.600 2.730 1759.860 3.050 ;
        RECT 1762.820 2.730 1763.080 3.050 ;
        RECT 1762.880 2.400 1763.020 2.730 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 967.450 1587.360 967.770 1587.420 ;
        RECT 971.590 1587.360 971.910 1587.420 ;
        RECT 967.450 1587.220 971.910 1587.360 ;
        RECT 967.450 1587.160 967.770 1587.220 ;
        RECT 971.590 1587.160 971.910 1587.220 ;
        RECT 971.590 51.920 971.910 51.980 ;
        RECT 1780.730 51.920 1781.050 51.980 ;
        RECT 971.590 51.780 1781.050 51.920 ;
        RECT 971.590 51.720 971.910 51.780 ;
        RECT 1780.730 51.720 1781.050 51.780 ;
      LAYER via ;
        RECT 967.480 1587.160 967.740 1587.420 ;
        RECT 971.620 1587.160 971.880 1587.420 ;
        RECT 971.620 51.720 971.880 51.980 ;
        RECT 1780.760 51.720 1781.020 51.980 ;
      LAYER met2 ;
        RECT 967.340 1600.380 967.620 1604.000 ;
        RECT 967.340 1600.000 967.680 1600.380 ;
        RECT 967.540 1587.450 967.680 1600.000 ;
        RECT 967.480 1587.130 967.740 1587.450 ;
        RECT 971.620 1587.130 971.880 1587.450 ;
        RECT 971.680 52.010 971.820 1587.130 ;
        RECT 971.620 51.690 971.880 52.010 ;
        RECT 1780.760 51.690 1781.020 52.010 ;
        RECT 1780.820 2.400 1780.960 51.690 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 973.430 1588.380 973.750 1588.440 ;
        RECT 978.950 1588.380 979.270 1588.440 ;
        RECT 973.430 1588.240 979.270 1588.380 ;
        RECT 973.430 1588.180 973.750 1588.240 ;
        RECT 978.950 1588.180 979.270 1588.240 ;
        RECT 978.950 51.580 979.270 51.640 ;
        RECT 1794.070 51.580 1794.390 51.640 ;
        RECT 978.950 51.440 1794.390 51.580 ;
        RECT 978.950 51.380 979.270 51.440 ;
        RECT 1794.070 51.380 1794.390 51.440 ;
        RECT 1794.070 2.960 1794.390 3.020 ;
        RECT 1798.670 2.960 1798.990 3.020 ;
        RECT 1794.070 2.820 1798.990 2.960 ;
        RECT 1794.070 2.760 1794.390 2.820 ;
        RECT 1798.670 2.760 1798.990 2.820 ;
      LAYER via ;
        RECT 973.460 1588.180 973.720 1588.440 ;
        RECT 978.980 1588.180 979.240 1588.440 ;
        RECT 978.980 51.380 979.240 51.640 ;
        RECT 1794.100 51.380 1794.360 51.640 ;
        RECT 1794.100 2.760 1794.360 3.020 ;
        RECT 1798.700 2.760 1798.960 3.020 ;
      LAYER met2 ;
        RECT 973.320 1600.380 973.600 1604.000 ;
        RECT 973.320 1600.000 973.660 1600.380 ;
        RECT 973.520 1588.470 973.660 1600.000 ;
        RECT 973.460 1588.150 973.720 1588.470 ;
        RECT 978.980 1588.150 979.240 1588.470 ;
        RECT 979.040 51.670 979.180 1588.150 ;
        RECT 978.980 51.350 979.240 51.670 ;
        RECT 1794.100 51.350 1794.360 51.670 ;
        RECT 1794.160 3.050 1794.300 51.350 ;
        RECT 1794.100 2.730 1794.360 3.050 ;
        RECT 1798.700 2.730 1798.960 3.050 ;
        RECT 1798.760 2.400 1798.900 2.730 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 979.300 1600.450 979.580 1604.000 ;
        RECT 978.580 1600.310 979.580 1600.450 ;
        RECT 978.580 54.245 978.720 1600.310 ;
        RECT 979.300 1600.000 979.580 1600.310 ;
        RECT 978.510 53.875 978.790 54.245 ;
        RECT 1814.790 53.875 1815.070 54.245 ;
        RECT 1814.860 3.130 1815.000 53.875 ;
        RECT 1814.860 2.990 1816.840 3.130 ;
        RECT 1816.700 2.400 1816.840 2.990 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
      LAYER via2 ;
        RECT 978.510 53.920 978.790 54.200 ;
        RECT 1814.790 53.920 1815.070 54.200 ;
      LAYER met3 ;
        RECT 978.485 54.210 978.815 54.225 ;
        RECT 1814.765 54.210 1815.095 54.225 ;
        RECT 978.485 53.910 1815.095 54.210 ;
        RECT 978.485 53.895 978.815 53.910 ;
        RECT 1814.765 53.895 1815.095 53.910 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1828.570 15.880 1828.890 15.940 ;
        RECT 1834.550 15.880 1834.870 15.940 ;
        RECT 1828.570 15.740 1834.870 15.880 ;
        RECT 1828.570 15.680 1828.890 15.740 ;
        RECT 1834.550 15.680 1834.870 15.740 ;
      LAYER via ;
        RECT 1828.600 15.680 1828.860 15.940 ;
        RECT 1834.580 15.680 1834.840 15.940 ;
      LAYER met2 ;
        RECT 985.740 1600.380 986.020 1604.000 ;
        RECT 985.740 1600.000 986.080 1600.380 ;
        RECT 985.940 1589.570 986.080 1600.000 ;
        RECT 985.480 1589.430 986.080 1589.570 ;
        RECT 985.480 53.565 985.620 1589.430 ;
        RECT 985.410 53.195 985.690 53.565 ;
        RECT 1828.590 53.195 1828.870 53.565 ;
        RECT 1828.660 15.970 1828.800 53.195 ;
        RECT 1828.600 15.650 1828.860 15.970 ;
        RECT 1834.580 15.650 1834.840 15.970 ;
        RECT 1834.640 2.400 1834.780 15.650 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
      LAYER via2 ;
        RECT 985.410 53.240 985.690 53.520 ;
        RECT 1828.590 53.240 1828.870 53.520 ;
      LAYER met3 ;
        RECT 985.385 53.530 985.715 53.545 ;
        RECT 1828.565 53.530 1828.895 53.545 ;
        RECT 985.385 53.230 1828.895 53.530 ;
        RECT 985.385 53.215 985.715 53.230 ;
        RECT 1828.565 53.215 1828.895 53.230 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1849.270 2.960 1849.590 3.020 ;
        RECT 1852.030 2.960 1852.350 3.020 ;
        RECT 1849.270 2.820 1852.350 2.960 ;
        RECT 1849.270 2.760 1849.590 2.820 ;
        RECT 1852.030 2.760 1852.350 2.820 ;
      LAYER via ;
        RECT 1849.300 2.760 1849.560 3.020 ;
        RECT 1852.060 2.760 1852.320 3.020 ;
      LAYER met2 ;
        RECT 991.720 1600.450 992.000 1604.000 ;
        RECT 991.720 1600.310 992.980 1600.450 ;
        RECT 991.720 1600.000 992.000 1600.310 ;
        RECT 992.840 52.885 992.980 1600.310 ;
        RECT 992.770 52.515 993.050 52.885 ;
        RECT 1849.290 52.515 1849.570 52.885 ;
        RECT 1849.360 3.050 1849.500 52.515 ;
        RECT 1849.300 2.730 1849.560 3.050 ;
        RECT 1852.060 2.730 1852.320 3.050 ;
        RECT 1852.120 2.400 1852.260 2.730 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
      LAYER via2 ;
        RECT 992.770 52.560 993.050 52.840 ;
        RECT 1849.290 52.560 1849.570 52.840 ;
      LAYER met3 ;
        RECT 992.745 52.850 993.075 52.865 ;
        RECT 1849.265 52.850 1849.595 52.865 ;
        RECT 992.745 52.550 1849.595 52.850 ;
        RECT 992.745 52.535 993.075 52.550 ;
        RECT 1849.265 52.535 1849.595 52.550 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 998.160 1600.450 998.440 1604.000 ;
        RECT 998.160 1600.310 999.420 1600.450 ;
        RECT 998.160 1600.000 998.440 1600.310 ;
        RECT 999.280 52.205 999.420 1600.310 ;
        RECT 999.210 51.835 999.490 52.205 ;
        RECT 1870.450 51.835 1870.730 52.205 ;
        RECT 1870.520 3.130 1870.660 51.835 ;
        RECT 1870.060 2.990 1870.660 3.130 ;
        RECT 1870.060 2.400 1870.200 2.990 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
      LAYER via2 ;
        RECT 999.210 51.880 999.490 52.160 ;
        RECT 1870.450 51.880 1870.730 52.160 ;
      LAYER met3 ;
        RECT 999.185 52.170 999.515 52.185 ;
        RECT 1870.425 52.170 1870.755 52.185 ;
        RECT 999.185 51.870 1870.755 52.170 ;
        RECT 999.185 51.855 999.515 51.870 ;
        RECT 1870.425 51.855 1870.755 51.870 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 638.625 18.105 638.795 19.635 ;
      LAYER mcon ;
        RECT 638.625 19.465 638.795 19.635 ;
      LAYER met1 ;
        RECT 608.650 1590.420 608.970 1590.480 ;
        RECT 612.790 1590.420 613.110 1590.480 ;
        RECT 608.650 1590.280 613.110 1590.420 ;
        RECT 608.650 1590.220 608.970 1590.280 ;
        RECT 612.790 1590.220 613.110 1590.280 ;
        RECT 638.565 19.620 638.855 19.665 ;
        RECT 746.190 19.620 746.510 19.680 ;
        RECT 638.565 19.480 746.510 19.620 ;
        RECT 638.565 19.435 638.855 19.480 ;
        RECT 746.190 19.420 746.510 19.480 ;
        RECT 638.565 18.260 638.855 18.305 ;
        RECT 617.020 18.120 638.855 18.260 ;
        RECT 612.790 17.580 613.110 17.640 ;
        RECT 617.020 17.580 617.160 18.120 ;
        RECT 638.565 18.075 638.855 18.120 ;
        RECT 612.790 17.440 617.160 17.580 ;
        RECT 612.790 17.380 613.110 17.440 ;
      LAYER via ;
        RECT 608.680 1590.220 608.940 1590.480 ;
        RECT 612.820 1590.220 613.080 1590.480 ;
        RECT 746.220 19.420 746.480 19.680 ;
        RECT 612.820 17.380 613.080 17.640 ;
      LAYER met2 ;
        RECT 608.540 1600.380 608.820 1604.000 ;
        RECT 608.540 1600.000 608.880 1600.380 ;
        RECT 608.740 1590.510 608.880 1600.000 ;
        RECT 608.680 1590.190 608.940 1590.510 ;
        RECT 612.820 1590.190 613.080 1590.510 ;
        RECT 612.880 17.670 613.020 1590.190 ;
        RECT 746.220 19.390 746.480 19.710 ;
        RECT 612.820 17.350 613.080 17.670 ;
        RECT 746.280 2.400 746.420 19.390 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1883.770 2.960 1884.090 3.020 ;
        RECT 1887.910 2.960 1888.230 3.020 ;
        RECT 1883.770 2.820 1888.230 2.960 ;
        RECT 1883.770 2.760 1884.090 2.820 ;
        RECT 1887.910 2.760 1888.230 2.820 ;
      LAYER via ;
        RECT 1883.800 2.760 1884.060 3.020 ;
        RECT 1887.940 2.760 1888.200 3.020 ;
      LAYER met2 ;
        RECT 1004.140 1600.450 1004.420 1604.000 ;
        RECT 1004.140 1600.310 1005.860 1600.450 ;
        RECT 1004.140 1600.000 1004.420 1600.310 ;
        RECT 1005.720 1588.210 1005.860 1600.310 ;
        RECT 1005.720 1588.070 1006.780 1588.210 ;
        RECT 1006.640 51.525 1006.780 1588.070 ;
        RECT 1006.570 51.155 1006.850 51.525 ;
        RECT 1883.790 51.155 1884.070 51.525 ;
        RECT 1883.860 3.050 1884.000 51.155 ;
        RECT 1883.800 2.730 1884.060 3.050 ;
        RECT 1887.940 2.730 1888.200 3.050 ;
        RECT 1888.000 2.400 1888.140 2.730 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
      LAYER via2 ;
        RECT 1006.570 51.200 1006.850 51.480 ;
        RECT 1883.790 51.200 1884.070 51.480 ;
      LAYER met3 ;
        RECT 1006.545 51.490 1006.875 51.505 ;
        RECT 1883.765 51.490 1884.095 51.505 ;
        RECT 1006.545 51.190 1884.095 51.490 ;
        RECT 1006.545 51.175 1006.875 51.190 ;
        RECT 1883.765 51.175 1884.095 51.190 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1010.690 1593.480 1011.010 1593.540 ;
        RECT 1013.450 1593.480 1013.770 1593.540 ;
        RECT 1010.690 1593.340 1013.770 1593.480 ;
        RECT 1010.690 1593.280 1011.010 1593.340 ;
        RECT 1013.450 1593.280 1013.770 1593.340 ;
        RECT 1013.450 75.040 1013.770 75.100 ;
        RECT 1904.470 75.040 1904.790 75.100 ;
        RECT 1013.450 74.900 1904.790 75.040 ;
        RECT 1013.450 74.840 1013.770 74.900 ;
        RECT 1904.470 74.840 1904.790 74.900 ;
      LAYER via ;
        RECT 1010.720 1593.280 1010.980 1593.540 ;
        RECT 1013.480 1593.280 1013.740 1593.540 ;
        RECT 1013.480 74.840 1013.740 75.100 ;
        RECT 1904.500 74.840 1904.760 75.100 ;
      LAYER met2 ;
        RECT 1010.580 1600.380 1010.860 1604.000 ;
        RECT 1010.580 1600.000 1010.920 1600.380 ;
        RECT 1010.780 1593.570 1010.920 1600.000 ;
        RECT 1010.720 1593.250 1010.980 1593.570 ;
        RECT 1013.480 1593.250 1013.740 1593.570 ;
        RECT 1013.540 75.130 1013.680 1593.250 ;
        RECT 1013.480 74.810 1013.740 75.130 ;
        RECT 1904.500 74.810 1904.760 75.130 ;
        RECT 1904.560 3.130 1904.700 74.810 ;
        RECT 1904.560 2.990 1906.080 3.130 ;
        RECT 1905.940 2.400 1906.080 2.990 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1016.670 1590.080 1016.990 1590.140 ;
        RECT 1019.430 1590.080 1019.750 1590.140 ;
        RECT 1016.670 1589.940 1019.750 1590.080 ;
        RECT 1016.670 1589.880 1016.990 1589.940 ;
        RECT 1019.430 1589.880 1019.750 1589.940 ;
        RECT 1019.430 74.700 1019.750 74.760 ;
        RECT 1918.270 74.700 1918.590 74.760 ;
        RECT 1019.430 74.560 1918.590 74.700 ;
        RECT 1019.430 74.500 1019.750 74.560 ;
        RECT 1918.270 74.500 1918.590 74.560 ;
      LAYER via ;
        RECT 1016.700 1589.880 1016.960 1590.140 ;
        RECT 1019.460 1589.880 1019.720 1590.140 ;
        RECT 1019.460 74.500 1019.720 74.760 ;
        RECT 1918.300 74.500 1918.560 74.760 ;
      LAYER met2 ;
        RECT 1016.560 1600.380 1016.840 1604.000 ;
        RECT 1016.560 1600.000 1016.900 1600.380 ;
        RECT 1016.760 1590.170 1016.900 1600.000 ;
        RECT 1016.700 1589.850 1016.960 1590.170 ;
        RECT 1019.460 1589.850 1019.720 1590.170 ;
        RECT 1019.520 74.790 1019.660 1589.850 ;
        RECT 1019.460 74.470 1019.720 74.790 ;
        RECT 1918.300 74.470 1918.560 74.790 ;
        RECT 1918.360 16.730 1918.500 74.470 ;
        RECT 1918.360 16.590 1923.560 16.730 ;
        RECT 1923.420 2.400 1923.560 16.590 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1023.110 1587.360 1023.430 1587.420 ;
        RECT 1027.250 1587.360 1027.570 1587.420 ;
        RECT 1023.110 1587.220 1027.570 1587.360 ;
        RECT 1023.110 1587.160 1023.430 1587.220 ;
        RECT 1027.250 1587.160 1027.570 1587.220 ;
        RECT 1027.250 74.360 1027.570 74.420 ;
        RECT 1938.970 74.360 1939.290 74.420 ;
        RECT 1027.250 74.220 1939.290 74.360 ;
        RECT 1027.250 74.160 1027.570 74.220 ;
        RECT 1938.970 74.160 1939.290 74.220 ;
      LAYER via ;
        RECT 1023.140 1587.160 1023.400 1587.420 ;
        RECT 1027.280 1587.160 1027.540 1587.420 ;
        RECT 1027.280 74.160 1027.540 74.420 ;
        RECT 1939.000 74.160 1939.260 74.420 ;
      LAYER met2 ;
        RECT 1023.000 1600.380 1023.280 1604.000 ;
        RECT 1023.000 1600.000 1023.340 1600.380 ;
        RECT 1023.200 1587.450 1023.340 1600.000 ;
        RECT 1023.140 1587.130 1023.400 1587.450 ;
        RECT 1027.280 1587.130 1027.540 1587.450 ;
        RECT 1027.340 74.450 1027.480 1587.130 ;
        RECT 1027.280 74.130 1027.540 74.450 ;
        RECT 1939.000 74.130 1939.260 74.450 ;
        RECT 1939.060 16.730 1939.200 74.130 ;
        RECT 1939.060 16.590 1941.500 16.730 ;
        RECT 1941.360 2.400 1941.500 16.590 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1029.090 1587.360 1029.410 1587.420 ;
        RECT 1033.690 1587.360 1034.010 1587.420 ;
        RECT 1029.090 1587.220 1034.010 1587.360 ;
        RECT 1029.090 1587.160 1029.410 1587.220 ;
        RECT 1033.690 1587.160 1034.010 1587.220 ;
        RECT 1034.150 73.680 1034.470 73.740 ;
        RECT 1952.770 73.680 1953.090 73.740 ;
        RECT 1034.150 73.540 1953.090 73.680 ;
        RECT 1034.150 73.480 1034.470 73.540 ;
        RECT 1952.770 73.480 1953.090 73.540 ;
        RECT 1952.770 18.600 1953.090 18.660 ;
        RECT 1959.210 18.600 1959.530 18.660 ;
        RECT 1952.770 18.460 1959.530 18.600 ;
        RECT 1952.770 18.400 1953.090 18.460 ;
        RECT 1959.210 18.400 1959.530 18.460 ;
      LAYER via ;
        RECT 1029.120 1587.160 1029.380 1587.420 ;
        RECT 1033.720 1587.160 1033.980 1587.420 ;
        RECT 1034.180 73.480 1034.440 73.740 ;
        RECT 1952.800 73.480 1953.060 73.740 ;
        RECT 1952.800 18.400 1953.060 18.660 ;
        RECT 1959.240 18.400 1959.500 18.660 ;
      LAYER met2 ;
        RECT 1028.980 1600.380 1029.260 1604.000 ;
        RECT 1028.980 1600.000 1029.320 1600.380 ;
        RECT 1029.180 1587.450 1029.320 1600.000 ;
        RECT 1029.120 1587.130 1029.380 1587.450 ;
        RECT 1033.720 1587.130 1033.980 1587.450 ;
        RECT 1033.780 1579.370 1033.920 1587.130 ;
        RECT 1033.780 1579.230 1034.380 1579.370 ;
        RECT 1034.240 73.770 1034.380 1579.230 ;
        RECT 1034.180 73.450 1034.440 73.770 ;
        RECT 1952.800 73.450 1953.060 73.770 ;
        RECT 1952.860 18.690 1953.000 73.450 ;
        RECT 1952.800 18.370 1953.060 18.690 ;
        RECT 1959.240 18.370 1959.500 18.690 ;
        RECT 1959.300 2.400 1959.440 18.370 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1035.070 1587.360 1035.390 1587.420 ;
        RECT 1040.130 1587.360 1040.450 1587.420 ;
        RECT 1035.070 1587.220 1040.450 1587.360 ;
        RECT 1035.070 1587.160 1035.390 1587.220 ;
        RECT 1040.130 1587.160 1040.450 1587.220 ;
        RECT 1040.590 56.000 1040.910 56.060 ;
        RECT 1973.470 56.000 1973.790 56.060 ;
        RECT 1040.590 55.860 1973.790 56.000 ;
        RECT 1040.590 55.800 1040.910 55.860 ;
        RECT 1973.470 55.800 1973.790 55.860 ;
        RECT 1973.470 2.960 1973.790 3.020 ;
        RECT 1977.150 2.960 1977.470 3.020 ;
        RECT 1973.470 2.820 1977.470 2.960 ;
        RECT 1973.470 2.760 1973.790 2.820 ;
        RECT 1977.150 2.760 1977.470 2.820 ;
      LAYER via ;
        RECT 1035.100 1587.160 1035.360 1587.420 ;
        RECT 1040.160 1587.160 1040.420 1587.420 ;
        RECT 1040.620 55.800 1040.880 56.060 ;
        RECT 1973.500 55.800 1973.760 56.060 ;
        RECT 1973.500 2.760 1973.760 3.020 ;
        RECT 1977.180 2.760 1977.440 3.020 ;
      LAYER met2 ;
        RECT 1034.960 1600.380 1035.240 1604.000 ;
        RECT 1034.960 1600.000 1035.300 1600.380 ;
        RECT 1035.160 1587.450 1035.300 1600.000 ;
        RECT 1035.100 1587.130 1035.360 1587.450 ;
        RECT 1040.160 1587.130 1040.420 1587.450 ;
        RECT 1040.220 1579.370 1040.360 1587.130 ;
        RECT 1040.220 1579.230 1040.820 1579.370 ;
        RECT 1040.680 56.090 1040.820 1579.230 ;
        RECT 1040.620 55.770 1040.880 56.090 ;
        RECT 1973.500 55.770 1973.760 56.090 ;
        RECT 1973.560 3.050 1973.700 55.770 ;
        RECT 1973.500 2.730 1973.760 3.050 ;
        RECT 1977.180 2.730 1977.440 3.050 ;
        RECT 1977.240 2.400 1977.380 2.730 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1039.210 1590.420 1039.530 1590.480 ;
        RECT 1041.510 1590.420 1041.830 1590.480 ;
        RECT 1039.210 1590.280 1041.830 1590.420 ;
        RECT 1039.210 1590.220 1039.530 1590.280 ;
        RECT 1041.510 1590.220 1041.830 1590.280 ;
        RECT 1040.130 56.340 1040.450 56.400 ;
        RECT 1994.170 56.340 1994.490 56.400 ;
        RECT 1040.130 56.200 1994.490 56.340 ;
        RECT 1040.130 56.140 1040.450 56.200 ;
        RECT 1994.170 56.140 1994.490 56.200 ;
      LAYER via ;
        RECT 1039.240 1590.220 1039.500 1590.480 ;
        RECT 1041.540 1590.220 1041.800 1590.480 ;
        RECT 1040.160 56.140 1040.420 56.400 ;
        RECT 1994.200 56.140 1994.460 56.400 ;
      LAYER met2 ;
        RECT 1041.400 1600.380 1041.680 1604.000 ;
        RECT 1041.400 1600.000 1041.740 1600.380 ;
        RECT 1041.600 1590.510 1041.740 1600.000 ;
        RECT 1039.240 1590.190 1039.500 1590.510 ;
        RECT 1041.540 1590.190 1041.800 1590.510 ;
        RECT 1039.300 1578.690 1039.440 1590.190 ;
        RECT 1039.300 1578.550 1040.360 1578.690 ;
        RECT 1040.220 56.430 1040.360 1578.550 ;
        RECT 1040.160 56.110 1040.420 56.430 ;
        RECT 1994.200 56.110 1994.460 56.430 ;
        RECT 1994.260 3.130 1994.400 56.110 ;
        RECT 1994.260 2.990 1995.320 3.130 ;
        RECT 1995.180 2.400 1995.320 2.990 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1047.950 56.680 1048.270 56.740 ;
        RECT 2007.970 56.680 2008.290 56.740 ;
        RECT 1047.950 56.540 2008.290 56.680 ;
        RECT 1047.950 56.480 1048.270 56.540 ;
        RECT 2007.970 56.480 2008.290 56.540 ;
        RECT 2007.970 2.960 2008.290 3.020 ;
        RECT 2012.570 2.960 2012.890 3.020 ;
        RECT 2007.970 2.820 2012.890 2.960 ;
        RECT 2007.970 2.760 2008.290 2.820 ;
        RECT 2012.570 2.760 2012.890 2.820 ;
      LAYER via ;
        RECT 1047.980 56.480 1048.240 56.740 ;
        RECT 2008.000 56.480 2008.260 56.740 ;
        RECT 2008.000 2.760 2008.260 3.020 ;
        RECT 2012.600 2.760 2012.860 3.020 ;
      LAYER met2 ;
        RECT 1047.380 1600.450 1047.660 1604.000 ;
        RECT 1047.380 1600.310 1048.180 1600.450 ;
        RECT 1047.380 1600.000 1047.660 1600.310 ;
        RECT 1048.040 56.770 1048.180 1600.310 ;
        RECT 1047.980 56.450 1048.240 56.770 ;
        RECT 2008.000 56.450 2008.260 56.770 ;
        RECT 2008.060 3.050 2008.200 56.450 ;
        RECT 2008.000 2.730 2008.260 3.050 ;
        RECT 2012.600 2.730 2012.860 3.050 ;
        RECT 2012.660 2.400 2012.800 2.730 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1054.850 57.020 1055.170 57.080 ;
        RECT 2028.670 57.020 2028.990 57.080 ;
        RECT 1054.850 56.880 2028.990 57.020 ;
        RECT 1054.850 56.820 1055.170 56.880 ;
        RECT 2028.670 56.820 2028.990 56.880 ;
        RECT 2028.670 2.960 2028.990 3.020 ;
        RECT 2030.510 2.960 2030.830 3.020 ;
        RECT 2028.670 2.820 2030.830 2.960 ;
        RECT 2028.670 2.760 2028.990 2.820 ;
        RECT 2030.510 2.760 2030.830 2.820 ;
      LAYER via ;
        RECT 1054.880 56.820 1055.140 57.080 ;
        RECT 2028.700 56.820 2028.960 57.080 ;
        RECT 2028.700 2.760 2028.960 3.020 ;
        RECT 2030.540 2.760 2030.800 3.020 ;
      LAYER met2 ;
        RECT 1053.820 1600.450 1054.100 1604.000 ;
        RECT 1053.820 1600.310 1055.080 1600.450 ;
        RECT 1053.820 1600.000 1054.100 1600.310 ;
        RECT 1054.940 57.110 1055.080 1600.310 ;
        RECT 1054.880 56.790 1055.140 57.110 ;
        RECT 2028.700 56.790 2028.960 57.110 ;
        RECT 2028.760 3.050 2028.900 56.790 ;
        RECT 2028.700 2.730 2028.960 3.050 ;
        RECT 2030.540 2.730 2030.800 3.050 ;
        RECT 2030.600 2.400 2030.740 2.730 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1061.750 57.360 1062.070 57.420 ;
        RECT 2042.470 57.360 2042.790 57.420 ;
        RECT 1061.750 57.220 2042.790 57.360 ;
        RECT 1061.750 57.160 1062.070 57.220 ;
        RECT 2042.470 57.160 2042.790 57.220 ;
        RECT 2042.470 18.260 2042.790 18.320 ;
        RECT 2048.450 18.260 2048.770 18.320 ;
        RECT 2042.470 18.120 2048.770 18.260 ;
        RECT 2042.470 18.060 2042.790 18.120 ;
        RECT 2048.450 18.060 2048.770 18.120 ;
      LAYER via ;
        RECT 1061.780 57.160 1062.040 57.420 ;
        RECT 2042.500 57.160 2042.760 57.420 ;
        RECT 2042.500 18.060 2042.760 18.320 ;
        RECT 2048.480 18.060 2048.740 18.320 ;
      LAYER met2 ;
        RECT 1059.800 1600.450 1060.080 1604.000 ;
        RECT 1059.800 1600.310 1061.520 1600.450 ;
        RECT 1059.800 1600.000 1060.080 1600.310 ;
        RECT 1061.380 1580.050 1061.520 1600.310 ;
        RECT 1061.380 1579.910 1061.980 1580.050 ;
        RECT 1061.840 57.450 1061.980 1579.910 ;
        RECT 1061.780 57.130 1062.040 57.450 ;
        RECT 2042.500 57.130 2042.760 57.450 ;
        RECT 2042.560 18.350 2042.700 57.130 ;
        RECT 2042.500 18.030 2042.760 18.350 ;
        RECT 2048.480 18.030 2048.740 18.350 ;
        RECT 2048.540 2.400 2048.680 18.030 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 637.705 15.895 637.875 17.595 ;
        RECT 639.545 15.895 639.715 16.235 ;
        RECT 637.705 15.725 639.715 15.895 ;
        RECT 744.885 15.045 745.055 16.235 ;
      LAYER mcon ;
        RECT 637.705 17.425 637.875 17.595 ;
        RECT 639.545 16.065 639.715 16.235 ;
        RECT 744.885 16.065 745.055 16.235 ;
      LAYER met1 ;
        RECT 614.630 1589.740 614.950 1589.800 ;
        RECT 620.610 1589.740 620.930 1589.800 ;
        RECT 614.630 1589.600 620.930 1589.740 ;
        RECT 614.630 1589.540 614.950 1589.600 ;
        RECT 620.610 1589.540 620.930 1589.600 ;
        RECT 621.530 17.580 621.850 17.640 ;
        RECT 637.645 17.580 637.935 17.625 ;
        RECT 621.530 17.440 637.935 17.580 ;
        RECT 621.530 17.380 621.850 17.440 ;
        RECT 637.645 17.395 637.935 17.440 ;
        RECT 639.485 16.220 639.775 16.265 ;
        RECT 744.825 16.220 745.115 16.265 ;
        RECT 639.485 16.080 745.115 16.220 ;
        RECT 639.485 16.035 639.775 16.080 ;
        RECT 744.825 16.035 745.115 16.080 ;
        RECT 744.825 15.200 745.115 15.245 ;
        RECT 763.670 15.200 763.990 15.260 ;
        RECT 744.825 15.060 763.990 15.200 ;
        RECT 744.825 15.015 745.115 15.060 ;
        RECT 763.670 15.000 763.990 15.060 ;
      LAYER via ;
        RECT 614.660 1589.540 614.920 1589.800 ;
        RECT 620.640 1589.540 620.900 1589.800 ;
        RECT 621.560 17.380 621.820 17.640 ;
        RECT 763.700 15.000 763.960 15.260 ;
      LAYER met2 ;
        RECT 614.520 1600.380 614.800 1604.000 ;
        RECT 614.520 1600.000 614.860 1600.380 ;
        RECT 614.720 1589.830 614.860 1600.000 ;
        RECT 614.660 1589.510 614.920 1589.830 ;
        RECT 620.640 1589.510 620.900 1589.830 ;
        RECT 620.700 18.090 620.840 1589.510 ;
        RECT 620.700 17.950 621.760 18.090 ;
        RECT 621.620 17.670 621.760 17.950 ;
        RECT 621.560 17.350 621.820 17.670 ;
        RECT 763.700 14.970 763.960 15.290 ;
        RECT 763.760 2.400 763.900 14.970 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1066.350 1590.080 1066.670 1590.140 ;
        RECT 1068.190 1590.080 1068.510 1590.140 ;
        RECT 1066.350 1589.940 1068.510 1590.080 ;
        RECT 1066.350 1589.880 1066.670 1589.940 ;
        RECT 1068.190 1589.880 1068.510 1589.940 ;
        RECT 1068.190 57.700 1068.510 57.760 ;
        RECT 2063.170 57.700 2063.490 57.760 ;
        RECT 1068.190 57.560 2063.490 57.700 ;
        RECT 1068.190 57.500 1068.510 57.560 ;
        RECT 2063.170 57.500 2063.490 57.560 ;
        RECT 2063.170 2.960 2063.490 3.020 ;
        RECT 2066.390 2.960 2066.710 3.020 ;
        RECT 2063.170 2.820 2066.710 2.960 ;
        RECT 2063.170 2.760 2063.490 2.820 ;
        RECT 2066.390 2.760 2066.710 2.820 ;
      LAYER via ;
        RECT 1066.380 1589.880 1066.640 1590.140 ;
        RECT 1068.220 1589.880 1068.480 1590.140 ;
        RECT 1068.220 57.500 1068.480 57.760 ;
        RECT 2063.200 57.500 2063.460 57.760 ;
        RECT 2063.200 2.760 2063.460 3.020 ;
        RECT 2066.420 2.760 2066.680 3.020 ;
      LAYER met2 ;
        RECT 1066.240 1600.380 1066.520 1604.000 ;
        RECT 1066.240 1600.000 1066.580 1600.380 ;
        RECT 1066.440 1590.170 1066.580 1600.000 ;
        RECT 1066.380 1589.850 1066.640 1590.170 ;
        RECT 1068.220 1589.850 1068.480 1590.170 ;
        RECT 1068.280 57.790 1068.420 1589.850 ;
        RECT 1068.220 57.470 1068.480 57.790 ;
        RECT 2063.200 57.470 2063.460 57.790 ;
        RECT 2063.260 3.050 2063.400 57.470 ;
        RECT 2063.200 2.730 2063.460 3.050 ;
        RECT 2066.420 2.730 2066.680 3.050 ;
        RECT 2066.480 2.400 2066.620 2.730 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1072.330 1593.480 1072.650 1593.540 ;
        RECT 1075.550 1593.480 1075.870 1593.540 ;
        RECT 1072.330 1593.340 1075.870 1593.480 ;
        RECT 1072.330 1593.280 1072.650 1593.340 ;
        RECT 1075.550 1593.280 1075.870 1593.340 ;
        RECT 1075.550 58.040 1075.870 58.100 ;
        RECT 2084.330 58.040 2084.650 58.100 ;
        RECT 1075.550 57.900 2084.650 58.040 ;
        RECT 1075.550 57.840 1075.870 57.900 ;
        RECT 2084.330 57.840 2084.650 57.900 ;
      LAYER via ;
        RECT 1072.360 1593.280 1072.620 1593.540 ;
        RECT 1075.580 1593.280 1075.840 1593.540 ;
        RECT 1075.580 57.840 1075.840 58.100 ;
        RECT 2084.360 57.840 2084.620 58.100 ;
      LAYER met2 ;
        RECT 1072.220 1600.380 1072.500 1604.000 ;
        RECT 1072.220 1600.000 1072.560 1600.380 ;
        RECT 1072.420 1593.570 1072.560 1600.000 ;
        RECT 1072.360 1593.250 1072.620 1593.570 ;
        RECT 1075.580 1593.250 1075.840 1593.570 ;
        RECT 1075.640 58.130 1075.780 1593.250 ;
        RECT 1075.580 57.810 1075.840 58.130 ;
        RECT 2084.360 57.810 2084.620 58.130 ;
        RECT 2084.420 2.400 2084.560 57.810 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1078.770 1590.080 1079.090 1590.140 ;
        RECT 1081.990 1590.080 1082.310 1590.140 ;
        RECT 1078.770 1589.940 1082.310 1590.080 ;
        RECT 1078.770 1589.880 1079.090 1589.940 ;
        RECT 1081.990 1589.880 1082.310 1589.940 ;
        RECT 1081.990 58.380 1082.310 58.440 ;
        RECT 2097.670 58.380 2097.990 58.440 ;
        RECT 1081.990 58.240 2097.990 58.380 ;
        RECT 1081.990 58.180 1082.310 58.240 ;
        RECT 2097.670 58.180 2097.990 58.240 ;
        RECT 2097.670 2.960 2097.990 3.020 ;
        RECT 2101.810 2.960 2102.130 3.020 ;
        RECT 2097.670 2.820 2102.130 2.960 ;
        RECT 2097.670 2.760 2097.990 2.820 ;
        RECT 2101.810 2.760 2102.130 2.820 ;
      LAYER via ;
        RECT 1078.800 1589.880 1079.060 1590.140 ;
        RECT 1082.020 1589.880 1082.280 1590.140 ;
        RECT 1082.020 58.180 1082.280 58.440 ;
        RECT 2097.700 58.180 2097.960 58.440 ;
        RECT 2097.700 2.760 2097.960 3.020 ;
        RECT 2101.840 2.760 2102.100 3.020 ;
      LAYER met2 ;
        RECT 1078.660 1600.380 1078.940 1604.000 ;
        RECT 1078.660 1600.000 1079.000 1600.380 ;
        RECT 1078.860 1590.170 1079.000 1600.000 ;
        RECT 1078.800 1589.850 1079.060 1590.170 ;
        RECT 1082.020 1589.850 1082.280 1590.170 ;
        RECT 1082.080 58.470 1082.220 1589.850 ;
        RECT 1082.020 58.150 1082.280 58.470 ;
        RECT 2097.700 58.150 2097.960 58.470 ;
        RECT 2097.760 3.050 2097.900 58.150 ;
        RECT 2097.700 2.730 2097.960 3.050 ;
        RECT 2101.840 2.730 2102.100 3.050 ;
        RECT 2101.900 2.400 2102.040 2.730 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1084.750 1590.080 1085.070 1590.140 ;
        RECT 1089.350 1590.080 1089.670 1590.140 ;
        RECT 1084.750 1589.940 1089.670 1590.080 ;
        RECT 1084.750 1589.880 1085.070 1589.940 ;
        RECT 1089.350 1589.880 1089.670 1589.940 ;
        RECT 1089.350 62.120 1089.670 62.180 ;
        RECT 2118.370 62.120 2118.690 62.180 ;
        RECT 1089.350 61.980 2118.690 62.120 ;
        RECT 1089.350 61.920 1089.670 61.980 ;
        RECT 2118.370 61.920 2118.690 61.980 ;
        RECT 2118.370 2.960 2118.690 3.020 ;
        RECT 2119.750 2.960 2120.070 3.020 ;
        RECT 2118.370 2.820 2120.070 2.960 ;
        RECT 2118.370 2.760 2118.690 2.820 ;
        RECT 2119.750 2.760 2120.070 2.820 ;
      LAYER via ;
        RECT 1084.780 1589.880 1085.040 1590.140 ;
        RECT 1089.380 1589.880 1089.640 1590.140 ;
        RECT 1089.380 61.920 1089.640 62.180 ;
        RECT 2118.400 61.920 2118.660 62.180 ;
        RECT 2118.400 2.760 2118.660 3.020 ;
        RECT 2119.780 2.760 2120.040 3.020 ;
      LAYER met2 ;
        RECT 1084.640 1600.380 1084.920 1604.000 ;
        RECT 1084.640 1600.000 1084.980 1600.380 ;
        RECT 1084.840 1590.170 1084.980 1600.000 ;
        RECT 1084.780 1589.850 1085.040 1590.170 ;
        RECT 1089.380 1589.850 1089.640 1590.170 ;
        RECT 1089.440 62.210 1089.580 1589.850 ;
        RECT 1089.380 61.890 1089.640 62.210 ;
        RECT 2118.400 61.890 2118.660 62.210 ;
        RECT 2118.460 3.050 2118.600 61.890 ;
        RECT 2118.400 2.730 2118.660 3.050 ;
        RECT 2119.780 2.730 2120.040 3.050 ;
        RECT 2119.840 2.400 2119.980 2.730 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1090.730 1590.080 1091.050 1590.140 ;
        RECT 1095.790 1590.080 1096.110 1590.140 ;
        RECT 1090.730 1589.940 1096.110 1590.080 ;
        RECT 1090.730 1589.880 1091.050 1589.940 ;
        RECT 1095.790 1589.880 1096.110 1589.940 ;
        RECT 1095.790 61.780 1096.110 61.840 ;
        RECT 2132.170 61.780 2132.490 61.840 ;
        RECT 1095.790 61.640 2132.490 61.780 ;
        RECT 1095.790 61.580 1096.110 61.640 ;
        RECT 2132.170 61.580 2132.490 61.640 ;
        RECT 2132.170 2.960 2132.490 3.020 ;
        RECT 2137.690 2.960 2138.010 3.020 ;
        RECT 2132.170 2.820 2138.010 2.960 ;
        RECT 2132.170 2.760 2132.490 2.820 ;
        RECT 2137.690 2.760 2138.010 2.820 ;
      LAYER via ;
        RECT 1090.760 1589.880 1091.020 1590.140 ;
        RECT 1095.820 1589.880 1096.080 1590.140 ;
        RECT 1095.820 61.580 1096.080 61.840 ;
        RECT 2132.200 61.580 2132.460 61.840 ;
        RECT 2132.200 2.760 2132.460 3.020 ;
        RECT 2137.720 2.760 2137.980 3.020 ;
      LAYER met2 ;
        RECT 1090.620 1600.380 1090.900 1604.000 ;
        RECT 1090.620 1600.000 1090.960 1600.380 ;
        RECT 1090.820 1590.170 1090.960 1600.000 ;
        RECT 1090.760 1589.850 1091.020 1590.170 ;
        RECT 1095.820 1589.850 1096.080 1590.170 ;
        RECT 1095.880 61.870 1096.020 1589.850 ;
        RECT 1095.820 61.550 1096.080 61.870 ;
        RECT 2132.200 61.550 2132.460 61.870 ;
        RECT 2132.260 3.050 2132.400 61.550 ;
        RECT 2132.200 2.730 2132.460 3.050 ;
        RECT 2137.720 2.730 2137.980 3.050 ;
        RECT 2137.780 2.400 2137.920 2.730 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1097.170 1590.080 1097.490 1590.140 ;
        RECT 1102.690 1590.080 1103.010 1590.140 ;
        RECT 1097.170 1589.940 1103.010 1590.080 ;
        RECT 1097.170 1589.880 1097.490 1589.940 ;
        RECT 1102.690 1589.880 1103.010 1589.940 ;
        RECT 1102.690 61.440 1103.010 61.500 ;
        RECT 2152.870 61.440 2153.190 61.500 ;
        RECT 1102.690 61.300 2153.190 61.440 ;
        RECT 1102.690 61.240 1103.010 61.300 ;
        RECT 2152.870 61.240 2153.190 61.300 ;
        RECT 2152.870 2.960 2153.190 3.020 ;
        RECT 2155.630 2.960 2155.950 3.020 ;
        RECT 2152.870 2.820 2155.950 2.960 ;
        RECT 2152.870 2.760 2153.190 2.820 ;
        RECT 2155.630 2.760 2155.950 2.820 ;
      LAYER via ;
        RECT 1097.200 1589.880 1097.460 1590.140 ;
        RECT 1102.720 1589.880 1102.980 1590.140 ;
        RECT 1102.720 61.240 1102.980 61.500 ;
        RECT 2152.900 61.240 2153.160 61.500 ;
        RECT 2152.900 2.760 2153.160 3.020 ;
        RECT 2155.660 2.760 2155.920 3.020 ;
      LAYER met2 ;
        RECT 1097.060 1600.380 1097.340 1604.000 ;
        RECT 1097.060 1600.000 1097.400 1600.380 ;
        RECT 1097.260 1590.170 1097.400 1600.000 ;
        RECT 1097.200 1589.850 1097.460 1590.170 ;
        RECT 1102.720 1589.850 1102.980 1590.170 ;
        RECT 1102.780 61.530 1102.920 1589.850 ;
        RECT 1102.720 61.210 1102.980 61.530 ;
        RECT 2152.900 61.210 2153.160 61.530 ;
        RECT 2152.960 3.050 2153.100 61.210 ;
        RECT 2152.900 2.730 2153.160 3.050 ;
        RECT 2155.660 2.730 2155.920 3.050 ;
        RECT 2155.720 2.400 2155.860 2.730 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1103.150 61.100 1103.470 61.160 ;
        RECT 2166.670 61.100 2166.990 61.160 ;
        RECT 1103.150 60.960 2166.990 61.100 ;
        RECT 1103.150 60.900 1103.470 60.960 ;
        RECT 2166.670 60.900 2166.990 60.960 ;
        RECT 2166.670 17.580 2166.990 17.640 ;
        RECT 2173.110 17.580 2173.430 17.640 ;
        RECT 2166.670 17.440 2173.430 17.580 ;
        RECT 2166.670 17.380 2166.990 17.440 ;
        RECT 2173.110 17.380 2173.430 17.440 ;
      LAYER via ;
        RECT 1103.180 60.900 1103.440 61.160 ;
        RECT 2166.700 60.900 2166.960 61.160 ;
        RECT 2166.700 17.380 2166.960 17.640 ;
        RECT 2173.140 17.380 2173.400 17.640 ;
      LAYER met2 ;
        RECT 1103.040 1600.380 1103.320 1604.000 ;
        RECT 1103.040 1600.000 1103.380 1600.380 ;
        RECT 1103.240 61.190 1103.380 1600.000 ;
        RECT 1103.180 60.870 1103.440 61.190 ;
        RECT 2166.700 60.870 2166.960 61.190 ;
        RECT 2166.760 17.670 2166.900 60.870 ;
        RECT 2166.700 17.350 2166.960 17.670 ;
        RECT 2173.140 17.350 2173.400 17.670 ;
        RECT 2173.200 2.400 2173.340 17.350 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1109.590 60.760 1109.910 60.820 ;
        RECT 2187.370 60.760 2187.690 60.820 ;
        RECT 1109.590 60.620 2187.690 60.760 ;
        RECT 1109.590 60.560 1109.910 60.620 ;
        RECT 2187.370 60.560 2187.690 60.620 ;
        RECT 2187.370 2.960 2187.690 3.020 ;
        RECT 2191.050 2.960 2191.370 3.020 ;
        RECT 2187.370 2.820 2191.370 2.960 ;
        RECT 2187.370 2.760 2187.690 2.820 ;
        RECT 2191.050 2.760 2191.370 2.820 ;
      LAYER via ;
        RECT 1109.620 60.560 1109.880 60.820 ;
        RECT 2187.400 60.560 2187.660 60.820 ;
        RECT 2187.400 2.760 2187.660 3.020 ;
        RECT 2191.080 2.760 2191.340 3.020 ;
      LAYER met2 ;
        RECT 1109.480 1600.380 1109.760 1604.000 ;
        RECT 1109.480 1600.000 1109.820 1600.380 ;
        RECT 1109.680 60.850 1109.820 1600.000 ;
        RECT 1109.620 60.530 1109.880 60.850 ;
        RECT 2187.400 60.530 2187.660 60.850 ;
        RECT 2187.460 3.050 2187.600 60.530 ;
        RECT 2187.400 2.730 2187.660 3.050 ;
        RECT 2191.080 2.730 2191.340 3.050 ;
        RECT 2191.140 2.400 2191.280 2.730 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1116.950 60.420 1117.270 60.480 ;
        RECT 2208.070 60.420 2208.390 60.480 ;
        RECT 1116.950 60.280 2208.390 60.420 ;
        RECT 1116.950 60.220 1117.270 60.280 ;
        RECT 2208.070 60.220 2208.390 60.280 ;
      LAYER via ;
        RECT 1116.980 60.220 1117.240 60.480 ;
        RECT 2208.100 60.220 2208.360 60.480 ;
      LAYER met2 ;
        RECT 1115.460 1600.450 1115.740 1604.000 ;
        RECT 1115.460 1600.310 1117.180 1600.450 ;
        RECT 1115.460 1600.000 1115.740 1600.310 ;
        RECT 1117.040 60.510 1117.180 1600.310 ;
        RECT 1116.980 60.190 1117.240 60.510 ;
        RECT 2208.100 60.190 2208.360 60.510 ;
        RECT 2208.160 17.410 2208.300 60.190 ;
        RECT 2208.160 17.270 2209.220 17.410 ;
        RECT 2209.080 2.400 2209.220 17.270 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1123.390 60.080 1123.710 60.140 ;
        RECT 2221.870 60.080 2222.190 60.140 ;
        RECT 1123.390 59.940 2222.190 60.080 ;
        RECT 1123.390 59.880 1123.710 59.940 ;
        RECT 2221.870 59.880 2222.190 59.940 ;
      LAYER via ;
        RECT 1123.420 59.880 1123.680 60.140 ;
        RECT 2221.900 59.880 2222.160 60.140 ;
      LAYER met2 ;
        RECT 1121.900 1600.450 1122.180 1604.000 ;
        RECT 1121.900 1600.310 1122.700 1600.450 ;
        RECT 1121.900 1600.000 1122.180 1600.310 ;
        RECT 1122.560 1580.050 1122.700 1600.310 ;
        RECT 1122.560 1579.910 1123.620 1580.050 ;
        RECT 1123.480 60.170 1123.620 1579.910 ;
        RECT 1123.420 59.850 1123.680 60.170 ;
        RECT 2221.900 59.850 2222.160 60.170 ;
        RECT 2221.960 17.410 2222.100 59.850 ;
        RECT 2221.960 17.270 2227.160 17.410 ;
        RECT 2227.020 2.400 2227.160 17.270 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 746.265 1588.905 746.435 1591.795 ;
      LAYER mcon ;
        RECT 746.265 1591.625 746.435 1591.795 ;
      LAYER met1 ;
        RECT 621.070 1591.780 621.390 1591.840 ;
        RECT 746.205 1591.780 746.495 1591.825 ;
        RECT 621.070 1591.640 746.495 1591.780 ;
        RECT 621.070 1591.580 621.390 1591.640 ;
        RECT 746.205 1591.595 746.495 1591.640 ;
        RECT 769.190 1589.740 769.510 1589.800 ;
        RECT 759.620 1589.600 769.510 1589.740 ;
        RECT 759.620 1589.400 759.760 1589.600 ;
        RECT 769.190 1589.540 769.510 1589.600 ;
        RECT 755.480 1589.260 759.760 1589.400 ;
        RECT 746.205 1589.060 746.495 1589.105 ;
        RECT 755.480 1589.060 755.620 1589.260 ;
        RECT 746.205 1588.920 755.620 1589.060 ;
        RECT 746.205 1588.875 746.495 1588.920 ;
        RECT 769.190 20.300 769.510 20.360 ;
        RECT 781.610 20.300 781.930 20.360 ;
        RECT 769.190 20.160 781.930 20.300 ;
        RECT 769.190 20.100 769.510 20.160 ;
        RECT 781.610 20.100 781.930 20.160 ;
      LAYER via ;
        RECT 621.100 1591.580 621.360 1591.840 ;
        RECT 769.220 1589.540 769.480 1589.800 ;
        RECT 769.220 20.100 769.480 20.360 ;
        RECT 781.640 20.100 781.900 20.360 ;
      LAYER met2 ;
        RECT 620.960 1600.380 621.240 1604.000 ;
        RECT 620.960 1600.000 621.300 1600.380 ;
        RECT 621.160 1591.870 621.300 1600.000 ;
        RECT 621.100 1591.550 621.360 1591.870 ;
        RECT 769.220 1589.510 769.480 1589.830 ;
        RECT 769.280 20.390 769.420 1589.510 ;
        RECT 769.220 20.070 769.480 20.390 ;
        RECT 781.640 20.070 781.900 20.390 ;
        RECT 781.700 2.400 781.840 20.070 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1130.290 59.740 1130.610 59.800 ;
        RECT 2242.570 59.740 2242.890 59.800 ;
        RECT 1130.290 59.600 2242.890 59.740 ;
        RECT 1130.290 59.540 1130.610 59.600 ;
        RECT 2242.570 59.540 2242.890 59.600 ;
      LAYER via ;
        RECT 1130.320 59.540 1130.580 59.800 ;
        RECT 2242.600 59.540 2242.860 59.800 ;
      LAYER met2 ;
        RECT 1127.880 1600.450 1128.160 1604.000 ;
        RECT 1127.880 1600.310 1129.140 1600.450 ;
        RECT 1127.880 1600.000 1128.160 1600.310 ;
        RECT 1129.000 1580.050 1129.140 1600.310 ;
        RECT 1129.000 1579.910 1130.520 1580.050 ;
        RECT 1130.380 59.830 1130.520 1579.910 ;
        RECT 1130.320 59.510 1130.580 59.830 ;
        RECT 2242.600 59.510 2242.860 59.830 ;
        RECT 2242.660 17.410 2242.800 59.510 ;
        RECT 2242.660 17.270 2245.100 17.410 ;
        RECT 2244.960 2.400 2245.100 17.270 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1136.805 1449.165 1136.975 1497.275 ;
        RECT 1136.805 786.505 1136.975 821.015 ;
        RECT 1136.805 689.605 1136.975 724.455 ;
        RECT 1136.805 593.045 1136.975 627.895 ;
        RECT 1136.805 496.485 1136.975 531.335 ;
        RECT 1136.805 386.325 1136.975 434.775 ;
        RECT 1136.805 255.085 1136.975 289.595 ;
        RECT 1136.805 59.245 1136.975 96.475 ;
      LAYER mcon ;
        RECT 1136.805 1497.105 1136.975 1497.275 ;
        RECT 1136.805 820.845 1136.975 821.015 ;
        RECT 1136.805 724.285 1136.975 724.455 ;
        RECT 1136.805 627.725 1136.975 627.895 ;
        RECT 1136.805 531.165 1136.975 531.335 ;
        RECT 1136.805 434.605 1136.975 434.775 ;
        RECT 1136.805 289.425 1136.975 289.595 ;
        RECT 1136.805 96.305 1136.975 96.475 ;
      LAYER met1 ;
        RECT 1136.730 1497.260 1137.050 1497.320 ;
        RECT 1136.535 1497.120 1137.050 1497.260 ;
        RECT 1136.730 1497.060 1137.050 1497.120 ;
        RECT 1136.745 1449.320 1137.035 1449.365 ;
        RECT 1137.190 1449.320 1137.510 1449.380 ;
        RECT 1136.745 1449.180 1137.510 1449.320 ;
        RECT 1136.745 1449.135 1137.035 1449.180 ;
        RECT 1137.190 1449.120 1137.510 1449.180 ;
        RECT 1136.270 1414.640 1136.590 1414.700 ;
        RECT 1137.190 1414.640 1137.510 1414.700 ;
        RECT 1136.270 1414.500 1137.510 1414.640 ;
        RECT 1136.270 1414.440 1136.590 1414.500 ;
        RECT 1137.190 1414.440 1137.510 1414.500 ;
        RECT 1136.270 1318.080 1136.590 1318.140 ;
        RECT 1137.190 1318.080 1137.510 1318.140 ;
        RECT 1136.270 1317.940 1137.510 1318.080 ;
        RECT 1136.270 1317.880 1136.590 1317.940 ;
        RECT 1137.190 1317.880 1137.510 1317.940 ;
        RECT 1136.270 1221.520 1136.590 1221.580 ;
        RECT 1137.190 1221.520 1137.510 1221.580 ;
        RECT 1136.270 1221.380 1137.510 1221.520 ;
        RECT 1136.270 1221.320 1136.590 1221.380 ;
        RECT 1137.190 1221.320 1137.510 1221.380 ;
        RECT 1136.270 1124.960 1136.590 1125.020 ;
        RECT 1137.190 1124.960 1137.510 1125.020 ;
        RECT 1136.270 1124.820 1137.510 1124.960 ;
        RECT 1136.270 1124.760 1136.590 1124.820 ;
        RECT 1137.190 1124.760 1137.510 1124.820 ;
        RECT 1136.270 1028.400 1136.590 1028.460 ;
        RECT 1137.190 1028.400 1137.510 1028.460 ;
        RECT 1136.270 1028.260 1137.510 1028.400 ;
        RECT 1136.270 1028.200 1136.590 1028.260 ;
        RECT 1137.190 1028.200 1137.510 1028.260 ;
        RECT 1136.270 931.840 1136.590 931.900 ;
        RECT 1137.190 931.840 1137.510 931.900 ;
        RECT 1136.270 931.700 1137.510 931.840 ;
        RECT 1136.270 931.640 1136.590 931.700 ;
        RECT 1137.190 931.640 1137.510 931.700 ;
        RECT 1135.810 869.620 1136.130 869.680 ;
        RECT 1137.190 869.620 1137.510 869.680 ;
        RECT 1135.810 869.480 1137.510 869.620 ;
        RECT 1135.810 869.420 1136.130 869.480 ;
        RECT 1137.190 869.420 1137.510 869.480 ;
        RECT 1136.270 835.280 1136.590 835.340 ;
        RECT 1137.190 835.280 1137.510 835.340 ;
        RECT 1136.270 835.140 1137.510 835.280 ;
        RECT 1136.270 835.080 1136.590 835.140 ;
        RECT 1137.190 835.080 1137.510 835.140 ;
        RECT 1136.730 821.000 1137.050 821.060 ;
        RECT 1136.535 820.860 1137.050 821.000 ;
        RECT 1136.730 820.800 1137.050 820.860 ;
        RECT 1136.730 786.660 1137.050 786.720 ;
        RECT 1136.535 786.520 1137.050 786.660 ;
        RECT 1136.730 786.460 1137.050 786.520 ;
        RECT 1136.270 738.380 1136.590 738.440 ;
        RECT 1137.190 738.380 1137.510 738.440 ;
        RECT 1136.270 738.240 1137.510 738.380 ;
        RECT 1136.270 738.180 1136.590 738.240 ;
        RECT 1137.190 738.180 1137.510 738.240 ;
        RECT 1136.730 724.440 1137.050 724.500 ;
        RECT 1136.535 724.300 1137.050 724.440 ;
        RECT 1136.730 724.240 1137.050 724.300 ;
        RECT 1136.730 689.760 1137.050 689.820 ;
        RECT 1136.535 689.620 1137.050 689.760 ;
        RECT 1136.730 689.560 1137.050 689.620 ;
        RECT 1136.270 641.820 1136.590 641.880 ;
        RECT 1137.190 641.820 1137.510 641.880 ;
        RECT 1136.270 641.680 1137.510 641.820 ;
        RECT 1136.270 641.620 1136.590 641.680 ;
        RECT 1137.190 641.620 1137.510 641.680 ;
        RECT 1136.730 627.880 1137.050 627.940 ;
        RECT 1136.535 627.740 1137.050 627.880 ;
        RECT 1136.730 627.680 1137.050 627.740 ;
        RECT 1136.730 593.200 1137.050 593.260 ;
        RECT 1136.535 593.060 1137.050 593.200 ;
        RECT 1136.730 593.000 1137.050 593.060 ;
        RECT 1136.270 545.260 1136.590 545.320 ;
        RECT 1137.190 545.260 1137.510 545.320 ;
        RECT 1136.270 545.120 1137.510 545.260 ;
        RECT 1136.270 545.060 1136.590 545.120 ;
        RECT 1137.190 545.060 1137.510 545.120 ;
        RECT 1136.730 531.320 1137.050 531.380 ;
        RECT 1136.535 531.180 1137.050 531.320 ;
        RECT 1136.730 531.120 1137.050 531.180 ;
        RECT 1136.730 496.640 1137.050 496.700 ;
        RECT 1136.535 496.500 1137.050 496.640 ;
        RECT 1136.730 496.440 1137.050 496.500 ;
        RECT 1136.270 448.700 1136.590 448.760 ;
        RECT 1137.190 448.700 1137.510 448.760 ;
        RECT 1136.270 448.560 1137.510 448.700 ;
        RECT 1136.270 448.500 1136.590 448.560 ;
        RECT 1137.190 448.500 1137.510 448.560 ;
        RECT 1136.730 434.760 1137.050 434.820 ;
        RECT 1136.535 434.620 1137.050 434.760 ;
        RECT 1136.730 434.560 1137.050 434.620 ;
        RECT 1136.745 386.480 1137.035 386.525 ;
        RECT 1137.190 386.480 1137.510 386.540 ;
        RECT 1136.745 386.340 1137.510 386.480 ;
        RECT 1136.745 386.295 1137.035 386.340 ;
        RECT 1137.190 386.280 1137.510 386.340 ;
        RECT 1136.745 289.580 1137.035 289.625 ;
        RECT 1137.190 289.580 1137.510 289.640 ;
        RECT 1136.745 289.440 1137.510 289.580 ;
        RECT 1136.745 289.395 1137.035 289.440 ;
        RECT 1137.190 289.380 1137.510 289.440 ;
        RECT 1136.730 255.240 1137.050 255.300 ;
        RECT 1136.535 255.100 1137.050 255.240 ;
        RECT 1136.730 255.040 1137.050 255.100 ;
        RECT 1136.270 158.680 1136.590 158.740 ;
        RECT 1137.190 158.680 1137.510 158.740 ;
        RECT 1136.270 158.540 1137.510 158.680 ;
        RECT 1136.270 158.480 1136.590 158.540 ;
        RECT 1137.190 158.480 1137.510 158.540 ;
        RECT 1136.730 96.460 1137.050 96.520 ;
        RECT 1136.535 96.320 1137.050 96.460 ;
        RECT 1136.730 96.260 1137.050 96.320 ;
        RECT 1136.745 59.400 1137.035 59.445 ;
        RECT 2256.370 59.400 2256.690 59.460 ;
        RECT 1136.745 59.260 2256.690 59.400 ;
        RECT 1136.745 59.215 1137.035 59.260 ;
        RECT 2256.370 59.200 2256.690 59.260 ;
        RECT 2256.370 17.580 2256.690 17.640 ;
        RECT 2262.350 17.580 2262.670 17.640 ;
        RECT 2256.370 17.440 2262.670 17.580 ;
        RECT 2256.370 17.380 2256.690 17.440 ;
        RECT 2262.350 17.380 2262.670 17.440 ;
      LAYER via ;
        RECT 1136.760 1497.060 1137.020 1497.320 ;
        RECT 1137.220 1449.120 1137.480 1449.380 ;
        RECT 1136.300 1414.440 1136.560 1414.700 ;
        RECT 1137.220 1414.440 1137.480 1414.700 ;
        RECT 1136.300 1317.880 1136.560 1318.140 ;
        RECT 1137.220 1317.880 1137.480 1318.140 ;
        RECT 1136.300 1221.320 1136.560 1221.580 ;
        RECT 1137.220 1221.320 1137.480 1221.580 ;
        RECT 1136.300 1124.760 1136.560 1125.020 ;
        RECT 1137.220 1124.760 1137.480 1125.020 ;
        RECT 1136.300 1028.200 1136.560 1028.460 ;
        RECT 1137.220 1028.200 1137.480 1028.460 ;
        RECT 1136.300 931.640 1136.560 931.900 ;
        RECT 1137.220 931.640 1137.480 931.900 ;
        RECT 1135.840 869.420 1136.100 869.680 ;
        RECT 1137.220 869.420 1137.480 869.680 ;
        RECT 1136.300 835.080 1136.560 835.340 ;
        RECT 1137.220 835.080 1137.480 835.340 ;
        RECT 1136.760 820.800 1137.020 821.060 ;
        RECT 1136.760 786.460 1137.020 786.720 ;
        RECT 1136.300 738.180 1136.560 738.440 ;
        RECT 1137.220 738.180 1137.480 738.440 ;
        RECT 1136.760 724.240 1137.020 724.500 ;
        RECT 1136.760 689.560 1137.020 689.820 ;
        RECT 1136.300 641.620 1136.560 641.880 ;
        RECT 1137.220 641.620 1137.480 641.880 ;
        RECT 1136.760 627.680 1137.020 627.940 ;
        RECT 1136.760 593.000 1137.020 593.260 ;
        RECT 1136.300 545.060 1136.560 545.320 ;
        RECT 1137.220 545.060 1137.480 545.320 ;
        RECT 1136.760 531.120 1137.020 531.380 ;
        RECT 1136.760 496.440 1137.020 496.700 ;
        RECT 1136.300 448.500 1136.560 448.760 ;
        RECT 1137.220 448.500 1137.480 448.760 ;
        RECT 1136.760 434.560 1137.020 434.820 ;
        RECT 1137.220 386.280 1137.480 386.540 ;
        RECT 1137.220 289.380 1137.480 289.640 ;
        RECT 1136.760 255.040 1137.020 255.300 ;
        RECT 1136.300 158.480 1136.560 158.740 ;
        RECT 1137.220 158.480 1137.480 158.740 ;
        RECT 1136.760 96.260 1137.020 96.520 ;
        RECT 2256.400 59.200 2256.660 59.460 ;
        RECT 2256.400 17.380 2256.660 17.640 ;
        RECT 2262.380 17.380 2262.640 17.640 ;
      LAYER met2 ;
        RECT 1134.320 1600.450 1134.600 1604.000 ;
        RECT 1134.320 1600.310 1135.120 1600.450 ;
        RECT 1134.320 1600.000 1134.600 1600.310 ;
        RECT 1134.980 1569.850 1135.120 1600.310 ;
        RECT 1134.980 1569.710 1136.500 1569.850 ;
        RECT 1136.360 1510.690 1136.500 1569.710 ;
        RECT 1136.360 1510.550 1136.960 1510.690 ;
        RECT 1136.820 1497.350 1136.960 1510.550 ;
        RECT 1136.760 1497.030 1137.020 1497.350 ;
        RECT 1137.220 1449.090 1137.480 1449.410 ;
        RECT 1137.280 1414.730 1137.420 1449.090 ;
        RECT 1136.300 1414.410 1136.560 1414.730 ;
        RECT 1137.220 1414.410 1137.480 1414.730 ;
        RECT 1136.360 1414.130 1136.500 1414.410 ;
        RECT 1136.360 1413.990 1136.960 1414.130 ;
        RECT 1136.820 1366.530 1136.960 1413.990 ;
        RECT 1136.820 1366.390 1137.420 1366.530 ;
        RECT 1137.280 1318.170 1137.420 1366.390 ;
        RECT 1136.300 1317.850 1136.560 1318.170 ;
        RECT 1137.220 1317.850 1137.480 1318.170 ;
        RECT 1136.360 1317.570 1136.500 1317.850 ;
        RECT 1136.360 1317.430 1136.960 1317.570 ;
        RECT 1136.820 1269.970 1136.960 1317.430 ;
        RECT 1136.820 1269.830 1137.420 1269.970 ;
        RECT 1137.280 1221.610 1137.420 1269.830 ;
        RECT 1136.300 1221.290 1136.560 1221.610 ;
        RECT 1137.220 1221.290 1137.480 1221.610 ;
        RECT 1136.360 1221.010 1136.500 1221.290 ;
        RECT 1136.360 1220.870 1136.960 1221.010 ;
        RECT 1136.820 1173.410 1136.960 1220.870 ;
        RECT 1136.820 1173.270 1137.420 1173.410 ;
        RECT 1137.280 1125.050 1137.420 1173.270 ;
        RECT 1136.300 1124.730 1136.560 1125.050 ;
        RECT 1137.220 1124.730 1137.480 1125.050 ;
        RECT 1136.360 1124.450 1136.500 1124.730 ;
        RECT 1136.360 1124.310 1136.960 1124.450 ;
        RECT 1136.820 1076.850 1136.960 1124.310 ;
        RECT 1136.820 1076.710 1137.420 1076.850 ;
        RECT 1137.280 1028.490 1137.420 1076.710 ;
        RECT 1136.300 1028.170 1136.560 1028.490 ;
        RECT 1137.220 1028.170 1137.480 1028.490 ;
        RECT 1136.360 1027.890 1136.500 1028.170 ;
        RECT 1136.360 1027.750 1136.960 1027.890 ;
        RECT 1136.820 980.290 1136.960 1027.750 ;
        RECT 1136.820 980.150 1137.420 980.290 ;
        RECT 1137.280 931.930 1137.420 980.150 ;
        RECT 1136.300 931.610 1136.560 931.930 ;
        RECT 1137.220 931.610 1137.480 931.930 ;
        RECT 1136.360 931.330 1136.500 931.610 ;
        RECT 1136.360 931.190 1136.960 931.330 ;
        RECT 1136.820 917.845 1136.960 931.190 ;
        RECT 1135.830 917.475 1136.110 917.845 ;
        RECT 1136.750 917.475 1137.030 917.845 ;
        RECT 1135.900 869.710 1136.040 917.475 ;
        RECT 1135.840 869.390 1136.100 869.710 ;
        RECT 1137.220 869.390 1137.480 869.710 ;
        RECT 1137.280 835.370 1137.420 869.390 ;
        RECT 1136.300 835.050 1136.560 835.370 ;
        RECT 1137.220 835.050 1137.480 835.370 ;
        RECT 1136.360 834.770 1136.500 835.050 ;
        RECT 1136.360 834.630 1136.960 834.770 ;
        RECT 1136.820 821.090 1136.960 834.630 ;
        RECT 1136.760 820.770 1137.020 821.090 ;
        RECT 1136.760 786.430 1137.020 786.750 ;
        RECT 1136.820 772.890 1136.960 786.430 ;
        RECT 1136.820 772.750 1137.420 772.890 ;
        RECT 1137.280 738.470 1137.420 772.750 ;
        RECT 1136.300 738.210 1136.560 738.470 ;
        RECT 1136.300 738.150 1136.960 738.210 ;
        RECT 1137.220 738.150 1137.480 738.470 ;
        RECT 1136.360 738.070 1136.960 738.150 ;
        RECT 1136.820 724.530 1136.960 738.070 ;
        RECT 1136.760 724.210 1137.020 724.530 ;
        RECT 1136.760 689.530 1137.020 689.850 ;
        RECT 1136.820 676.330 1136.960 689.530 ;
        RECT 1136.820 676.190 1137.420 676.330 ;
        RECT 1137.280 641.910 1137.420 676.190 ;
        RECT 1136.300 641.650 1136.560 641.910 ;
        RECT 1136.300 641.590 1136.960 641.650 ;
        RECT 1137.220 641.590 1137.480 641.910 ;
        RECT 1136.360 641.510 1136.960 641.590 ;
        RECT 1136.820 627.970 1136.960 641.510 ;
        RECT 1136.760 627.650 1137.020 627.970 ;
        RECT 1136.760 592.970 1137.020 593.290 ;
        RECT 1136.820 579.770 1136.960 592.970 ;
        RECT 1136.820 579.630 1137.420 579.770 ;
        RECT 1137.280 545.350 1137.420 579.630 ;
        RECT 1136.300 545.090 1136.560 545.350 ;
        RECT 1136.300 545.030 1136.960 545.090 ;
        RECT 1137.220 545.030 1137.480 545.350 ;
        RECT 1136.360 544.950 1136.960 545.030 ;
        RECT 1136.820 531.410 1136.960 544.950 ;
        RECT 1136.760 531.090 1137.020 531.410 ;
        RECT 1136.760 496.410 1137.020 496.730 ;
        RECT 1136.820 483.210 1136.960 496.410 ;
        RECT 1136.820 483.070 1137.420 483.210 ;
        RECT 1137.280 448.790 1137.420 483.070 ;
        RECT 1136.300 448.530 1136.560 448.790 ;
        RECT 1136.300 448.470 1136.960 448.530 ;
        RECT 1137.220 448.470 1137.480 448.790 ;
        RECT 1136.360 448.390 1136.960 448.470 ;
        RECT 1136.820 434.850 1136.960 448.390 ;
        RECT 1136.760 434.530 1137.020 434.850 ;
        RECT 1137.220 386.250 1137.480 386.570 ;
        RECT 1137.280 351.290 1137.420 386.250 ;
        RECT 1136.820 351.150 1137.420 351.290 ;
        RECT 1136.820 303.690 1136.960 351.150 ;
        RECT 1136.820 303.550 1137.420 303.690 ;
        RECT 1137.280 289.670 1137.420 303.550 ;
        RECT 1137.220 289.350 1137.480 289.670 ;
        RECT 1136.760 255.010 1137.020 255.330 ;
        RECT 1136.820 207.130 1136.960 255.010 ;
        RECT 1136.820 206.990 1137.420 207.130 ;
        RECT 1137.280 158.850 1137.420 206.990 ;
        RECT 1136.360 158.770 1137.420 158.850 ;
        RECT 1136.300 158.710 1137.480 158.770 ;
        RECT 1136.300 158.450 1136.560 158.710 ;
        RECT 1137.220 158.450 1137.480 158.710 ;
        RECT 1136.360 158.295 1136.500 158.450 ;
        RECT 1137.280 110.685 1137.420 158.450 ;
        RECT 1137.210 110.315 1137.490 110.685 ;
        RECT 1136.750 96.715 1137.030 97.085 ;
        RECT 1136.820 96.550 1136.960 96.715 ;
        RECT 1136.760 96.230 1137.020 96.550 ;
        RECT 2256.400 59.170 2256.660 59.490 ;
        RECT 2256.460 17.670 2256.600 59.170 ;
        RECT 2256.400 17.350 2256.660 17.670 ;
        RECT 2262.380 17.350 2262.640 17.670 ;
        RECT 2262.440 2.400 2262.580 17.350 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
      LAYER via2 ;
        RECT 1135.830 917.520 1136.110 917.800 ;
        RECT 1136.750 917.520 1137.030 917.800 ;
        RECT 1137.210 110.360 1137.490 110.640 ;
        RECT 1136.750 96.760 1137.030 97.040 ;
      LAYER met3 ;
        RECT 1135.805 917.810 1136.135 917.825 ;
        RECT 1136.725 917.810 1137.055 917.825 ;
        RECT 1135.805 917.510 1137.055 917.810 ;
        RECT 1135.805 917.495 1136.135 917.510 ;
        RECT 1136.725 917.495 1137.055 917.510 ;
        RECT 1136.470 110.650 1136.850 110.660 ;
        RECT 1137.185 110.650 1137.515 110.665 ;
        RECT 1136.470 110.350 1137.515 110.650 ;
        RECT 1136.470 110.340 1136.850 110.350 ;
        RECT 1137.185 110.335 1137.515 110.350 ;
        RECT 1136.725 97.060 1137.055 97.065 ;
        RECT 1136.470 97.050 1137.055 97.060 ;
        RECT 1136.470 96.750 1137.280 97.050 ;
        RECT 1136.470 96.740 1137.055 96.750 ;
        RECT 1136.725 96.735 1137.055 96.740 ;
      LAYER via3 ;
        RECT 1136.500 110.340 1136.820 110.660 ;
        RECT 1136.500 96.740 1136.820 97.060 ;
      LAYER met4 ;
        RECT 1136.495 110.335 1136.825 110.665 ;
        RECT 1136.510 97.065 1136.810 110.335 ;
        RECT 1136.495 96.735 1136.825 97.065 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1140.410 1590.080 1140.730 1590.140 ;
        RECT 1144.090 1590.080 1144.410 1590.140 ;
        RECT 1140.410 1589.940 1144.410 1590.080 ;
        RECT 1140.410 1589.880 1140.730 1589.940 ;
        RECT 1144.090 1589.880 1144.410 1589.940 ;
        RECT 1144.090 59.060 1144.410 59.120 ;
        RECT 2277.070 59.060 2277.390 59.120 ;
        RECT 1144.090 58.920 2277.390 59.060 ;
        RECT 1144.090 58.860 1144.410 58.920 ;
        RECT 2277.070 58.860 2277.390 58.920 ;
        RECT 2277.070 2.960 2277.390 3.020 ;
        RECT 2280.290 2.960 2280.610 3.020 ;
        RECT 2277.070 2.820 2280.610 2.960 ;
        RECT 2277.070 2.760 2277.390 2.820 ;
        RECT 2280.290 2.760 2280.610 2.820 ;
      LAYER via ;
        RECT 1140.440 1589.880 1140.700 1590.140 ;
        RECT 1144.120 1589.880 1144.380 1590.140 ;
        RECT 1144.120 58.860 1144.380 59.120 ;
        RECT 2277.100 58.860 2277.360 59.120 ;
        RECT 2277.100 2.760 2277.360 3.020 ;
        RECT 2280.320 2.760 2280.580 3.020 ;
      LAYER met2 ;
        RECT 1140.300 1600.380 1140.580 1604.000 ;
        RECT 1140.300 1600.000 1140.640 1600.380 ;
        RECT 1140.500 1590.170 1140.640 1600.000 ;
        RECT 1140.440 1589.850 1140.700 1590.170 ;
        RECT 1144.120 1589.850 1144.380 1590.170 ;
        RECT 1144.180 59.150 1144.320 1589.850 ;
        RECT 1144.120 58.830 1144.380 59.150 ;
        RECT 2277.100 58.830 2277.360 59.150 ;
        RECT 2277.160 3.050 2277.300 58.830 ;
        RECT 2277.100 2.730 2277.360 3.050 ;
        RECT 2280.320 2.730 2280.580 3.050 ;
        RECT 2280.380 2.400 2280.520 2.730 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1146.390 1590.080 1146.710 1590.140 ;
        RECT 1151.450 1590.080 1151.770 1590.140 ;
        RECT 1146.390 1589.940 1151.770 1590.080 ;
        RECT 1146.390 1589.880 1146.710 1589.940 ;
        RECT 1151.450 1589.880 1151.770 1589.940 ;
        RECT 1151.450 58.720 1151.770 58.780 ;
        RECT 2298.230 58.720 2298.550 58.780 ;
        RECT 1151.450 58.580 2298.550 58.720 ;
        RECT 1151.450 58.520 1151.770 58.580 ;
        RECT 2298.230 58.520 2298.550 58.580 ;
      LAYER via ;
        RECT 1146.420 1589.880 1146.680 1590.140 ;
        RECT 1151.480 1589.880 1151.740 1590.140 ;
        RECT 1151.480 58.520 1151.740 58.780 ;
        RECT 2298.260 58.520 2298.520 58.780 ;
      LAYER met2 ;
        RECT 1146.280 1600.380 1146.560 1604.000 ;
        RECT 1146.280 1600.000 1146.620 1600.380 ;
        RECT 1146.480 1590.170 1146.620 1600.000 ;
        RECT 1146.420 1589.850 1146.680 1590.170 ;
        RECT 1151.480 1589.850 1151.740 1590.170 ;
        RECT 1151.540 58.810 1151.680 1589.850 ;
        RECT 1151.480 58.490 1151.740 58.810 ;
        RECT 2298.260 58.490 2298.520 58.810 ;
        RECT 2298.320 2.400 2298.460 58.490 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1152.830 1576.820 1153.150 1576.880 ;
        RECT 1157.430 1576.820 1157.750 1576.880 ;
        RECT 1152.830 1576.680 1157.750 1576.820 ;
        RECT 1152.830 1576.620 1153.150 1576.680 ;
        RECT 1157.430 1576.620 1157.750 1576.680 ;
        RECT 2311.570 2.960 2311.890 3.020 ;
        RECT 2316.170 2.960 2316.490 3.020 ;
        RECT 2311.570 2.820 2316.490 2.960 ;
        RECT 2311.570 2.760 2311.890 2.820 ;
        RECT 2316.170 2.760 2316.490 2.820 ;
      LAYER via ;
        RECT 1152.860 1576.620 1153.120 1576.880 ;
        RECT 1157.460 1576.620 1157.720 1576.880 ;
        RECT 2311.600 2.760 2311.860 3.020 ;
        RECT 2316.200 2.760 2316.460 3.020 ;
      LAYER met2 ;
        RECT 1152.720 1600.380 1153.000 1604.000 ;
        RECT 1152.720 1600.000 1153.060 1600.380 ;
        RECT 1152.920 1576.910 1153.060 1600.000 ;
        RECT 1152.860 1576.590 1153.120 1576.910 ;
        RECT 1157.460 1576.590 1157.720 1576.910 ;
        RECT 1157.520 61.725 1157.660 1576.590 ;
        RECT 1157.450 61.355 1157.730 61.725 ;
        RECT 2311.590 61.355 2311.870 61.725 ;
        RECT 2311.660 3.050 2311.800 61.355 ;
        RECT 2311.600 2.730 2311.860 3.050 ;
        RECT 2316.200 2.730 2316.460 3.050 ;
        RECT 2316.260 2.400 2316.400 2.730 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
      LAYER via2 ;
        RECT 1157.450 61.400 1157.730 61.680 ;
        RECT 2311.590 61.400 2311.870 61.680 ;
      LAYER met3 ;
        RECT 1157.425 61.690 1157.755 61.705 ;
        RECT 2311.565 61.690 2311.895 61.705 ;
        RECT 1157.425 61.390 2311.895 61.690 ;
        RECT 1157.425 61.375 1157.755 61.390 ;
        RECT 2311.565 61.375 2311.895 61.390 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1153.290 1600.960 1153.610 1601.020 ;
        RECT 1157.430 1600.960 1157.750 1601.020 ;
        RECT 1153.290 1600.820 1157.750 1600.960 ;
        RECT 1153.290 1600.760 1153.610 1600.820 ;
        RECT 1157.430 1600.760 1157.750 1600.820 ;
        RECT 1152.830 1535.340 1153.150 1535.400 ;
        RECT 1157.890 1535.340 1158.210 1535.400 ;
        RECT 1152.830 1535.200 1158.210 1535.340 ;
        RECT 1152.830 1535.140 1153.150 1535.200 ;
        RECT 1157.890 1535.140 1158.210 1535.200 ;
        RECT 2332.270 2.960 2332.590 3.020 ;
        RECT 2334.110 2.960 2334.430 3.020 ;
        RECT 2332.270 2.820 2334.430 2.960 ;
        RECT 2332.270 2.760 2332.590 2.820 ;
        RECT 2334.110 2.760 2334.430 2.820 ;
      LAYER via ;
        RECT 1153.320 1600.760 1153.580 1601.020 ;
        RECT 1157.460 1600.760 1157.720 1601.020 ;
        RECT 1152.860 1535.140 1153.120 1535.400 ;
        RECT 1157.920 1535.140 1158.180 1535.400 ;
        RECT 2332.300 2.760 2332.560 3.020 ;
        RECT 2334.140 2.760 2334.400 3.020 ;
      LAYER met2 ;
        RECT 1158.700 1601.130 1158.980 1604.000 ;
        RECT 1157.520 1601.050 1158.980 1601.130 ;
        RECT 1153.320 1600.730 1153.580 1601.050 ;
        RECT 1157.460 1600.990 1158.980 1601.050 ;
        RECT 1157.460 1600.730 1157.720 1600.990 ;
        RECT 1153.380 1569.170 1153.520 1600.730 ;
        RECT 1158.700 1600.000 1158.980 1600.990 ;
        RECT 1152.920 1569.030 1153.520 1569.170 ;
        RECT 1152.920 1535.430 1153.060 1569.030 ;
        RECT 1152.860 1535.110 1153.120 1535.430 ;
        RECT 1157.920 1535.110 1158.180 1535.430 ;
        RECT 1157.980 61.045 1158.120 1535.110 ;
        RECT 1157.910 60.675 1158.190 61.045 ;
        RECT 2332.290 60.675 2332.570 61.045 ;
        RECT 2332.360 3.050 2332.500 60.675 ;
        RECT 2332.300 2.730 2332.560 3.050 ;
        RECT 2334.140 2.730 2334.400 3.050 ;
        RECT 2334.200 2.400 2334.340 2.730 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
      LAYER via2 ;
        RECT 1157.910 60.720 1158.190 61.000 ;
        RECT 2332.290 60.720 2332.570 61.000 ;
      LAYER met3 ;
        RECT 1157.885 61.010 1158.215 61.025 ;
        RECT 2332.265 61.010 2332.595 61.025 ;
        RECT 1157.885 60.710 2332.595 61.010 ;
        RECT 1157.885 60.695 1158.215 60.710 ;
        RECT 2332.265 60.695 2332.595 60.710 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1159.270 1590.080 1159.590 1590.140 ;
        RECT 1165.250 1590.080 1165.570 1590.140 ;
        RECT 1159.270 1589.940 1165.570 1590.080 ;
        RECT 1159.270 1589.880 1159.590 1589.940 ;
        RECT 1165.250 1589.880 1165.570 1589.940 ;
        RECT 1159.270 1535.340 1159.590 1535.400 ;
        RECT 1165.250 1535.340 1165.570 1535.400 ;
        RECT 1159.270 1535.200 1165.570 1535.340 ;
        RECT 1159.270 1535.140 1159.590 1535.200 ;
        RECT 1165.250 1535.140 1165.570 1535.200 ;
        RECT 2346.070 2.960 2346.390 3.020 ;
        RECT 2351.590 2.960 2351.910 3.020 ;
        RECT 2346.070 2.820 2351.910 2.960 ;
        RECT 2346.070 2.760 2346.390 2.820 ;
        RECT 2351.590 2.760 2351.910 2.820 ;
      LAYER via ;
        RECT 1159.300 1589.880 1159.560 1590.140 ;
        RECT 1165.280 1589.880 1165.540 1590.140 ;
        RECT 1159.300 1535.140 1159.560 1535.400 ;
        RECT 1165.280 1535.140 1165.540 1535.400 ;
        RECT 2346.100 2.760 2346.360 3.020 ;
        RECT 2351.620 2.760 2351.880 3.020 ;
      LAYER met2 ;
        RECT 1165.140 1600.380 1165.420 1604.000 ;
        RECT 1165.140 1600.000 1165.480 1600.380 ;
        RECT 1165.340 1590.170 1165.480 1600.000 ;
        RECT 1159.300 1589.850 1159.560 1590.170 ;
        RECT 1165.280 1589.850 1165.540 1590.170 ;
        RECT 1159.360 1535.430 1159.500 1589.850 ;
        RECT 1159.300 1535.110 1159.560 1535.430 ;
        RECT 1165.280 1535.110 1165.540 1535.430 ;
        RECT 1165.340 60.365 1165.480 1535.110 ;
        RECT 1165.270 59.995 1165.550 60.365 ;
        RECT 2346.090 59.995 2346.370 60.365 ;
        RECT 2346.160 3.050 2346.300 59.995 ;
        RECT 2346.100 2.730 2346.360 3.050 ;
        RECT 2351.620 2.730 2351.880 3.050 ;
        RECT 2351.680 2.400 2351.820 2.730 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
      LAYER via2 ;
        RECT 1165.270 60.040 1165.550 60.320 ;
        RECT 2346.090 60.040 2346.370 60.320 ;
      LAYER met3 ;
        RECT 1165.245 60.330 1165.575 60.345 ;
        RECT 2346.065 60.330 2346.395 60.345 ;
        RECT 1165.245 60.030 2346.395 60.330 ;
        RECT 1165.245 60.015 1165.575 60.030 ;
        RECT 2346.065 60.015 2346.395 60.030 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1170.385 1304.325 1170.555 1352.095 ;
        RECT 1169.005 1041.845 1169.175 1083.155 ;
        RECT 1170.845 758.965 1171.015 807.075 ;
        RECT 1170.845 620.925 1171.015 710.515 ;
        RECT 1171.305 572.985 1171.475 596.955 ;
        RECT 1170.845 524.365 1171.015 572.475 ;
        RECT 1170.845 476.085 1171.015 500.395 ;
        RECT 1170.845 435.285 1171.015 458.915 ;
        RECT 1170.845 379.525 1171.015 427.635 ;
        RECT 1170.385 289.085 1170.555 331.075 ;
        RECT 1170.385 193.205 1170.555 234.515 ;
      LAYER mcon ;
        RECT 1170.385 1351.925 1170.555 1352.095 ;
        RECT 1169.005 1082.985 1169.175 1083.155 ;
        RECT 1170.845 806.905 1171.015 807.075 ;
        RECT 1170.845 710.345 1171.015 710.515 ;
        RECT 1171.305 596.785 1171.475 596.955 ;
        RECT 1170.845 572.305 1171.015 572.475 ;
        RECT 1170.845 500.225 1171.015 500.395 ;
        RECT 1170.845 458.745 1171.015 458.915 ;
        RECT 1170.845 427.465 1171.015 427.635 ;
        RECT 1170.385 330.905 1170.555 331.075 ;
        RECT 1170.385 234.345 1170.555 234.515 ;
      LAYER met1 ;
        RECT 1166.630 1590.080 1166.950 1590.140 ;
        RECT 1171.230 1590.080 1171.550 1590.140 ;
        RECT 1166.630 1589.940 1171.550 1590.080 ;
        RECT 1166.630 1589.880 1166.950 1589.940 ;
        RECT 1171.230 1589.880 1171.550 1589.940 ;
        RECT 1166.630 1559.140 1166.950 1559.200 ;
        RECT 1171.690 1559.140 1172.010 1559.200 ;
        RECT 1166.630 1559.000 1172.010 1559.140 ;
        RECT 1166.630 1558.940 1166.950 1559.000 ;
        RECT 1171.690 1558.940 1172.010 1559.000 ;
        RECT 1171.230 1497.600 1171.550 1497.660 ;
        RECT 1171.690 1497.600 1172.010 1497.660 ;
        RECT 1171.230 1497.460 1172.010 1497.600 ;
        RECT 1171.230 1497.400 1171.550 1497.460 ;
        RECT 1171.690 1497.400 1172.010 1497.460 ;
        RECT 1169.850 1435.380 1170.170 1435.440 ;
        RECT 1170.310 1435.380 1170.630 1435.440 ;
        RECT 1169.850 1435.240 1170.630 1435.380 ;
        RECT 1169.850 1435.180 1170.170 1435.240 ;
        RECT 1170.310 1435.180 1170.630 1435.240 ;
        RECT 1170.325 1352.080 1170.615 1352.125 ;
        RECT 1170.770 1352.080 1171.090 1352.140 ;
        RECT 1170.325 1351.940 1171.090 1352.080 ;
        RECT 1170.325 1351.895 1170.615 1351.940 ;
        RECT 1170.770 1351.880 1171.090 1351.940 ;
        RECT 1170.310 1304.480 1170.630 1304.540 ;
        RECT 1170.115 1304.340 1170.630 1304.480 ;
        RECT 1170.310 1304.280 1170.630 1304.340 ;
        RECT 1170.310 1256.200 1170.630 1256.260 ;
        RECT 1170.770 1256.200 1171.090 1256.260 ;
        RECT 1170.310 1256.060 1171.090 1256.200 ;
        RECT 1170.310 1256.000 1170.630 1256.060 ;
        RECT 1170.770 1256.000 1171.090 1256.060 ;
        RECT 1170.310 1200.780 1170.630 1200.840 ;
        RECT 1170.770 1200.780 1171.090 1200.840 ;
        RECT 1170.310 1200.640 1171.090 1200.780 ;
        RECT 1170.310 1200.580 1170.630 1200.640 ;
        RECT 1170.770 1200.580 1171.090 1200.640 ;
        RECT 1170.310 1173.040 1170.630 1173.300 ;
        RECT 1170.400 1172.560 1170.540 1173.040 ;
        RECT 1170.770 1172.560 1171.090 1172.620 ;
        RECT 1170.400 1172.420 1171.090 1172.560 ;
        RECT 1170.770 1172.360 1171.090 1172.420 ;
        RECT 1170.770 1125.300 1171.090 1125.360 ;
        RECT 1170.400 1125.160 1171.090 1125.300 ;
        RECT 1170.400 1124.680 1170.540 1125.160 ;
        RECT 1170.770 1125.100 1171.090 1125.160 ;
        RECT 1170.310 1124.420 1170.630 1124.680 ;
        RECT 1168.930 1083.140 1169.250 1083.200 ;
        RECT 1168.735 1083.000 1169.250 1083.140 ;
        RECT 1168.930 1082.940 1169.250 1083.000 ;
        RECT 1168.930 1042.000 1169.250 1042.060 ;
        RECT 1168.735 1041.860 1169.250 1042.000 ;
        RECT 1168.930 1041.800 1169.250 1041.860 ;
        RECT 1168.930 1017.860 1169.250 1017.920 ;
        RECT 1171.690 1017.860 1172.010 1017.920 ;
        RECT 1168.930 1017.720 1172.010 1017.860 ;
        RECT 1168.930 1017.660 1169.250 1017.720 ;
        RECT 1171.690 1017.660 1172.010 1017.720 ;
        RECT 1170.770 814.200 1171.090 814.260 ;
        RECT 1171.690 814.200 1172.010 814.260 ;
        RECT 1170.770 814.060 1172.010 814.200 ;
        RECT 1170.770 814.000 1171.090 814.060 ;
        RECT 1171.690 814.000 1172.010 814.060 ;
        RECT 1170.770 807.060 1171.090 807.120 ;
        RECT 1170.575 806.920 1171.090 807.060 ;
        RECT 1170.770 806.860 1171.090 806.920 ;
        RECT 1170.770 759.120 1171.090 759.180 ;
        RECT 1170.575 758.980 1171.090 759.120 ;
        RECT 1170.770 758.920 1171.090 758.980 ;
        RECT 1170.770 724.580 1171.090 724.840 ;
        RECT 1170.860 724.100 1171.000 724.580 ;
        RECT 1171.230 724.100 1171.550 724.160 ;
        RECT 1170.860 723.960 1171.550 724.100 ;
        RECT 1171.230 723.900 1171.550 723.960 ;
        RECT 1170.785 710.500 1171.075 710.545 ;
        RECT 1171.230 710.500 1171.550 710.560 ;
        RECT 1170.785 710.360 1171.550 710.500 ;
        RECT 1170.785 710.315 1171.075 710.360 ;
        RECT 1171.230 710.300 1171.550 710.360 ;
        RECT 1170.785 621.080 1171.075 621.125 ;
        RECT 1171.230 621.080 1171.550 621.140 ;
        RECT 1170.785 620.940 1171.550 621.080 ;
        RECT 1170.785 620.895 1171.075 620.940 ;
        RECT 1171.230 620.880 1171.550 620.940 ;
        RECT 1171.230 596.940 1171.550 597.000 ;
        RECT 1171.035 596.800 1171.550 596.940 ;
        RECT 1171.230 596.740 1171.550 596.800 ;
        RECT 1170.310 573.140 1170.630 573.200 ;
        RECT 1171.245 573.140 1171.535 573.185 ;
        RECT 1170.310 573.000 1171.535 573.140 ;
        RECT 1170.310 572.940 1170.630 573.000 ;
        RECT 1171.245 572.955 1171.535 573.000 ;
        RECT 1170.770 572.460 1171.090 572.520 ;
        RECT 1170.575 572.320 1171.090 572.460 ;
        RECT 1170.770 572.260 1171.090 572.320 ;
        RECT 1170.785 524.520 1171.075 524.565 ;
        RECT 1171.230 524.520 1171.550 524.580 ;
        RECT 1170.785 524.380 1171.550 524.520 ;
        RECT 1170.785 524.335 1171.075 524.380 ;
        RECT 1171.230 524.320 1171.550 524.380 ;
        RECT 1170.785 500.380 1171.075 500.425 ;
        RECT 1171.230 500.380 1171.550 500.440 ;
        RECT 1170.785 500.240 1171.550 500.380 ;
        RECT 1170.785 500.195 1171.075 500.240 ;
        RECT 1171.230 500.180 1171.550 500.240 ;
        RECT 1170.770 476.240 1171.090 476.300 ;
        RECT 1170.575 476.100 1171.090 476.240 ;
        RECT 1170.770 476.040 1171.090 476.100 ;
        RECT 1170.770 458.900 1171.090 458.960 ;
        RECT 1170.575 458.760 1171.090 458.900 ;
        RECT 1170.770 458.700 1171.090 458.760 ;
        RECT 1170.785 435.440 1171.075 435.485 ;
        RECT 1171.690 435.440 1172.010 435.500 ;
        RECT 1170.785 435.300 1172.010 435.440 ;
        RECT 1170.785 435.255 1171.075 435.300 ;
        RECT 1171.690 435.240 1172.010 435.300 ;
        RECT 1170.785 427.620 1171.075 427.665 ;
        RECT 1171.230 427.620 1171.550 427.680 ;
        RECT 1170.785 427.480 1171.550 427.620 ;
        RECT 1170.785 427.435 1171.075 427.480 ;
        RECT 1171.230 427.420 1171.550 427.480 ;
        RECT 1170.770 379.680 1171.090 379.740 ;
        RECT 1170.575 379.540 1171.090 379.680 ;
        RECT 1170.770 379.480 1171.090 379.540 ;
        RECT 1170.310 338.200 1170.630 338.260 ;
        RECT 1171.230 338.200 1171.550 338.260 ;
        RECT 1170.310 338.060 1171.550 338.200 ;
        RECT 1170.310 338.000 1170.630 338.060 ;
        RECT 1171.230 338.000 1171.550 338.060 ;
        RECT 1170.310 331.060 1170.630 331.120 ;
        RECT 1170.115 330.920 1170.630 331.060 ;
        RECT 1170.310 330.860 1170.630 330.920 ;
        RECT 1170.325 289.240 1170.615 289.285 ;
        RECT 1171.230 289.240 1171.550 289.300 ;
        RECT 1170.325 289.100 1171.550 289.240 ;
        RECT 1170.325 289.055 1170.615 289.100 ;
        RECT 1171.230 289.040 1171.550 289.100 ;
        RECT 1170.310 241.640 1170.630 241.700 ;
        RECT 1171.230 241.640 1171.550 241.700 ;
        RECT 1170.310 241.500 1171.550 241.640 ;
        RECT 1170.310 241.440 1170.630 241.500 ;
        RECT 1171.230 241.440 1171.550 241.500 ;
        RECT 1170.310 234.500 1170.630 234.560 ;
        RECT 1170.115 234.360 1170.630 234.500 ;
        RECT 1170.310 234.300 1170.630 234.360 ;
        RECT 1170.310 193.360 1170.630 193.420 ;
        RECT 1170.115 193.220 1170.630 193.360 ;
        RECT 1170.310 193.160 1170.630 193.220 ;
        RECT 1171.690 96.460 1172.010 96.520 ;
        RECT 1173.070 96.460 1173.390 96.520 ;
        RECT 1171.690 96.320 1173.390 96.460 ;
        RECT 1171.690 96.260 1172.010 96.320 ;
        RECT 1173.070 96.260 1173.390 96.320 ;
      LAYER via ;
        RECT 1166.660 1589.880 1166.920 1590.140 ;
        RECT 1171.260 1589.880 1171.520 1590.140 ;
        RECT 1166.660 1558.940 1166.920 1559.200 ;
        RECT 1171.720 1558.940 1171.980 1559.200 ;
        RECT 1171.260 1497.400 1171.520 1497.660 ;
        RECT 1171.720 1497.400 1171.980 1497.660 ;
        RECT 1169.880 1435.180 1170.140 1435.440 ;
        RECT 1170.340 1435.180 1170.600 1435.440 ;
        RECT 1170.800 1351.880 1171.060 1352.140 ;
        RECT 1170.340 1304.280 1170.600 1304.540 ;
        RECT 1170.340 1256.000 1170.600 1256.260 ;
        RECT 1170.800 1256.000 1171.060 1256.260 ;
        RECT 1170.340 1200.580 1170.600 1200.840 ;
        RECT 1170.800 1200.580 1171.060 1200.840 ;
        RECT 1170.340 1173.040 1170.600 1173.300 ;
        RECT 1170.800 1172.360 1171.060 1172.620 ;
        RECT 1170.800 1125.100 1171.060 1125.360 ;
        RECT 1170.340 1124.420 1170.600 1124.680 ;
        RECT 1168.960 1082.940 1169.220 1083.200 ;
        RECT 1168.960 1041.800 1169.220 1042.060 ;
        RECT 1168.960 1017.660 1169.220 1017.920 ;
        RECT 1171.720 1017.660 1171.980 1017.920 ;
        RECT 1170.800 814.000 1171.060 814.260 ;
        RECT 1171.720 814.000 1171.980 814.260 ;
        RECT 1170.800 806.860 1171.060 807.120 ;
        RECT 1170.800 758.920 1171.060 759.180 ;
        RECT 1170.800 724.580 1171.060 724.840 ;
        RECT 1171.260 723.900 1171.520 724.160 ;
        RECT 1171.260 710.300 1171.520 710.560 ;
        RECT 1171.260 620.880 1171.520 621.140 ;
        RECT 1171.260 596.740 1171.520 597.000 ;
        RECT 1170.340 572.940 1170.600 573.200 ;
        RECT 1170.800 572.260 1171.060 572.520 ;
        RECT 1171.260 524.320 1171.520 524.580 ;
        RECT 1171.260 500.180 1171.520 500.440 ;
        RECT 1170.800 476.040 1171.060 476.300 ;
        RECT 1170.800 458.700 1171.060 458.960 ;
        RECT 1171.720 435.240 1171.980 435.500 ;
        RECT 1171.260 427.420 1171.520 427.680 ;
        RECT 1170.800 379.480 1171.060 379.740 ;
        RECT 1170.340 338.000 1170.600 338.260 ;
        RECT 1171.260 338.000 1171.520 338.260 ;
        RECT 1170.340 330.860 1170.600 331.120 ;
        RECT 1171.260 289.040 1171.520 289.300 ;
        RECT 1170.340 241.440 1170.600 241.700 ;
        RECT 1171.260 241.440 1171.520 241.700 ;
        RECT 1170.340 234.300 1170.600 234.560 ;
        RECT 1170.340 193.160 1170.600 193.420 ;
        RECT 1171.720 96.260 1171.980 96.520 ;
        RECT 1173.100 96.260 1173.360 96.520 ;
      LAYER met2 ;
        RECT 1171.120 1600.380 1171.400 1604.000 ;
        RECT 1171.120 1600.000 1171.460 1600.380 ;
        RECT 1171.320 1590.170 1171.460 1600.000 ;
        RECT 1166.660 1589.850 1166.920 1590.170 ;
        RECT 1171.260 1589.850 1171.520 1590.170 ;
        RECT 1166.720 1559.230 1166.860 1589.850 ;
        RECT 1166.660 1558.910 1166.920 1559.230 ;
        RECT 1171.720 1558.910 1171.980 1559.230 ;
        RECT 1171.780 1497.690 1171.920 1558.910 ;
        RECT 1171.260 1497.370 1171.520 1497.690 ;
        RECT 1171.720 1497.370 1171.980 1497.690 ;
        RECT 1171.320 1483.605 1171.460 1497.370 ;
        RECT 1169.870 1483.235 1170.150 1483.605 ;
        RECT 1171.250 1483.235 1171.530 1483.605 ;
        RECT 1169.940 1435.470 1170.080 1483.235 ;
        RECT 1169.880 1435.150 1170.140 1435.470 ;
        RECT 1170.340 1435.150 1170.600 1435.470 ;
        RECT 1170.400 1418.210 1170.540 1435.150 ;
        RECT 1170.400 1418.070 1171.000 1418.210 ;
        RECT 1170.860 1352.170 1171.000 1418.070 ;
        RECT 1170.800 1351.850 1171.060 1352.170 ;
        RECT 1170.340 1304.250 1170.600 1304.570 ;
        RECT 1170.400 1256.290 1170.540 1304.250 ;
        RECT 1170.340 1255.970 1170.600 1256.290 ;
        RECT 1170.800 1255.970 1171.060 1256.290 ;
        RECT 1170.860 1200.870 1171.000 1255.970 ;
        RECT 1170.340 1200.550 1170.600 1200.870 ;
        RECT 1170.800 1200.550 1171.060 1200.870 ;
        RECT 1170.400 1173.330 1170.540 1200.550 ;
        RECT 1170.340 1173.010 1170.600 1173.330 ;
        RECT 1170.800 1172.330 1171.060 1172.650 ;
        RECT 1170.860 1125.390 1171.000 1172.330 ;
        RECT 1170.800 1125.070 1171.060 1125.390 ;
        RECT 1170.340 1124.390 1170.600 1124.710 ;
        RECT 1170.400 1089.885 1170.540 1124.390 ;
        RECT 1168.950 1089.515 1169.230 1089.885 ;
        RECT 1170.330 1089.515 1170.610 1089.885 ;
        RECT 1169.020 1083.230 1169.160 1089.515 ;
        RECT 1168.960 1082.910 1169.220 1083.230 ;
        RECT 1168.960 1041.770 1169.220 1042.090 ;
        RECT 1169.020 1017.950 1169.160 1041.770 ;
        RECT 1168.960 1017.630 1169.220 1017.950 ;
        RECT 1171.720 1017.630 1171.980 1017.950 ;
        RECT 1171.780 893.250 1171.920 1017.630 ;
        RECT 1170.860 893.110 1171.920 893.250 ;
        RECT 1170.860 869.565 1171.000 893.110 ;
        RECT 1170.790 869.195 1171.070 869.565 ;
        RECT 1171.710 869.195 1171.990 869.565 ;
        RECT 1171.780 814.290 1171.920 869.195 ;
        RECT 1170.800 813.970 1171.060 814.290 ;
        RECT 1171.720 813.970 1171.980 814.290 ;
        RECT 1170.860 807.150 1171.000 813.970 ;
        RECT 1170.800 806.830 1171.060 807.150 ;
        RECT 1170.800 758.890 1171.060 759.210 ;
        RECT 1170.860 724.870 1171.000 758.890 ;
        RECT 1170.800 724.550 1171.060 724.870 ;
        RECT 1171.260 723.870 1171.520 724.190 ;
        RECT 1171.320 710.590 1171.460 723.870 ;
        RECT 1171.260 710.270 1171.520 710.590 ;
        RECT 1171.260 620.850 1171.520 621.170 ;
        RECT 1171.320 597.030 1171.460 620.850 ;
        RECT 1171.260 596.710 1171.520 597.030 ;
        RECT 1170.340 572.970 1170.600 573.230 ;
        RECT 1170.340 572.910 1171.000 572.970 ;
        RECT 1170.400 572.830 1171.000 572.910 ;
        RECT 1170.860 572.550 1171.000 572.830 ;
        RECT 1170.800 572.230 1171.060 572.550 ;
        RECT 1171.260 524.290 1171.520 524.610 ;
        RECT 1171.320 500.470 1171.460 524.290 ;
        RECT 1171.260 500.150 1171.520 500.470 ;
        RECT 1170.800 476.010 1171.060 476.330 ;
        RECT 1170.860 458.990 1171.000 476.010 ;
        RECT 1170.800 458.670 1171.060 458.990 ;
        RECT 1171.720 435.210 1171.980 435.530 ;
        RECT 1171.780 434.930 1171.920 435.210 ;
        RECT 1171.320 434.790 1171.920 434.930 ;
        RECT 1171.320 427.710 1171.460 434.790 ;
        RECT 1171.260 427.390 1171.520 427.710 ;
        RECT 1170.800 379.450 1171.060 379.770 ;
        RECT 1170.860 352.650 1171.000 379.450 ;
        RECT 1170.860 352.510 1171.460 352.650 ;
        RECT 1171.320 338.290 1171.460 352.510 ;
        RECT 1170.340 337.970 1170.600 338.290 ;
        RECT 1171.260 337.970 1171.520 338.290 ;
        RECT 1170.400 331.150 1170.540 337.970 ;
        RECT 1170.340 330.830 1170.600 331.150 ;
        RECT 1171.260 289.010 1171.520 289.330 ;
        RECT 1171.320 241.730 1171.460 289.010 ;
        RECT 1170.340 241.410 1170.600 241.730 ;
        RECT 1171.260 241.410 1171.520 241.730 ;
        RECT 1170.400 234.590 1170.540 241.410 ;
        RECT 1170.340 234.270 1170.600 234.590 ;
        RECT 1170.340 193.130 1170.600 193.450 ;
        RECT 1170.400 158.170 1170.540 193.130 ;
        RECT 1170.400 158.030 1171.460 158.170 ;
        RECT 1171.320 110.570 1171.460 158.030 ;
        RECT 1171.320 110.430 1171.920 110.570 ;
        RECT 1171.780 96.550 1171.920 110.430 ;
        RECT 1171.720 96.230 1171.980 96.550 ;
        RECT 1173.100 96.230 1173.360 96.550 ;
        RECT 1173.160 59.685 1173.300 96.230 ;
        RECT 1173.090 59.315 1173.370 59.685 ;
        RECT 2366.790 59.315 2367.070 59.685 ;
        RECT 2366.860 3.130 2367.000 59.315 ;
        RECT 2366.860 2.990 2369.300 3.130 ;
        RECT 2369.160 2.960 2369.300 2.990 ;
        RECT 2369.160 2.820 2369.760 2.960 ;
        RECT 2369.620 2.400 2369.760 2.820 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
      LAYER via2 ;
        RECT 1169.870 1483.280 1170.150 1483.560 ;
        RECT 1171.250 1483.280 1171.530 1483.560 ;
        RECT 1168.950 1089.560 1169.230 1089.840 ;
        RECT 1170.330 1089.560 1170.610 1089.840 ;
        RECT 1170.790 869.240 1171.070 869.520 ;
        RECT 1171.710 869.240 1171.990 869.520 ;
        RECT 1173.090 59.360 1173.370 59.640 ;
        RECT 2366.790 59.360 2367.070 59.640 ;
      LAYER met3 ;
        RECT 1169.845 1483.570 1170.175 1483.585 ;
        RECT 1171.225 1483.570 1171.555 1483.585 ;
        RECT 1169.845 1483.270 1171.555 1483.570 ;
        RECT 1169.845 1483.255 1170.175 1483.270 ;
        RECT 1171.225 1483.255 1171.555 1483.270 ;
        RECT 1168.925 1089.850 1169.255 1089.865 ;
        RECT 1170.305 1089.850 1170.635 1089.865 ;
        RECT 1168.925 1089.550 1170.635 1089.850 ;
        RECT 1168.925 1089.535 1169.255 1089.550 ;
        RECT 1170.305 1089.535 1170.635 1089.550 ;
        RECT 1170.765 869.530 1171.095 869.545 ;
        RECT 1171.685 869.530 1172.015 869.545 ;
        RECT 1170.765 869.230 1172.015 869.530 ;
        RECT 1170.765 869.215 1171.095 869.230 ;
        RECT 1171.685 869.215 1172.015 869.230 ;
        RECT 1173.065 59.650 1173.395 59.665 ;
        RECT 2366.765 59.650 2367.095 59.665 ;
        RECT 1173.065 59.350 2367.095 59.650 ;
        RECT 1173.065 59.335 1173.395 59.350 ;
        RECT 2366.765 59.335 2367.095 59.350 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1178.130 1600.960 1178.450 1601.020 ;
        RECT 1177.300 1600.820 1178.450 1600.960 ;
        RECT 1177.300 1599.660 1177.440 1600.820 ;
        RECT 1178.130 1600.760 1178.450 1600.820 ;
        RECT 1177.210 1599.400 1177.530 1599.660 ;
        RECT 1173.070 1579.880 1173.390 1579.940 ;
        RECT 1177.210 1579.880 1177.530 1579.940 ;
        RECT 1173.070 1579.740 1177.530 1579.880 ;
        RECT 1173.070 1579.680 1173.390 1579.740 ;
        RECT 1177.210 1579.680 1177.530 1579.740 ;
        RECT 1173.070 1535.340 1173.390 1535.400 ;
        RECT 1179.050 1535.340 1179.370 1535.400 ;
        RECT 1173.070 1535.200 1179.370 1535.340 ;
        RECT 1173.070 1535.140 1173.390 1535.200 ;
        RECT 1179.050 1535.140 1179.370 1535.200 ;
      LAYER via ;
        RECT 1178.160 1600.760 1178.420 1601.020 ;
        RECT 1177.240 1599.400 1177.500 1599.660 ;
        RECT 1173.100 1579.680 1173.360 1579.940 ;
        RECT 1177.240 1579.680 1177.500 1579.940 ;
        RECT 1173.100 1535.140 1173.360 1535.400 ;
        RECT 1179.080 1535.140 1179.340 1535.400 ;
      LAYER met2 ;
        RECT 1177.560 1601.130 1177.840 1604.000 ;
        RECT 1177.560 1601.050 1178.360 1601.130 ;
        RECT 1177.560 1600.990 1178.420 1601.050 ;
        RECT 1177.560 1600.000 1177.840 1600.990 ;
        RECT 1178.160 1600.730 1178.420 1600.990 ;
        RECT 1177.240 1599.370 1177.500 1599.690 ;
        RECT 1177.300 1579.970 1177.440 1599.370 ;
        RECT 1173.100 1579.650 1173.360 1579.970 ;
        RECT 1177.240 1579.650 1177.500 1579.970 ;
        RECT 1173.160 1535.430 1173.300 1579.650 ;
        RECT 1173.100 1535.110 1173.360 1535.430 ;
        RECT 1179.080 1535.110 1179.340 1535.430 ;
        RECT 1179.140 59.005 1179.280 1535.110 ;
        RECT 1179.070 58.635 1179.350 59.005 ;
        RECT 2387.950 58.635 2388.230 59.005 ;
        RECT 2388.020 17.410 2388.160 58.635 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.400 2387.700 17.270 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
      LAYER via2 ;
        RECT 1179.070 58.680 1179.350 58.960 ;
        RECT 2387.950 58.680 2388.230 58.960 ;
      LAYER met3 ;
        RECT 1179.045 58.970 1179.375 58.985 ;
        RECT 2387.925 58.970 2388.255 58.985 ;
        RECT 1179.045 58.670 2388.255 58.970 ;
        RECT 1179.045 58.655 1179.375 58.670 ;
        RECT 2387.925 58.655 2388.255 58.670 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1179.970 1579.880 1180.290 1579.940 ;
        RECT 1182.270 1579.880 1182.590 1579.940 ;
        RECT 1179.970 1579.740 1182.590 1579.880 ;
        RECT 1179.970 1579.680 1180.290 1579.740 ;
        RECT 1182.270 1579.680 1182.590 1579.740 ;
        RECT 1179.970 1535.340 1180.290 1535.400 ;
        RECT 1186.410 1535.340 1186.730 1535.400 ;
        RECT 1179.970 1535.200 1186.730 1535.340 ;
        RECT 1179.970 1535.140 1180.290 1535.200 ;
        RECT 1186.410 1535.140 1186.730 1535.200 ;
      LAYER via ;
        RECT 1180.000 1579.680 1180.260 1579.940 ;
        RECT 1182.300 1579.680 1182.560 1579.940 ;
        RECT 1180.000 1535.140 1180.260 1535.400 ;
        RECT 1186.440 1535.140 1186.700 1535.400 ;
      LAYER met2 ;
        RECT 1183.540 1600.450 1183.820 1604.000 ;
        RECT 1182.360 1600.310 1183.820 1600.450 ;
        RECT 1182.360 1579.970 1182.500 1600.310 ;
        RECT 1183.540 1600.000 1183.820 1600.310 ;
        RECT 1180.000 1579.650 1180.260 1579.970 ;
        RECT 1182.300 1579.650 1182.560 1579.970 ;
        RECT 1180.060 1535.430 1180.200 1579.650 ;
        RECT 1180.000 1535.110 1180.260 1535.430 ;
        RECT 1186.440 1535.110 1186.700 1535.430 ;
        RECT 1186.500 58.325 1186.640 1535.110 ;
        RECT 1186.430 57.955 1186.710 58.325 ;
        RECT 2401.290 57.955 2401.570 58.325 ;
        RECT 2401.360 17.410 2401.500 57.955 ;
        RECT 2401.360 17.270 2405.640 17.410 ;
        RECT 2405.500 2.400 2405.640 17.270 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
      LAYER via2 ;
        RECT 1186.430 58.000 1186.710 58.280 ;
        RECT 2401.290 58.000 2401.570 58.280 ;
      LAYER met3 ;
        RECT 1186.405 58.290 1186.735 58.305 ;
        RECT 2401.265 58.290 2401.595 58.305 ;
        RECT 1186.405 57.990 2401.595 58.290 ;
        RECT 1186.405 57.975 1186.735 57.990 ;
        RECT 2401.265 57.975 2401.595 57.990 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 626.940 1600.380 627.220 1604.000 ;
        RECT 626.940 1600.000 627.280 1600.380 ;
        RECT 627.140 20.130 627.280 1600.000 ;
        RECT 626.680 19.990 627.280 20.130 ;
        RECT 626.680 16.165 626.820 19.990 ;
        RECT 626.610 15.795 626.890 16.165 ;
        RECT 799.570 15.795 799.850 16.165 ;
        RECT 799.640 2.400 799.780 15.795 ;
        RECT 799.430 -4.800 799.990 2.400 ;
      LAYER via2 ;
        RECT 626.610 15.840 626.890 16.120 ;
        RECT 799.570 15.840 799.850 16.120 ;
      LAYER met3 ;
        RECT 626.585 16.130 626.915 16.145 ;
        RECT 799.545 16.130 799.875 16.145 ;
        RECT 626.585 15.830 799.875 16.130 ;
        RECT 626.585 15.815 626.915 15.830 ;
        RECT 799.545 15.815 799.875 15.830 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 637.245 19.805 639.255 19.975 ;
      LAYER mcon ;
        RECT 639.085 19.805 639.255 19.975 ;
      LAYER met1 ;
        RECT 573.690 1590.420 574.010 1590.480 ;
        RECT 578.290 1590.420 578.610 1590.480 ;
        RECT 573.690 1590.280 578.610 1590.420 ;
        RECT 573.690 1590.220 574.010 1590.280 ;
        RECT 578.290 1590.220 578.610 1590.280 ;
        RECT 578.290 19.960 578.610 20.020 ;
        RECT 637.185 19.960 637.475 20.005 ;
        RECT 578.290 19.820 637.475 19.960 ;
        RECT 578.290 19.760 578.610 19.820 ;
        RECT 637.185 19.775 637.475 19.820 ;
        RECT 639.025 19.960 639.315 20.005 ;
        RECT 644.990 19.960 645.310 20.020 ;
        RECT 639.025 19.820 645.310 19.960 ;
        RECT 639.025 19.775 639.315 19.820 ;
        RECT 644.990 19.760 645.310 19.820 ;
      LAYER via ;
        RECT 573.720 1590.220 573.980 1590.480 ;
        RECT 578.320 1590.220 578.580 1590.480 ;
        RECT 578.320 19.760 578.580 20.020 ;
        RECT 645.020 19.760 645.280 20.020 ;
      LAYER met2 ;
        RECT 573.580 1600.380 573.860 1604.000 ;
        RECT 573.580 1600.000 573.920 1600.380 ;
        RECT 573.780 1590.510 573.920 1600.000 ;
        RECT 573.720 1590.190 573.980 1590.510 ;
        RECT 578.320 1590.190 578.580 1590.510 ;
        RECT 578.380 20.050 578.520 1590.190 ;
        RECT 578.320 19.730 578.580 20.050 ;
        RECT 645.020 19.730 645.280 20.050 ;
        RECT 645.080 2.400 645.220 19.730 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1187.330 1579.880 1187.650 1579.940 ;
        RECT 1190.550 1579.880 1190.870 1579.940 ;
        RECT 1187.330 1579.740 1190.870 1579.880 ;
        RECT 1187.330 1579.680 1187.650 1579.740 ;
        RECT 1190.550 1579.680 1190.870 1579.740 ;
        RECT 1187.330 1510.860 1187.650 1510.920 ;
        RECT 1191.930 1510.860 1192.250 1510.920 ;
        RECT 1187.330 1510.720 1192.250 1510.860 ;
        RECT 1187.330 1510.660 1187.650 1510.720 ;
        RECT 1191.930 1510.660 1192.250 1510.720 ;
        RECT 1191.930 72.660 1192.250 72.720 ;
        RECT 2428.870 72.660 2429.190 72.720 ;
        RECT 1191.930 72.520 2429.190 72.660 ;
        RECT 1191.930 72.460 1192.250 72.520 ;
        RECT 2428.870 72.460 2429.190 72.520 ;
      LAYER via ;
        RECT 1187.360 1579.680 1187.620 1579.940 ;
        RECT 1190.580 1579.680 1190.840 1579.940 ;
        RECT 1187.360 1510.660 1187.620 1510.920 ;
        RECT 1191.960 1510.660 1192.220 1510.920 ;
        RECT 1191.960 72.460 1192.220 72.720 ;
        RECT 2428.900 72.460 2429.160 72.720 ;
      LAYER met2 ;
        RECT 1191.820 1600.450 1192.100 1604.000 ;
        RECT 1190.640 1600.310 1192.100 1600.450 ;
        RECT 1190.640 1579.970 1190.780 1600.310 ;
        RECT 1191.820 1600.000 1192.100 1600.310 ;
        RECT 1187.360 1579.650 1187.620 1579.970 ;
        RECT 1190.580 1579.650 1190.840 1579.970 ;
        RECT 1187.420 1510.950 1187.560 1579.650 ;
        RECT 1187.360 1510.630 1187.620 1510.950 ;
        RECT 1191.960 1510.630 1192.220 1510.950 ;
        RECT 1192.020 1448.810 1192.160 1510.630 ;
        RECT 1192.020 1448.670 1192.620 1448.810 ;
        RECT 1192.480 134.370 1192.620 1448.670 ;
        RECT 1192.020 134.230 1192.620 134.370 ;
        RECT 1192.020 72.750 1192.160 134.230 ;
        RECT 1191.960 72.430 1192.220 72.750 ;
        RECT 2428.900 72.430 2429.160 72.750 ;
        RECT 2428.960 2.400 2429.100 72.430 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1193.770 1579.880 1194.090 1579.940 ;
        RECT 1196.530 1579.880 1196.850 1579.940 ;
        RECT 1193.770 1579.740 1196.850 1579.880 ;
        RECT 1193.770 1579.680 1194.090 1579.740 ;
        RECT 1196.530 1579.680 1196.850 1579.740 ;
        RECT 1193.770 1535.000 1194.090 1535.060 ;
        RECT 1200.210 1535.000 1200.530 1535.060 ;
        RECT 1193.770 1534.860 1200.530 1535.000 ;
        RECT 1193.770 1534.800 1194.090 1534.860 ;
        RECT 1200.210 1534.800 1200.530 1534.860 ;
        RECT 1200.210 63.480 1200.530 63.540 ;
        RECT 2442.670 63.480 2442.990 63.540 ;
        RECT 1200.210 63.340 2442.990 63.480 ;
        RECT 1200.210 63.280 1200.530 63.340 ;
        RECT 2442.670 63.280 2442.990 63.340 ;
      LAYER via ;
        RECT 1193.800 1579.680 1194.060 1579.940 ;
        RECT 1196.560 1579.680 1196.820 1579.940 ;
        RECT 1193.800 1534.800 1194.060 1535.060 ;
        RECT 1200.240 1534.800 1200.500 1535.060 ;
        RECT 1200.240 63.280 1200.500 63.540 ;
        RECT 2442.700 63.280 2442.960 63.540 ;
      LAYER met2 ;
        RECT 1197.800 1600.450 1198.080 1604.000 ;
        RECT 1196.620 1600.310 1198.080 1600.450 ;
        RECT 1196.620 1579.970 1196.760 1600.310 ;
        RECT 1197.800 1600.000 1198.080 1600.310 ;
        RECT 1193.800 1579.650 1194.060 1579.970 ;
        RECT 1196.560 1579.650 1196.820 1579.970 ;
        RECT 1193.860 1535.090 1194.000 1579.650 ;
        RECT 1193.800 1534.770 1194.060 1535.090 ;
        RECT 1200.240 1534.770 1200.500 1535.090 ;
        RECT 1200.300 63.570 1200.440 1534.770 ;
        RECT 1200.240 63.250 1200.500 63.570 ;
        RECT 2442.700 63.250 2442.960 63.570 ;
        RECT 2442.760 17.410 2442.900 63.250 ;
        RECT 2442.760 17.270 2447.040 17.410 ;
        RECT 2446.900 2.400 2447.040 17.270 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1202.510 1594.160 1202.830 1594.220 ;
        RECT 1204.350 1594.160 1204.670 1594.220 ;
        RECT 1202.510 1594.020 1204.670 1594.160 ;
        RECT 1202.510 1593.960 1202.830 1594.020 ;
        RECT 1204.350 1593.960 1204.670 1594.020 ;
        RECT 1202.510 1587.020 1202.830 1587.080 ;
        RECT 1206.190 1587.020 1206.510 1587.080 ;
        RECT 1202.510 1586.880 1206.510 1587.020 ;
        RECT 1202.510 1586.820 1202.830 1586.880 ;
        RECT 1206.190 1586.820 1206.510 1586.880 ;
        RECT 1205.730 63.820 1206.050 63.880 ;
        RECT 2463.370 63.820 2463.690 63.880 ;
        RECT 1205.730 63.680 2463.690 63.820 ;
        RECT 1205.730 63.620 1206.050 63.680 ;
        RECT 2463.370 63.620 2463.690 63.680 ;
      LAYER via ;
        RECT 1202.540 1593.960 1202.800 1594.220 ;
        RECT 1204.380 1593.960 1204.640 1594.220 ;
        RECT 1202.540 1586.820 1202.800 1587.080 ;
        RECT 1206.220 1586.820 1206.480 1587.080 ;
        RECT 1205.760 63.620 1206.020 63.880 ;
        RECT 2463.400 63.620 2463.660 63.880 ;
      LAYER met2 ;
        RECT 1204.240 1600.380 1204.520 1604.000 ;
        RECT 1204.240 1600.000 1204.580 1600.380 ;
        RECT 1204.440 1594.250 1204.580 1600.000 ;
        RECT 1202.540 1593.930 1202.800 1594.250 ;
        RECT 1204.380 1593.930 1204.640 1594.250 ;
        RECT 1202.600 1587.110 1202.740 1593.930 ;
        RECT 1202.540 1586.790 1202.800 1587.110 ;
        RECT 1206.220 1586.790 1206.480 1587.110 ;
        RECT 1206.280 1390.330 1206.420 1586.790 ;
        RECT 1205.820 1390.190 1206.420 1390.330 ;
        RECT 1205.820 63.910 1205.960 1390.190 ;
        RECT 1205.760 63.590 1206.020 63.910 ;
        RECT 2463.400 63.590 2463.660 63.910 ;
        RECT 2463.460 3.130 2463.600 63.590 ;
        RECT 2463.460 2.990 2464.520 3.130 ;
        RECT 2464.380 2.960 2464.520 2.990 ;
        RECT 2464.380 2.820 2464.980 2.960 ;
        RECT 2464.840 2.400 2464.980 2.820 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1213.165 1442.025 1213.335 1490.475 ;
        RECT 1212.705 814.385 1212.875 862.495 ;
        RECT 1212.705 717.825 1212.875 765.935 ;
        RECT 1212.705 620.925 1212.875 669.375 ;
        RECT 1212.705 524.365 1212.875 572.475 ;
        RECT 1212.705 427.805 1212.875 475.915 ;
        RECT 1212.705 331.245 1212.875 379.355 ;
        RECT 1212.705 234.685 1212.875 282.795 ;
        RECT 1212.705 138.125 1212.875 186.235 ;
      LAYER mcon ;
        RECT 1213.165 1490.305 1213.335 1490.475 ;
        RECT 1212.705 862.325 1212.875 862.495 ;
        RECT 1212.705 765.765 1212.875 765.935 ;
        RECT 1212.705 669.205 1212.875 669.375 ;
        RECT 1212.705 572.305 1212.875 572.475 ;
        RECT 1212.705 475.745 1212.875 475.915 ;
        RECT 1212.705 379.185 1212.875 379.355 ;
        RECT 1212.705 282.625 1212.875 282.795 ;
        RECT 1212.705 186.065 1212.875 186.235 ;
      LAYER met1 ;
        RECT 1208.030 1594.160 1208.350 1594.220 ;
        RECT 1210.330 1594.160 1210.650 1594.220 ;
        RECT 1208.030 1594.020 1210.650 1594.160 ;
        RECT 1208.030 1593.960 1208.350 1594.020 ;
        RECT 1210.330 1593.960 1210.650 1594.020 ;
        RECT 1208.030 1570.700 1208.350 1570.760 ;
        RECT 1213.090 1570.700 1213.410 1570.760 ;
        RECT 1208.030 1570.560 1213.410 1570.700 ;
        RECT 1208.030 1570.500 1208.350 1570.560 ;
        RECT 1213.090 1570.500 1213.410 1570.560 ;
        RECT 1213.090 1490.460 1213.410 1490.520 ;
        RECT 1212.895 1490.320 1213.410 1490.460 ;
        RECT 1213.090 1490.260 1213.410 1490.320 ;
        RECT 1213.090 1442.180 1213.410 1442.240 ;
        RECT 1212.895 1442.040 1213.410 1442.180 ;
        RECT 1213.090 1441.980 1213.410 1442.040 ;
        RECT 1212.630 1352.420 1212.950 1352.480 ;
        RECT 1213.090 1352.420 1213.410 1352.480 ;
        RECT 1212.630 1352.280 1213.410 1352.420 ;
        RECT 1212.630 1352.220 1212.950 1352.280 ;
        RECT 1213.090 1352.220 1213.410 1352.280 ;
        RECT 1211.710 1200.780 1212.030 1200.840 ;
        RECT 1212.630 1200.780 1212.950 1200.840 ;
        RECT 1211.710 1200.640 1212.950 1200.780 ;
        RECT 1211.710 1200.580 1212.030 1200.640 ;
        RECT 1212.630 1200.580 1212.950 1200.640 ;
        RECT 1211.710 1104.220 1212.030 1104.280 ;
        RECT 1212.630 1104.220 1212.950 1104.280 ;
        RECT 1211.710 1104.080 1212.950 1104.220 ;
        RECT 1211.710 1104.020 1212.030 1104.080 ;
        RECT 1212.630 1104.020 1212.950 1104.080 ;
        RECT 1211.710 1055.600 1212.030 1055.660 ;
        RECT 1212.630 1055.600 1212.950 1055.660 ;
        RECT 1211.710 1055.460 1212.950 1055.600 ;
        RECT 1211.710 1055.400 1212.030 1055.460 ;
        RECT 1212.630 1055.400 1212.950 1055.460 ;
        RECT 1211.710 959.040 1212.030 959.100 ;
        RECT 1212.630 959.040 1212.950 959.100 ;
        RECT 1211.710 958.900 1212.950 959.040 ;
        RECT 1211.710 958.840 1212.030 958.900 ;
        RECT 1212.630 958.840 1212.950 958.900 ;
        RECT 1212.630 862.480 1212.950 862.540 ;
        RECT 1212.435 862.340 1212.950 862.480 ;
        RECT 1212.630 862.280 1212.950 862.340 ;
        RECT 1212.630 814.540 1212.950 814.600 ;
        RECT 1212.435 814.400 1212.950 814.540 ;
        RECT 1212.630 814.340 1212.950 814.400 ;
        RECT 1212.630 765.920 1212.950 765.980 ;
        RECT 1212.435 765.780 1212.950 765.920 ;
        RECT 1212.630 765.720 1212.950 765.780 ;
        RECT 1212.630 717.980 1212.950 718.040 ;
        RECT 1212.435 717.840 1212.950 717.980 ;
        RECT 1212.630 717.780 1212.950 717.840 ;
        RECT 1212.630 669.360 1212.950 669.420 ;
        RECT 1212.435 669.220 1212.950 669.360 ;
        RECT 1212.630 669.160 1212.950 669.220 ;
        RECT 1212.630 621.080 1212.950 621.140 ;
        RECT 1212.435 620.940 1212.950 621.080 ;
        RECT 1212.630 620.880 1212.950 620.940 ;
        RECT 1212.630 572.460 1212.950 572.520 ;
        RECT 1212.435 572.320 1212.950 572.460 ;
        RECT 1212.630 572.260 1212.950 572.320 ;
        RECT 1212.630 524.520 1212.950 524.580 ;
        RECT 1212.435 524.380 1212.950 524.520 ;
        RECT 1212.630 524.320 1212.950 524.380 ;
        RECT 1212.630 475.900 1212.950 475.960 ;
        RECT 1212.435 475.760 1212.950 475.900 ;
        RECT 1212.630 475.700 1212.950 475.760 ;
        RECT 1212.630 427.960 1212.950 428.020 ;
        RECT 1212.435 427.820 1212.950 427.960 ;
        RECT 1212.630 427.760 1212.950 427.820 ;
        RECT 1212.630 379.340 1212.950 379.400 ;
        RECT 1212.435 379.200 1212.950 379.340 ;
        RECT 1212.630 379.140 1212.950 379.200 ;
        RECT 1212.630 331.400 1212.950 331.460 ;
        RECT 1212.435 331.260 1212.950 331.400 ;
        RECT 1212.630 331.200 1212.950 331.260 ;
        RECT 1212.630 282.780 1212.950 282.840 ;
        RECT 1212.435 282.640 1212.950 282.780 ;
        RECT 1212.630 282.580 1212.950 282.640 ;
        RECT 1212.630 234.840 1212.950 234.900 ;
        RECT 1212.435 234.700 1212.950 234.840 ;
        RECT 1212.630 234.640 1212.950 234.700 ;
        RECT 1212.630 186.220 1212.950 186.280 ;
        RECT 1212.435 186.080 1212.950 186.220 ;
        RECT 1212.630 186.020 1212.950 186.080 ;
        RECT 1212.630 138.280 1212.950 138.340 ;
        RECT 1212.435 138.140 1212.950 138.280 ;
        RECT 1212.630 138.080 1212.950 138.140 ;
        RECT 1212.170 64.160 1212.490 64.220 ;
        RECT 2477.170 64.160 2477.490 64.220 ;
        RECT 1212.170 64.020 2477.490 64.160 ;
        RECT 1212.170 63.960 1212.490 64.020 ;
        RECT 2477.170 63.960 2477.490 64.020 ;
        RECT 2477.170 2.960 2477.490 3.020 ;
        RECT 2482.690 2.960 2483.010 3.020 ;
        RECT 2477.170 2.820 2483.010 2.960 ;
        RECT 2477.170 2.760 2477.490 2.820 ;
        RECT 2482.690 2.760 2483.010 2.820 ;
      LAYER via ;
        RECT 1208.060 1593.960 1208.320 1594.220 ;
        RECT 1210.360 1593.960 1210.620 1594.220 ;
        RECT 1208.060 1570.500 1208.320 1570.760 ;
        RECT 1213.120 1570.500 1213.380 1570.760 ;
        RECT 1213.120 1490.260 1213.380 1490.520 ;
        RECT 1213.120 1441.980 1213.380 1442.240 ;
        RECT 1212.660 1352.220 1212.920 1352.480 ;
        RECT 1213.120 1352.220 1213.380 1352.480 ;
        RECT 1211.740 1200.580 1212.000 1200.840 ;
        RECT 1212.660 1200.580 1212.920 1200.840 ;
        RECT 1211.740 1104.020 1212.000 1104.280 ;
        RECT 1212.660 1104.020 1212.920 1104.280 ;
        RECT 1211.740 1055.400 1212.000 1055.660 ;
        RECT 1212.660 1055.400 1212.920 1055.660 ;
        RECT 1211.740 958.840 1212.000 959.100 ;
        RECT 1212.660 958.840 1212.920 959.100 ;
        RECT 1212.660 862.280 1212.920 862.540 ;
        RECT 1212.660 814.340 1212.920 814.600 ;
        RECT 1212.660 765.720 1212.920 765.980 ;
        RECT 1212.660 717.780 1212.920 718.040 ;
        RECT 1212.660 669.160 1212.920 669.420 ;
        RECT 1212.660 620.880 1212.920 621.140 ;
        RECT 1212.660 572.260 1212.920 572.520 ;
        RECT 1212.660 524.320 1212.920 524.580 ;
        RECT 1212.660 475.700 1212.920 475.960 ;
        RECT 1212.660 427.760 1212.920 428.020 ;
        RECT 1212.660 379.140 1212.920 379.400 ;
        RECT 1212.660 331.200 1212.920 331.460 ;
        RECT 1212.660 282.580 1212.920 282.840 ;
        RECT 1212.660 234.640 1212.920 234.900 ;
        RECT 1212.660 186.020 1212.920 186.280 ;
        RECT 1212.660 138.080 1212.920 138.340 ;
        RECT 1212.200 63.960 1212.460 64.220 ;
        RECT 2477.200 63.960 2477.460 64.220 ;
        RECT 2477.200 2.760 2477.460 3.020 ;
        RECT 2482.720 2.760 2482.980 3.020 ;
      LAYER met2 ;
        RECT 1210.220 1600.380 1210.500 1604.000 ;
        RECT 1210.220 1600.000 1210.560 1600.380 ;
        RECT 1210.420 1594.250 1210.560 1600.000 ;
        RECT 1208.060 1593.930 1208.320 1594.250 ;
        RECT 1210.360 1593.930 1210.620 1594.250 ;
        RECT 1208.120 1570.790 1208.260 1593.930 ;
        RECT 1208.060 1570.470 1208.320 1570.790 ;
        RECT 1213.120 1570.470 1213.380 1570.790 ;
        RECT 1213.180 1490.550 1213.320 1570.470 ;
        RECT 1213.120 1490.230 1213.380 1490.550 ;
        RECT 1213.120 1441.950 1213.380 1442.270 ;
        RECT 1213.180 1352.510 1213.320 1441.950 ;
        RECT 1212.660 1352.190 1212.920 1352.510 ;
        RECT 1213.120 1352.190 1213.380 1352.510 ;
        RECT 1212.720 1249.005 1212.860 1352.190 ;
        RECT 1211.730 1248.635 1212.010 1249.005 ;
        RECT 1212.650 1248.635 1212.930 1249.005 ;
        RECT 1211.800 1200.870 1211.940 1248.635 ;
        RECT 1211.740 1200.550 1212.000 1200.870 ;
        RECT 1212.660 1200.550 1212.920 1200.870 ;
        RECT 1212.720 1152.445 1212.860 1200.550 ;
        RECT 1211.730 1152.075 1212.010 1152.445 ;
        RECT 1212.650 1152.075 1212.930 1152.445 ;
        RECT 1211.800 1104.310 1211.940 1152.075 ;
        RECT 1211.740 1103.990 1212.000 1104.310 ;
        RECT 1212.660 1103.990 1212.920 1104.310 ;
        RECT 1212.720 1055.690 1212.860 1103.990 ;
        RECT 1211.740 1055.370 1212.000 1055.690 ;
        RECT 1212.660 1055.370 1212.920 1055.690 ;
        RECT 1211.800 1007.605 1211.940 1055.370 ;
        RECT 1211.730 1007.235 1212.010 1007.605 ;
        RECT 1212.650 1007.235 1212.930 1007.605 ;
        RECT 1212.720 959.130 1212.860 1007.235 ;
        RECT 1211.740 958.810 1212.000 959.130 ;
        RECT 1212.660 958.810 1212.920 959.130 ;
        RECT 1211.800 911.045 1211.940 958.810 ;
        RECT 1211.730 910.675 1212.010 911.045 ;
        RECT 1212.650 910.675 1212.930 911.045 ;
        RECT 1212.720 862.570 1212.860 910.675 ;
        RECT 1212.660 862.250 1212.920 862.570 ;
        RECT 1212.660 814.310 1212.920 814.630 ;
        RECT 1212.720 766.010 1212.860 814.310 ;
        RECT 1212.660 765.690 1212.920 766.010 ;
        RECT 1212.660 717.750 1212.920 718.070 ;
        RECT 1212.720 669.450 1212.860 717.750 ;
        RECT 1212.660 669.130 1212.920 669.450 ;
        RECT 1212.660 620.850 1212.920 621.170 ;
        RECT 1212.720 572.550 1212.860 620.850 ;
        RECT 1212.660 572.230 1212.920 572.550 ;
        RECT 1212.660 524.290 1212.920 524.610 ;
        RECT 1212.720 475.990 1212.860 524.290 ;
        RECT 1212.660 475.670 1212.920 475.990 ;
        RECT 1212.660 427.730 1212.920 428.050 ;
        RECT 1212.720 379.430 1212.860 427.730 ;
        RECT 1212.660 379.110 1212.920 379.430 ;
        RECT 1212.660 331.170 1212.920 331.490 ;
        RECT 1212.720 282.870 1212.860 331.170 ;
        RECT 1212.660 282.550 1212.920 282.870 ;
        RECT 1212.660 234.610 1212.920 234.930 ;
        RECT 1212.720 186.310 1212.860 234.610 ;
        RECT 1212.660 185.990 1212.920 186.310 ;
        RECT 1212.660 138.050 1212.920 138.370 ;
        RECT 1212.720 113.970 1212.860 138.050 ;
        RECT 1211.800 113.830 1212.860 113.970 ;
        RECT 1211.800 96.290 1211.940 113.830 ;
        RECT 1211.800 96.150 1212.400 96.290 ;
        RECT 1212.260 64.250 1212.400 96.150 ;
        RECT 1212.200 63.930 1212.460 64.250 ;
        RECT 2477.200 63.930 2477.460 64.250 ;
        RECT 2477.260 3.050 2477.400 63.930 ;
        RECT 2477.200 2.730 2477.460 3.050 ;
        RECT 2482.720 2.730 2482.980 3.050 ;
        RECT 2482.780 2.400 2482.920 2.730 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
      LAYER via2 ;
        RECT 1211.730 1248.680 1212.010 1248.960 ;
        RECT 1212.650 1248.680 1212.930 1248.960 ;
        RECT 1211.730 1152.120 1212.010 1152.400 ;
        RECT 1212.650 1152.120 1212.930 1152.400 ;
        RECT 1211.730 1007.280 1212.010 1007.560 ;
        RECT 1212.650 1007.280 1212.930 1007.560 ;
        RECT 1211.730 910.720 1212.010 911.000 ;
        RECT 1212.650 910.720 1212.930 911.000 ;
      LAYER met3 ;
        RECT 1211.705 1248.970 1212.035 1248.985 ;
        RECT 1212.625 1248.970 1212.955 1248.985 ;
        RECT 1211.705 1248.670 1212.955 1248.970 ;
        RECT 1211.705 1248.655 1212.035 1248.670 ;
        RECT 1212.625 1248.655 1212.955 1248.670 ;
        RECT 1211.705 1152.410 1212.035 1152.425 ;
        RECT 1212.625 1152.410 1212.955 1152.425 ;
        RECT 1211.705 1152.110 1212.955 1152.410 ;
        RECT 1211.705 1152.095 1212.035 1152.110 ;
        RECT 1212.625 1152.095 1212.955 1152.110 ;
        RECT 1211.705 1007.570 1212.035 1007.585 ;
        RECT 1212.625 1007.570 1212.955 1007.585 ;
        RECT 1211.705 1007.270 1212.955 1007.570 ;
        RECT 1211.705 1007.255 1212.035 1007.270 ;
        RECT 1212.625 1007.255 1212.955 1007.270 ;
        RECT 1211.705 911.010 1212.035 911.025 ;
        RECT 1212.625 911.010 1212.955 911.025 ;
        RECT 1211.705 910.710 1212.955 911.010 ;
        RECT 1211.705 910.695 1212.035 910.710 ;
        RECT 1212.625 910.695 1212.955 910.710 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1219.605 1442.025 1219.775 1490.475 ;
        RECT 1219.145 1386.945 1219.315 1394.255 ;
        RECT 1219.145 758.965 1219.315 807.075 ;
        RECT 1219.145 620.925 1219.315 669.035 ;
        RECT 1219.145 565.845 1219.315 613.955 ;
      LAYER mcon ;
        RECT 1219.605 1490.305 1219.775 1490.475 ;
        RECT 1219.145 1394.085 1219.315 1394.255 ;
        RECT 1219.145 806.905 1219.315 807.075 ;
        RECT 1219.145 668.865 1219.315 669.035 ;
        RECT 1219.145 613.785 1219.315 613.955 ;
      LAYER met1 ;
        RECT 1214.470 1579.880 1214.790 1579.940 ;
        RECT 1215.390 1579.880 1215.710 1579.940 ;
        RECT 1214.470 1579.740 1215.710 1579.880 ;
        RECT 1214.470 1579.680 1214.790 1579.740 ;
        RECT 1215.390 1579.680 1215.710 1579.740 ;
        RECT 1214.470 1534.320 1214.790 1534.380 ;
        RECT 1219.530 1534.320 1219.850 1534.380 ;
        RECT 1214.470 1534.180 1219.850 1534.320 ;
        RECT 1214.470 1534.120 1214.790 1534.180 ;
        RECT 1219.530 1534.120 1219.850 1534.180 ;
        RECT 1219.530 1490.460 1219.850 1490.520 ;
        RECT 1219.335 1490.320 1219.850 1490.460 ;
        RECT 1219.530 1490.260 1219.850 1490.320 ;
        RECT 1219.070 1442.180 1219.390 1442.240 ;
        RECT 1219.545 1442.180 1219.835 1442.225 ;
        RECT 1219.070 1442.040 1219.835 1442.180 ;
        RECT 1219.070 1441.980 1219.390 1442.040 ;
        RECT 1219.545 1441.995 1219.835 1442.040 ;
        RECT 1219.070 1394.240 1219.390 1394.300 ;
        RECT 1218.875 1394.100 1219.390 1394.240 ;
        RECT 1219.070 1394.040 1219.390 1394.100 ;
        RECT 1219.070 1387.100 1219.390 1387.160 ;
        RECT 1218.875 1386.960 1219.390 1387.100 ;
        RECT 1219.070 1386.900 1219.390 1386.960 ;
        RECT 1219.070 1345.960 1219.390 1346.020 ;
        RECT 1218.700 1345.820 1219.390 1345.960 ;
        RECT 1218.700 1345.340 1218.840 1345.820 ;
        RECT 1219.070 1345.760 1219.390 1345.820 ;
        RECT 1218.610 1345.080 1218.930 1345.340 ;
        RECT 1218.150 1249.060 1218.470 1249.120 ;
        RECT 1219.070 1249.060 1219.390 1249.120 ;
        RECT 1218.150 1248.920 1219.390 1249.060 ;
        RECT 1218.150 1248.860 1218.470 1248.920 ;
        RECT 1219.070 1248.860 1219.390 1248.920 ;
        RECT 1218.150 1152.500 1218.470 1152.560 ;
        RECT 1219.070 1152.500 1219.390 1152.560 ;
        RECT 1218.150 1152.360 1219.390 1152.500 ;
        RECT 1218.150 1152.300 1218.470 1152.360 ;
        RECT 1219.070 1152.300 1219.390 1152.360 ;
        RECT 1218.610 1055.940 1218.930 1056.000 ;
        RECT 1219.070 1055.940 1219.390 1056.000 ;
        RECT 1218.610 1055.800 1219.390 1055.940 ;
        RECT 1218.610 1055.740 1218.930 1055.800 ;
        RECT 1219.070 1055.740 1219.390 1055.800 ;
        RECT 1218.610 959.380 1218.930 959.440 ;
        RECT 1219.070 959.380 1219.390 959.440 ;
        RECT 1218.610 959.240 1219.390 959.380 ;
        RECT 1218.610 959.180 1218.930 959.240 ;
        RECT 1219.070 959.180 1219.390 959.240 ;
        RECT 1218.610 862.820 1218.930 862.880 ;
        RECT 1219.070 862.820 1219.390 862.880 ;
        RECT 1218.610 862.680 1219.390 862.820 ;
        RECT 1218.610 862.620 1218.930 862.680 ;
        RECT 1219.070 862.620 1219.390 862.680 ;
        RECT 1219.070 862.140 1219.390 862.200 ;
        RECT 1219.530 862.140 1219.850 862.200 ;
        RECT 1219.070 862.000 1219.850 862.140 ;
        RECT 1219.070 861.940 1219.390 862.000 ;
        RECT 1219.530 861.940 1219.850 862.000 ;
        RECT 1219.070 807.060 1219.390 807.120 ;
        RECT 1218.875 806.920 1219.390 807.060 ;
        RECT 1219.070 806.860 1219.390 806.920 ;
        RECT 1219.070 759.120 1219.390 759.180 ;
        RECT 1218.875 758.980 1219.390 759.120 ;
        RECT 1219.070 758.920 1219.390 758.980 ;
        RECT 1218.150 717.980 1218.470 718.040 ;
        RECT 1219.070 717.980 1219.390 718.040 ;
        RECT 1218.150 717.840 1219.390 717.980 ;
        RECT 1218.150 717.780 1218.470 717.840 ;
        RECT 1219.070 717.780 1219.390 717.840 ;
        RECT 1218.150 669.700 1218.470 669.760 ;
        RECT 1219.070 669.700 1219.390 669.760 ;
        RECT 1218.150 669.560 1219.390 669.700 ;
        RECT 1218.150 669.500 1218.470 669.560 ;
        RECT 1219.070 669.500 1219.390 669.560 ;
        RECT 1219.070 669.020 1219.390 669.080 ;
        RECT 1218.875 668.880 1219.390 669.020 ;
        RECT 1219.070 668.820 1219.390 668.880 ;
        RECT 1219.070 621.080 1219.390 621.140 ;
        RECT 1218.875 620.940 1219.390 621.080 ;
        RECT 1219.070 620.880 1219.390 620.940 ;
        RECT 1219.070 613.940 1219.390 614.000 ;
        RECT 1218.875 613.800 1219.390 613.940 ;
        RECT 1219.070 613.740 1219.390 613.800 ;
        RECT 1219.070 566.000 1219.390 566.060 ;
        RECT 1218.875 565.860 1219.390 566.000 ;
        RECT 1219.070 565.800 1219.390 565.860 ;
        RECT 1219.070 524.860 1219.390 524.920 ;
        RECT 1218.240 524.720 1219.390 524.860 ;
        RECT 1218.240 524.580 1218.380 524.720 ;
        RECT 1219.070 524.660 1219.390 524.720 ;
        RECT 1218.150 524.320 1218.470 524.580 ;
        RECT 1218.150 476.240 1218.470 476.300 ;
        RECT 1219.070 476.240 1219.390 476.300 ;
        RECT 1218.150 476.100 1219.390 476.240 ;
        RECT 1218.150 476.040 1218.470 476.100 ;
        RECT 1219.070 476.040 1219.390 476.100 ;
        RECT 1218.150 379.680 1218.470 379.740 ;
        RECT 1219.070 379.680 1219.390 379.740 ;
        RECT 1218.150 379.540 1219.390 379.680 ;
        RECT 1218.150 379.480 1218.470 379.540 ;
        RECT 1219.070 379.480 1219.390 379.540 ;
        RECT 1218.150 283.120 1218.470 283.180 ;
        RECT 1219.070 283.120 1219.390 283.180 ;
        RECT 1218.150 282.980 1219.390 283.120 ;
        RECT 1218.150 282.920 1218.470 282.980 ;
        RECT 1219.070 282.920 1219.390 282.980 ;
        RECT 1218.150 186.560 1218.470 186.620 ;
        RECT 1219.070 186.560 1219.390 186.620 ;
        RECT 1218.150 186.420 1219.390 186.560 ;
        RECT 1218.150 186.360 1218.470 186.420 ;
        RECT 1219.070 186.360 1219.390 186.420 ;
        RECT 1218.610 90.000 1218.930 90.060 ;
        RECT 1219.070 90.000 1219.390 90.060 ;
        RECT 1218.610 89.860 1219.390 90.000 ;
        RECT 1218.610 89.800 1218.930 89.860 ;
        RECT 1219.070 89.800 1219.390 89.860 ;
        RECT 1219.070 64.500 1219.390 64.560 ;
        RECT 2497.870 64.500 2498.190 64.560 ;
        RECT 1219.070 64.360 2498.190 64.500 ;
        RECT 1219.070 64.300 1219.390 64.360 ;
        RECT 2497.870 64.300 2498.190 64.360 ;
        RECT 2497.870 2.960 2498.190 3.020 ;
        RECT 2500.630 2.960 2500.950 3.020 ;
        RECT 2497.870 2.820 2500.950 2.960 ;
        RECT 2497.870 2.760 2498.190 2.820 ;
        RECT 2500.630 2.760 2500.950 2.820 ;
      LAYER via ;
        RECT 1214.500 1579.680 1214.760 1579.940 ;
        RECT 1215.420 1579.680 1215.680 1579.940 ;
        RECT 1214.500 1534.120 1214.760 1534.380 ;
        RECT 1219.560 1534.120 1219.820 1534.380 ;
        RECT 1219.560 1490.260 1219.820 1490.520 ;
        RECT 1219.100 1441.980 1219.360 1442.240 ;
        RECT 1219.100 1394.040 1219.360 1394.300 ;
        RECT 1219.100 1386.900 1219.360 1387.160 ;
        RECT 1219.100 1345.760 1219.360 1346.020 ;
        RECT 1218.640 1345.080 1218.900 1345.340 ;
        RECT 1218.180 1248.860 1218.440 1249.120 ;
        RECT 1219.100 1248.860 1219.360 1249.120 ;
        RECT 1218.180 1152.300 1218.440 1152.560 ;
        RECT 1219.100 1152.300 1219.360 1152.560 ;
        RECT 1218.640 1055.740 1218.900 1056.000 ;
        RECT 1219.100 1055.740 1219.360 1056.000 ;
        RECT 1218.640 959.180 1218.900 959.440 ;
        RECT 1219.100 959.180 1219.360 959.440 ;
        RECT 1218.640 862.620 1218.900 862.880 ;
        RECT 1219.100 862.620 1219.360 862.880 ;
        RECT 1219.100 861.940 1219.360 862.200 ;
        RECT 1219.560 861.940 1219.820 862.200 ;
        RECT 1219.100 806.860 1219.360 807.120 ;
        RECT 1219.100 758.920 1219.360 759.180 ;
        RECT 1218.180 717.780 1218.440 718.040 ;
        RECT 1219.100 717.780 1219.360 718.040 ;
        RECT 1218.180 669.500 1218.440 669.760 ;
        RECT 1219.100 669.500 1219.360 669.760 ;
        RECT 1219.100 668.820 1219.360 669.080 ;
        RECT 1219.100 620.880 1219.360 621.140 ;
        RECT 1219.100 613.740 1219.360 614.000 ;
        RECT 1219.100 565.800 1219.360 566.060 ;
        RECT 1219.100 524.660 1219.360 524.920 ;
        RECT 1218.180 524.320 1218.440 524.580 ;
        RECT 1218.180 476.040 1218.440 476.300 ;
        RECT 1219.100 476.040 1219.360 476.300 ;
        RECT 1218.180 379.480 1218.440 379.740 ;
        RECT 1219.100 379.480 1219.360 379.740 ;
        RECT 1218.180 282.920 1218.440 283.180 ;
        RECT 1219.100 282.920 1219.360 283.180 ;
        RECT 1218.180 186.360 1218.440 186.620 ;
        RECT 1219.100 186.360 1219.360 186.620 ;
        RECT 1218.640 89.800 1218.900 90.060 ;
        RECT 1219.100 89.800 1219.360 90.060 ;
        RECT 1219.100 64.300 1219.360 64.560 ;
        RECT 2497.900 64.300 2498.160 64.560 ;
        RECT 2497.900 2.760 2498.160 3.020 ;
        RECT 2500.660 2.760 2500.920 3.020 ;
      LAYER met2 ;
        RECT 1216.660 1600.450 1216.940 1604.000 ;
        RECT 1215.480 1600.310 1216.940 1600.450 ;
        RECT 1215.480 1579.970 1215.620 1600.310 ;
        RECT 1216.660 1600.000 1216.940 1600.310 ;
        RECT 1214.500 1579.650 1214.760 1579.970 ;
        RECT 1215.420 1579.650 1215.680 1579.970 ;
        RECT 1214.560 1534.410 1214.700 1579.650 ;
        RECT 1214.500 1534.090 1214.760 1534.410 ;
        RECT 1219.560 1534.090 1219.820 1534.410 ;
        RECT 1219.620 1490.550 1219.760 1534.090 ;
        RECT 1219.560 1490.230 1219.820 1490.550 ;
        RECT 1219.100 1441.950 1219.360 1442.270 ;
        RECT 1219.160 1394.330 1219.300 1441.950 ;
        RECT 1219.100 1394.010 1219.360 1394.330 ;
        RECT 1219.100 1386.870 1219.360 1387.190 ;
        RECT 1219.160 1346.050 1219.300 1386.870 ;
        RECT 1219.100 1345.730 1219.360 1346.050 ;
        RECT 1218.640 1345.050 1218.900 1345.370 ;
        RECT 1218.700 1322.330 1218.840 1345.050 ;
        RECT 1218.240 1322.190 1218.840 1322.330 ;
        RECT 1218.240 1249.150 1218.380 1322.190 ;
        RECT 1218.180 1248.830 1218.440 1249.150 ;
        RECT 1219.100 1248.830 1219.360 1249.150 ;
        RECT 1219.160 1225.090 1219.300 1248.830 ;
        RECT 1218.240 1224.950 1219.300 1225.090 ;
        RECT 1218.240 1152.590 1218.380 1224.950 ;
        RECT 1218.180 1152.270 1218.440 1152.590 ;
        RECT 1219.100 1152.270 1219.360 1152.590 ;
        RECT 1219.160 1104.050 1219.300 1152.270 ;
        RECT 1218.700 1103.910 1219.300 1104.050 ;
        RECT 1218.700 1056.030 1218.840 1103.910 ;
        RECT 1218.640 1055.710 1218.900 1056.030 ;
        RECT 1219.100 1055.710 1219.360 1056.030 ;
        RECT 1219.160 1031.290 1219.300 1055.710 ;
        RECT 1218.700 1031.150 1219.300 1031.290 ;
        RECT 1218.700 959.470 1218.840 1031.150 ;
        RECT 1218.640 959.150 1218.900 959.470 ;
        RECT 1219.100 959.150 1219.360 959.470 ;
        RECT 1219.160 910.930 1219.300 959.150 ;
        RECT 1218.700 910.790 1219.300 910.930 ;
        RECT 1218.700 862.910 1218.840 910.790 ;
        RECT 1218.640 862.590 1218.900 862.910 ;
        RECT 1219.100 862.590 1219.360 862.910 ;
        RECT 1219.160 862.230 1219.300 862.590 ;
        RECT 1219.100 861.910 1219.360 862.230 ;
        RECT 1219.560 861.910 1219.820 862.230 ;
        RECT 1219.620 814.370 1219.760 861.910 ;
        RECT 1219.160 814.230 1219.760 814.370 ;
        RECT 1219.160 807.150 1219.300 814.230 ;
        RECT 1219.100 806.830 1219.360 807.150 ;
        RECT 1219.100 758.890 1219.360 759.210 ;
        RECT 1219.160 718.070 1219.300 758.890 ;
        RECT 1218.180 717.750 1218.440 718.070 ;
        RECT 1219.100 717.750 1219.360 718.070 ;
        RECT 1218.240 669.790 1218.380 717.750 ;
        RECT 1218.180 669.470 1218.440 669.790 ;
        RECT 1219.100 669.470 1219.360 669.790 ;
        RECT 1219.160 669.110 1219.300 669.470 ;
        RECT 1219.100 668.790 1219.360 669.110 ;
        RECT 1219.100 620.850 1219.360 621.170 ;
        RECT 1219.160 614.030 1219.300 620.850 ;
        RECT 1219.100 613.710 1219.360 614.030 ;
        RECT 1219.100 565.770 1219.360 566.090 ;
        RECT 1219.160 524.950 1219.300 565.770 ;
        RECT 1219.100 524.630 1219.360 524.950 ;
        RECT 1218.180 524.290 1218.440 524.610 ;
        RECT 1218.240 476.330 1218.380 524.290 ;
        RECT 1218.180 476.010 1218.440 476.330 ;
        RECT 1219.100 476.010 1219.360 476.330 ;
        RECT 1219.160 451.250 1219.300 476.010 ;
        RECT 1218.240 451.110 1219.300 451.250 ;
        RECT 1218.240 379.770 1218.380 451.110 ;
        RECT 1218.180 379.450 1218.440 379.770 ;
        RECT 1219.100 379.450 1219.360 379.770 ;
        RECT 1219.160 355.370 1219.300 379.450 ;
        RECT 1218.240 355.230 1219.300 355.370 ;
        RECT 1218.240 283.210 1218.380 355.230 ;
        RECT 1218.180 282.890 1218.440 283.210 ;
        RECT 1219.100 282.890 1219.360 283.210 ;
        RECT 1219.160 234.445 1219.300 282.890 ;
        RECT 1218.170 234.075 1218.450 234.445 ;
        RECT 1219.090 234.075 1219.370 234.445 ;
        RECT 1218.240 186.650 1218.380 234.075 ;
        RECT 1218.180 186.330 1218.440 186.650 ;
        RECT 1219.100 186.330 1219.360 186.650 ;
        RECT 1219.160 137.770 1219.300 186.330 ;
        RECT 1218.700 137.630 1219.300 137.770 ;
        RECT 1218.700 90.090 1218.840 137.630 ;
        RECT 1218.640 89.770 1218.900 90.090 ;
        RECT 1219.100 89.770 1219.360 90.090 ;
        RECT 1219.160 64.590 1219.300 89.770 ;
        RECT 1219.100 64.270 1219.360 64.590 ;
        RECT 2497.900 64.270 2498.160 64.590 ;
        RECT 2497.960 3.050 2498.100 64.270 ;
        RECT 2497.900 2.730 2498.160 3.050 ;
        RECT 2500.660 2.730 2500.920 3.050 ;
        RECT 2500.720 2.400 2500.860 2.730 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
      LAYER via2 ;
        RECT 1218.170 234.120 1218.450 234.400 ;
        RECT 1219.090 234.120 1219.370 234.400 ;
      LAYER met3 ;
        RECT 1218.145 234.410 1218.475 234.425 ;
        RECT 1219.065 234.410 1219.395 234.425 ;
        RECT 1218.145 234.110 1219.395 234.410 ;
        RECT 1218.145 234.095 1218.475 234.110 ;
        RECT 1219.065 234.095 1219.395 234.110 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1221.830 1481.620 1222.150 1481.680 ;
        RECT 1226.890 1481.620 1227.210 1481.680 ;
        RECT 1221.830 1481.480 1227.210 1481.620 ;
        RECT 1221.830 1481.420 1222.150 1481.480 ;
        RECT 1226.890 1481.420 1227.210 1481.480 ;
        RECT 1226.890 64.840 1227.210 64.900 ;
        RECT 2511.670 64.840 2511.990 64.900 ;
        RECT 1226.890 64.700 2511.990 64.840 ;
        RECT 1226.890 64.640 1227.210 64.700 ;
        RECT 2511.670 64.640 2511.990 64.700 ;
        RECT 2511.670 17.580 2511.990 17.640 ;
        RECT 2518.110 17.580 2518.430 17.640 ;
        RECT 2511.670 17.440 2518.430 17.580 ;
        RECT 2511.670 17.380 2511.990 17.440 ;
        RECT 2518.110 17.380 2518.430 17.440 ;
      LAYER via ;
        RECT 1221.860 1481.420 1222.120 1481.680 ;
        RECT 1226.920 1481.420 1227.180 1481.680 ;
        RECT 1226.920 64.640 1227.180 64.900 ;
        RECT 2511.700 64.640 2511.960 64.900 ;
        RECT 2511.700 17.380 2511.960 17.640 ;
        RECT 2518.140 17.380 2518.400 17.640 ;
      LAYER met2 ;
        RECT 1222.640 1601.130 1222.920 1604.000 ;
        RECT 1221.920 1600.990 1222.920 1601.130 ;
        RECT 1221.920 1481.710 1222.060 1600.990 ;
        RECT 1222.640 1600.000 1222.920 1600.990 ;
        RECT 1221.860 1481.390 1222.120 1481.710 ;
        RECT 1226.920 1481.390 1227.180 1481.710 ;
        RECT 1226.980 64.930 1227.120 1481.390 ;
        RECT 1226.920 64.610 1227.180 64.930 ;
        RECT 2511.700 64.610 2511.960 64.930 ;
        RECT 2511.760 17.670 2511.900 64.610 ;
        RECT 2511.700 17.350 2511.960 17.670 ;
        RECT 2518.140 17.350 2518.400 17.670 ;
        RECT 2518.200 2.400 2518.340 17.350 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1228.730 1594.160 1229.050 1594.220 ;
        RECT 1229.190 1594.160 1229.510 1594.220 ;
        RECT 1228.730 1594.020 1229.510 1594.160 ;
        RECT 1228.730 1593.960 1229.050 1594.020 ;
        RECT 1229.190 1593.960 1229.510 1594.020 ;
        RECT 1228.730 1473.120 1229.050 1473.180 ;
        RECT 1233.790 1473.120 1234.110 1473.180 ;
        RECT 1228.730 1472.980 1234.110 1473.120 ;
        RECT 1228.730 1472.920 1229.050 1472.980 ;
        RECT 1233.790 1472.920 1234.110 1472.980 ;
        RECT 1233.790 65.180 1234.110 65.240 ;
        RECT 2532.370 65.180 2532.690 65.240 ;
        RECT 1233.790 65.040 2532.690 65.180 ;
        RECT 1233.790 64.980 1234.110 65.040 ;
        RECT 2532.370 64.980 2532.690 65.040 ;
        RECT 2532.370 2.960 2532.690 3.020 ;
        RECT 2536.050 2.960 2536.370 3.020 ;
        RECT 2532.370 2.820 2536.370 2.960 ;
        RECT 2532.370 2.760 2532.690 2.820 ;
        RECT 2536.050 2.760 2536.370 2.820 ;
      LAYER via ;
        RECT 1228.760 1593.960 1229.020 1594.220 ;
        RECT 1229.220 1593.960 1229.480 1594.220 ;
        RECT 1228.760 1472.920 1229.020 1473.180 ;
        RECT 1233.820 1472.920 1234.080 1473.180 ;
        RECT 1233.820 64.980 1234.080 65.240 ;
        RECT 2532.400 64.980 2532.660 65.240 ;
        RECT 2532.400 2.760 2532.660 3.020 ;
        RECT 2536.080 2.760 2536.340 3.020 ;
      LAYER met2 ;
        RECT 1229.080 1600.380 1229.360 1604.000 ;
        RECT 1229.080 1600.000 1229.420 1600.380 ;
        RECT 1229.280 1594.250 1229.420 1600.000 ;
        RECT 1228.760 1593.930 1229.020 1594.250 ;
        RECT 1229.220 1593.930 1229.480 1594.250 ;
        RECT 1228.820 1473.210 1228.960 1593.930 ;
        RECT 1228.760 1472.890 1229.020 1473.210 ;
        RECT 1233.820 1472.890 1234.080 1473.210 ;
        RECT 1233.880 65.270 1234.020 1472.890 ;
        RECT 1233.820 64.950 1234.080 65.270 ;
        RECT 2532.400 64.950 2532.660 65.270 ;
        RECT 2532.460 3.050 2532.600 64.950 ;
        RECT 2532.400 2.730 2532.660 3.050 ;
        RECT 2536.080 2.730 2536.340 3.050 ;
        RECT 2536.140 2.400 2536.280 2.730 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1235.170 1536.700 1235.490 1536.760 ;
        RECT 1240.690 1536.700 1241.010 1536.760 ;
        RECT 1235.170 1536.560 1241.010 1536.700 ;
        RECT 1235.170 1536.500 1235.490 1536.560 ;
        RECT 1240.690 1536.500 1241.010 1536.560 ;
        RECT 1240.690 68.920 1241.010 68.980 ;
        RECT 2553.070 68.920 2553.390 68.980 ;
        RECT 1240.690 68.780 2553.390 68.920 ;
        RECT 1240.690 68.720 1241.010 68.780 ;
        RECT 2553.070 68.720 2553.390 68.780 ;
        RECT 2553.070 2.960 2553.390 3.020 ;
        RECT 2553.990 2.960 2554.310 3.020 ;
        RECT 2553.070 2.820 2554.310 2.960 ;
        RECT 2553.070 2.760 2553.390 2.820 ;
        RECT 2553.990 2.760 2554.310 2.820 ;
      LAYER via ;
        RECT 1235.200 1536.500 1235.460 1536.760 ;
        RECT 1240.720 1536.500 1240.980 1536.760 ;
        RECT 1240.720 68.720 1240.980 68.980 ;
        RECT 2553.100 68.720 2553.360 68.980 ;
        RECT 2553.100 2.760 2553.360 3.020 ;
        RECT 2554.020 2.760 2554.280 3.020 ;
      LAYER met2 ;
        RECT 1235.060 1600.380 1235.340 1604.000 ;
        RECT 1235.060 1600.000 1235.400 1600.380 ;
        RECT 1235.260 1536.790 1235.400 1600.000 ;
        RECT 1235.200 1536.470 1235.460 1536.790 ;
        RECT 1240.720 1536.470 1240.980 1536.790 ;
        RECT 1240.780 69.010 1240.920 1536.470 ;
        RECT 1240.720 68.690 1240.980 69.010 ;
        RECT 2553.100 68.690 2553.360 69.010 ;
        RECT 2553.160 3.050 2553.300 68.690 ;
        RECT 2553.100 2.730 2553.360 3.050 ;
        RECT 2554.020 2.730 2554.280 3.050 ;
        RECT 2554.080 2.400 2554.220 2.730 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1235.630 1600.960 1235.950 1601.020 ;
        RECT 1240.230 1600.960 1240.550 1601.020 ;
        RECT 1235.630 1600.820 1240.550 1600.960 ;
        RECT 1235.630 1600.760 1235.950 1600.820 ;
        RECT 1240.230 1600.760 1240.550 1600.820 ;
        RECT 1236.090 1473.120 1236.410 1473.180 ;
        RECT 1240.230 1473.120 1240.550 1473.180 ;
        RECT 1236.090 1472.980 1240.550 1473.120 ;
        RECT 1236.090 1472.920 1236.410 1472.980 ;
        RECT 1240.230 1472.920 1240.550 1472.980 ;
        RECT 1240.230 68.580 1240.550 68.640 ;
        RECT 2566.870 68.580 2567.190 68.640 ;
        RECT 1240.230 68.440 2567.190 68.580 ;
        RECT 1240.230 68.380 1240.550 68.440 ;
        RECT 2566.870 68.380 2567.190 68.440 ;
        RECT 2566.870 2.960 2567.190 3.020 ;
        RECT 2571.930 2.960 2572.250 3.020 ;
        RECT 2566.870 2.820 2572.250 2.960 ;
        RECT 2566.870 2.760 2567.190 2.820 ;
        RECT 2571.930 2.760 2572.250 2.820 ;
      LAYER via ;
        RECT 1235.660 1600.760 1235.920 1601.020 ;
        RECT 1240.260 1600.760 1240.520 1601.020 ;
        RECT 1236.120 1472.920 1236.380 1473.180 ;
        RECT 1240.260 1472.920 1240.520 1473.180 ;
        RECT 1240.260 68.380 1240.520 68.640 ;
        RECT 2566.900 68.380 2567.160 68.640 ;
        RECT 2566.900 2.760 2567.160 3.020 ;
        RECT 2571.960 2.760 2572.220 3.020 ;
      LAYER met2 ;
        RECT 1241.500 1601.130 1241.780 1604.000 ;
        RECT 1240.320 1601.050 1241.780 1601.130 ;
        RECT 1235.660 1600.730 1235.920 1601.050 ;
        RECT 1240.260 1600.990 1241.780 1601.050 ;
        RECT 1240.260 1600.730 1240.520 1600.990 ;
        RECT 1235.720 1535.170 1235.860 1600.730 ;
        RECT 1241.500 1600.000 1241.780 1600.990 ;
        RECT 1235.720 1535.030 1236.320 1535.170 ;
        RECT 1236.180 1473.210 1236.320 1535.030 ;
        RECT 1236.120 1472.890 1236.380 1473.210 ;
        RECT 1240.260 1472.890 1240.520 1473.210 ;
        RECT 1240.320 68.670 1240.460 1472.890 ;
        RECT 1240.260 68.350 1240.520 68.670 ;
        RECT 2566.900 68.350 2567.160 68.670 ;
        RECT 2566.960 3.050 2567.100 68.350 ;
        RECT 2566.900 2.730 2567.160 3.050 ;
        RECT 2571.960 2.730 2572.220 3.050 ;
        RECT 2572.020 2.400 2572.160 2.730 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1242.530 1558.120 1242.850 1558.180 ;
        RECT 1247.130 1558.120 1247.450 1558.180 ;
        RECT 1242.530 1557.980 1247.450 1558.120 ;
        RECT 1242.530 1557.920 1242.850 1557.980 ;
        RECT 1247.130 1557.920 1247.450 1557.980 ;
        RECT 1242.530 1473.120 1242.850 1473.180 ;
        RECT 1247.590 1473.120 1247.910 1473.180 ;
        RECT 1242.530 1472.980 1247.910 1473.120 ;
        RECT 1242.530 1472.920 1242.850 1472.980 ;
        RECT 1247.590 1472.920 1247.910 1472.980 ;
        RECT 1247.590 68.240 1247.910 68.300 ;
        RECT 2587.570 68.240 2587.890 68.300 ;
        RECT 1247.590 68.100 2587.890 68.240 ;
        RECT 1247.590 68.040 1247.910 68.100 ;
        RECT 2587.570 68.040 2587.890 68.100 ;
      LAYER via ;
        RECT 1242.560 1557.920 1242.820 1558.180 ;
        RECT 1247.160 1557.920 1247.420 1558.180 ;
        RECT 1242.560 1472.920 1242.820 1473.180 ;
        RECT 1247.620 1472.920 1247.880 1473.180 ;
        RECT 1247.620 68.040 1247.880 68.300 ;
        RECT 2587.600 68.040 2587.860 68.300 ;
      LAYER met2 ;
        RECT 1247.480 1600.380 1247.760 1604.000 ;
        RECT 1247.480 1600.000 1247.820 1600.380 ;
        RECT 1247.680 1597.220 1247.820 1600.000 ;
        RECT 1247.220 1597.080 1247.820 1597.220 ;
        RECT 1247.220 1558.210 1247.360 1597.080 ;
        RECT 1242.560 1557.890 1242.820 1558.210 ;
        RECT 1247.160 1557.890 1247.420 1558.210 ;
        RECT 1242.620 1473.210 1242.760 1557.890 ;
        RECT 1242.560 1472.890 1242.820 1473.210 ;
        RECT 1247.620 1472.890 1247.880 1473.210 ;
        RECT 1247.680 68.330 1247.820 1472.890 ;
        RECT 1247.620 68.010 1247.880 68.330 ;
        RECT 2587.600 68.010 2587.860 68.330 ;
        RECT 2587.660 3.130 2587.800 68.010 ;
        RECT 2587.660 2.990 2589.640 3.130 ;
        RECT 2589.500 2.400 2589.640 2.990 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 662.545 20.145 662.715 21.335 ;
        RECT 768.345 20.485 769.895 20.655 ;
        RECT 786.745 20.145 786.915 20.995 ;
      LAYER mcon ;
        RECT 662.545 21.165 662.715 21.335 ;
        RECT 786.745 20.825 786.915 20.995 ;
        RECT 769.725 20.485 769.895 20.655 ;
      LAYER met1 ;
        RECT 635.330 1588.720 635.650 1588.780 ;
        RECT 640.850 1588.720 641.170 1588.780 ;
        RECT 635.330 1588.580 641.170 1588.720 ;
        RECT 635.330 1588.520 635.650 1588.580 ;
        RECT 640.850 1588.520 641.170 1588.580 ;
        RECT 662.485 21.320 662.775 21.365 ;
        RECT 662.485 21.180 681.560 21.320 ;
        RECT 662.485 21.135 662.775 21.180 ;
        RECT 681.420 20.980 681.560 21.180 ;
        RECT 786.685 20.980 786.975 21.025 ;
        RECT 681.420 20.840 728.480 20.980 ;
        RECT 728.340 20.640 728.480 20.840 ;
        RECT 785.840 20.840 786.975 20.980 ;
        RECT 768.285 20.640 768.575 20.685 ;
        RECT 728.340 20.500 768.575 20.640 ;
        RECT 768.285 20.455 768.575 20.500 ;
        RECT 769.665 20.640 769.955 20.685 ;
        RECT 785.840 20.640 785.980 20.840 ;
        RECT 786.685 20.795 786.975 20.840 ;
        RECT 769.665 20.500 785.980 20.640 ;
        RECT 769.665 20.455 769.955 20.500 ;
        RECT 640.850 20.300 641.170 20.360 ;
        RECT 662.485 20.300 662.775 20.345 ;
        RECT 640.850 20.160 662.775 20.300 ;
        RECT 640.850 20.100 641.170 20.160 ;
        RECT 662.485 20.115 662.775 20.160 ;
        RECT 786.685 20.300 786.975 20.345 ;
        RECT 823.470 20.300 823.790 20.360 ;
        RECT 786.685 20.160 823.790 20.300 ;
        RECT 786.685 20.115 786.975 20.160 ;
        RECT 823.470 20.100 823.790 20.160 ;
      LAYER via ;
        RECT 635.360 1588.520 635.620 1588.780 ;
        RECT 640.880 1588.520 641.140 1588.780 ;
        RECT 640.880 20.100 641.140 20.360 ;
        RECT 823.500 20.100 823.760 20.360 ;
      LAYER met2 ;
        RECT 635.220 1600.380 635.500 1604.000 ;
        RECT 635.220 1600.000 635.560 1600.380 ;
        RECT 635.420 1588.810 635.560 1600.000 ;
        RECT 635.360 1588.490 635.620 1588.810 ;
        RECT 640.880 1588.490 641.140 1588.810 ;
        RECT 640.940 20.390 641.080 1588.490 ;
        RECT 640.880 20.070 641.140 20.390 ;
        RECT 823.500 20.070 823.760 20.390 ;
        RECT 823.560 2.400 823.700 20.070 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1249.430 1558.120 1249.750 1558.180 ;
        RECT 1253.110 1558.120 1253.430 1558.180 ;
        RECT 1249.430 1557.980 1253.430 1558.120 ;
        RECT 1249.430 1557.920 1249.750 1557.980 ;
        RECT 1253.110 1557.920 1253.430 1557.980 ;
        RECT 1249.430 1481.620 1249.750 1481.680 ;
        RECT 1254.490 1481.620 1254.810 1481.680 ;
        RECT 1249.430 1481.480 1254.810 1481.620 ;
        RECT 1249.430 1481.420 1249.750 1481.480 ;
        RECT 1254.490 1481.420 1254.810 1481.480 ;
        RECT 1254.490 67.900 1254.810 67.960 ;
        RECT 2601.370 67.900 2601.690 67.960 ;
        RECT 1254.490 67.760 2601.690 67.900 ;
        RECT 1254.490 67.700 1254.810 67.760 ;
        RECT 2601.370 67.700 2601.690 67.760 ;
        RECT 2601.370 17.580 2601.690 17.640 ;
        RECT 2607.350 17.580 2607.670 17.640 ;
        RECT 2601.370 17.440 2607.670 17.580 ;
        RECT 2601.370 17.380 2601.690 17.440 ;
        RECT 2607.350 17.380 2607.670 17.440 ;
      LAYER via ;
        RECT 1249.460 1557.920 1249.720 1558.180 ;
        RECT 1253.140 1557.920 1253.400 1558.180 ;
        RECT 1249.460 1481.420 1249.720 1481.680 ;
        RECT 1254.520 1481.420 1254.780 1481.680 ;
        RECT 1254.520 67.700 1254.780 67.960 ;
        RECT 2601.400 67.700 2601.660 67.960 ;
        RECT 2601.400 17.380 2601.660 17.640 ;
        RECT 2607.380 17.380 2607.640 17.640 ;
      LAYER met2 ;
        RECT 1253.460 1600.380 1253.740 1604.000 ;
        RECT 1253.460 1600.000 1253.800 1600.380 ;
        RECT 1253.660 1597.220 1253.800 1600.000 ;
        RECT 1253.200 1597.080 1253.800 1597.220 ;
        RECT 1253.200 1558.210 1253.340 1597.080 ;
        RECT 1249.460 1557.890 1249.720 1558.210 ;
        RECT 1253.140 1557.890 1253.400 1558.210 ;
        RECT 1249.520 1481.710 1249.660 1557.890 ;
        RECT 1249.460 1481.390 1249.720 1481.710 ;
        RECT 1254.520 1481.390 1254.780 1481.710 ;
        RECT 1254.580 67.990 1254.720 1481.390 ;
        RECT 1254.520 67.670 1254.780 67.990 ;
        RECT 2601.400 67.670 2601.660 67.990 ;
        RECT 2601.460 17.670 2601.600 67.670 ;
        RECT 2601.400 17.350 2601.660 17.670 ;
        RECT 2607.380 17.350 2607.640 17.670 ;
        RECT 2607.440 2.400 2607.580 17.350 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1256.405 1534.505 1256.575 1547.935 ;
        RECT 1256.405 1486.225 1256.575 1497.275 ;
      LAYER mcon ;
        RECT 1256.405 1547.765 1256.575 1547.935 ;
        RECT 1256.405 1497.105 1256.575 1497.275 ;
      LAYER met1 ;
        RECT 1256.345 1547.920 1256.635 1547.965 ;
        RECT 1258.630 1547.920 1258.950 1547.980 ;
        RECT 1256.345 1547.780 1258.950 1547.920 ;
        RECT 1256.345 1547.735 1256.635 1547.780 ;
        RECT 1258.630 1547.720 1258.950 1547.780 ;
        RECT 1256.330 1534.660 1256.650 1534.720 ;
        RECT 1256.135 1534.520 1256.650 1534.660 ;
        RECT 1256.330 1534.460 1256.650 1534.520 ;
        RECT 1256.330 1497.260 1256.650 1497.320 ;
        RECT 1256.135 1497.120 1256.650 1497.260 ;
        RECT 1256.330 1497.060 1256.650 1497.120 ;
        RECT 1256.345 1486.380 1256.635 1486.425 ;
        RECT 1260.930 1486.380 1261.250 1486.440 ;
        RECT 1256.345 1486.240 1261.250 1486.380 ;
        RECT 1256.345 1486.195 1256.635 1486.240 ;
        RECT 1260.930 1486.180 1261.250 1486.240 ;
        RECT 1260.930 67.560 1261.250 67.620 ;
        RECT 2622.070 67.560 2622.390 67.620 ;
        RECT 1260.930 67.420 2622.390 67.560 ;
        RECT 1260.930 67.360 1261.250 67.420 ;
        RECT 2622.070 67.360 2622.390 67.420 ;
        RECT 2622.070 2.960 2622.390 3.020 ;
        RECT 2625.290 2.960 2625.610 3.020 ;
        RECT 2622.070 2.820 2625.610 2.960 ;
        RECT 2622.070 2.760 2622.390 2.820 ;
        RECT 2625.290 2.760 2625.610 2.820 ;
      LAYER via ;
        RECT 1258.660 1547.720 1258.920 1547.980 ;
        RECT 1256.360 1534.460 1256.620 1534.720 ;
        RECT 1256.360 1497.060 1256.620 1497.320 ;
        RECT 1260.960 1486.180 1261.220 1486.440 ;
        RECT 1260.960 67.360 1261.220 67.620 ;
        RECT 2622.100 67.360 2622.360 67.620 ;
        RECT 2622.100 2.760 2622.360 3.020 ;
        RECT 2625.320 2.760 2625.580 3.020 ;
      LAYER met2 ;
        RECT 1259.900 1600.450 1260.180 1604.000 ;
        RECT 1258.720 1600.310 1260.180 1600.450 ;
        RECT 1258.720 1548.010 1258.860 1600.310 ;
        RECT 1259.900 1600.000 1260.180 1600.310 ;
        RECT 1258.660 1547.690 1258.920 1548.010 ;
        RECT 1256.360 1534.430 1256.620 1534.750 ;
        RECT 1256.420 1497.350 1256.560 1534.430 ;
        RECT 1256.360 1497.030 1256.620 1497.350 ;
        RECT 1260.960 1486.150 1261.220 1486.470 ;
        RECT 1261.020 67.650 1261.160 1486.150 ;
        RECT 1260.960 67.330 1261.220 67.650 ;
        RECT 2622.100 67.330 2622.360 67.650 ;
        RECT 2622.160 3.050 2622.300 67.330 ;
        RECT 2622.100 2.730 2622.360 3.050 ;
        RECT 2625.320 2.730 2625.580 3.050 ;
        RECT 2625.380 2.400 2625.520 2.730 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1263.690 1473.120 1264.010 1473.180 ;
        RECT 1268.290 1473.120 1268.610 1473.180 ;
        RECT 1263.690 1472.980 1268.610 1473.120 ;
        RECT 1263.690 1472.920 1264.010 1472.980 ;
        RECT 1268.290 1472.920 1268.610 1472.980 ;
        RECT 1268.290 67.220 1268.610 67.280 ;
        RECT 2642.770 67.220 2643.090 67.280 ;
        RECT 1268.290 67.080 2643.090 67.220 ;
        RECT 1268.290 67.020 1268.610 67.080 ;
        RECT 2642.770 67.020 2643.090 67.080 ;
      LAYER via ;
        RECT 1263.720 1472.920 1263.980 1473.180 ;
        RECT 1268.320 1472.920 1268.580 1473.180 ;
        RECT 1268.320 67.020 1268.580 67.280 ;
        RECT 2642.800 67.020 2643.060 67.280 ;
      LAYER met2 ;
        RECT 1265.880 1600.450 1266.160 1604.000 ;
        RECT 1264.700 1600.310 1266.160 1600.450 ;
        RECT 1264.700 1546.165 1264.840 1600.310 ;
        RECT 1265.880 1600.000 1266.160 1600.310 ;
        RECT 1264.630 1545.795 1264.910 1546.165 ;
        RECT 1263.710 1545.115 1263.990 1545.485 ;
        RECT 1263.780 1473.210 1263.920 1545.115 ;
        RECT 1263.720 1472.890 1263.980 1473.210 ;
        RECT 1268.320 1472.890 1268.580 1473.210 ;
        RECT 1268.380 67.310 1268.520 1472.890 ;
        RECT 1268.320 66.990 1268.580 67.310 ;
        RECT 2642.800 66.990 2643.060 67.310 ;
        RECT 2642.860 2.960 2643.000 66.990 ;
        RECT 2642.860 2.820 2643.460 2.960 ;
        RECT 2643.320 2.400 2643.460 2.820 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
      LAYER via2 ;
        RECT 1264.630 1545.840 1264.910 1546.120 ;
        RECT 1263.710 1545.160 1263.990 1545.440 ;
      LAYER met3 ;
        RECT 1264.605 1546.130 1264.935 1546.145 ;
        RECT 1263.470 1545.830 1264.935 1546.130 ;
        RECT 1263.470 1545.465 1263.770 1545.830 ;
        RECT 1264.605 1545.815 1264.935 1545.830 ;
        RECT 1263.470 1545.150 1264.015 1545.465 ;
        RECT 1263.685 1545.135 1264.015 1545.150 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1270.205 1497.445 1270.375 1545.555 ;
      LAYER mcon ;
        RECT 1270.205 1545.385 1270.375 1545.555 ;
      LAYER met1 ;
        RECT 1270.130 1545.540 1270.450 1545.600 ;
        RECT 1269.935 1545.400 1270.450 1545.540 ;
        RECT 1270.130 1545.340 1270.450 1545.400 ;
        RECT 1270.145 1497.600 1270.435 1497.645 ;
        RECT 1275.190 1497.600 1275.510 1497.660 ;
        RECT 1270.145 1497.460 1275.510 1497.600 ;
        RECT 1270.145 1497.415 1270.435 1497.460 ;
        RECT 1275.190 1497.400 1275.510 1497.460 ;
        RECT 1275.190 66.880 1275.510 66.940 ;
        RECT 2656.570 66.880 2656.890 66.940 ;
        RECT 1275.190 66.740 2656.890 66.880 ;
        RECT 1275.190 66.680 1275.510 66.740 ;
        RECT 2656.570 66.680 2656.890 66.740 ;
        RECT 2656.570 2.960 2656.890 3.020 ;
        RECT 2661.170 2.960 2661.490 3.020 ;
        RECT 2656.570 2.820 2661.490 2.960 ;
        RECT 2656.570 2.760 2656.890 2.820 ;
        RECT 2661.170 2.760 2661.490 2.820 ;
      LAYER via ;
        RECT 1270.160 1545.340 1270.420 1545.600 ;
        RECT 1275.220 1497.400 1275.480 1497.660 ;
        RECT 1275.220 66.680 1275.480 66.940 ;
        RECT 2656.600 66.680 2656.860 66.940 ;
        RECT 2656.600 2.760 2656.860 3.020 ;
        RECT 2661.200 2.760 2661.460 3.020 ;
      LAYER met2 ;
        RECT 1272.320 1600.450 1272.600 1604.000 ;
        RECT 1270.680 1600.310 1272.600 1600.450 ;
        RECT 1270.680 1546.050 1270.820 1600.310 ;
        RECT 1272.320 1600.000 1272.600 1600.310 ;
        RECT 1270.220 1545.910 1270.820 1546.050 ;
        RECT 1270.220 1545.630 1270.360 1545.910 ;
        RECT 1270.160 1545.310 1270.420 1545.630 ;
        RECT 1275.220 1497.370 1275.480 1497.690 ;
        RECT 1275.280 66.970 1275.420 1497.370 ;
        RECT 1275.220 66.650 1275.480 66.970 ;
        RECT 2656.600 66.650 2656.860 66.970 ;
        RECT 2656.660 3.050 2656.800 66.650 ;
        RECT 2656.600 2.730 2656.860 3.050 ;
        RECT 2661.200 2.730 2661.460 3.050 ;
        RECT 2661.260 2.400 2661.400 2.730 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1279.790 1600.960 1280.110 1601.020 ;
        RECT 1281.630 1600.960 1281.950 1601.020 ;
        RECT 1279.790 1600.820 1281.950 1600.960 ;
        RECT 1279.790 1600.760 1280.110 1600.820 ;
        RECT 1281.630 1600.760 1281.950 1600.820 ;
        RECT 1281.630 66.540 1281.950 66.600 ;
        RECT 2677.270 66.540 2677.590 66.600 ;
        RECT 1281.630 66.400 2677.590 66.540 ;
        RECT 1281.630 66.340 1281.950 66.400 ;
        RECT 2677.270 66.340 2677.590 66.400 ;
      LAYER via ;
        RECT 1279.820 1600.760 1280.080 1601.020 ;
        RECT 1281.660 1600.760 1281.920 1601.020 ;
        RECT 1281.660 66.340 1281.920 66.600 ;
        RECT 2677.300 66.340 2677.560 66.600 ;
      LAYER met2 ;
        RECT 1278.300 1601.130 1278.580 1604.000 ;
        RECT 1278.300 1601.050 1280.020 1601.130 ;
        RECT 1278.300 1600.990 1280.080 1601.050 ;
        RECT 1278.300 1600.000 1278.580 1600.990 ;
        RECT 1279.820 1600.730 1280.080 1600.990 ;
        RECT 1281.660 1600.730 1281.920 1601.050 ;
        RECT 1281.720 66.630 1281.860 1600.730 ;
        RECT 1281.660 66.310 1281.920 66.630 ;
        RECT 2677.300 66.310 2677.560 66.630 ;
        RECT 2677.360 3.130 2677.500 66.310 ;
        RECT 2677.360 2.990 2678.420 3.130 ;
        RECT 2678.280 2.960 2678.420 2.990 ;
        RECT 2678.280 2.820 2678.880 2.960 ;
        RECT 2678.740 2.400 2678.880 2.820 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1284.850 1580.560 1285.170 1580.620 ;
        RECT 1288.990 1580.560 1289.310 1580.620 ;
        RECT 1284.850 1580.420 1289.310 1580.560 ;
        RECT 1284.850 1580.360 1285.170 1580.420 ;
        RECT 1288.990 1580.360 1289.310 1580.420 ;
        RECT 1288.990 66.200 1289.310 66.260 ;
        RECT 2691.070 66.200 2691.390 66.260 ;
        RECT 1288.990 66.060 2691.390 66.200 ;
        RECT 1288.990 66.000 1289.310 66.060 ;
        RECT 2691.070 66.000 2691.390 66.060 ;
        RECT 2691.070 2.960 2691.390 3.020 ;
        RECT 2696.590 2.960 2696.910 3.020 ;
        RECT 2691.070 2.820 2696.910 2.960 ;
        RECT 2691.070 2.760 2691.390 2.820 ;
        RECT 2696.590 2.760 2696.910 2.820 ;
      LAYER via ;
        RECT 1284.880 1580.360 1285.140 1580.620 ;
        RECT 1289.020 1580.360 1289.280 1580.620 ;
        RECT 1289.020 66.000 1289.280 66.260 ;
        RECT 2691.100 66.000 2691.360 66.260 ;
        RECT 2691.100 2.760 2691.360 3.020 ;
        RECT 2696.620 2.760 2696.880 3.020 ;
      LAYER met2 ;
        RECT 1284.740 1600.380 1285.020 1604.000 ;
        RECT 1284.740 1600.000 1285.080 1600.380 ;
        RECT 1284.940 1580.650 1285.080 1600.000 ;
        RECT 1284.880 1580.330 1285.140 1580.650 ;
        RECT 1289.020 1580.330 1289.280 1580.650 ;
        RECT 1289.080 66.290 1289.220 1580.330 ;
        RECT 1289.020 65.970 1289.280 66.290 ;
        RECT 2691.100 65.970 2691.360 66.290 ;
        RECT 2691.160 3.050 2691.300 65.970 ;
        RECT 2691.100 2.730 2691.360 3.050 ;
        RECT 2696.620 2.730 2696.880 3.050 ;
        RECT 2696.680 2.400 2696.820 2.730 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1295.965 65.705 1296.135 113.815 ;
      LAYER mcon ;
        RECT 1295.965 113.645 1296.135 113.815 ;
      LAYER met1 ;
        RECT 1295.890 113.800 1296.210 113.860 ;
        RECT 1295.695 113.660 1296.210 113.800 ;
        RECT 1295.890 113.600 1296.210 113.660 ;
        RECT 1295.905 65.860 1296.195 65.905 ;
        RECT 2711.770 65.860 2712.090 65.920 ;
        RECT 1295.905 65.720 2712.090 65.860 ;
        RECT 1295.905 65.675 1296.195 65.720 ;
        RECT 2711.770 65.660 2712.090 65.720 ;
        RECT 2711.770 2.960 2712.090 3.020 ;
        RECT 2714.530 2.960 2714.850 3.020 ;
        RECT 2711.770 2.820 2714.850 2.960 ;
        RECT 2711.770 2.760 2712.090 2.820 ;
        RECT 2714.530 2.760 2714.850 2.820 ;
      LAYER via ;
        RECT 1295.920 113.600 1296.180 113.860 ;
        RECT 2711.800 65.660 2712.060 65.920 ;
        RECT 2711.800 2.760 2712.060 3.020 ;
        RECT 2714.560 2.760 2714.820 3.020 ;
      LAYER met2 ;
        RECT 1290.720 1601.130 1291.000 1604.000 ;
        RECT 1290.000 1600.990 1291.000 1601.130 ;
        RECT 1290.000 1597.050 1290.140 1600.990 ;
        RECT 1290.720 1600.000 1291.000 1600.990 ;
        RECT 1290.000 1596.910 1290.600 1597.050 ;
        RECT 1290.460 1535.340 1290.600 1596.910 ;
        RECT 1290.460 1535.200 1291.060 1535.340 ;
        RECT 1290.920 1486.890 1291.060 1535.200 ;
        RECT 1290.920 1486.750 1296.120 1486.890 ;
        RECT 1295.980 113.890 1296.120 1486.750 ;
        RECT 1295.920 113.570 1296.180 113.890 ;
        RECT 2711.800 65.630 2712.060 65.950 ;
        RECT 2711.860 3.050 2712.000 65.630 ;
        RECT 2711.800 2.730 2712.060 3.050 ;
        RECT 2714.560 2.730 2714.820 3.050 ;
        RECT 2714.620 2.400 2714.760 2.730 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1301.945 65.365 1302.115 131.155 ;
      LAYER mcon ;
        RECT 1301.945 130.985 1302.115 131.155 ;
      LAYER met1 ;
        RECT 1297.730 1510.520 1298.050 1510.580 ;
        RECT 1302.330 1510.520 1302.650 1510.580 ;
        RECT 1297.730 1510.380 1302.650 1510.520 ;
        RECT 1297.730 1510.320 1298.050 1510.380 ;
        RECT 1302.330 1510.320 1302.650 1510.380 ;
        RECT 1301.410 952.240 1301.730 952.300 ;
        RECT 1302.330 952.240 1302.650 952.300 ;
        RECT 1301.410 952.100 1302.650 952.240 ;
        RECT 1301.410 952.040 1301.730 952.100 ;
        RECT 1302.330 952.040 1302.650 952.100 ;
        RECT 1301.885 131.140 1302.175 131.185 ;
        RECT 1302.330 131.140 1302.650 131.200 ;
        RECT 1301.885 131.000 1302.650 131.140 ;
        RECT 1301.885 130.955 1302.175 131.000 ;
        RECT 1302.330 130.940 1302.650 131.000 ;
        RECT 1301.885 65.520 1302.175 65.565 ;
        RECT 2732.470 65.520 2732.790 65.580 ;
        RECT 1301.885 65.380 2732.790 65.520 ;
        RECT 1301.885 65.335 1302.175 65.380 ;
        RECT 2732.470 65.320 2732.790 65.380 ;
      LAYER via ;
        RECT 1297.760 1510.320 1298.020 1510.580 ;
        RECT 1302.360 1510.320 1302.620 1510.580 ;
        RECT 1301.440 952.040 1301.700 952.300 ;
        RECT 1302.360 952.040 1302.620 952.300 ;
        RECT 1302.360 130.940 1302.620 131.200 ;
        RECT 2732.500 65.320 2732.760 65.580 ;
      LAYER met2 ;
        RECT 1297.160 1600.450 1297.440 1604.000 ;
        RECT 1297.160 1600.310 1297.960 1600.450 ;
        RECT 1297.160 1600.000 1297.440 1600.310 ;
        RECT 1297.820 1510.610 1297.960 1600.310 ;
        RECT 1297.760 1510.290 1298.020 1510.610 ;
        RECT 1302.360 1510.290 1302.620 1510.610 ;
        RECT 1302.420 952.330 1302.560 1510.290 ;
        RECT 1301.440 952.010 1301.700 952.330 ;
        RECT 1302.360 952.010 1302.620 952.330 ;
        RECT 1301.500 904.245 1301.640 952.010 ;
        RECT 1301.430 903.875 1301.710 904.245 ;
        RECT 1302.350 903.875 1302.630 904.245 ;
        RECT 1302.420 131.230 1302.560 903.875 ;
        RECT 1302.360 130.910 1302.620 131.230 ;
        RECT 2732.500 65.290 2732.760 65.610 ;
        RECT 2732.560 2.400 2732.700 65.290 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
      LAYER via2 ;
        RECT 1301.430 903.920 1301.710 904.200 ;
        RECT 1302.350 903.920 1302.630 904.200 ;
      LAYER met3 ;
        RECT 1301.405 904.210 1301.735 904.225 ;
        RECT 1302.325 904.210 1302.655 904.225 ;
        RECT 1301.405 903.910 1302.655 904.210 ;
        RECT 1301.405 903.895 1301.735 903.910 ;
        RECT 1302.325 903.895 1302.655 903.910 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2746.270 2.960 2746.590 3.020 ;
        RECT 2750.410 2.960 2750.730 3.020 ;
        RECT 2746.270 2.820 2750.730 2.960 ;
        RECT 2746.270 2.760 2746.590 2.820 ;
        RECT 2750.410 2.760 2750.730 2.820 ;
      LAYER via ;
        RECT 2746.300 2.760 2746.560 3.020 ;
        RECT 2750.440 2.760 2750.700 3.020 ;
      LAYER met2 ;
        RECT 1303.140 1601.130 1303.420 1604.000 ;
        RECT 1302.420 1600.990 1303.420 1601.130 ;
        RECT 1302.420 1597.050 1302.560 1600.990 ;
        RECT 1303.140 1600.000 1303.420 1600.990 ;
        RECT 1302.420 1596.910 1303.020 1597.050 ;
        RECT 1302.880 68.525 1303.020 1596.910 ;
        RECT 1302.810 68.155 1303.090 68.525 ;
        RECT 2746.290 68.155 2746.570 68.525 ;
        RECT 2746.360 3.050 2746.500 68.155 ;
        RECT 2746.300 2.730 2746.560 3.050 ;
        RECT 2750.440 2.730 2750.700 3.050 ;
        RECT 2750.500 2.400 2750.640 2.730 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
      LAYER via2 ;
        RECT 1302.810 68.200 1303.090 68.480 ;
        RECT 2746.290 68.200 2746.570 68.480 ;
      LAYER met3 ;
        RECT 1302.785 68.490 1303.115 68.505 ;
        RECT 2746.265 68.490 2746.595 68.505 ;
        RECT 1302.785 68.190 2746.595 68.490 ;
        RECT 1302.785 68.175 1303.115 68.190 ;
        RECT 2746.265 68.175 2746.595 68.190 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1304.170 1600.960 1304.490 1601.020 ;
        RECT 1307.850 1600.960 1308.170 1601.020 ;
        RECT 1304.170 1600.820 1308.170 1600.960 ;
        RECT 1304.170 1600.760 1304.490 1600.820 ;
        RECT 1307.850 1600.760 1308.170 1600.820 ;
      LAYER via ;
        RECT 1304.200 1600.760 1304.460 1601.020 ;
        RECT 1307.880 1600.760 1308.140 1601.020 ;
      LAYER met2 ;
        RECT 1309.120 1601.130 1309.400 1604.000 ;
        RECT 1307.940 1601.050 1309.400 1601.130 ;
        RECT 1304.200 1600.730 1304.460 1601.050 ;
        RECT 1307.880 1600.990 1309.400 1601.050 ;
        RECT 1307.880 1600.730 1308.140 1600.990 ;
        RECT 1304.260 1535.340 1304.400 1600.730 ;
        RECT 1309.120 1600.000 1309.400 1600.990 ;
        RECT 1304.260 1535.200 1304.860 1535.340 ;
        RECT 1304.720 1486.890 1304.860 1535.200 ;
        RECT 1304.720 1486.750 1309.920 1486.890 ;
        RECT 1309.780 67.845 1309.920 1486.750 ;
        RECT 1309.710 67.475 1309.990 67.845 ;
        RECT 2766.990 67.475 2767.270 67.845 ;
        RECT 2767.060 3.130 2767.200 67.475 ;
        RECT 2767.060 2.990 2768.120 3.130 ;
        RECT 2767.980 2.400 2768.120 2.990 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
      LAYER via2 ;
        RECT 1309.710 67.520 1309.990 67.800 ;
        RECT 2766.990 67.520 2767.270 67.800 ;
      LAYER met3 ;
        RECT 1309.685 67.810 1310.015 67.825 ;
        RECT 2766.965 67.810 2767.295 67.825 ;
        RECT 1309.685 67.510 2767.295 67.810 ;
        RECT 1309.685 67.495 1310.015 67.510 ;
        RECT 2766.965 67.495 2767.295 67.510 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 738.445 1586.865 738.615 1591.115 ;
        RECT 758.685 1587.205 758.855 1590.775 ;
        RECT 806.065 15.725 806.235 37.315 ;
      LAYER mcon ;
        RECT 738.445 1590.945 738.615 1591.115 ;
        RECT 758.685 1590.605 758.855 1590.775 ;
        RECT 806.065 37.145 806.235 37.315 ;
      LAYER met1 ;
        RECT 641.310 1591.100 641.630 1591.160 ;
        RECT 738.385 1591.100 738.675 1591.145 ;
        RECT 641.310 1590.960 738.675 1591.100 ;
        RECT 641.310 1590.900 641.630 1590.960 ;
        RECT 738.385 1590.915 738.675 1590.960 ;
        RECT 758.625 1590.760 758.915 1590.805 ;
        RECT 782.990 1590.760 783.310 1590.820 ;
        RECT 758.625 1590.620 783.310 1590.760 ;
        RECT 758.625 1590.575 758.915 1590.620 ;
        RECT 782.990 1590.560 783.310 1590.620 ;
        RECT 758.625 1587.360 758.915 1587.405 ;
        RECT 745.360 1587.220 758.915 1587.360 ;
        RECT 738.385 1587.020 738.675 1587.065 ;
        RECT 745.360 1587.020 745.500 1587.220 ;
        RECT 758.625 1587.175 758.915 1587.220 ;
        RECT 738.385 1586.880 745.500 1587.020 ;
        RECT 738.385 1586.835 738.675 1586.880 ;
        RECT 782.990 37.300 783.310 37.360 ;
        RECT 806.005 37.300 806.295 37.345 ;
        RECT 782.990 37.160 806.295 37.300 ;
        RECT 782.990 37.100 783.310 37.160 ;
        RECT 806.005 37.115 806.295 37.160 ;
        RECT 806.005 15.880 806.295 15.925 ;
        RECT 840.950 15.880 841.270 15.940 ;
        RECT 806.005 15.740 841.270 15.880 ;
        RECT 806.005 15.695 806.295 15.740 ;
        RECT 840.950 15.680 841.270 15.740 ;
      LAYER via ;
        RECT 641.340 1590.900 641.600 1591.160 ;
        RECT 783.020 1590.560 783.280 1590.820 ;
        RECT 783.020 37.100 783.280 37.360 ;
        RECT 840.980 15.680 841.240 15.940 ;
      LAYER met2 ;
        RECT 641.200 1600.380 641.480 1604.000 ;
        RECT 641.200 1600.000 641.540 1600.380 ;
        RECT 641.400 1591.190 641.540 1600.000 ;
        RECT 641.340 1590.870 641.600 1591.190 ;
        RECT 783.020 1590.530 783.280 1590.850 ;
        RECT 783.080 37.390 783.220 1590.530 ;
        RECT 783.020 37.070 783.280 37.390 ;
        RECT 840.980 15.650 841.240 15.970 ;
        RECT 841.040 2.400 841.180 15.650 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.530 1563.900 1311.850 1563.960 ;
        RECT 1313.830 1563.900 1314.150 1563.960 ;
        RECT 1311.530 1563.760 1314.150 1563.900 ;
        RECT 1311.530 1563.700 1311.850 1563.760 ;
        RECT 1313.830 1563.700 1314.150 1563.760 ;
        RECT 1311.530 1530.240 1311.850 1530.300 ;
        RECT 1316.130 1530.240 1316.450 1530.300 ;
        RECT 1311.530 1530.100 1316.450 1530.240 ;
        RECT 1311.530 1530.040 1311.850 1530.100 ;
        RECT 1316.130 1530.040 1316.450 1530.100 ;
        RECT 2780.770 2.960 2781.090 3.020 ;
        RECT 2785.830 2.960 2786.150 3.020 ;
        RECT 2780.770 2.820 2786.150 2.960 ;
        RECT 2780.770 2.760 2781.090 2.820 ;
        RECT 2785.830 2.760 2786.150 2.820 ;
      LAYER via ;
        RECT 1311.560 1563.700 1311.820 1563.960 ;
        RECT 1313.860 1563.700 1314.120 1563.960 ;
        RECT 1311.560 1530.040 1311.820 1530.300 ;
        RECT 1316.160 1530.040 1316.420 1530.300 ;
        RECT 2780.800 2.760 2781.060 3.020 ;
        RECT 2785.860 2.760 2786.120 3.020 ;
      LAYER met2 ;
        RECT 1315.560 1600.450 1315.840 1604.000 ;
        RECT 1313.920 1600.310 1315.840 1600.450 ;
        RECT 1313.920 1563.990 1314.060 1600.310 ;
        RECT 1315.560 1600.000 1315.840 1600.310 ;
        RECT 1311.560 1563.670 1311.820 1563.990 ;
        RECT 1313.860 1563.670 1314.120 1563.990 ;
        RECT 1311.620 1530.330 1311.760 1563.670 ;
        RECT 1311.560 1530.010 1311.820 1530.330 ;
        RECT 1316.160 1530.010 1316.420 1530.330 ;
        RECT 1316.220 67.165 1316.360 1530.010 ;
        RECT 1316.150 66.795 1316.430 67.165 ;
        RECT 2780.790 66.795 2781.070 67.165 ;
        RECT 2780.860 3.050 2781.000 66.795 ;
        RECT 2780.800 2.730 2781.060 3.050 ;
        RECT 2785.860 2.730 2786.120 3.050 ;
        RECT 2785.920 2.400 2786.060 2.730 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
      LAYER via2 ;
        RECT 1316.150 66.840 1316.430 67.120 ;
        RECT 2780.790 66.840 2781.070 67.120 ;
      LAYER met3 ;
        RECT 1316.125 67.130 1316.455 67.145 ;
        RECT 2780.765 67.130 2781.095 67.145 ;
        RECT 1316.125 66.830 2781.095 67.130 ;
        RECT 1316.125 66.815 1316.455 66.830 ;
        RECT 2780.765 66.815 2781.095 66.830 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1323.105 1324.725 1323.275 1373.175 ;
        RECT 1323.105 928.285 1323.275 962.795 ;
        RECT 1323.105 800.445 1323.275 848.555 ;
        RECT 1323.105 510.765 1323.275 558.535 ;
        RECT 1323.105 414.205 1323.275 461.975 ;
        RECT 1323.105 221.425 1323.275 268.855 ;
      LAYER mcon ;
        RECT 1323.105 1373.005 1323.275 1373.175 ;
        RECT 1323.105 962.625 1323.275 962.795 ;
        RECT 1323.105 848.385 1323.275 848.555 ;
        RECT 1323.105 558.365 1323.275 558.535 ;
        RECT 1323.105 461.805 1323.275 461.975 ;
        RECT 1323.105 268.685 1323.275 268.855 ;
      LAYER met1 ;
        RECT 1317.970 1600.960 1318.290 1601.020 ;
        RECT 1320.270 1600.960 1320.590 1601.020 ;
        RECT 1317.970 1600.820 1320.590 1600.960 ;
        RECT 1317.970 1600.760 1318.290 1600.820 ;
        RECT 1320.270 1600.760 1320.590 1600.820 ;
        RECT 1322.570 1421.440 1322.890 1421.500 ;
        RECT 1323.490 1421.440 1323.810 1421.500 ;
        RECT 1322.570 1421.300 1323.810 1421.440 ;
        RECT 1322.570 1421.240 1322.890 1421.300 ;
        RECT 1323.490 1421.240 1323.810 1421.300 ;
        RECT 1323.045 1373.160 1323.335 1373.205 ;
        RECT 1323.490 1373.160 1323.810 1373.220 ;
        RECT 1323.045 1373.020 1323.810 1373.160 ;
        RECT 1323.045 1372.975 1323.335 1373.020 ;
        RECT 1323.490 1372.960 1323.810 1373.020 ;
        RECT 1323.030 1324.880 1323.350 1324.940 ;
        RECT 1322.835 1324.740 1323.350 1324.880 ;
        RECT 1323.030 1324.680 1323.350 1324.740 ;
        RECT 1323.030 962.780 1323.350 962.840 ;
        RECT 1322.835 962.640 1323.350 962.780 ;
        RECT 1323.030 962.580 1323.350 962.640 ;
        RECT 1323.030 928.440 1323.350 928.500 ;
        RECT 1322.835 928.300 1323.350 928.440 ;
        RECT 1323.030 928.240 1323.350 928.300 ;
        RECT 1323.030 848.540 1323.350 848.600 ;
        RECT 1322.835 848.400 1323.350 848.540 ;
        RECT 1323.030 848.340 1323.350 848.400 ;
        RECT 1323.030 800.600 1323.350 800.660 ;
        RECT 1322.835 800.460 1323.350 800.600 ;
        RECT 1323.030 800.400 1323.350 800.460 ;
        RECT 1322.570 752.320 1322.890 752.380 ;
        RECT 1323.030 752.320 1323.350 752.380 ;
        RECT 1322.570 752.180 1323.350 752.320 ;
        RECT 1322.570 752.120 1322.890 752.180 ;
        RECT 1323.030 752.120 1323.350 752.180 ;
        RECT 1322.570 704.040 1322.890 704.100 ;
        RECT 1323.030 704.040 1323.350 704.100 ;
        RECT 1322.570 703.900 1323.350 704.040 ;
        RECT 1322.570 703.840 1322.890 703.900 ;
        RECT 1323.030 703.840 1323.350 703.900 ;
        RECT 1322.570 655.760 1322.890 655.820 ;
        RECT 1323.030 655.760 1323.350 655.820 ;
        RECT 1322.570 655.620 1323.350 655.760 ;
        RECT 1322.570 655.560 1322.890 655.620 ;
        RECT 1323.030 655.560 1323.350 655.620 ;
        RECT 1322.570 607.480 1322.890 607.540 ;
        RECT 1323.030 607.480 1323.350 607.540 ;
        RECT 1322.570 607.340 1323.350 607.480 ;
        RECT 1322.570 607.280 1322.890 607.340 ;
        RECT 1323.030 607.280 1323.350 607.340 ;
        RECT 1322.570 559.200 1322.890 559.260 ;
        RECT 1323.030 559.200 1323.350 559.260 ;
        RECT 1322.570 559.060 1323.350 559.200 ;
        RECT 1322.570 559.000 1322.890 559.060 ;
        RECT 1323.030 559.000 1323.350 559.060 ;
        RECT 1323.030 558.520 1323.350 558.580 ;
        RECT 1322.835 558.380 1323.350 558.520 ;
        RECT 1323.030 558.320 1323.350 558.380 ;
        RECT 1323.030 510.920 1323.350 510.980 ;
        RECT 1322.835 510.780 1323.350 510.920 ;
        RECT 1323.030 510.720 1323.350 510.780 ;
        RECT 1322.570 462.640 1322.890 462.700 ;
        RECT 1323.030 462.640 1323.350 462.700 ;
        RECT 1322.570 462.500 1323.350 462.640 ;
        RECT 1322.570 462.440 1322.890 462.500 ;
        RECT 1323.030 462.440 1323.350 462.500 ;
        RECT 1323.030 461.960 1323.350 462.020 ;
        RECT 1322.835 461.820 1323.350 461.960 ;
        RECT 1323.030 461.760 1323.350 461.820 ;
        RECT 1323.030 414.360 1323.350 414.420 ;
        RECT 1322.835 414.220 1323.350 414.360 ;
        RECT 1323.030 414.160 1323.350 414.220 ;
        RECT 1322.570 366.080 1322.890 366.140 ;
        RECT 1323.030 366.080 1323.350 366.140 ;
        RECT 1322.570 365.940 1323.350 366.080 ;
        RECT 1322.570 365.880 1322.890 365.940 ;
        RECT 1323.030 365.880 1323.350 365.940 ;
        RECT 1323.030 268.840 1323.350 268.900 ;
        RECT 1322.835 268.700 1323.350 268.840 ;
        RECT 1323.030 268.640 1323.350 268.700 ;
        RECT 1323.030 221.580 1323.350 221.640 ;
        RECT 1322.835 221.440 1323.350 221.580 ;
        RECT 1323.030 221.380 1323.350 221.440 ;
        RECT 1322.110 166.160 1322.430 166.220 ;
        RECT 1323.030 166.160 1323.350 166.220 ;
        RECT 1322.110 166.020 1323.350 166.160 ;
        RECT 1322.110 165.960 1322.430 166.020 ;
        RECT 1323.030 165.960 1323.350 166.020 ;
        RECT 1322.110 124.340 1322.430 124.400 ;
        RECT 1323.490 124.340 1323.810 124.400 ;
        RECT 1322.110 124.200 1323.810 124.340 ;
        RECT 1322.110 124.140 1322.430 124.200 ;
        RECT 1323.490 124.140 1323.810 124.200 ;
      LAYER via ;
        RECT 1318.000 1600.760 1318.260 1601.020 ;
        RECT 1320.300 1600.760 1320.560 1601.020 ;
        RECT 1322.600 1421.240 1322.860 1421.500 ;
        RECT 1323.520 1421.240 1323.780 1421.500 ;
        RECT 1323.520 1372.960 1323.780 1373.220 ;
        RECT 1323.060 1324.680 1323.320 1324.940 ;
        RECT 1323.060 962.580 1323.320 962.840 ;
        RECT 1323.060 928.240 1323.320 928.500 ;
        RECT 1323.060 848.340 1323.320 848.600 ;
        RECT 1323.060 800.400 1323.320 800.660 ;
        RECT 1322.600 752.120 1322.860 752.380 ;
        RECT 1323.060 752.120 1323.320 752.380 ;
        RECT 1322.600 703.840 1322.860 704.100 ;
        RECT 1323.060 703.840 1323.320 704.100 ;
        RECT 1322.600 655.560 1322.860 655.820 ;
        RECT 1323.060 655.560 1323.320 655.820 ;
        RECT 1322.600 607.280 1322.860 607.540 ;
        RECT 1323.060 607.280 1323.320 607.540 ;
        RECT 1322.600 559.000 1322.860 559.260 ;
        RECT 1323.060 559.000 1323.320 559.260 ;
        RECT 1323.060 558.320 1323.320 558.580 ;
        RECT 1323.060 510.720 1323.320 510.980 ;
        RECT 1322.600 462.440 1322.860 462.700 ;
        RECT 1323.060 462.440 1323.320 462.700 ;
        RECT 1323.060 461.760 1323.320 462.020 ;
        RECT 1323.060 414.160 1323.320 414.420 ;
        RECT 1322.600 365.880 1322.860 366.140 ;
        RECT 1323.060 365.880 1323.320 366.140 ;
        RECT 1323.060 268.640 1323.320 268.900 ;
        RECT 1323.060 221.380 1323.320 221.640 ;
        RECT 1322.140 165.960 1322.400 166.220 ;
        RECT 1323.060 165.960 1323.320 166.220 ;
        RECT 1322.140 124.140 1322.400 124.400 ;
        RECT 1323.520 124.140 1323.780 124.400 ;
      LAYER met2 ;
        RECT 1321.540 1601.130 1321.820 1604.000 ;
        RECT 1320.360 1601.050 1321.820 1601.130 ;
        RECT 1318.000 1600.730 1318.260 1601.050 ;
        RECT 1320.300 1600.990 1321.820 1601.050 ;
        RECT 1320.300 1600.730 1320.560 1600.990 ;
        RECT 1318.060 1535.170 1318.200 1600.730 ;
        RECT 1321.540 1600.000 1321.820 1600.990 ;
        RECT 1318.060 1535.030 1318.660 1535.170 ;
        RECT 1318.520 1470.005 1318.660 1535.030 ;
        RECT 1318.450 1469.635 1318.730 1470.005 ;
        RECT 1323.510 1469.635 1323.790 1470.005 ;
        RECT 1323.580 1421.530 1323.720 1469.635 ;
        RECT 1322.600 1421.210 1322.860 1421.530 ;
        RECT 1323.520 1421.210 1323.780 1421.530 ;
        RECT 1322.660 1373.445 1322.800 1421.210 ;
        RECT 1322.590 1373.075 1322.870 1373.445 ;
        RECT 1323.510 1373.075 1323.790 1373.445 ;
        RECT 1323.520 1372.930 1323.780 1373.075 ;
        RECT 1323.060 1324.650 1323.320 1324.970 ;
        RECT 1323.120 962.870 1323.260 1324.650 ;
        RECT 1323.060 962.550 1323.320 962.870 ;
        RECT 1323.060 928.210 1323.320 928.530 ;
        RECT 1323.120 904.130 1323.260 928.210 ;
        RECT 1323.120 903.990 1323.720 904.130 ;
        RECT 1323.580 849.050 1323.720 903.990 ;
        RECT 1323.120 848.910 1323.720 849.050 ;
        RECT 1323.120 848.630 1323.260 848.910 ;
        RECT 1323.060 848.310 1323.320 848.630 ;
        RECT 1323.060 800.370 1323.320 800.690 ;
        RECT 1323.120 800.090 1323.260 800.370 ;
        RECT 1322.660 799.950 1323.260 800.090 ;
        RECT 1322.660 752.410 1322.800 799.950 ;
        RECT 1322.600 752.090 1322.860 752.410 ;
        RECT 1323.060 752.090 1323.320 752.410 ;
        RECT 1323.120 751.810 1323.260 752.090 ;
        RECT 1322.660 751.670 1323.260 751.810 ;
        RECT 1322.660 704.130 1322.800 751.670 ;
        RECT 1322.600 703.810 1322.860 704.130 ;
        RECT 1323.060 703.810 1323.320 704.130 ;
        RECT 1323.120 703.530 1323.260 703.810 ;
        RECT 1322.660 703.390 1323.260 703.530 ;
        RECT 1322.660 655.850 1322.800 703.390 ;
        RECT 1322.600 655.530 1322.860 655.850 ;
        RECT 1323.060 655.530 1323.320 655.850 ;
        RECT 1323.120 655.250 1323.260 655.530 ;
        RECT 1322.660 655.110 1323.260 655.250 ;
        RECT 1322.660 607.570 1322.800 655.110 ;
        RECT 1322.600 607.250 1322.860 607.570 ;
        RECT 1323.060 607.250 1323.320 607.570 ;
        RECT 1323.120 606.970 1323.260 607.250 ;
        RECT 1322.660 606.830 1323.260 606.970 ;
        RECT 1322.660 559.290 1322.800 606.830 ;
        RECT 1322.600 558.970 1322.860 559.290 ;
        RECT 1323.060 558.970 1323.320 559.290 ;
        RECT 1323.120 558.610 1323.260 558.970 ;
        RECT 1323.060 558.290 1323.320 558.610 ;
        RECT 1323.060 510.690 1323.320 511.010 ;
        RECT 1323.120 510.410 1323.260 510.690 ;
        RECT 1322.660 510.270 1323.260 510.410 ;
        RECT 1322.660 462.730 1322.800 510.270 ;
        RECT 1322.600 462.410 1322.860 462.730 ;
        RECT 1323.060 462.410 1323.320 462.730 ;
        RECT 1323.120 462.050 1323.260 462.410 ;
        RECT 1323.060 461.730 1323.320 462.050 ;
        RECT 1323.060 414.130 1323.320 414.450 ;
        RECT 1323.120 413.850 1323.260 414.130 ;
        RECT 1322.660 413.710 1323.260 413.850 ;
        RECT 1322.660 366.170 1322.800 413.710 ;
        RECT 1322.600 365.850 1322.860 366.170 ;
        RECT 1323.060 365.850 1323.320 366.170 ;
        RECT 1323.120 268.930 1323.260 365.850 ;
        RECT 1323.060 268.610 1323.320 268.930 ;
        RECT 1323.060 221.350 1323.320 221.670 ;
        RECT 1323.120 166.250 1323.260 221.350 ;
        RECT 1322.140 165.930 1322.400 166.250 ;
        RECT 1323.060 165.930 1323.320 166.250 ;
        RECT 1322.200 124.430 1322.340 165.930 ;
        RECT 1322.140 124.110 1322.400 124.430 ;
        RECT 1323.520 124.110 1323.780 124.430 ;
        RECT 1323.580 76.005 1323.720 124.110 ;
        RECT 1323.510 75.635 1323.790 76.005 ;
        RECT 1325.810 74.955 1326.090 75.325 ;
        RECT 1325.880 66.485 1326.020 74.955 ;
        RECT 1325.810 66.115 1326.090 66.485 ;
        RECT 2801.490 66.115 2801.770 66.485 ;
        RECT 2801.560 3.130 2801.700 66.115 ;
        RECT 2801.560 2.990 2804.000 3.130 ;
        RECT 2803.860 2.400 2804.000 2.990 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
      LAYER via2 ;
        RECT 1318.450 1469.680 1318.730 1469.960 ;
        RECT 1323.510 1469.680 1323.790 1469.960 ;
        RECT 1322.590 1373.120 1322.870 1373.400 ;
        RECT 1323.510 1373.120 1323.790 1373.400 ;
        RECT 1323.510 75.680 1323.790 75.960 ;
        RECT 1325.810 75.000 1326.090 75.280 ;
        RECT 1325.810 66.160 1326.090 66.440 ;
        RECT 2801.490 66.160 2801.770 66.440 ;
      LAYER met3 ;
        RECT 1318.425 1469.970 1318.755 1469.985 ;
        RECT 1323.485 1469.970 1323.815 1469.985 ;
        RECT 1318.425 1469.670 1323.815 1469.970 ;
        RECT 1318.425 1469.655 1318.755 1469.670 ;
        RECT 1323.485 1469.655 1323.815 1469.670 ;
        RECT 1322.565 1373.410 1322.895 1373.425 ;
        RECT 1323.485 1373.410 1323.815 1373.425 ;
        RECT 1322.565 1373.110 1323.815 1373.410 ;
        RECT 1322.565 1373.095 1322.895 1373.110 ;
        RECT 1323.485 1373.095 1323.815 1373.110 ;
        RECT 1323.485 75.655 1323.815 75.985 ;
        RECT 1323.500 75.290 1323.800 75.655 ;
        RECT 1325.785 75.290 1326.115 75.305 ;
        RECT 1323.500 74.990 1326.115 75.290 ;
        RECT 1325.785 74.975 1326.115 74.990 ;
        RECT 1325.785 66.450 1326.115 66.465 ;
        RECT 2801.465 66.450 2801.795 66.465 ;
        RECT 1325.785 66.150 2801.795 66.450 ;
        RECT 1325.785 66.135 1326.115 66.150 ;
        RECT 2801.465 66.135 2801.795 66.150 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1329.085 1463.105 1329.255 1510.875 ;
        RECT 1330.005 1090.125 1330.175 1152.515 ;
        RECT 1330.005 848.725 1330.175 896.835 ;
        RECT 1330.005 752.165 1330.175 800.275 ;
        RECT 1330.005 655.605 1330.175 703.715 ;
        RECT 1330.005 559.045 1330.175 607.155 ;
        RECT 1330.005 462.485 1330.175 510.595 ;
        RECT 1330.005 365.925 1330.175 414.035 ;
      LAYER mcon ;
        RECT 1329.085 1510.705 1329.255 1510.875 ;
        RECT 1330.005 1152.345 1330.175 1152.515 ;
        RECT 1330.005 896.665 1330.175 896.835 ;
        RECT 1330.005 800.105 1330.175 800.275 ;
        RECT 1330.005 703.545 1330.175 703.715 ;
        RECT 1330.005 606.985 1330.175 607.155 ;
        RECT 1330.005 510.425 1330.175 510.595 ;
        RECT 1330.005 413.865 1330.175 414.035 ;
      LAYER met1 ;
        RECT 1329.010 1510.860 1329.330 1510.920 ;
        RECT 1328.815 1510.720 1329.330 1510.860 ;
        RECT 1329.010 1510.660 1329.330 1510.720 ;
        RECT 1329.025 1463.260 1329.315 1463.305 ;
        RECT 1329.470 1463.260 1329.790 1463.320 ;
        RECT 1329.025 1463.120 1329.790 1463.260 ;
        RECT 1329.025 1463.075 1329.315 1463.120 ;
        RECT 1329.470 1463.060 1329.790 1463.120 ;
        RECT 1329.470 1462.380 1329.790 1462.640 ;
        RECT 1329.560 1462.240 1329.700 1462.380 ;
        RECT 1329.930 1462.240 1330.250 1462.300 ;
        RECT 1329.560 1462.100 1330.250 1462.240 ;
        RECT 1329.930 1462.040 1330.250 1462.100 ;
        RECT 1329.930 1152.500 1330.250 1152.560 ;
        RECT 1329.735 1152.360 1330.250 1152.500 ;
        RECT 1329.930 1152.300 1330.250 1152.360 ;
        RECT 1329.930 1090.280 1330.250 1090.340 ;
        RECT 1329.735 1090.140 1330.250 1090.280 ;
        RECT 1329.930 1090.080 1330.250 1090.140 ;
        RECT 1329.930 904.780 1330.250 905.040 ;
        RECT 1330.020 904.360 1330.160 904.780 ;
        RECT 1329.930 904.100 1330.250 904.360 ;
        RECT 1329.930 896.820 1330.250 896.880 ;
        RECT 1329.735 896.680 1330.250 896.820 ;
        RECT 1329.930 896.620 1330.250 896.680 ;
        RECT 1329.930 848.880 1330.250 848.940 ;
        RECT 1329.735 848.740 1330.250 848.880 ;
        RECT 1329.930 848.680 1330.250 848.740 ;
        RECT 1329.930 800.260 1330.250 800.320 ;
        RECT 1329.735 800.120 1330.250 800.260 ;
        RECT 1329.930 800.060 1330.250 800.120 ;
        RECT 1329.930 752.320 1330.250 752.380 ;
        RECT 1329.735 752.180 1330.250 752.320 ;
        RECT 1329.930 752.120 1330.250 752.180 ;
        RECT 1329.930 703.700 1330.250 703.760 ;
        RECT 1329.735 703.560 1330.250 703.700 ;
        RECT 1329.930 703.500 1330.250 703.560 ;
        RECT 1329.930 655.760 1330.250 655.820 ;
        RECT 1329.735 655.620 1330.250 655.760 ;
        RECT 1329.930 655.560 1330.250 655.620 ;
        RECT 1329.930 607.140 1330.250 607.200 ;
        RECT 1329.735 607.000 1330.250 607.140 ;
        RECT 1329.930 606.940 1330.250 607.000 ;
        RECT 1329.930 559.200 1330.250 559.260 ;
        RECT 1329.735 559.060 1330.250 559.200 ;
        RECT 1329.930 559.000 1330.250 559.060 ;
        RECT 1329.930 510.580 1330.250 510.640 ;
        RECT 1329.735 510.440 1330.250 510.580 ;
        RECT 1329.930 510.380 1330.250 510.440 ;
        RECT 1329.930 462.640 1330.250 462.700 ;
        RECT 1329.735 462.500 1330.250 462.640 ;
        RECT 1329.930 462.440 1330.250 462.500 ;
        RECT 1329.930 414.020 1330.250 414.080 ;
        RECT 1329.735 413.880 1330.250 414.020 ;
        RECT 1329.930 413.820 1330.250 413.880 ;
        RECT 1329.930 366.080 1330.250 366.140 ;
        RECT 1329.735 365.940 1330.250 366.080 ;
        RECT 1329.930 365.880 1330.250 365.940 ;
        RECT 2815.270 17.580 2815.590 17.640 ;
        RECT 2821.710 17.580 2822.030 17.640 ;
        RECT 2815.270 17.440 2822.030 17.580 ;
        RECT 2815.270 17.380 2815.590 17.440 ;
        RECT 2821.710 17.380 2822.030 17.440 ;
      LAYER via ;
        RECT 1329.040 1510.660 1329.300 1510.920 ;
        RECT 1329.500 1463.060 1329.760 1463.320 ;
        RECT 1329.500 1462.380 1329.760 1462.640 ;
        RECT 1329.960 1462.040 1330.220 1462.300 ;
        RECT 1329.960 1152.300 1330.220 1152.560 ;
        RECT 1329.960 1090.080 1330.220 1090.340 ;
        RECT 1329.960 904.780 1330.220 905.040 ;
        RECT 1329.960 904.100 1330.220 904.360 ;
        RECT 1329.960 896.620 1330.220 896.880 ;
        RECT 1329.960 848.680 1330.220 848.940 ;
        RECT 1329.960 800.060 1330.220 800.320 ;
        RECT 1329.960 752.120 1330.220 752.380 ;
        RECT 1329.960 703.500 1330.220 703.760 ;
        RECT 1329.960 655.560 1330.220 655.820 ;
        RECT 1329.960 606.940 1330.220 607.200 ;
        RECT 1329.960 559.000 1330.220 559.260 ;
        RECT 1329.960 510.380 1330.220 510.640 ;
        RECT 1329.960 462.440 1330.220 462.700 ;
        RECT 1329.960 413.820 1330.220 414.080 ;
        RECT 1329.960 365.880 1330.220 366.140 ;
        RECT 2815.300 17.380 2815.560 17.640 ;
        RECT 2821.740 17.380 2822.000 17.640 ;
      LAYER met2 ;
        RECT 1327.980 1600.450 1328.260 1604.000 ;
        RECT 1326.800 1600.310 1328.260 1600.450 ;
        RECT 1326.800 1573.365 1326.940 1600.310 ;
        RECT 1327.980 1600.000 1328.260 1600.310 ;
        RECT 1326.730 1572.995 1327.010 1573.365 ;
        RECT 1329.030 1572.995 1329.310 1573.365 ;
        RECT 1329.100 1510.950 1329.240 1572.995 ;
        RECT 1329.040 1510.630 1329.300 1510.950 ;
        RECT 1329.500 1463.030 1329.760 1463.350 ;
        RECT 1329.560 1462.670 1329.700 1463.030 ;
        RECT 1329.500 1462.350 1329.760 1462.670 ;
        RECT 1329.960 1462.010 1330.220 1462.330 ;
        RECT 1330.020 1152.590 1330.160 1462.010 ;
        RECT 1329.960 1152.270 1330.220 1152.590 ;
        RECT 1329.960 1090.050 1330.220 1090.370 ;
        RECT 1330.020 905.070 1330.160 1090.050 ;
        RECT 1329.960 904.750 1330.220 905.070 ;
        RECT 1329.960 904.070 1330.220 904.390 ;
        RECT 1330.020 896.910 1330.160 904.070 ;
        RECT 1329.960 896.590 1330.220 896.910 ;
        RECT 1329.960 848.650 1330.220 848.970 ;
        RECT 1330.020 800.350 1330.160 848.650 ;
        RECT 1329.960 800.030 1330.220 800.350 ;
        RECT 1329.960 752.090 1330.220 752.410 ;
        RECT 1330.020 703.790 1330.160 752.090 ;
        RECT 1329.960 703.470 1330.220 703.790 ;
        RECT 1329.960 655.530 1330.220 655.850 ;
        RECT 1330.020 607.230 1330.160 655.530 ;
        RECT 1329.960 606.910 1330.220 607.230 ;
        RECT 1329.960 558.970 1330.220 559.290 ;
        RECT 1330.020 510.670 1330.160 558.970 ;
        RECT 1329.960 510.350 1330.220 510.670 ;
        RECT 1329.960 462.410 1330.220 462.730 ;
        RECT 1330.020 414.110 1330.160 462.410 ;
        RECT 1329.960 413.790 1330.220 414.110 ;
        RECT 1329.960 365.850 1330.220 366.170 ;
        RECT 1330.020 179.250 1330.160 365.850 ;
        RECT 1330.020 179.110 1330.620 179.250 ;
        RECT 1330.480 65.805 1330.620 179.110 ;
        RECT 1330.410 65.435 1330.690 65.805 ;
        RECT 2815.290 65.435 2815.570 65.805 ;
        RECT 2815.360 17.670 2815.500 65.435 ;
        RECT 2815.300 17.350 2815.560 17.670 ;
        RECT 2821.740 17.350 2822.000 17.670 ;
        RECT 2821.800 2.400 2821.940 17.350 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
      LAYER via2 ;
        RECT 1326.730 1573.040 1327.010 1573.320 ;
        RECT 1329.030 1573.040 1329.310 1573.320 ;
        RECT 1330.410 65.480 1330.690 65.760 ;
        RECT 2815.290 65.480 2815.570 65.760 ;
      LAYER met3 ;
        RECT 1326.705 1573.330 1327.035 1573.345 ;
        RECT 1329.005 1573.330 1329.335 1573.345 ;
        RECT 1326.705 1573.030 1329.335 1573.330 ;
        RECT 1326.705 1573.015 1327.035 1573.030 ;
        RECT 1329.005 1573.015 1329.335 1573.030 ;
        RECT 1330.385 65.770 1330.715 65.785 ;
        RECT 2815.265 65.770 2815.595 65.785 ;
        RECT 1330.385 65.470 2815.595 65.770 ;
        RECT 1330.385 65.455 1330.715 65.470 ;
        RECT 2815.265 65.455 2815.595 65.470 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1335.525 1497.105 1335.695 1518.015 ;
        RECT 1335.985 1414.485 1336.155 1438.795 ;
        RECT 1336.445 848.725 1336.615 896.835 ;
        RECT 1336.445 752.165 1336.615 800.275 ;
        RECT 1336.445 655.605 1336.615 703.715 ;
        RECT 1336.905 559.045 1337.075 607.155 ;
        RECT 1336.445 462.485 1336.615 510.595 ;
        RECT 1336.445 365.925 1336.615 414.035 ;
        RECT 1336.445 269.025 1336.615 317.475 ;
        RECT 1336.445 178.925 1336.615 220.575 ;
      LAYER mcon ;
        RECT 1335.525 1517.845 1335.695 1518.015 ;
        RECT 1335.985 1438.625 1336.155 1438.795 ;
        RECT 1336.445 896.665 1336.615 896.835 ;
        RECT 1336.445 800.105 1336.615 800.275 ;
        RECT 1336.445 703.545 1336.615 703.715 ;
        RECT 1336.905 606.985 1337.075 607.155 ;
        RECT 1336.445 510.425 1336.615 510.595 ;
        RECT 1336.445 413.865 1336.615 414.035 ;
        RECT 1336.445 317.305 1336.615 317.475 ;
        RECT 1336.445 220.405 1336.615 220.575 ;
      LAYER met1 ;
        RECT 1332.690 1531.940 1333.010 1532.000 ;
        RECT 1335.450 1531.940 1335.770 1532.000 ;
        RECT 1332.690 1531.800 1335.770 1531.940 ;
        RECT 1332.690 1531.740 1333.010 1531.800 ;
        RECT 1335.450 1531.740 1335.770 1531.800 ;
        RECT 1335.450 1518.000 1335.770 1518.060 ;
        RECT 1335.255 1517.860 1335.770 1518.000 ;
        RECT 1335.450 1517.800 1335.770 1517.860 ;
        RECT 1335.450 1497.260 1335.770 1497.320 ;
        RECT 1335.255 1497.120 1335.770 1497.260 ;
        RECT 1335.450 1497.060 1335.770 1497.120 ;
        RECT 1335.910 1438.780 1336.230 1438.840 ;
        RECT 1335.715 1438.640 1336.230 1438.780 ;
        RECT 1335.910 1438.580 1336.230 1438.640 ;
        RECT 1335.925 1414.640 1336.215 1414.685 ;
        RECT 1336.370 1414.640 1336.690 1414.700 ;
        RECT 1335.925 1414.500 1336.690 1414.640 ;
        RECT 1335.925 1414.455 1336.215 1414.500 ;
        RECT 1336.370 1414.440 1336.690 1414.500 ;
        RECT 1336.370 932.180 1336.690 932.240 ;
        RECT 1335.540 932.040 1336.690 932.180 ;
        RECT 1335.540 931.900 1335.680 932.040 ;
        RECT 1336.370 931.980 1336.690 932.040 ;
        RECT 1335.450 931.640 1335.770 931.900 ;
        RECT 1336.370 896.820 1336.690 896.880 ;
        RECT 1336.175 896.680 1336.690 896.820 ;
        RECT 1336.370 896.620 1336.690 896.680 ;
        RECT 1336.370 848.880 1336.690 848.940 ;
        RECT 1336.175 848.740 1336.690 848.880 ;
        RECT 1336.370 848.680 1336.690 848.740 ;
        RECT 1336.370 800.260 1336.690 800.320 ;
        RECT 1336.175 800.120 1336.690 800.260 ;
        RECT 1336.370 800.060 1336.690 800.120 ;
        RECT 1336.370 752.320 1336.690 752.380 ;
        RECT 1336.175 752.180 1336.690 752.320 ;
        RECT 1336.370 752.120 1336.690 752.180 ;
        RECT 1336.370 703.700 1336.690 703.760 ;
        RECT 1336.175 703.560 1336.690 703.700 ;
        RECT 1336.370 703.500 1336.690 703.560 ;
        RECT 1336.370 655.760 1336.690 655.820 ;
        RECT 1336.175 655.620 1336.690 655.760 ;
        RECT 1336.370 655.560 1336.690 655.620 ;
        RECT 1336.370 607.140 1336.690 607.200 ;
        RECT 1336.845 607.140 1337.135 607.185 ;
        RECT 1336.370 607.000 1337.135 607.140 ;
        RECT 1336.370 606.940 1336.690 607.000 ;
        RECT 1336.845 606.955 1337.135 607.000 ;
        RECT 1336.370 559.200 1336.690 559.260 ;
        RECT 1336.845 559.200 1337.135 559.245 ;
        RECT 1336.370 559.060 1337.135 559.200 ;
        RECT 1336.370 559.000 1336.690 559.060 ;
        RECT 1336.845 559.015 1337.135 559.060 ;
        RECT 1336.370 510.580 1336.690 510.640 ;
        RECT 1336.175 510.440 1336.690 510.580 ;
        RECT 1336.370 510.380 1336.690 510.440 ;
        RECT 1336.370 462.640 1336.690 462.700 ;
        RECT 1336.175 462.500 1336.690 462.640 ;
        RECT 1336.370 462.440 1336.690 462.500 ;
        RECT 1336.370 414.020 1336.690 414.080 ;
        RECT 1336.175 413.880 1336.690 414.020 ;
        RECT 1336.370 413.820 1336.690 413.880 ;
        RECT 1336.370 366.080 1336.690 366.140 ;
        RECT 1336.175 365.940 1336.690 366.080 ;
        RECT 1336.370 365.880 1336.690 365.940 ;
        RECT 1336.370 317.460 1336.690 317.520 ;
        RECT 1336.175 317.320 1336.690 317.460 ;
        RECT 1336.370 317.260 1336.690 317.320 ;
        RECT 1336.370 269.180 1336.690 269.240 ;
        RECT 1336.175 269.040 1336.690 269.180 ;
        RECT 1336.370 268.980 1336.690 269.040 ;
        RECT 1336.370 220.560 1336.690 220.620 ;
        RECT 1336.175 220.420 1336.690 220.560 ;
        RECT 1336.370 220.360 1336.690 220.420 ;
        RECT 1336.385 179.080 1336.675 179.125 ;
        RECT 1336.830 179.080 1337.150 179.140 ;
        RECT 1336.385 178.940 1337.150 179.080 ;
        RECT 1336.385 178.895 1336.675 178.940 ;
        RECT 1336.830 178.880 1337.150 178.940 ;
      LAYER via ;
        RECT 1332.720 1531.740 1332.980 1532.000 ;
        RECT 1335.480 1531.740 1335.740 1532.000 ;
        RECT 1335.480 1517.800 1335.740 1518.060 ;
        RECT 1335.480 1497.060 1335.740 1497.320 ;
        RECT 1335.940 1438.580 1336.200 1438.840 ;
        RECT 1336.400 1414.440 1336.660 1414.700 ;
        RECT 1336.400 931.980 1336.660 932.240 ;
        RECT 1335.480 931.640 1335.740 931.900 ;
        RECT 1336.400 896.620 1336.660 896.880 ;
        RECT 1336.400 848.680 1336.660 848.940 ;
        RECT 1336.400 800.060 1336.660 800.320 ;
        RECT 1336.400 752.120 1336.660 752.380 ;
        RECT 1336.400 703.500 1336.660 703.760 ;
        RECT 1336.400 655.560 1336.660 655.820 ;
        RECT 1336.400 606.940 1336.660 607.200 ;
        RECT 1336.400 559.000 1336.660 559.260 ;
        RECT 1336.400 510.380 1336.660 510.640 ;
        RECT 1336.400 462.440 1336.660 462.700 ;
        RECT 1336.400 413.820 1336.660 414.080 ;
        RECT 1336.400 365.880 1336.660 366.140 ;
        RECT 1336.400 317.260 1336.660 317.520 ;
        RECT 1336.400 268.980 1336.660 269.240 ;
        RECT 1336.400 220.360 1336.660 220.620 ;
        RECT 1336.860 178.880 1337.120 179.140 ;
      LAYER met2 ;
        RECT 1333.960 1600.450 1334.240 1604.000 ;
        RECT 1332.780 1600.310 1334.240 1600.450 ;
        RECT 1332.780 1532.030 1332.920 1600.310 ;
        RECT 1333.960 1600.000 1334.240 1600.310 ;
        RECT 1332.720 1531.710 1332.980 1532.030 ;
        RECT 1335.480 1531.710 1335.740 1532.030 ;
        RECT 1335.540 1518.090 1335.680 1531.710 ;
        RECT 1335.480 1517.770 1335.740 1518.090 ;
        RECT 1335.480 1497.030 1335.740 1497.350 ;
        RECT 1335.540 1469.890 1335.680 1497.030 ;
        RECT 1335.540 1469.750 1336.140 1469.890 ;
        RECT 1336.000 1438.870 1336.140 1469.750 ;
        RECT 1335.940 1438.550 1336.200 1438.870 ;
        RECT 1336.400 1414.410 1336.660 1414.730 ;
        RECT 1336.460 932.270 1336.600 1414.410 ;
        RECT 1336.400 931.950 1336.660 932.270 ;
        RECT 1335.480 931.610 1335.740 931.930 ;
        RECT 1335.540 904.245 1335.680 931.610 ;
        RECT 1335.470 903.875 1335.750 904.245 ;
        RECT 1336.390 903.875 1336.670 904.245 ;
        RECT 1336.460 896.910 1336.600 903.875 ;
        RECT 1336.400 896.590 1336.660 896.910 ;
        RECT 1336.400 848.650 1336.660 848.970 ;
        RECT 1336.460 800.350 1336.600 848.650 ;
        RECT 1336.400 800.030 1336.660 800.350 ;
        RECT 1336.400 752.090 1336.660 752.410 ;
        RECT 1336.460 703.790 1336.600 752.090 ;
        RECT 1336.400 703.470 1336.660 703.790 ;
        RECT 1336.400 655.530 1336.660 655.850 ;
        RECT 1336.460 607.230 1336.600 655.530 ;
        RECT 1336.400 606.910 1336.660 607.230 ;
        RECT 1336.400 558.970 1336.660 559.290 ;
        RECT 1336.460 510.670 1336.600 558.970 ;
        RECT 1336.400 510.350 1336.660 510.670 ;
        RECT 1336.400 462.410 1336.660 462.730 ;
        RECT 1336.460 414.110 1336.600 462.410 ;
        RECT 1336.400 413.790 1336.660 414.110 ;
        RECT 1336.400 365.850 1336.660 366.170 ;
        RECT 1336.460 317.550 1336.600 365.850 ;
        RECT 1336.400 317.230 1336.660 317.550 ;
        RECT 1336.400 268.950 1336.660 269.270 ;
        RECT 1336.460 220.650 1336.600 268.950 ;
        RECT 1336.400 220.330 1336.660 220.650 ;
        RECT 1336.860 178.850 1337.120 179.170 ;
        RECT 1336.920 65.125 1337.060 178.850 ;
        RECT 1336.850 64.755 1337.130 65.125 ;
        RECT 2835.990 64.755 2836.270 65.125 ;
        RECT 2836.060 17.410 2836.200 64.755 ;
        RECT 2836.060 17.270 2839.420 17.410 ;
        RECT 2839.280 2.400 2839.420 17.270 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
      LAYER via2 ;
        RECT 1335.470 903.920 1335.750 904.200 ;
        RECT 1336.390 903.920 1336.670 904.200 ;
        RECT 1336.850 64.800 1337.130 65.080 ;
        RECT 2835.990 64.800 2836.270 65.080 ;
      LAYER met3 ;
        RECT 1335.445 904.210 1335.775 904.225 ;
        RECT 1336.365 904.210 1336.695 904.225 ;
        RECT 1335.445 903.910 1336.695 904.210 ;
        RECT 1335.445 903.895 1335.775 903.910 ;
        RECT 1336.365 903.895 1336.695 903.910 ;
        RECT 1336.825 65.090 1337.155 65.105 ;
        RECT 2835.965 65.090 2836.295 65.105 ;
        RECT 1336.825 64.790 2836.295 65.090 ;
        RECT 1336.825 64.775 1337.155 64.790 ;
        RECT 2835.965 64.775 2836.295 64.790 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1343.345 1338.665 1343.515 1366.375 ;
        RECT 1343.345 565.845 1343.515 613.955 ;
        RECT 1342.885 469.285 1343.055 517.395 ;
      LAYER mcon ;
        RECT 1343.345 1366.205 1343.515 1366.375 ;
        RECT 1343.345 613.785 1343.515 613.955 ;
        RECT 1342.885 517.225 1343.055 517.395 ;
      LAYER met1 ;
        RECT 1339.130 1573.420 1339.450 1573.480 ;
        RECT 1340.510 1573.420 1340.830 1573.480 ;
        RECT 1339.130 1573.280 1340.830 1573.420 ;
        RECT 1339.130 1573.220 1339.450 1573.280 ;
        RECT 1340.510 1573.220 1340.830 1573.280 ;
        RECT 1339.130 1497.600 1339.450 1497.660 ;
        RECT 1343.730 1497.600 1344.050 1497.660 ;
        RECT 1339.130 1497.460 1344.050 1497.600 ;
        RECT 1339.130 1497.400 1339.450 1497.460 ;
        RECT 1343.730 1497.400 1344.050 1497.460 ;
        RECT 1343.270 1366.360 1343.590 1366.420 ;
        RECT 1343.075 1366.220 1343.590 1366.360 ;
        RECT 1343.270 1366.160 1343.590 1366.220 ;
        RECT 1343.270 1338.820 1343.590 1338.880 ;
        RECT 1343.075 1338.680 1343.590 1338.820 ;
        RECT 1343.270 1338.620 1343.590 1338.680 ;
        RECT 1343.270 1221.520 1343.590 1221.580 ;
        RECT 1344.190 1221.520 1344.510 1221.580 ;
        RECT 1343.270 1221.380 1344.510 1221.520 ;
        RECT 1343.270 1221.320 1343.590 1221.380 ;
        RECT 1344.190 1221.320 1344.510 1221.380 ;
        RECT 1343.270 1124.960 1343.590 1125.020 ;
        RECT 1344.190 1124.960 1344.510 1125.020 ;
        RECT 1343.270 1124.820 1344.510 1124.960 ;
        RECT 1343.270 1124.760 1343.590 1124.820 ;
        RECT 1344.190 1124.760 1344.510 1124.820 ;
        RECT 1343.270 1028.400 1343.590 1028.460 ;
        RECT 1344.190 1028.400 1344.510 1028.460 ;
        RECT 1343.270 1028.260 1344.510 1028.400 ;
        RECT 1343.270 1028.200 1343.590 1028.260 ;
        RECT 1344.190 1028.200 1344.510 1028.260 ;
        RECT 1343.270 931.840 1343.590 931.900 ;
        RECT 1344.190 931.840 1344.510 931.900 ;
        RECT 1343.270 931.700 1344.510 931.840 ;
        RECT 1343.270 931.640 1343.590 931.700 ;
        RECT 1344.190 931.640 1344.510 931.700 ;
        RECT 1343.270 738.380 1343.590 738.440 ;
        RECT 1344.190 738.380 1344.510 738.440 ;
        RECT 1343.270 738.240 1344.510 738.380 ;
        RECT 1343.270 738.180 1343.590 738.240 ;
        RECT 1344.190 738.180 1344.510 738.240 ;
        RECT 1343.270 641.820 1343.590 641.880 ;
        RECT 1344.190 641.820 1344.510 641.880 ;
        RECT 1343.270 641.680 1344.510 641.820 ;
        RECT 1343.270 641.620 1343.590 641.680 ;
        RECT 1344.190 641.620 1344.510 641.680 ;
        RECT 1343.270 613.940 1343.590 614.000 ;
        RECT 1343.075 613.800 1343.590 613.940 ;
        RECT 1343.270 613.740 1343.590 613.800 ;
        RECT 1343.285 566.000 1343.575 566.045 ;
        RECT 1344.190 566.000 1344.510 566.060 ;
        RECT 1343.285 565.860 1344.510 566.000 ;
        RECT 1343.285 565.815 1343.575 565.860 ;
        RECT 1344.190 565.800 1344.510 565.860 ;
        RECT 1343.270 545.260 1343.590 545.320 ;
        RECT 1344.190 545.260 1344.510 545.320 ;
        RECT 1343.270 545.120 1344.510 545.260 ;
        RECT 1343.270 545.060 1343.590 545.120 ;
        RECT 1344.190 545.060 1344.510 545.120 ;
        RECT 1342.825 517.380 1343.115 517.425 ;
        RECT 1343.270 517.380 1343.590 517.440 ;
        RECT 1342.825 517.240 1343.590 517.380 ;
        RECT 1342.825 517.195 1343.115 517.240 ;
        RECT 1343.270 517.180 1343.590 517.240 ;
        RECT 1342.810 469.440 1343.130 469.500 ;
        RECT 1342.615 469.300 1343.130 469.440 ;
        RECT 1342.810 469.240 1343.130 469.300 ;
        RECT 1343.270 352.140 1343.590 352.200 ;
        RECT 1344.190 352.140 1344.510 352.200 ;
        RECT 1343.270 352.000 1344.510 352.140 ;
        RECT 1343.270 351.940 1343.590 352.000 ;
        RECT 1344.190 351.940 1344.510 352.000 ;
      LAYER via ;
        RECT 1339.160 1573.220 1339.420 1573.480 ;
        RECT 1340.540 1573.220 1340.800 1573.480 ;
        RECT 1339.160 1497.400 1339.420 1497.660 ;
        RECT 1343.760 1497.400 1344.020 1497.660 ;
        RECT 1343.300 1366.160 1343.560 1366.420 ;
        RECT 1343.300 1338.620 1343.560 1338.880 ;
        RECT 1343.300 1221.320 1343.560 1221.580 ;
        RECT 1344.220 1221.320 1344.480 1221.580 ;
        RECT 1343.300 1124.760 1343.560 1125.020 ;
        RECT 1344.220 1124.760 1344.480 1125.020 ;
        RECT 1343.300 1028.200 1343.560 1028.460 ;
        RECT 1344.220 1028.200 1344.480 1028.460 ;
        RECT 1343.300 931.640 1343.560 931.900 ;
        RECT 1344.220 931.640 1344.480 931.900 ;
        RECT 1343.300 738.180 1343.560 738.440 ;
        RECT 1344.220 738.180 1344.480 738.440 ;
        RECT 1343.300 641.620 1343.560 641.880 ;
        RECT 1344.220 641.620 1344.480 641.880 ;
        RECT 1343.300 613.740 1343.560 614.000 ;
        RECT 1344.220 565.800 1344.480 566.060 ;
        RECT 1343.300 545.060 1343.560 545.320 ;
        RECT 1344.220 545.060 1344.480 545.320 ;
        RECT 1343.300 517.180 1343.560 517.440 ;
        RECT 1342.840 469.240 1343.100 469.500 ;
        RECT 1343.300 351.940 1343.560 352.200 ;
        RECT 1344.220 351.940 1344.480 352.200 ;
      LAYER met2 ;
        RECT 1340.400 1600.380 1340.680 1604.000 ;
        RECT 1340.400 1600.000 1340.740 1600.380 ;
        RECT 1340.600 1573.510 1340.740 1600.000 ;
        RECT 1339.160 1573.190 1339.420 1573.510 ;
        RECT 1340.540 1573.190 1340.800 1573.510 ;
        RECT 1339.220 1497.690 1339.360 1573.190 ;
        RECT 1339.160 1497.370 1339.420 1497.690 ;
        RECT 1343.760 1497.370 1344.020 1497.690 ;
        RECT 1343.820 1386.930 1343.960 1497.370 ;
        RECT 1343.360 1386.790 1343.960 1386.930 ;
        RECT 1343.360 1366.450 1343.500 1386.790 ;
        RECT 1343.300 1366.130 1343.560 1366.450 ;
        RECT 1343.300 1338.590 1343.560 1338.910 ;
        RECT 1343.360 1292.410 1343.500 1338.590 ;
        RECT 1343.360 1292.270 1344.420 1292.410 ;
        RECT 1344.280 1221.610 1344.420 1292.270 ;
        RECT 1343.300 1221.290 1343.560 1221.610 ;
        RECT 1344.220 1221.290 1344.480 1221.610 ;
        RECT 1343.360 1195.850 1343.500 1221.290 ;
        RECT 1343.360 1195.710 1344.420 1195.850 ;
        RECT 1344.280 1125.050 1344.420 1195.710 ;
        RECT 1343.300 1124.730 1343.560 1125.050 ;
        RECT 1344.220 1124.730 1344.480 1125.050 ;
        RECT 1343.360 1099.970 1343.500 1124.730 ;
        RECT 1343.360 1099.830 1344.420 1099.970 ;
        RECT 1344.280 1028.490 1344.420 1099.830 ;
        RECT 1343.300 1028.170 1343.560 1028.490 ;
        RECT 1344.220 1028.170 1344.480 1028.490 ;
        RECT 1343.360 1003.410 1343.500 1028.170 ;
        RECT 1343.360 1003.270 1344.420 1003.410 ;
        RECT 1344.280 931.930 1344.420 1003.270 ;
        RECT 1343.300 931.610 1343.560 931.930 ;
        RECT 1344.220 931.610 1344.480 931.930 ;
        RECT 1343.360 883.730 1343.500 931.610 ;
        RECT 1343.360 883.590 1343.960 883.730 ;
        RECT 1343.820 883.050 1343.960 883.590 ;
        RECT 1342.900 882.910 1343.960 883.050 ;
        RECT 1342.900 810.970 1343.040 882.910 ;
        RECT 1342.900 810.830 1344.420 810.970 ;
        RECT 1344.280 738.470 1344.420 810.830 ;
        RECT 1343.300 738.150 1343.560 738.470 ;
        RECT 1344.220 738.150 1344.480 738.470 ;
        RECT 1343.360 693.330 1343.500 738.150 ;
        RECT 1343.360 693.190 1343.960 693.330 ;
        RECT 1343.820 689.930 1343.960 693.190 ;
        RECT 1343.820 689.790 1344.420 689.930 ;
        RECT 1344.280 641.910 1344.420 689.790 ;
        RECT 1343.300 641.590 1343.560 641.910 ;
        RECT 1344.220 641.590 1344.480 641.910 ;
        RECT 1343.360 614.030 1343.500 641.590 ;
        RECT 1343.300 613.710 1343.560 614.030 ;
        RECT 1344.220 565.770 1344.480 566.090 ;
        RECT 1344.280 545.350 1344.420 565.770 ;
        RECT 1343.300 545.030 1343.560 545.350 ;
        RECT 1344.220 545.030 1344.480 545.350 ;
        RECT 1343.360 517.470 1343.500 545.030 ;
        RECT 1343.300 517.150 1343.560 517.470 ;
        RECT 1342.840 469.210 1343.100 469.530 ;
        RECT 1342.900 424.050 1343.040 469.210 ;
        RECT 1342.900 423.910 1344.420 424.050 ;
        RECT 1344.280 352.230 1344.420 423.910 ;
        RECT 1343.300 351.910 1343.560 352.230 ;
        RECT 1344.220 351.910 1344.480 352.230 ;
        RECT 1343.360 283.120 1343.500 351.910 ;
        RECT 1342.900 282.980 1343.500 283.120 ;
        RECT 1342.900 133.690 1343.040 282.980 ;
        RECT 1342.900 133.550 1344.420 133.690 ;
        RECT 1344.280 75.325 1344.420 133.550 ;
        RECT 1344.210 74.955 1344.490 75.325 ;
        RECT 2856.690 74.955 2856.970 75.325 ;
        RECT 2856.760 17.410 2856.900 74.955 ;
        RECT 2856.760 17.270 2857.360 17.410 ;
        RECT 2857.220 2.400 2857.360 17.270 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
      LAYER via2 ;
        RECT 1344.210 75.000 1344.490 75.280 ;
        RECT 2856.690 75.000 2856.970 75.280 ;
      LAYER met3 ;
        RECT 1344.185 75.290 1344.515 75.305 ;
        RECT 2856.665 75.290 2856.995 75.305 ;
        RECT 1344.185 74.990 2856.995 75.290 ;
        RECT 1344.185 74.975 1344.515 74.990 ;
        RECT 2856.665 74.975 2856.995 74.990 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.030 1594.160 1346.350 1594.220 ;
        RECT 1346.950 1594.160 1347.270 1594.220 ;
        RECT 1346.030 1594.020 1347.270 1594.160 ;
        RECT 1346.030 1593.960 1346.350 1594.020 ;
        RECT 1346.950 1593.960 1347.270 1594.020 ;
      LAYER via ;
        RECT 1346.060 1593.960 1346.320 1594.220 ;
        RECT 1346.980 1593.960 1347.240 1594.220 ;
      LAYER met2 ;
        RECT 1346.380 1600.450 1346.660 1604.000 ;
        RECT 1346.380 1600.310 1347.180 1600.450 ;
        RECT 1346.380 1600.000 1346.660 1600.310 ;
        RECT 1347.040 1594.250 1347.180 1600.310 ;
        RECT 1346.060 1593.930 1346.320 1594.250 ;
        RECT 1346.980 1593.930 1347.240 1594.250 ;
        RECT 1346.120 1558.970 1346.260 1593.930 ;
        RECT 1346.120 1558.830 1351.780 1558.970 ;
        RECT 1351.640 74.645 1351.780 1558.830 ;
        RECT 1351.570 74.275 1351.850 74.645 ;
        RECT 2870.490 74.275 2870.770 74.645 ;
        RECT 2870.560 17.410 2870.700 74.275 ;
        RECT 2870.560 17.270 2875.300 17.410 ;
        RECT 2875.160 2.400 2875.300 17.270 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
      LAYER via2 ;
        RECT 1351.570 74.320 1351.850 74.600 ;
        RECT 2870.490 74.320 2870.770 74.600 ;
      LAYER met3 ;
        RECT 1351.545 74.610 1351.875 74.625 ;
        RECT 2870.465 74.610 2870.795 74.625 ;
        RECT 1351.545 74.310 2870.795 74.610 ;
        RECT 1351.545 74.295 1351.875 74.310 ;
        RECT 2870.465 74.295 2870.795 74.310 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1357.605 1467.525 1357.775 1497.275 ;
      LAYER mcon ;
        RECT 1357.605 1497.105 1357.775 1497.275 ;
      LAYER met1 ;
        RECT 1353.850 1545.880 1354.170 1545.940 ;
        RECT 1357.530 1545.880 1357.850 1545.940 ;
        RECT 1353.850 1545.740 1357.850 1545.880 ;
        RECT 1353.850 1545.680 1354.170 1545.740 ;
        RECT 1357.530 1545.680 1357.850 1545.740 ;
        RECT 1357.530 1497.260 1357.850 1497.320 ;
        RECT 1357.335 1497.120 1357.850 1497.260 ;
        RECT 1357.530 1497.060 1357.850 1497.120 ;
        RECT 1357.530 1467.680 1357.850 1467.740 ;
        RECT 1357.335 1467.540 1357.850 1467.680 ;
        RECT 1357.530 1467.480 1357.850 1467.540 ;
      LAYER via ;
        RECT 1353.880 1545.680 1354.140 1545.940 ;
        RECT 1357.560 1545.680 1357.820 1545.940 ;
        RECT 1357.560 1497.060 1357.820 1497.320 ;
        RECT 1357.560 1467.480 1357.820 1467.740 ;
      LAYER met2 ;
        RECT 1352.820 1600.450 1353.100 1604.000 ;
        RECT 1352.820 1600.310 1354.080 1600.450 ;
        RECT 1352.820 1600.000 1353.100 1600.310 ;
        RECT 1353.940 1545.970 1354.080 1600.310 ;
        RECT 1353.880 1545.650 1354.140 1545.970 ;
        RECT 1357.560 1545.650 1357.820 1545.970 ;
        RECT 1357.620 1497.350 1357.760 1545.650 ;
        RECT 1357.560 1497.030 1357.820 1497.350 ;
        RECT 1357.560 1467.450 1357.820 1467.770 ;
        RECT 1357.620 73.285 1357.760 1467.450 ;
        RECT 1357.550 72.915 1357.830 73.285 ;
        RECT 2891.190 72.915 2891.470 73.285 ;
        RECT 2891.260 3.130 2891.400 72.915 ;
        RECT 2891.260 2.990 2893.240 3.130 ;
        RECT 2893.100 2.400 2893.240 2.990 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
      LAYER via2 ;
        RECT 1357.550 72.960 1357.830 73.240 ;
        RECT 2891.190 72.960 2891.470 73.240 ;
      LAYER met3 ;
        RECT 1357.525 73.250 1357.855 73.265 ;
        RECT 2891.165 73.250 2891.495 73.265 ;
        RECT 1357.525 72.950 2891.495 73.250 ;
        RECT 1357.525 72.935 1357.855 72.950 ;
        RECT 2891.165 72.935 2891.495 72.950 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1358.450 1597.220 1358.770 1597.280 ;
        RECT 1359.370 1597.220 1359.690 1597.280 ;
        RECT 1358.450 1597.080 1359.690 1597.220 ;
        RECT 1358.450 1597.020 1358.770 1597.080 ;
        RECT 1359.370 1597.020 1359.690 1597.080 ;
        RECT 1352.470 1580.220 1352.790 1580.280 ;
        RECT 1358.450 1580.220 1358.770 1580.280 ;
        RECT 1352.470 1580.080 1358.770 1580.220 ;
        RECT 1352.470 1580.020 1352.790 1580.080 ;
        RECT 1358.450 1580.020 1358.770 1580.080 ;
        RECT 1352.470 1535.340 1352.790 1535.400 ;
        RECT 1357.990 1535.340 1358.310 1535.400 ;
        RECT 1352.470 1535.200 1358.310 1535.340 ;
        RECT 1352.470 1535.140 1352.790 1535.200 ;
        RECT 1357.990 1535.140 1358.310 1535.200 ;
        RECT 2904.970 17.580 2905.290 17.640 ;
        RECT 2910.950 17.580 2911.270 17.640 ;
        RECT 2904.970 17.440 2911.270 17.580 ;
        RECT 2904.970 17.380 2905.290 17.440 ;
        RECT 2910.950 17.380 2911.270 17.440 ;
      LAYER via ;
        RECT 1358.480 1597.020 1358.740 1597.280 ;
        RECT 1359.400 1597.020 1359.660 1597.280 ;
        RECT 1352.500 1580.020 1352.760 1580.280 ;
        RECT 1358.480 1580.020 1358.740 1580.280 ;
        RECT 1352.500 1535.140 1352.760 1535.400 ;
        RECT 1358.020 1535.140 1358.280 1535.400 ;
        RECT 2905.000 17.380 2905.260 17.640 ;
        RECT 2910.980 17.380 2911.240 17.640 ;
      LAYER met2 ;
        RECT 1358.800 1600.450 1359.080 1604.000 ;
        RECT 1358.800 1600.310 1359.600 1600.450 ;
        RECT 1358.800 1600.000 1359.080 1600.310 ;
        RECT 1359.460 1597.310 1359.600 1600.310 ;
        RECT 1358.480 1596.990 1358.740 1597.310 ;
        RECT 1359.400 1596.990 1359.660 1597.310 ;
        RECT 1358.540 1580.310 1358.680 1596.990 ;
        RECT 1352.500 1579.990 1352.760 1580.310 ;
        RECT 1358.480 1579.990 1358.740 1580.310 ;
        RECT 1352.560 1535.430 1352.700 1579.990 ;
        RECT 1352.500 1535.110 1352.760 1535.430 ;
        RECT 1358.020 1535.110 1358.280 1535.430 ;
        RECT 1358.080 72.605 1358.220 1535.110 ;
        RECT 1358.010 72.235 1358.290 72.605 ;
        RECT 2904.990 72.235 2905.270 72.605 ;
        RECT 2905.060 17.670 2905.200 72.235 ;
        RECT 2905.000 17.350 2905.260 17.670 ;
        RECT 2910.980 17.350 2911.240 17.670 ;
        RECT 2911.040 2.400 2911.180 17.350 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 1358.010 72.280 1358.290 72.560 ;
        RECT 2904.990 72.280 2905.270 72.560 ;
      LAYER met3 ;
        RECT 1357.985 72.570 1358.315 72.585 ;
        RECT 2904.965 72.570 2905.295 72.585 ;
        RECT 1357.985 72.270 2905.295 72.570 ;
        RECT 1357.985 72.255 1358.315 72.270 ;
        RECT 2904.965 72.255 2905.295 72.270 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 647.640 1600.380 647.920 1604.000 ;
        RECT 647.640 1600.000 647.980 1600.380 ;
        RECT 647.840 20.245 647.980 1600.000 ;
        RECT 647.770 19.875 648.050 20.245 ;
        RECT 858.910 19.875 859.190 20.245 ;
        RECT 858.980 2.400 859.120 19.875 ;
        RECT 858.770 -4.800 859.330 2.400 ;
      LAYER via2 ;
        RECT 647.770 19.920 648.050 20.200 ;
        RECT 858.910 19.920 859.190 20.200 ;
      LAYER met3 ;
        RECT 647.745 20.210 648.075 20.225 ;
        RECT 858.885 20.210 859.215 20.225 ;
        RECT 647.745 19.910 859.215 20.210 ;
        RECT 647.745 19.895 648.075 19.910 ;
        RECT 858.885 19.895 859.215 19.910 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 653.620 1600.450 653.900 1604.000 ;
        RECT 653.620 1600.310 654.880 1600.450 ;
        RECT 653.620 1600.000 653.900 1600.310 ;
        RECT 654.740 19.565 654.880 1600.310 ;
        RECT 654.670 19.195 654.950 19.565 ;
        RECT 876.850 19.195 877.130 19.565 ;
        RECT 876.920 2.400 877.060 19.195 ;
        RECT 876.710 -4.800 877.270 2.400 ;
      LAYER via2 ;
        RECT 654.670 19.240 654.950 19.520 ;
        RECT 876.850 19.240 877.130 19.520 ;
      LAYER met3 ;
        RECT 654.645 19.530 654.975 19.545 ;
        RECT 876.825 19.530 877.155 19.545 ;
        RECT 654.645 19.230 877.155 19.530 ;
        RECT 654.645 19.215 654.975 19.230 ;
        RECT 876.825 19.215 877.155 19.230 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 660.060 1600.450 660.340 1604.000 ;
        RECT 660.060 1600.310 661.320 1600.450 ;
        RECT 660.060 1600.000 660.340 1600.310 ;
        RECT 661.180 1590.250 661.320 1600.310 ;
        RECT 661.180 1590.110 661.780 1590.250 ;
        RECT 661.640 18.885 661.780 1590.110 ;
        RECT 661.570 18.515 661.850 18.885 ;
        RECT 894.790 18.515 895.070 18.885 ;
        RECT 894.860 2.400 895.000 18.515 ;
        RECT 894.650 -4.800 895.210 2.400 ;
      LAYER via2 ;
        RECT 661.570 18.560 661.850 18.840 ;
        RECT 894.790 18.560 895.070 18.840 ;
      LAYER met3 ;
        RECT 661.545 18.850 661.875 18.865 ;
        RECT 894.765 18.850 895.095 18.865 ;
        RECT 661.545 18.550 895.095 18.850 ;
        RECT 661.545 18.535 661.875 18.550 ;
        RECT 894.765 18.535 895.095 18.550 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 812.045 16.065 812.215 17.935 ;
      LAYER mcon ;
        RECT 812.045 17.765 812.215 17.935 ;
      LAYER met1 ;
        RECT 667.530 1592.460 667.850 1592.520 ;
        RECT 789.890 1592.460 790.210 1592.520 ;
        RECT 667.530 1592.320 790.210 1592.460 ;
        RECT 667.530 1592.260 667.850 1592.320 ;
        RECT 789.890 1592.260 790.210 1592.320 ;
        RECT 811.985 17.920 812.275 17.965 ;
        RECT 823.930 17.920 824.250 17.980 ;
        RECT 811.985 17.780 824.250 17.920 ;
        RECT 811.985 17.735 812.275 17.780 ;
        RECT 823.930 17.720 824.250 17.780 ;
        RECT 824.390 16.900 824.710 16.960 ;
        RECT 912.710 16.900 913.030 16.960 ;
        RECT 824.390 16.760 913.030 16.900 ;
        RECT 824.390 16.700 824.710 16.760 ;
        RECT 912.710 16.700 913.030 16.760 ;
        RECT 789.890 16.560 790.210 16.620 ;
        RECT 789.890 16.420 794.260 16.560 ;
        RECT 789.890 16.360 790.210 16.420 ;
        RECT 794.120 16.220 794.260 16.420 ;
        RECT 811.985 16.220 812.275 16.265 ;
        RECT 794.120 16.080 812.275 16.220 ;
        RECT 811.985 16.035 812.275 16.080 ;
      LAYER via ;
        RECT 667.560 1592.260 667.820 1592.520 ;
        RECT 789.920 1592.260 790.180 1592.520 ;
        RECT 823.960 17.720 824.220 17.980 ;
        RECT 824.420 16.700 824.680 16.960 ;
        RECT 912.740 16.700 913.000 16.960 ;
        RECT 789.920 16.360 790.180 16.620 ;
      LAYER met2 ;
        RECT 666.040 1600.450 666.320 1604.000 ;
        RECT 666.040 1600.310 667.760 1600.450 ;
        RECT 666.040 1600.000 666.320 1600.310 ;
        RECT 667.620 1592.550 667.760 1600.310 ;
        RECT 667.560 1592.230 667.820 1592.550 ;
        RECT 789.920 1592.230 790.180 1592.550 ;
        RECT 789.980 16.650 790.120 1592.230 ;
        RECT 823.960 17.690 824.220 18.010 ;
        RECT 824.020 17.410 824.160 17.690 ;
        RECT 824.020 17.270 824.620 17.410 ;
        RECT 824.480 16.990 824.620 17.270 ;
        RECT 824.420 16.670 824.680 16.990 ;
        RECT 912.740 16.670 913.000 16.990 ;
        RECT 789.920 16.330 790.180 16.650 ;
        RECT 912.800 2.400 912.940 16.670 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 824.005 16.745 824.175 20.315 ;
      LAYER mcon ;
        RECT 824.005 20.145 824.175 20.315 ;
      LAYER met1 ;
        RECT 672.590 1593.140 672.910 1593.200 ;
        RECT 796.790 1593.140 797.110 1593.200 ;
        RECT 672.590 1593.000 797.110 1593.140 ;
        RECT 672.590 1592.940 672.910 1593.000 ;
        RECT 796.790 1592.940 797.110 1593.000 ;
        RECT 823.945 20.300 824.235 20.345 ;
        RECT 930.190 20.300 930.510 20.360 ;
        RECT 823.945 20.160 930.510 20.300 ;
        RECT 823.945 20.115 824.235 20.160 ;
        RECT 930.190 20.100 930.510 20.160 ;
        RECT 796.790 16.900 797.110 16.960 ;
        RECT 823.945 16.900 824.235 16.945 ;
        RECT 796.790 16.760 824.235 16.900 ;
        RECT 796.790 16.700 797.110 16.760 ;
        RECT 823.945 16.715 824.235 16.760 ;
      LAYER via ;
        RECT 672.620 1592.940 672.880 1593.200 ;
        RECT 796.820 1592.940 797.080 1593.200 ;
        RECT 930.220 20.100 930.480 20.360 ;
        RECT 796.820 16.700 797.080 16.960 ;
      LAYER met2 ;
        RECT 672.480 1600.380 672.760 1604.000 ;
        RECT 672.480 1600.000 672.820 1600.380 ;
        RECT 672.680 1593.230 672.820 1600.000 ;
        RECT 672.620 1592.910 672.880 1593.230 ;
        RECT 796.820 1592.910 797.080 1593.230 ;
        RECT 796.880 16.990 797.020 1592.910 ;
        RECT 930.220 20.070 930.480 20.390 ;
        RECT 796.820 16.670 797.080 16.990 ;
        RECT 930.280 2.400 930.420 20.070 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 810.205 15.895 810.375 16.575 ;
        RECT 812.505 15.895 812.675 16.235 ;
        RECT 810.205 15.725 812.675 15.895 ;
        RECT 817.105 14.195 817.275 16.235 ;
        RECT 817.105 14.025 818.655 14.195 ;
      LAYER mcon ;
        RECT 810.205 16.405 810.375 16.575 ;
        RECT 812.505 16.065 812.675 16.235 ;
        RECT 817.105 16.065 817.275 16.235 ;
        RECT 818.485 14.025 818.655 14.195 ;
      LAYER met1 ;
        RECT 678.570 1593.820 678.890 1593.880 ;
        RECT 797.250 1593.820 797.570 1593.880 ;
        RECT 678.570 1593.680 797.570 1593.820 ;
        RECT 678.570 1593.620 678.890 1593.680 ;
        RECT 797.250 1593.620 797.570 1593.680 ;
        RECT 797.250 16.560 797.570 16.620 ;
        RECT 810.145 16.560 810.435 16.605 ;
        RECT 797.250 16.420 810.435 16.560 ;
        RECT 797.250 16.360 797.570 16.420 ;
        RECT 810.145 16.375 810.435 16.420 ;
        RECT 812.445 16.220 812.735 16.265 ;
        RECT 817.045 16.220 817.335 16.265 ;
        RECT 812.445 16.080 817.335 16.220 ;
        RECT 812.445 16.035 812.735 16.080 ;
        RECT 817.045 16.035 817.335 16.080 ;
        RECT 818.425 14.180 818.715 14.225 ;
        RECT 948.130 14.180 948.450 14.240 ;
        RECT 818.425 14.040 948.450 14.180 ;
        RECT 818.425 13.995 818.715 14.040 ;
        RECT 948.130 13.980 948.450 14.040 ;
      LAYER via ;
        RECT 678.600 1593.620 678.860 1593.880 ;
        RECT 797.280 1593.620 797.540 1593.880 ;
        RECT 797.280 16.360 797.540 16.620 ;
        RECT 948.160 13.980 948.420 14.240 ;
      LAYER met2 ;
        RECT 678.460 1600.380 678.740 1604.000 ;
        RECT 678.460 1600.000 678.800 1600.380 ;
        RECT 678.660 1593.910 678.800 1600.000 ;
        RECT 678.600 1593.590 678.860 1593.910 ;
        RECT 797.280 1593.590 797.540 1593.910 ;
        RECT 797.340 16.650 797.480 1593.590 ;
        RECT 797.280 16.330 797.540 16.650 ;
        RECT 948.160 13.950 948.420 14.270 ;
        RECT 948.220 2.400 948.360 13.950 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 744.425 15.045 744.595 17.595 ;
      LAYER mcon ;
        RECT 744.425 17.425 744.595 17.595 ;
      LAYER met1 ;
        RECT 685.010 1590.080 685.330 1590.140 ;
        RECT 689.610 1590.080 689.930 1590.140 ;
        RECT 685.010 1589.940 689.930 1590.080 ;
        RECT 685.010 1589.880 685.330 1589.940 ;
        RECT 689.610 1589.880 689.930 1589.940 ;
        RECT 744.365 17.580 744.655 17.625 ;
        RECT 966.070 17.580 966.390 17.640 ;
        RECT 744.365 17.440 966.390 17.580 ;
        RECT 744.365 17.395 744.655 17.440 ;
        RECT 966.070 17.380 966.390 17.440 ;
        RECT 689.610 15.200 689.930 15.260 ;
        RECT 744.365 15.200 744.655 15.245 ;
        RECT 689.610 15.060 693.060 15.200 ;
        RECT 689.610 15.000 689.930 15.060 ;
        RECT 692.920 14.860 693.060 15.060 ;
        RECT 734.320 15.060 744.655 15.200 ;
        RECT 734.320 14.860 734.460 15.060 ;
        RECT 744.365 15.015 744.655 15.060 ;
        RECT 692.920 14.720 734.460 14.860 ;
      LAYER via ;
        RECT 685.040 1589.880 685.300 1590.140 ;
        RECT 689.640 1589.880 689.900 1590.140 ;
        RECT 966.100 17.380 966.360 17.640 ;
        RECT 689.640 15.000 689.900 15.260 ;
      LAYER met2 ;
        RECT 684.900 1600.380 685.180 1604.000 ;
        RECT 684.900 1600.000 685.240 1600.380 ;
        RECT 685.100 1590.170 685.240 1600.000 ;
        RECT 685.040 1589.850 685.300 1590.170 ;
        RECT 689.640 1589.850 689.900 1590.170 ;
        RECT 689.700 15.290 689.840 1589.850 ;
        RECT 966.100 17.350 966.360 17.670 ;
        RECT 689.640 14.970 689.900 15.290 ;
        RECT 966.160 2.400 966.300 17.350 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 709.465 1586.525 709.635 1588.395 ;
        RECT 728.325 1586.525 728.495 1588.735 ;
        RECT 733.845 1588.565 734.015 1589.755 ;
        RECT 759.145 1588.905 759.315 1589.755 ;
      LAYER mcon ;
        RECT 733.845 1589.585 734.015 1589.755 ;
        RECT 759.145 1589.585 759.315 1589.755 ;
        RECT 728.325 1588.565 728.495 1588.735 ;
        RECT 709.465 1588.225 709.635 1588.395 ;
      LAYER met1 ;
        RECT 733.785 1589.740 734.075 1589.785 ;
        RECT 759.085 1589.740 759.375 1589.785 ;
        RECT 733.785 1589.600 759.375 1589.740 ;
        RECT 733.785 1589.555 734.075 1589.600 ;
        RECT 759.085 1589.555 759.375 1589.600 ;
        RECT 759.085 1589.060 759.375 1589.105 ;
        RECT 803.690 1589.060 804.010 1589.120 ;
        RECT 759.085 1588.920 804.010 1589.060 ;
        RECT 759.085 1588.875 759.375 1588.920 ;
        RECT 803.690 1588.860 804.010 1588.920 ;
        RECT 728.265 1588.720 728.555 1588.765 ;
        RECT 733.785 1588.720 734.075 1588.765 ;
        RECT 728.265 1588.580 734.075 1588.720 ;
        RECT 728.265 1588.535 728.555 1588.580 ;
        RECT 733.785 1588.535 734.075 1588.580 ;
        RECT 690.990 1588.380 691.310 1588.440 ;
        RECT 709.405 1588.380 709.695 1588.425 ;
        RECT 690.990 1588.240 709.695 1588.380 ;
        RECT 690.990 1588.180 691.310 1588.240 ;
        RECT 709.405 1588.195 709.695 1588.240 ;
        RECT 709.405 1586.680 709.695 1586.725 ;
        RECT 728.265 1586.680 728.555 1586.725 ;
        RECT 709.405 1586.540 728.555 1586.680 ;
        RECT 709.405 1586.495 709.695 1586.540 ;
        RECT 728.265 1586.495 728.555 1586.540 ;
        RECT 817.950 14.860 818.270 14.920 ;
        RECT 984.010 14.860 984.330 14.920 ;
        RECT 817.950 14.720 984.330 14.860 ;
        RECT 817.950 14.660 818.270 14.720 ;
        RECT 984.010 14.660 984.330 14.720 ;
        RECT 803.690 14.180 804.010 14.240 ;
        RECT 817.950 14.180 818.270 14.240 ;
        RECT 803.690 14.040 818.270 14.180 ;
        RECT 803.690 13.980 804.010 14.040 ;
        RECT 817.950 13.980 818.270 14.040 ;
      LAYER via ;
        RECT 803.720 1588.860 803.980 1589.120 ;
        RECT 691.020 1588.180 691.280 1588.440 ;
        RECT 817.980 14.660 818.240 14.920 ;
        RECT 984.040 14.660 984.300 14.920 ;
        RECT 803.720 13.980 803.980 14.240 ;
        RECT 817.980 13.980 818.240 14.240 ;
      LAYER met2 ;
        RECT 690.880 1600.380 691.160 1604.000 ;
        RECT 690.880 1600.000 691.220 1600.380 ;
        RECT 691.080 1588.470 691.220 1600.000 ;
        RECT 803.720 1588.830 803.980 1589.150 ;
        RECT 691.020 1588.150 691.280 1588.470 ;
        RECT 803.780 14.270 803.920 1588.830 ;
        RECT 817.980 14.630 818.240 14.950 ;
        RECT 984.040 14.630 984.300 14.950 ;
        RECT 818.040 14.270 818.180 14.630 ;
        RECT 803.720 13.950 803.980 14.270 ;
        RECT 817.980 13.950 818.240 14.270 ;
        RECT 984.100 2.400 984.240 14.630 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 1590.080 579.990 1590.140 ;
        RECT 585.650 1590.080 585.970 1590.140 ;
        RECT 579.670 1589.940 585.970 1590.080 ;
        RECT 579.670 1589.880 579.990 1589.940 ;
        RECT 585.650 1589.880 585.970 1589.940 ;
        RECT 586.110 14.860 586.430 14.920 ;
        RECT 662.930 14.860 663.250 14.920 ;
        RECT 586.110 14.720 663.250 14.860 ;
        RECT 586.110 14.660 586.430 14.720 ;
        RECT 662.930 14.660 663.250 14.720 ;
      LAYER via ;
        RECT 579.700 1589.880 579.960 1590.140 ;
        RECT 585.680 1589.880 585.940 1590.140 ;
        RECT 586.140 14.660 586.400 14.920 ;
        RECT 662.960 14.660 663.220 14.920 ;
      LAYER met2 ;
        RECT 579.560 1600.380 579.840 1604.000 ;
        RECT 579.560 1600.000 579.900 1600.380 ;
        RECT 579.760 1590.170 579.900 1600.000 ;
        RECT 579.700 1589.850 579.960 1590.170 ;
        RECT 585.680 1589.850 585.940 1590.170 ;
        RECT 585.740 24.890 585.880 1589.850 ;
        RECT 585.740 24.750 586.340 24.890 ;
        RECT 586.200 14.950 586.340 24.750 ;
        RECT 586.140 14.630 586.400 14.950 ;
        RECT 662.960 14.630 663.220 14.950 ;
        RECT 663.020 2.400 663.160 14.630 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 696.970 1588.040 697.290 1588.100 ;
        RECT 703.410 1588.040 703.730 1588.100 ;
        RECT 696.970 1587.900 703.730 1588.040 ;
        RECT 696.970 1587.840 697.290 1587.900 ;
        RECT 703.410 1587.840 703.730 1587.900 ;
        RECT 703.410 17.240 703.730 17.300 ;
        RECT 1001.950 17.240 1002.270 17.300 ;
        RECT 703.410 17.100 1002.270 17.240 ;
        RECT 703.410 17.040 703.730 17.100 ;
        RECT 1001.950 17.040 1002.270 17.100 ;
      LAYER via ;
        RECT 697.000 1587.840 697.260 1588.100 ;
        RECT 703.440 1587.840 703.700 1588.100 ;
        RECT 703.440 17.040 703.700 17.300 ;
        RECT 1001.980 17.040 1002.240 17.300 ;
      LAYER met2 ;
        RECT 696.860 1600.380 697.140 1604.000 ;
        RECT 696.860 1600.000 697.200 1600.380 ;
        RECT 697.060 1588.130 697.200 1600.000 ;
        RECT 697.000 1587.810 697.260 1588.130 ;
        RECT 703.440 1587.810 703.700 1588.130 ;
        RECT 703.500 17.330 703.640 1587.810 ;
        RECT 703.440 17.010 703.700 17.330 ;
        RECT 1001.980 17.010 1002.240 17.330 ;
        RECT 1002.040 2.400 1002.180 17.010 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 713.605 1589.585 713.775 1591.455 ;
        RECT 810.665 1545.725 810.835 1590.095 ;
        RECT 810.665 16.405 810.835 33.235 ;
      LAYER mcon ;
        RECT 713.605 1591.285 713.775 1591.455 ;
        RECT 810.665 1589.925 810.835 1590.095 ;
        RECT 810.665 33.065 810.835 33.235 ;
      LAYER met1 ;
        RECT 703.410 1591.440 703.730 1591.500 ;
        RECT 713.545 1591.440 713.835 1591.485 ;
        RECT 703.410 1591.300 713.835 1591.440 ;
        RECT 703.410 1591.240 703.730 1591.300 ;
        RECT 713.545 1591.255 713.835 1591.300 ;
        RECT 810.605 1590.080 810.895 1590.125 ;
        RECT 733.400 1589.940 810.895 1590.080 ;
        RECT 713.545 1589.740 713.835 1589.785 ;
        RECT 733.400 1589.740 733.540 1589.940 ;
        RECT 810.605 1589.895 810.895 1589.940 ;
        RECT 713.545 1589.600 733.540 1589.740 ;
        RECT 713.545 1589.555 713.835 1589.600 ;
        RECT 810.590 1545.880 810.910 1545.940 ;
        RECT 810.395 1545.740 810.910 1545.880 ;
        RECT 810.590 1545.680 810.910 1545.740 ;
        RECT 810.590 48.860 810.910 48.920 ;
        RECT 809.760 48.720 810.910 48.860 ;
        RECT 809.760 48.580 809.900 48.720 ;
        RECT 810.590 48.660 810.910 48.720 ;
        RECT 809.670 48.320 809.990 48.580 ;
        RECT 809.670 33.220 809.990 33.280 ;
        RECT 810.605 33.220 810.895 33.265 ;
        RECT 809.670 33.080 810.895 33.220 ;
        RECT 809.670 33.020 809.990 33.080 ;
        RECT 810.605 33.035 810.895 33.080 ;
        RECT 810.605 16.560 810.895 16.605 ;
        RECT 810.605 16.420 850.380 16.560 ;
        RECT 810.605 16.375 810.895 16.420 ;
        RECT 850.240 15.880 850.380 16.420 ;
        RECT 1019.430 15.880 1019.750 15.940 ;
        RECT 850.240 15.740 1019.750 15.880 ;
        RECT 1019.430 15.680 1019.750 15.740 ;
      LAYER via ;
        RECT 703.440 1591.240 703.700 1591.500 ;
        RECT 810.620 1545.680 810.880 1545.940 ;
        RECT 810.620 48.660 810.880 48.920 ;
        RECT 809.700 48.320 809.960 48.580 ;
        RECT 809.700 33.020 809.960 33.280 ;
        RECT 1019.460 15.680 1019.720 15.940 ;
      LAYER met2 ;
        RECT 703.300 1600.380 703.580 1604.000 ;
        RECT 703.300 1600.000 703.640 1600.380 ;
        RECT 703.500 1591.530 703.640 1600.000 ;
        RECT 703.440 1591.210 703.700 1591.530 ;
        RECT 810.620 1545.650 810.880 1545.970 ;
        RECT 810.680 48.950 810.820 1545.650 ;
        RECT 810.620 48.630 810.880 48.950 ;
        RECT 809.700 48.290 809.960 48.610 ;
        RECT 809.760 33.310 809.900 48.290 ;
        RECT 809.700 32.990 809.960 33.310 ;
        RECT 1019.460 15.650 1019.720 15.970 ;
        RECT 1019.520 2.400 1019.660 15.650 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 714.525 1593.325 714.695 1594.175 ;
        RECT 725.105 1588.225 725.275 1593.495 ;
      LAYER mcon ;
        RECT 714.525 1594.005 714.695 1594.175 ;
        RECT 725.105 1593.325 725.275 1593.495 ;
      LAYER met1 ;
        RECT 710.310 1594.160 710.630 1594.220 ;
        RECT 714.465 1594.160 714.755 1594.205 ;
        RECT 710.310 1594.020 714.755 1594.160 ;
        RECT 710.310 1593.960 710.630 1594.020 ;
        RECT 714.465 1593.975 714.755 1594.020 ;
        RECT 714.465 1593.480 714.755 1593.525 ;
        RECT 725.045 1593.480 725.335 1593.525 ;
        RECT 714.465 1593.340 725.335 1593.480 ;
        RECT 714.465 1593.295 714.755 1593.340 ;
        RECT 725.045 1593.295 725.335 1593.340 ;
        RECT 725.045 1588.380 725.335 1588.425 ;
        RECT 790.350 1588.380 790.670 1588.440 ;
        RECT 725.045 1588.240 790.670 1588.380 ;
        RECT 725.045 1588.195 725.335 1588.240 ;
        RECT 790.350 1588.180 790.670 1588.240 ;
      LAYER via ;
        RECT 710.340 1593.960 710.600 1594.220 ;
        RECT 790.380 1588.180 790.640 1588.440 ;
      LAYER met2 ;
        RECT 709.280 1600.450 709.560 1604.000 ;
        RECT 709.280 1600.310 710.540 1600.450 ;
        RECT 709.280 1600.000 709.560 1600.310 ;
        RECT 710.400 1594.250 710.540 1600.310 ;
        RECT 710.340 1593.930 710.600 1594.250 ;
        RECT 790.380 1588.150 790.640 1588.470 ;
        RECT 790.440 18.205 790.580 1588.150 ;
        RECT 790.370 17.835 790.650 18.205 ;
        RECT 1037.390 17.835 1037.670 18.205 ;
        RECT 1037.460 2.400 1037.600 17.835 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
      LAYER via2 ;
        RECT 790.370 17.880 790.650 18.160 ;
        RECT 1037.390 17.880 1037.670 18.160 ;
      LAYER met3 ;
        RECT 790.345 18.170 790.675 18.185 ;
        RECT 1037.365 18.170 1037.695 18.185 ;
        RECT 790.345 17.870 1037.695 18.170 ;
        RECT 790.345 17.855 790.675 17.870 ;
        RECT 1037.365 17.855 1037.695 17.870 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 845.165 16.065 845.335 17.935 ;
      LAYER mcon ;
        RECT 845.165 17.765 845.335 17.935 ;
      LAYER met1 ;
        RECT 845.105 17.920 845.395 17.965 ;
        RECT 1055.310 17.920 1055.630 17.980 ;
        RECT 845.105 17.780 1055.630 17.920 ;
        RECT 845.105 17.735 845.395 17.780 ;
        RECT 1055.310 17.720 1055.630 17.780 ;
        RECT 817.490 16.220 817.810 16.280 ;
        RECT 845.105 16.220 845.395 16.265 ;
        RECT 817.490 16.080 845.395 16.220 ;
        RECT 817.490 16.020 817.810 16.080 ;
        RECT 845.105 16.035 845.395 16.080 ;
      LAYER via ;
        RECT 1055.340 17.720 1055.600 17.980 ;
        RECT 817.520 16.020 817.780 16.280 ;
      LAYER met2 ;
        RECT 715.720 1600.380 716.000 1604.000 ;
        RECT 715.720 1600.000 716.060 1600.380 ;
        RECT 715.920 1590.365 716.060 1600.000 ;
        RECT 715.850 1589.995 716.130 1590.365 ;
        RECT 817.510 1589.995 817.790 1590.365 ;
        RECT 817.580 16.310 817.720 1589.995 ;
        RECT 1055.340 17.690 1055.600 18.010 ;
        RECT 817.520 15.990 817.780 16.310 ;
        RECT 1055.400 2.400 1055.540 17.690 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
      LAYER via2 ;
        RECT 715.850 1590.040 716.130 1590.320 ;
        RECT 817.510 1590.040 817.790 1590.320 ;
      LAYER met3 ;
        RECT 715.825 1590.330 716.155 1590.345 ;
        RECT 817.485 1590.330 817.815 1590.345 ;
        RECT 715.825 1590.030 817.815 1590.330 ;
        RECT 715.825 1590.015 716.155 1590.030 ;
        RECT 817.485 1590.015 817.815 1590.030 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 721.810 1588.040 722.130 1588.100 ;
        RECT 724.110 1588.040 724.430 1588.100 ;
        RECT 721.810 1587.900 724.430 1588.040 ;
        RECT 721.810 1587.840 722.130 1587.900 ;
        RECT 724.110 1587.840 724.430 1587.900 ;
      LAYER via ;
        RECT 721.840 1587.840 722.100 1588.100 ;
        RECT 724.140 1587.840 724.400 1588.100 ;
      LAYER met2 ;
        RECT 721.700 1600.380 721.980 1604.000 ;
        RECT 721.700 1600.000 722.040 1600.380 ;
        RECT 721.900 1588.130 722.040 1600.000 ;
        RECT 721.840 1587.810 722.100 1588.130 ;
        RECT 724.140 1587.810 724.400 1588.130 ;
        RECT 724.200 16.845 724.340 1587.810 ;
        RECT 724.130 16.475 724.410 16.845 ;
        RECT 1073.270 16.475 1073.550 16.845 ;
        RECT 1073.340 2.400 1073.480 16.475 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
      LAYER via2 ;
        RECT 724.130 16.520 724.410 16.800 ;
        RECT 1073.270 16.520 1073.550 16.800 ;
      LAYER met3 ;
        RECT 724.105 16.810 724.435 16.825 ;
        RECT 1073.245 16.810 1073.575 16.825 ;
        RECT 724.105 16.510 1073.575 16.810 ;
        RECT 724.105 16.495 724.435 16.510 ;
        RECT 1073.245 16.495 1073.575 16.510 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 740.285 1590.945 740.455 1593.495 ;
        RECT 752.245 1590.945 752.415 1592.135 ;
        RECT 770.185 1587.885 770.355 1592.135 ;
      LAYER mcon ;
        RECT 740.285 1593.325 740.455 1593.495 ;
        RECT 752.245 1591.965 752.415 1592.135 ;
        RECT 770.185 1591.965 770.355 1592.135 ;
      LAYER met1 ;
        RECT 728.250 1593.480 728.570 1593.540 ;
        RECT 740.225 1593.480 740.515 1593.525 ;
        RECT 728.250 1593.340 740.515 1593.480 ;
        RECT 728.250 1593.280 728.570 1593.340 ;
        RECT 740.225 1593.295 740.515 1593.340 ;
        RECT 752.185 1592.120 752.475 1592.165 ;
        RECT 770.125 1592.120 770.415 1592.165 ;
        RECT 752.185 1591.980 770.415 1592.120 ;
        RECT 752.185 1591.935 752.475 1591.980 ;
        RECT 770.125 1591.935 770.415 1591.980 ;
        RECT 740.225 1591.100 740.515 1591.145 ;
        RECT 752.185 1591.100 752.475 1591.145 ;
        RECT 740.225 1590.960 752.475 1591.100 ;
        RECT 740.225 1590.915 740.515 1590.960 ;
        RECT 752.185 1590.915 752.475 1590.960 ;
        RECT 770.125 1588.040 770.415 1588.085 ;
        RECT 830.830 1588.040 831.150 1588.100 ;
        RECT 770.125 1587.900 831.150 1588.040 ;
        RECT 770.125 1587.855 770.415 1587.900 ;
        RECT 830.830 1587.840 831.150 1587.900 ;
      LAYER via ;
        RECT 728.280 1593.280 728.540 1593.540 ;
        RECT 830.860 1587.840 831.120 1588.100 ;
      LAYER met2 ;
        RECT 728.140 1600.380 728.420 1604.000 ;
        RECT 728.140 1600.000 728.480 1600.380 ;
        RECT 728.340 1593.570 728.480 1600.000 ;
        RECT 728.280 1593.250 728.540 1593.570 ;
        RECT 830.860 1587.810 831.120 1588.130 ;
        RECT 830.920 1582.090 831.060 1587.810 ;
        RECT 830.920 1581.950 831.520 1582.090 ;
        RECT 831.380 17.525 831.520 1581.950 ;
        RECT 831.310 17.155 831.590 17.525 ;
        RECT 1090.750 17.155 1091.030 17.525 ;
        RECT 1090.820 2.400 1090.960 17.155 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
      LAYER via2 ;
        RECT 831.310 17.200 831.590 17.480 ;
        RECT 1090.750 17.200 1091.030 17.480 ;
      LAYER met3 ;
        RECT 831.285 17.490 831.615 17.505 ;
        RECT 1090.725 17.490 1091.055 17.505 ;
        RECT 831.285 17.190 1091.055 17.490 ;
        RECT 831.285 17.175 831.615 17.190 ;
        RECT 1090.725 17.175 1091.055 17.190 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 762.365 1589.245 762.535 1590.435 ;
        RECT 849.765 16.405 850.855 16.575 ;
        RECT 849.765 15.725 849.935 16.405 ;
      LAYER mcon ;
        RECT 762.365 1590.265 762.535 1590.435 ;
        RECT 850.685 16.405 850.855 16.575 ;
      LAYER met1 ;
        RECT 734.230 1590.420 734.550 1590.480 ;
        RECT 762.305 1590.420 762.595 1590.465 ;
        RECT 734.230 1590.280 762.595 1590.420 ;
        RECT 734.230 1590.220 734.550 1590.280 ;
        RECT 762.305 1590.235 762.595 1590.280 ;
        RECT 762.305 1589.400 762.595 1589.445 ;
        RECT 838.190 1589.400 838.510 1589.460 ;
        RECT 762.305 1589.260 838.510 1589.400 ;
        RECT 762.305 1589.215 762.595 1589.260 ;
        RECT 838.190 1589.200 838.510 1589.260 ;
        RECT 838.190 17.920 838.510 17.980 ;
        RECT 841.410 17.920 841.730 17.980 ;
        RECT 838.190 17.780 841.730 17.920 ;
        RECT 838.190 17.720 838.510 17.780 ;
        RECT 841.410 17.720 841.730 17.780 ;
        RECT 850.625 16.560 850.915 16.605 ;
        RECT 850.625 16.420 859.580 16.560 ;
        RECT 850.625 16.375 850.915 16.420 ;
        RECT 859.440 16.220 859.580 16.420 ;
        RECT 1108.670 16.220 1108.990 16.280 ;
        RECT 859.440 16.080 1108.990 16.220 ;
        RECT 1108.670 16.020 1108.990 16.080 ;
        RECT 841.410 15.880 841.730 15.940 ;
        RECT 849.705 15.880 849.995 15.925 ;
        RECT 841.410 15.740 849.995 15.880 ;
        RECT 841.410 15.680 841.730 15.740 ;
        RECT 849.705 15.695 849.995 15.740 ;
      LAYER via ;
        RECT 734.260 1590.220 734.520 1590.480 ;
        RECT 838.220 1589.200 838.480 1589.460 ;
        RECT 838.220 17.720 838.480 17.980 ;
        RECT 841.440 17.720 841.700 17.980 ;
        RECT 1108.700 16.020 1108.960 16.280 ;
        RECT 841.440 15.680 841.700 15.940 ;
      LAYER met2 ;
        RECT 734.120 1600.380 734.400 1604.000 ;
        RECT 734.120 1600.000 734.460 1600.380 ;
        RECT 734.320 1590.510 734.460 1600.000 ;
        RECT 734.260 1590.190 734.520 1590.510 ;
        RECT 838.220 1589.170 838.480 1589.490 ;
        RECT 838.280 18.010 838.420 1589.170 ;
        RECT 838.220 17.690 838.480 18.010 ;
        RECT 841.440 17.690 841.700 18.010 ;
        RECT 841.500 15.970 841.640 17.690 ;
        RECT 1108.700 15.990 1108.960 16.310 ;
        RECT 841.440 15.650 841.700 15.970 ;
        RECT 1108.760 2.400 1108.900 15.990 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 763.745 1591.285 763.915 1593.495 ;
        RECT 950.505 1588.905 950.675 1591.455 ;
        RECT 969.365 1538.925 969.535 1546.235 ;
        RECT 969.365 1442.025 969.535 1490.475 ;
        RECT 969.365 766.105 969.535 814.215 ;
        RECT 969.365 669.545 969.535 717.655 ;
        RECT 969.365 572.645 969.535 620.755 ;
        RECT 969.365 476.085 969.535 524.195 ;
        RECT 969.365 379.525 969.535 427.635 ;
        RECT 969.365 282.965 969.535 331.075 ;
        RECT 969.365 144.925 969.535 234.515 ;
        RECT 968.905 61.965 969.075 96.475 ;
      LAYER mcon ;
        RECT 763.745 1593.325 763.915 1593.495 ;
        RECT 950.505 1591.285 950.675 1591.455 ;
        RECT 969.365 1546.065 969.535 1546.235 ;
        RECT 969.365 1490.305 969.535 1490.475 ;
        RECT 969.365 814.045 969.535 814.215 ;
        RECT 969.365 717.485 969.535 717.655 ;
        RECT 969.365 620.585 969.535 620.755 ;
        RECT 969.365 524.025 969.535 524.195 ;
        RECT 969.365 427.465 969.535 427.635 ;
        RECT 969.365 330.905 969.535 331.075 ;
        RECT 969.365 234.345 969.535 234.515 ;
        RECT 968.905 96.305 969.075 96.475 ;
      LAYER met1 ;
        RECT 740.670 1593.480 740.990 1593.540 ;
        RECT 763.685 1593.480 763.975 1593.525 ;
        RECT 740.670 1593.340 763.975 1593.480 ;
        RECT 740.670 1593.280 740.990 1593.340 ;
        RECT 763.685 1593.295 763.975 1593.340 ;
        RECT 763.685 1591.440 763.975 1591.485 ;
        RECT 950.445 1591.440 950.735 1591.485 ;
        RECT 763.685 1591.300 950.735 1591.440 ;
        RECT 763.685 1591.255 763.975 1591.300 ;
        RECT 950.445 1591.255 950.735 1591.300 ;
        RECT 950.445 1589.060 950.735 1589.105 ;
        RECT 968.830 1589.060 969.150 1589.120 ;
        RECT 950.445 1588.920 969.150 1589.060 ;
        RECT 950.445 1588.875 950.735 1588.920 ;
        RECT 968.830 1588.860 969.150 1588.920 ;
        RECT 969.305 1546.220 969.595 1546.265 ;
        RECT 969.750 1546.220 970.070 1546.280 ;
        RECT 969.305 1546.080 970.070 1546.220 ;
        RECT 969.305 1546.035 969.595 1546.080 ;
        RECT 969.750 1546.020 970.070 1546.080 ;
        RECT 969.290 1539.080 969.610 1539.140 ;
        RECT 969.095 1538.940 969.610 1539.080 ;
        RECT 969.290 1538.880 969.610 1538.940 ;
        RECT 969.290 1490.460 969.610 1490.520 ;
        RECT 969.095 1490.320 969.610 1490.460 ;
        RECT 969.290 1490.260 969.610 1490.320 ;
        RECT 969.290 1442.180 969.610 1442.240 ;
        RECT 969.095 1442.040 969.610 1442.180 ;
        RECT 969.290 1441.980 969.610 1442.040 ;
        RECT 968.370 1345.620 968.690 1345.680 ;
        RECT 969.290 1345.620 969.610 1345.680 ;
        RECT 968.370 1345.480 969.610 1345.620 ;
        RECT 968.370 1345.420 968.690 1345.480 ;
        RECT 969.290 1345.420 969.610 1345.480 ;
        RECT 968.370 1249.060 968.690 1249.120 ;
        RECT 969.290 1249.060 969.610 1249.120 ;
        RECT 968.370 1248.920 969.610 1249.060 ;
        RECT 968.370 1248.860 968.690 1248.920 ;
        RECT 969.290 1248.860 969.610 1248.920 ;
        RECT 968.370 1152.500 968.690 1152.560 ;
        RECT 969.290 1152.500 969.610 1152.560 ;
        RECT 968.370 1152.360 969.610 1152.500 ;
        RECT 968.370 1152.300 968.690 1152.360 ;
        RECT 969.290 1152.300 969.610 1152.360 ;
        RECT 968.370 1007.320 968.690 1007.380 ;
        RECT 969.290 1007.320 969.610 1007.380 ;
        RECT 968.370 1007.180 969.610 1007.320 ;
        RECT 968.370 1007.120 968.690 1007.180 ;
        RECT 969.290 1007.120 969.610 1007.180 ;
        RECT 968.370 910.760 968.690 910.820 ;
        RECT 969.290 910.760 969.610 910.820 ;
        RECT 968.370 910.620 969.610 910.760 ;
        RECT 968.370 910.560 968.690 910.620 ;
        RECT 969.290 910.560 969.610 910.620 ;
        RECT 969.290 814.200 969.610 814.260 ;
        RECT 969.095 814.060 969.610 814.200 ;
        RECT 969.290 814.000 969.610 814.060 ;
        RECT 969.290 766.260 969.610 766.320 ;
        RECT 969.095 766.120 969.610 766.260 ;
        RECT 969.290 766.060 969.610 766.120 ;
        RECT 969.290 717.640 969.610 717.700 ;
        RECT 969.095 717.500 969.610 717.640 ;
        RECT 969.290 717.440 969.610 717.500 ;
        RECT 969.290 669.700 969.610 669.760 ;
        RECT 969.095 669.560 969.610 669.700 ;
        RECT 969.290 669.500 969.610 669.560 ;
        RECT 969.290 620.740 969.610 620.800 ;
        RECT 969.095 620.600 969.610 620.740 ;
        RECT 969.290 620.540 969.610 620.600 ;
        RECT 969.290 572.800 969.610 572.860 ;
        RECT 969.095 572.660 969.610 572.800 ;
        RECT 969.290 572.600 969.610 572.660 ;
        RECT 969.290 524.180 969.610 524.240 ;
        RECT 969.095 524.040 969.610 524.180 ;
        RECT 969.290 523.980 969.610 524.040 ;
        RECT 969.290 476.240 969.610 476.300 ;
        RECT 969.095 476.100 969.610 476.240 ;
        RECT 969.290 476.040 969.610 476.100 ;
        RECT 969.290 427.620 969.610 427.680 ;
        RECT 969.095 427.480 969.610 427.620 ;
        RECT 969.290 427.420 969.610 427.480 ;
        RECT 969.290 379.680 969.610 379.740 ;
        RECT 969.095 379.540 969.610 379.680 ;
        RECT 969.290 379.480 969.610 379.540 ;
        RECT 969.290 331.060 969.610 331.120 ;
        RECT 969.095 330.920 969.610 331.060 ;
        RECT 969.290 330.860 969.610 330.920 ;
        RECT 969.290 283.120 969.610 283.180 ;
        RECT 969.095 282.980 969.610 283.120 ;
        RECT 969.290 282.920 969.610 282.980 ;
        RECT 969.290 234.500 969.610 234.560 ;
        RECT 969.095 234.360 969.610 234.500 ;
        RECT 969.290 234.300 969.610 234.360 ;
        RECT 969.305 145.080 969.595 145.125 ;
        RECT 969.750 145.080 970.070 145.140 ;
        RECT 969.305 144.940 970.070 145.080 ;
        RECT 969.305 144.895 969.595 144.940 ;
        RECT 969.750 144.880 970.070 144.940 ;
        RECT 968.830 96.460 969.150 96.520 ;
        RECT 968.635 96.320 969.150 96.460 ;
        RECT 968.830 96.260 969.150 96.320 ;
        RECT 968.830 62.120 969.150 62.180 ;
        RECT 968.635 61.980 969.150 62.120 ;
        RECT 968.830 61.920 969.150 61.980 ;
        RECT 969.290 20.980 969.610 21.040 ;
        RECT 1126.610 20.980 1126.930 21.040 ;
        RECT 969.290 20.840 1126.930 20.980 ;
        RECT 969.290 20.780 969.610 20.840 ;
        RECT 1126.610 20.780 1126.930 20.840 ;
      LAYER via ;
        RECT 740.700 1593.280 740.960 1593.540 ;
        RECT 968.860 1588.860 969.120 1589.120 ;
        RECT 969.780 1546.020 970.040 1546.280 ;
        RECT 969.320 1538.880 969.580 1539.140 ;
        RECT 969.320 1490.260 969.580 1490.520 ;
        RECT 969.320 1441.980 969.580 1442.240 ;
        RECT 968.400 1345.420 968.660 1345.680 ;
        RECT 969.320 1345.420 969.580 1345.680 ;
        RECT 968.400 1248.860 968.660 1249.120 ;
        RECT 969.320 1248.860 969.580 1249.120 ;
        RECT 968.400 1152.300 968.660 1152.560 ;
        RECT 969.320 1152.300 969.580 1152.560 ;
        RECT 968.400 1007.120 968.660 1007.380 ;
        RECT 969.320 1007.120 969.580 1007.380 ;
        RECT 968.400 910.560 968.660 910.820 ;
        RECT 969.320 910.560 969.580 910.820 ;
        RECT 969.320 814.000 969.580 814.260 ;
        RECT 969.320 766.060 969.580 766.320 ;
        RECT 969.320 717.440 969.580 717.700 ;
        RECT 969.320 669.500 969.580 669.760 ;
        RECT 969.320 620.540 969.580 620.800 ;
        RECT 969.320 572.600 969.580 572.860 ;
        RECT 969.320 523.980 969.580 524.240 ;
        RECT 969.320 476.040 969.580 476.300 ;
        RECT 969.320 427.420 969.580 427.680 ;
        RECT 969.320 379.480 969.580 379.740 ;
        RECT 969.320 330.860 969.580 331.120 ;
        RECT 969.320 282.920 969.580 283.180 ;
        RECT 969.320 234.300 969.580 234.560 ;
        RECT 969.780 144.880 970.040 145.140 ;
        RECT 968.860 96.260 969.120 96.520 ;
        RECT 968.860 61.920 969.120 62.180 ;
        RECT 969.320 20.780 969.580 21.040 ;
        RECT 1126.640 20.780 1126.900 21.040 ;
      LAYER met2 ;
        RECT 740.560 1600.380 740.840 1604.000 ;
        RECT 740.560 1600.000 740.900 1600.380 ;
        RECT 740.760 1593.570 740.900 1600.000 ;
        RECT 740.700 1593.250 740.960 1593.570 ;
        RECT 968.860 1588.830 969.120 1589.150 ;
        RECT 968.920 1587.530 969.060 1588.830 ;
        RECT 968.920 1587.390 969.980 1587.530 ;
        RECT 969.840 1546.310 969.980 1587.390 ;
        RECT 969.780 1545.990 970.040 1546.310 ;
        RECT 969.320 1538.850 969.580 1539.170 ;
        RECT 969.380 1490.550 969.520 1538.850 ;
        RECT 969.320 1490.230 969.580 1490.550 ;
        RECT 969.320 1441.950 969.580 1442.270 ;
        RECT 969.380 1393.845 969.520 1441.950 ;
        RECT 968.390 1393.475 968.670 1393.845 ;
        RECT 969.310 1393.475 969.590 1393.845 ;
        RECT 968.460 1345.710 968.600 1393.475 ;
        RECT 968.400 1345.390 968.660 1345.710 ;
        RECT 969.320 1345.390 969.580 1345.710 ;
        RECT 969.380 1297.285 969.520 1345.390 ;
        RECT 968.390 1296.915 968.670 1297.285 ;
        RECT 969.310 1296.915 969.590 1297.285 ;
        RECT 968.460 1249.150 968.600 1296.915 ;
        RECT 968.400 1248.830 968.660 1249.150 ;
        RECT 969.320 1248.830 969.580 1249.150 ;
        RECT 969.380 1208.885 969.520 1248.830 ;
        RECT 969.310 1208.515 969.590 1208.885 ;
        RECT 969.310 1207.835 969.590 1208.205 ;
        RECT 969.380 1200.725 969.520 1207.835 ;
        RECT 968.390 1200.355 968.670 1200.725 ;
        RECT 969.310 1200.355 969.590 1200.725 ;
        RECT 968.460 1152.590 968.600 1200.355 ;
        RECT 968.400 1152.270 968.660 1152.590 ;
        RECT 969.320 1152.270 969.580 1152.590 ;
        RECT 969.380 1104.165 969.520 1152.270 ;
        RECT 968.390 1103.795 968.670 1104.165 ;
        RECT 969.310 1103.795 969.590 1104.165 ;
        RECT 968.460 1055.885 968.600 1103.795 ;
        RECT 968.390 1055.515 968.670 1055.885 ;
        RECT 969.310 1055.515 969.590 1055.885 ;
        RECT 969.380 1007.410 969.520 1055.515 ;
        RECT 968.400 1007.090 968.660 1007.410 ;
        RECT 969.320 1007.090 969.580 1007.410 ;
        RECT 968.460 959.325 968.600 1007.090 ;
        RECT 968.390 958.955 968.670 959.325 ;
        RECT 969.310 958.955 969.590 959.325 ;
        RECT 969.380 910.850 969.520 958.955 ;
        RECT 968.400 910.530 968.660 910.850 ;
        RECT 969.320 910.530 969.580 910.850 ;
        RECT 968.460 862.765 968.600 910.530 ;
        RECT 968.390 862.395 968.670 862.765 ;
        RECT 969.310 862.395 969.590 862.765 ;
        RECT 969.380 814.290 969.520 862.395 ;
        RECT 969.320 813.970 969.580 814.290 ;
        RECT 969.320 766.030 969.580 766.350 ;
        RECT 969.380 717.730 969.520 766.030 ;
        RECT 969.320 717.410 969.580 717.730 ;
        RECT 969.320 669.470 969.580 669.790 ;
        RECT 969.380 620.830 969.520 669.470 ;
        RECT 969.320 620.510 969.580 620.830 ;
        RECT 969.320 572.570 969.580 572.890 ;
        RECT 969.380 524.270 969.520 572.570 ;
        RECT 969.320 523.950 969.580 524.270 ;
        RECT 969.320 476.010 969.580 476.330 ;
        RECT 969.380 427.710 969.520 476.010 ;
        RECT 969.320 427.390 969.580 427.710 ;
        RECT 969.320 379.450 969.580 379.770 ;
        RECT 969.380 331.150 969.520 379.450 ;
        RECT 969.320 330.830 969.580 331.150 ;
        RECT 969.320 282.890 969.580 283.210 ;
        RECT 969.380 234.590 969.520 282.890 ;
        RECT 969.320 234.270 969.580 234.590 ;
        RECT 969.780 144.850 970.040 145.170 ;
        RECT 969.840 110.570 969.980 144.850 ;
        RECT 968.920 110.430 969.980 110.570 ;
        RECT 968.920 96.550 969.060 110.430 ;
        RECT 968.860 96.230 969.120 96.550 ;
        RECT 968.860 61.890 969.120 62.210 ;
        RECT 968.920 48.690 969.060 61.890 ;
        RECT 968.920 48.550 969.520 48.690 ;
        RECT 969.380 21.070 969.520 48.550 ;
        RECT 969.320 20.750 969.580 21.070 ;
        RECT 1126.640 20.750 1126.900 21.070 ;
        RECT 1126.700 2.400 1126.840 20.750 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
      LAYER via2 ;
        RECT 968.390 1393.520 968.670 1393.800 ;
        RECT 969.310 1393.520 969.590 1393.800 ;
        RECT 968.390 1296.960 968.670 1297.240 ;
        RECT 969.310 1296.960 969.590 1297.240 ;
        RECT 969.310 1208.560 969.590 1208.840 ;
        RECT 969.310 1207.880 969.590 1208.160 ;
        RECT 968.390 1200.400 968.670 1200.680 ;
        RECT 969.310 1200.400 969.590 1200.680 ;
        RECT 968.390 1103.840 968.670 1104.120 ;
        RECT 969.310 1103.840 969.590 1104.120 ;
        RECT 968.390 1055.560 968.670 1055.840 ;
        RECT 969.310 1055.560 969.590 1055.840 ;
        RECT 968.390 959.000 968.670 959.280 ;
        RECT 969.310 959.000 969.590 959.280 ;
        RECT 968.390 862.440 968.670 862.720 ;
        RECT 969.310 862.440 969.590 862.720 ;
      LAYER met3 ;
        RECT 968.365 1393.810 968.695 1393.825 ;
        RECT 969.285 1393.810 969.615 1393.825 ;
        RECT 968.365 1393.510 969.615 1393.810 ;
        RECT 968.365 1393.495 968.695 1393.510 ;
        RECT 969.285 1393.495 969.615 1393.510 ;
        RECT 968.365 1297.250 968.695 1297.265 ;
        RECT 969.285 1297.250 969.615 1297.265 ;
        RECT 968.365 1296.950 969.615 1297.250 ;
        RECT 968.365 1296.935 968.695 1296.950 ;
        RECT 969.285 1296.935 969.615 1296.950 ;
        RECT 969.285 1208.850 969.615 1208.865 ;
        RECT 969.285 1208.550 970.290 1208.850 ;
        RECT 969.285 1208.535 969.615 1208.550 ;
        RECT 969.285 1208.170 969.615 1208.185 ;
        RECT 969.990 1208.170 970.290 1208.550 ;
        RECT 969.285 1207.870 970.290 1208.170 ;
        RECT 969.285 1207.855 969.615 1207.870 ;
        RECT 968.365 1200.690 968.695 1200.705 ;
        RECT 969.285 1200.690 969.615 1200.705 ;
        RECT 968.365 1200.390 969.615 1200.690 ;
        RECT 968.365 1200.375 968.695 1200.390 ;
        RECT 969.285 1200.375 969.615 1200.390 ;
        RECT 968.365 1104.130 968.695 1104.145 ;
        RECT 969.285 1104.130 969.615 1104.145 ;
        RECT 968.365 1103.830 969.615 1104.130 ;
        RECT 968.365 1103.815 968.695 1103.830 ;
        RECT 969.285 1103.815 969.615 1103.830 ;
        RECT 968.365 1055.850 968.695 1055.865 ;
        RECT 969.285 1055.850 969.615 1055.865 ;
        RECT 968.365 1055.550 969.615 1055.850 ;
        RECT 968.365 1055.535 968.695 1055.550 ;
        RECT 969.285 1055.535 969.615 1055.550 ;
        RECT 968.365 959.290 968.695 959.305 ;
        RECT 969.285 959.290 969.615 959.305 ;
        RECT 968.365 958.990 969.615 959.290 ;
        RECT 968.365 958.975 968.695 958.990 ;
        RECT 969.285 958.975 969.615 958.990 ;
        RECT 968.365 862.730 968.695 862.745 ;
        RECT 969.285 862.730 969.615 862.745 ;
        RECT 968.365 862.430 969.615 862.730 ;
        RECT 968.365 862.415 968.695 862.430 ;
        RECT 969.285 862.415 969.615 862.430 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 766.505 1590.265 766.675 1591.795 ;
        RECT 990.065 1545.725 990.235 1589.415 ;
        RECT 1008.005 21.505 1008.175 35.275 ;
        RECT 1024.105 21.335 1024.275 21.675 ;
        RECT 1024.105 21.165 1027.035 21.335 ;
      LAYER mcon ;
        RECT 766.505 1591.625 766.675 1591.795 ;
        RECT 990.065 1589.245 990.235 1589.415 ;
        RECT 1008.005 35.105 1008.175 35.275 ;
        RECT 1024.105 21.505 1024.275 21.675 ;
        RECT 1026.865 21.165 1027.035 21.335 ;
      LAYER met1 ;
        RECT 746.650 1591.780 746.970 1591.840 ;
        RECT 766.445 1591.780 766.735 1591.825 ;
        RECT 746.650 1591.640 766.735 1591.780 ;
        RECT 746.650 1591.580 746.970 1591.640 ;
        RECT 766.445 1591.595 766.735 1591.640 ;
        RECT 766.445 1590.420 766.735 1590.465 ;
        RECT 766.445 1590.280 938.240 1590.420 ;
        RECT 766.445 1590.235 766.735 1590.280 ;
        RECT 938.100 1589.400 938.240 1590.280 ;
        RECT 990.005 1589.400 990.295 1589.445 ;
        RECT 938.100 1589.260 990.295 1589.400 ;
        RECT 990.005 1589.215 990.295 1589.260 ;
        RECT 989.990 1545.880 990.310 1545.940 ;
        RECT 989.795 1545.740 990.310 1545.880 ;
        RECT 989.990 1545.680 990.310 1545.740 ;
        RECT 989.990 35.260 990.310 35.320 ;
        RECT 1007.945 35.260 1008.235 35.305 ;
        RECT 989.990 35.120 1008.235 35.260 ;
        RECT 989.990 35.060 990.310 35.120 ;
        RECT 1007.945 35.075 1008.235 35.120 ;
        RECT 1007.945 21.660 1008.235 21.705 ;
        RECT 1024.045 21.660 1024.335 21.705 ;
        RECT 1007.945 21.520 1024.335 21.660 ;
        RECT 1007.945 21.475 1008.235 21.520 ;
        RECT 1024.045 21.475 1024.335 21.520 ;
        RECT 1026.805 21.320 1027.095 21.365 ;
        RECT 1026.805 21.180 1129.140 21.320 ;
        RECT 1026.805 21.135 1027.095 21.180 ;
        RECT 1129.000 20.980 1129.140 21.180 ;
        RECT 1144.550 20.980 1144.870 21.040 ;
        RECT 1129.000 20.840 1144.870 20.980 ;
        RECT 1144.550 20.780 1144.870 20.840 ;
      LAYER via ;
        RECT 746.680 1591.580 746.940 1591.840 ;
        RECT 990.020 1545.680 990.280 1545.940 ;
        RECT 990.020 35.060 990.280 35.320 ;
        RECT 1144.580 20.780 1144.840 21.040 ;
      LAYER met2 ;
        RECT 746.540 1600.380 746.820 1604.000 ;
        RECT 746.540 1600.000 746.880 1600.380 ;
        RECT 746.740 1591.870 746.880 1600.000 ;
        RECT 746.680 1591.550 746.940 1591.870 ;
        RECT 990.020 1545.650 990.280 1545.970 ;
        RECT 990.080 35.350 990.220 1545.650 ;
        RECT 990.020 35.030 990.280 35.350 ;
        RECT 1144.580 20.750 1144.840 21.070 ;
        RECT 1144.640 2.400 1144.780 20.750 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 764.205 1593.325 764.375 1594.175 ;
        RECT 786.285 1590.605 786.455 1593.495 ;
      LAYER mcon ;
        RECT 764.205 1594.005 764.375 1594.175 ;
        RECT 786.285 1593.325 786.455 1593.495 ;
      LAYER met1 ;
        RECT 754.010 1594.160 754.330 1594.220 ;
        RECT 764.145 1594.160 764.435 1594.205 ;
        RECT 754.010 1594.020 764.435 1594.160 ;
        RECT 754.010 1593.960 754.330 1594.020 ;
        RECT 764.145 1593.975 764.435 1594.020 ;
        RECT 764.145 1593.480 764.435 1593.525 ;
        RECT 786.225 1593.480 786.515 1593.525 ;
        RECT 764.145 1593.340 786.515 1593.480 ;
        RECT 764.145 1593.295 764.435 1593.340 ;
        RECT 786.225 1593.295 786.515 1593.340 ;
        RECT 786.225 1590.760 786.515 1590.805 ;
        RECT 786.225 1590.620 995.280 1590.760 ;
        RECT 786.225 1590.575 786.515 1590.620 ;
        RECT 995.140 1590.080 995.280 1590.620 ;
        RECT 1010.690 1590.080 1011.010 1590.140 ;
        RECT 995.140 1589.940 1011.010 1590.080 ;
        RECT 1010.690 1589.880 1011.010 1589.940 ;
        RECT 1162.490 21.660 1162.810 21.720 ;
        RECT 1026.420 21.520 1162.810 21.660 ;
        RECT 1010.690 21.320 1011.010 21.380 ;
        RECT 1026.420 21.320 1026.560 21.520 ;
        RECT 1162.490 21.460 1162.810 21.520 ;
        RECT 1010.690 21.180 1026.560 21.320 ;
        RECT 1010.690 21.120 1011.010 21.180 ;
      LAYER via ;
        RECT 754.040 1593.960 754.300 1594.220 ;
        RECT 1010.720 1589.880 1010.980 1590.140 ;
        RECT 1010.720 21.120 1010.980 21.380 ;
        RECT 1162.520 21.460 1162.780 21.720 ;
      LAYER met2 ;
        RECT 752.520 1600.450 752.800 1604.000 ;
        RECT 752.520 1600.310 754.240 1600.450 ;
        RECT 752.520 1600.000 752.800 1600.310 ;
        RECT 754.100 1594.250 754.240 1600.310 ;
        RECT 754.040 1593.930 754.300 1594.250 ;
        RECT 1010.720 1589.850 1010.980 1590.170 ;
        RECT 1010.780 21.410 1010.920 1589.850 ;
        RECT 1162.520 21.430 1162.780 21.750 ;
        RECT 1010.720 21.090 1010.980 21.410 ;
        RECT 1162.580 2.400 1162.720 21.430 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 585.650 1593.140 585.970 1593.200 ;
        RECT 666.150 1593.140 666.470 1593.200 ;
        RECT 585.650 1593.000 666.470 1593.140 ;
        RECT 585.650 1592.940 585.970 1593.000 ;
        RECT 666.150 1592.940 666.470 1593.000 ;
        RECT 666.150 17.580 666.470 17.640 ;
        RECT 680.410 17.580 680.730 17.640 ;
        RECT 666.150 17.440 680.730 17.580 ;
        RECT 666.150 17.380 666.470 17.440 ;
        RECT 680.410 17.380 680.730 17.440 ;
      LAYER via ;
        RECT 585.680 1592.940 585.940 1593.200 ;
        RECT 666.180 1592.940 666.440 1593.200 ;
        RECT 666.180 17.380 666.440 17.640 ;
        RECT 680.440 17.380 680.700 17.640 ;
      LAYER met2 ;
        RECT 585.540 1600.380 585.820 1604.000 ;
        RECT 585.540 1600.000 585.880 1600.380 ;
        RECT 585.740 1593.230 585.880 1600.000 ;
        RECT 585.680 1592.910 585.940 1593.230 ;
        RECT 666.180 1592.910 666.440 1593.230 ;
        RECT 666.240 17.670 666.380 1592.910 ;
        RECT 666.180 17.350 666.440 17.670 ;
        RECT 680.440 17.350 680.700 17.670 ;
        RECT 680.500 2.400 680.640 17.350 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 759.070 1587.360 759.390 1587.420 ;
        RECT 763.210 1587.360 763.530 1587.420 ;
        RECT 759.070 1587.220 763.530 1587.360 ;
        RECT 759.070 1587.160 759.390 1587.220 ;
        RECT 763.210 1587.160 763.530 1587.220 ;
        RECT 764.130 43.420 764.450 43.480 ;
        RECT 1179.970 43.420 1180.290 43.480 ;
        RECT 764.130 43.280 1180.290 43.420 ;
        RECT 764.130 43.220 764.450 43.280 ;
        RECT 1179.970 43.220 1180.290 43.280 ;
      LAYER via ;
        RECT 759.100 1587.160 759.360 1587.420 ;
        RECT 763.240 1587.160 763.500 1587.420 ;
        RECT 764.160 43.220 764.420 43.480 ;
        RECT 1180.000 43.220 1180.260 43.480 ;
      LAYER met2 ;
        RECT 758.960 1600.380 759.240 1604.000 ;
        RECT 758.960 1600.000 759.300 1600.380 ;
        RECT 759.160 1587.450 759.300 1600.000 ;
        RECT 759.100 1587.130 759.360 1587.450 ;
        RECT 763.240 1587.130 763.500 1587.450 ;
        RECT 763.300 1579.370 763.440 1587.130 ;
        RECT 763.300 1579.230 764.360 1579.370 ;
        RECT 764.220 43.510 764.360 1579.230 ;
        RECT 764.160 43.190 764.420 43.510 ;
        RECT 1180.000 43.190 1180.260 43.510 ;
        RECT 1180.060 2.400 1180.200 43.190 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 806.525 43.945 806.695 44.795 ;
        RECT 835.045 42.925 835.215 44.115 ;
        RECT 882.885 42.925 883.055 44.115 ;
        RECT 931.645 41.905 931.815 44.115 ;
        RECT 979.025 43.945 979.655 44.115 ;
        RECT 979.025 42.245 979.195 43.945 ;
      LAYER mcon ;
        RECT 806.525 44.625 806.695 44.795 ;
        RECT 835.045 43.945 835.215 44.115 ;
        RECT 882.885 43.945 883.055 44.115 ;
        RECT 931.645 43.945 931.815 44.115 ;
        RECT 979.485 43.945 979.655 44.115 ;
      LAYER met1 ;
        RECT 765.050 44.780 765.370 44.840 ;
        RECT 806.465 44.780 806.755 44.825 ;
        RECT 765.050 44.640 806.755 44.780 ;
        RECT 765.050 44.580 765.370 44.640 ;
        RECT 806.465 44.595 806.755 44.640 ;
        RECT 806.465 44.100 806.755 44.145 ;
        RECT 834.985 44.100 835.275 44.145 ;
        RECT 806.465 43.960 835.275 44.100 ;
        RECT 806.465 43.915 806.755 43.960 ;
        RECT 834.985 43.915 835.275 43.960 ;
        RECT 882.825 44.100 883.115 44.145 ;
        RECT 931.585 44.100 931.875 44.145 ;
        RECT 882.825 43.960 931.875 44.100 ;
        RECT 882.825 43.915 883.115 43.960 ;
        RECT 931.585 43.915 931.875 43.960 ;
        RECT 979.425 44.100 979.715 44.145 ;
        RECT 1028.170 44.100 1028.490 44.160 ;
        RECT 979.425 43.960 1028.490 44.100 ;
        RECT 979.425 43.915 979.715 43.960 ;
        RECT 1028.170 43.900 1028.490 43.960 ;
        RECT 1075.550 44.100 1075.870 44.160 ;
        RECT 1124.770 44.100 1125.090 44.160 ;
        RECT 1075.550 43.960 1125.090 44.100 ;
        RECT 1075.550 43.900 1075.870 43.960 ;
        RECT 1124.770 43.900 1125.090 43.960 ;
        RECT 834.985 43.080 835.275 43.125 ;
        RECT 882.825 43.080 883.115 43.125 ;
        RECT 834.985 42.940 883.115 43.080 ;
        RECT 834.985 42.895 835.275 42.940 ;
        RECT 882.825 42.895 883.115 42.940 ;
        RECT 978.965 42.400 979.255 42.445 ;
        RECT 951.900 42.260 979.255 42.400 ;
        RECT 931.585 42.060 931.875 42.105 ;
        RECT 951.900 42.060 952.040 42.260 ;
        RECT 978.965 42.215 979.255 42.260 ;
        RECT 931.585 41.920 952.040 42.060 ;
        RECT 931.585 41.875 931.875 41.920 ;
      LAYER via ;
        RECT 765.080 44.580 765.340 44.840 ;
        RECT 1028.200 43.900 1028.460 44.160 ;
        RECT 1075.580 43.900 1075.840 44.160 ;
        RECT 1124.800 43.900 1125.060 44.160 ;
      LAYER met2 ;
        RECT 764.940 1600.380 765.220 1604.000 ;
        RECT 764.940 1600.000 765.280 1600.380 ;
        RECT 765.140 44.870 765.280 1600.000 ;
        RECT 765.080 44.550 765.340 44.870 ;
        RECT 1028.200 44.045 1028.460 44.190 ;
        RECT 1075.580 44.045 1075.840 44.190 ;
        RECT 1124.800 44.045 1125.060 44.190 ;
        RECT 1028.190 43.675 1028.470 44.045 ;
        RECT 1075.570 43.675 1075.850 44.045 ;
        RECT 1124.790 43.675 1125.070 44.045 ;
        RECT 1197.930 43.675 1198.210 44.045 ;
        RECT 1198.000 2.400 1198.140 43.675 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
      LAYER via2 ;
        RECT 1028.190 43.720 1028.470 44.000 ;
        RECT 1075.570 43.720 1075.850 44.000 ;
        RECT 1124.790 43.720 1125.070 44.000 ;
        RECT 1197.930 43.720 1198.210 44.000 ;
      LAYER met3 ;
        RECT 1028.165 44.010 1028.495 44.025 ;
        RECT 1075.545 44.010 1075.875 44.025 ;
        RECT 1028.165 43.710 1075.875 44.010 ;
        RECT 1028.165 43.695 1028.495 43.710 ;
        RECT 1075.545 43.695 1075.875 43.710 ;
        RECT 1124.765 44.010 1125.095 44.025 ;
        RECT 1197.905 44.010 1198.235 44.025 ;
        RECT 1124.765 43.710 1198.235 44.010 ;
        RECT 1124.765 43.695 1125.095 43.710 ;
        RECT 1197.905 43.695 1198.235 43.710 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1194.305 43.265 1194.475 48.195 ;
      LAYER mcon ;
        RECT 1194.305 48.025 1194.475 48.195 ;
      LAYER met1 ;
        RECT 771.950 48.180 772.270 48.240 ;
        RECT 1194.245 48.180 1194.535 48.225 ;
        RECT 771.950 48.040 1194.535 48.180 ;
        RECT 771.950 47.980 772.270 48.040 ;
        RECT 1194.245 47.995 1194.535 48.040 ;
        RECT 1194.245 43.420 1194.535 43.465 ;
        RECT 1215.850 43.420 1216.170 43.480 ;
        RECT 1194.245 43.280 1216.170 43.420 ;
        RECT 1194.245 43.235 1194.535 43.280 ;
        RECT 1215.850 43.220 1216.170 43.280 ;
      LAYER via ;
        RECT 771.980 47.980 772.240 48.240 ;
        RECT 1215.880 43.220 1216.140 43.480 ;
      LAYER met2 ;
        RECT 771.380 1600.450 771.660 1604.000 ;
        RECT 771.380 1600.310 772.180 1600.450 ;
        RECT 771.380 1600.000 771.660 1600.310 ;
        RECT 772.040 48.270 772.180 1600.310 ;
        RECT 771.980 47.950 772.240 48.270 ;
        RECT 1215.880 43.190 1216.140 43.510 ;
        RECT 1215.940 2.400 1216.080 43.190 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1233.790 47.840 1234.110 47.900 ;
        RECT 1197.080 47.700 1234.110 47.840 ;
        RECT 778.390 47.500 778.710 47.560 ;
        RECT 1197.080 47.500 1197.220 47.700 ;
        RECT 1233.790 47.640 1234.110 47.700 ;
        RECT 778.390 47.360 1197.220 47.500 ;
        RECT 778.390 47.300 778.710 47.360 ;
      LAYER via ;
        RECT 778.420 47.300 778.680 47.560 ;
        RECT 1233.820 47.640 1234.080 47.900 ;
      LAYER met2 ;
        RECT 777.360 1600.450 777.640 1604.000 ;
        RECT 777.360 1600.310 778.620 1600.450 ;
        RECT 777.360 1600.000 777.640 1600.310 ;
        RECT 778.480 47.590 778.620 1600.310 ;
        RECT 1233.820 47.610 1234.080 47.930 ;
        RECT 778.420 47.270 778.680 47.590 ;
        RECT 1233.880 2.400 1234.020 47.610 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1197.065 46.665 1197.235 48.195 ;
      LAYER mcon ;
        RECT 1197.065 48.025 1197.235 48.195 ;
      LAYER met1 ;
        RECT 1197.005 48.180 1197.295 48.225 ;
        RECT 1251.730 48.180 1252.050 48.240 ;
        RECT 1197.005 48.040 1252.050 48.180 ;
        RECT 1197.005 47.995 1197.295 48.040 ;
        RECT 1251.730 47.980 1252.050 48.040 ;
        RECT 784.830 46.820 785.150 46.880 ;
        RECT 1197.005 46.820 1197.295 46.865 ;
        RECT 784.830 46.680 1197.295 46.820 ;
        RECT 784.830 46.620 785.150 46.680 ;
        RECT 1197.005 46.635 1197.295 46.680 ;
      LAYER via ;
        RECT 1251.760 47.980 1252.020 48.240 ;
        RECT 784.860 46.620 785.120 46.880 ;
      LAYER met2 ;
        RECT 783.800 1600.450 784.080 1604.000 ;
        RECT 783.800 1600.310 785.060 1600.450 ;
        RECT 783.800 1600.000 784.080 1600.310 ;
        RECT 784.920 46.910 785.060 1600.310 ;
        RECT 1251.760 47.950 1252.020 48.270 ;
        RECT 784.860 46.590 785.120 46.910 ;
        RECT 1251.820 2.400 1251.960 47.950 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1233.405 46.325 1233.575 47.515 ;
      LAYER mcon ;
        RECT 1233.405 47.345 1233.575 47.515 ;
      LAYER met1 ;
        RECT 1234.340 47.700 1248.740 47.840 ;
        RECT 1233.345 47.500 1233.635 47.545 ;
        RECT 1234.340 47.500 1234.480 47.700 ;
        RECT 1233.345 47.360 1234.480 47.500 ;
        RECT 1233.345 47.315 1233.635 47.360 ;
        RECT 1248.600 47.160 1248.740 47.700 ;
        RECT 1269.210 47.160 1269.530 47.220 ;
        RECT 1248.600 47.020 1269.530 47.160 ;
        RECT 1269.210 46.960 1269.530 47.020 ;
        RECT 792.650 46.480 792.970 46.540 ;
        RECT 1233.345 46.480 1233.635 46.525 ;
        RECT 792.650 46.340 1233.635 46.480 ;
        RECT 792.650 46.280 792.970 46.340 ;
        RECT 1233.345 46.295 1233.635 46.340 ;
      LAYER via ;
        RECT 1269.240 46.960 1269.500 47.220 ;
        RECT 792.680 46.280 792.940 46.540 ;
      LAYER met2 ;
        RECT 789.780 1600.450 790.060 1604.000 ;
        RECT 789.780 1600.310 791.500 1600.450 ;
        RECT 789.780 1600.000 790.060 1600.310 ;
        RECT 791.360 1580.050 791.500 1600.310 ;
        RECT 791.360 1579.910 792.880 1580.050 ;
        RECT 792.740 46.570 792.880 1579.910 ;
        RECT 1269.240 46.930 1269.500 47.250 ;
        RECT 792.680 46.250 792.940 46.570 ;
        RECT 1269.300 2.400 1269.440 46.930 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1002.945 1591.965 1003.115 1594.175 ;
        RECT 1024.565 1545.725 1024.735 1593.835 ;
        RECT 1023.645 379.525 1023.815 427.635 ;
        RECT 1024.565 282.965 1024.735 331.075 ;
        RECT 1024.565 186.405 1024.735 234.515 ;
        RECT 1024.565 89.845 1024.735 137.955 ;
        RECT 1025.945 21.845 1026.115 35.275 ;
        RECT 1220.525 21.845 1222.075 22.015 ;
      LAYER mcon ;
        RECT 1002.945 1594.005 1003.115 1594.175 ;
        RECT 1024.565 1593.665 1024.735 1593.835 ;
        RECT 1023.645 427.465 1023.815 427.635 ;
        RECT 1024.565 330.905 1024.735 331.075 ;
        RECT 1024.565 234.345 1024.735 234.515 ;
        RECT 1024.565 137.785 1024.735 137.955 ;
        RECT 1025.945 35.105 1026.115 35.275 ;
        RECT 1221.905 21.845 1222.075 22.015 ;
      LAYER met1 ;
        RECT 1002.885 1594.160 1003.175 1594.205 ;
        RECT 1002.885 1594.020 1004.480 1594.160 ;
        RECT 1002.885 1593.975 1003.175 1594.020 ;
        RECT 1004.340 1593.820 1004.480 1594.020 ;
        RECT 1024.505 1593.820 1024.795 1593.865 ;
        RECT 1004.340 1593.680 1024.795 1593.820 ;
        RECT 1024.505 1593.635 1024.795 1593.680 ;
        RECT 796.330 1592.120 796.650 1592.180 ;
        RECT 1002.885 1592.120 1003.175 1592.165 ;
        RECT 796.330 1591.980 1003.175 1592.120 ;
        RECT 796.330 1591.920 796.650 1591.980 ;
        RECT 1002.885 1591.935 1003.175 1591.980 ;
        RECT 1024.490 1545.880 1024.810 1545.940 ;
        RECT 1024.295 1545.740 1024.810 1545.880 ;
        RECT 1024.490 1545.680 1024.810 1545.740 ;
        RECT 1024.490 918.240 1024.810 918.300 ;
        RECT 1023.660 918.100 1024.810 918.240 ;
        RECT 1023.660 917.960 1023.800 918.100 ;
        RECT 1024.490 918.040 1024.810 918.100 ;
        RECT 1023.570 917.700 1023.890 917.960 ;
        RECT 1023.570 869.620 1023.890 869.680 ;
        RECT 1024.490 869.620 1024.810 869.680 ;
        RECT 1023.570 869.480 1024.810 869.620 ;
        RECT 1023.570 869.420 1023.890 869.480 ;
        RECT 1024.490 869.420 1024.810 869.480 ;
        RECT 1024.030 820.660 1024.350 820.720 ;
        RECT 1024.490 820.660 1024.810 820.720 ;
        RECT 1024.030 820.520 1024.810 820.660 ;
        RECT 1024.030 820.460 1024.350 820.520 ;
        RECT 1024.490 820.460 1024.810 820.520 ;
        RECT 1024.030 724.100 1024.350 724.160 ;
        RECT 1024.490 724.100 1024.810 724.160 ;
        RECT 1024.030 723.960 1024.810 724.100 ;
        RECT 1024.030 723.900 1024.350 723.960 ;
        RECT 1024.490 723.900 1024.810 723.960 ;
        RECT 1024.490 579.940 1024.810 580.000 ;
        RECT 1025.410 579.940 1025.730 580.000 ;
        RECT 1024.490 579.800 1025.730 579.940 ;
        RECT 1024.490 579.740 1024.810 579.800 ;
        RECT 1025.410 579.740 1025.730 579.800 ;
        RECT 1023.570 531.660 1023.890 531.720 ;
        RECT 1024.490 531.660 1024.810 531.720 ;
        RECT 1023.570 531.520 1024.810 531.660 ;
        RECT 1023.570 531.460 1023.890 531.520 ;
        RECT 1024.490 531.460 1024.810 531.520 ;
        RECT 1023.570 483.380 1023.890 483.440 ;
        RECT 1024.490 483.380 1024.810 483.440 ;
        RECT 1023.570 483.240 1024.810 483.380 ;
        RECT 1023.570 483.180 1023.890 483.240 ;
        RECT 1024.490 483.180 1024.810 483.240 ;
        RECT 1023.570 435.100 1023.890 435.160 ;
        RECT 1024.490 435.100 1024.810 435.160 ;
        RECT 1023.570 434.960 1024.810 435.100 ;
        RECT 1023.570 434.900 1023.890 434.960 ;
        RECT 1024.490 434.900 1024.810 434.960 ;
        RECT 1023.570 427.620 1023.890 427.680 ;
        RECT 1023.375 427.480 1023.890 427.620 ;
        RECT 1023.570 427.420 1023.890 427.480 ;
        RECT 1023.585 379.680 1023.875 379.725 ;
        RECT 1024.490 379.680 1024.810 379.740 ;
        RECT 1023.585 379.540 1024.810 379.680 ;
        RECT 1023.585 379.495 1023.875 379.540 ;
        RECT 1024.490 379.480 1024.810 379.540 ;
        RECT 1024.490 331.060 1024.810 331.120 ;
        RECT 1024.295 330.920 1024.810 331.060 ;
        RECT 1024.490 330.860 1024.810 330.920 ;
        RECT 1024.490 283.120 1024.810 283.180 ;
        RECT 1024.295 282.980 1024.810 283.120 ;
        RECT 1024.490 282.920 1024.810 282.980 ;
        RECT 1024.490 234.500 1024.810 234.560 ;
        RECT 1024.295 234.360 1024.810 234.500 ;
        RECT 1024.490 234.300 1024.810 234.360 ;
        RECT 1024.490 186.560 1024.810 186.620 ;
        RECT 1024.295 186.420 1024.810 186.560 ;
        RECT 1024.490 186.360 1024.810 186.420 ;
        RECT 1024.490 137.940 1024.810 138.000 ;
        RECT 1024.295 137.800 1024.810 137.940 ;
        RECT 1024.490 137.740 1024.810 137.800 ;
        RECT 1024.490 90.000 1024.810 90.060 ;
        RECT 1024.295 89.860 1024.810 90.000 ;
        RECT 1024.490 89.800 1024.810 89.860 ;
        RECT 1024.030 35.260 1024.350 35.320 ;
        RECT 1025.885 35.260 1026.175 35.305 ;
        RECT 1024.030 35.120 1026.175 35.260 ;
        RECT 1024.030 35.060 1024.350 35.120 ;
        RECT 1025.885 35.075 1026.175 35.120 ;
        RECT 1287.150 23.020 1287.470 23.080 ;
        RECT 1245.380 22.880 1287.470 23.020 ;
        RECT 1025.885 22.000 1026.175 22.045 ;
        RECT 1159.270 22.000 1159.590 22.060 ;
        RECT 1220.465 22.000 1220.755 22.045 ;
        RECT 1025.885 21.860 1159.590 22.000 ;
        RECT 1025.885 21.815 1026.175 21.860 ;
        RECT 1159.270 21.800 1159.590 21.860 ;
        RECT 1197.080 21.860 1220.755 22.000 ;
        RECT 1159.730 21.320 1160.050 21.380 ;
        RECT 1197.080 21.320 1197.220 21.860 ;
        RECT 1220.465 21.815 1220.755 21.860 ;
        RECT 1221.845 22.000 1222.135 22.045 ;
        RECT 1245.380 22.000 1245.520 22.880 ;
        RECT 1287.150 22.820 1287.470 22.880 ;
        RECT 1221.845 21.860 1245.520 22.000 ;
        RECT 1221.845 21.815 1222.135 21.860 ;
        RECT 1159.730 21.180 1197.220 21.320 ;
        RECT 1159.730 21.120 1160.050 21.180 ;
      LAYER via ;
        RECT 796.360 1591.920 796.620 1592.180 ;
        RECT 1024.520 1545.680 1024.780 1545.940 ;
        RECT 1024.520 918.040 1024.780 918.300 ;
        RECT 1023.600 917.700 1023.860 917.960 ;
        RECT 1023.600 869.420 1023.860 869.680 ;
        RECT 1024.520 869.420 1024.780 869.680 ;
        RECT 1024.060 820.460 1024.320 820.720 ;
        RECT 1024.520 820.460 1024.780 820.720 ;
        RECT 1024.060 723.900 1024.320 724.160 ;
        RECT 1024.520 723.900 1024.780 724.160 ;
        RECT 1024.520 579.740 1024.780 580.000 ;
        RECT 1025.440 579.740 1025.700 580.000 ;
        RECT 1023.600 531.460 1023.860 531.720 ;
        RECT 1024.520 531.460 1024.780 531.720 ;
        RECT 1023.600 483.180 1023.860 483.440 ;
        RECT 1024.520 483.180 1024.780 483.440 ;
        RECT 1023.600 434.900 1023.860 435.160 ;
        RECT 1024.520 434.900 1024.780 435.160 ;
        RECT 1023.600 427.420 1023.860 427.680 ;
        RECT 1024.520 379.480 1024.780 379.740 ;
        RECT 1024.520 330.860 1024.780 331.120 ;
        RECT 1024.520 282.920 1024.780 283.180 ;
        RECT 1024.520 234.300 1024.780 234.560 ;
        RECT 1024.520 186.360 1024.780 186.620 ;
        RECT 1024.520 137.740 1024.780 138.000 ;
        RECT 1024.520 89.800 1024.780 90.060 ;
        RECT 1024.060 35.060 1024.320 35.320 ;
        RECT 1159.300 21.800 1159.560 22.060 ;
        RECT 1159.760 21.120 1160.020 21.380 ;
        RECT 1287.180 22.820 1287.440 23.080 ;
      LAYER met2 ;
        RECT 796.220 1600.380 796.500 1604.000 ;
        RECT 796.220 1600.000 796.560 1600.380 ;
        RECT 796.420 1592.210 796.560 1600.000 ;
        RECT 796.360 1591.890 796.620 1592.210 ;
        RECT 1024.520 1545.650 1024.780 1545.970 ;
        RECT 1024.580 918.330 1024.720 1545.650 ;
        RECT 1024.520 918.010 1024.780 918.330 ;
        RECT 1023.600 917.670 1023.860 917.990 ;
        RECT 1023.660 869.710 1023.800 917.670 ;
        RECT 1023.600 869.390 1023.860 869.710 ;
        RECT 1024.520 869.390 1024.780 869.710 ;
        RECT 1024.580 820.750 1024.720 869.390 ;
        RECT 1024.060 820.430 1024.320 820.750 ;
        RECT 1024.520 820.430 1024.780 820.750 ;
        RECT 1024.120 773.685 1024.260 820.430 ;
        RECT 1024.050 773.315 1024.330 773.685 ;
        RECT 1024.510 772.635 1024.790 773.005 ;
        RECT 1024.580 724.190 1024.720 772.635 ;
        RECT 1024.060 723.870 1024.320 724.190 ;
        RECT 1024.520 723.870 1024.780 724.190 ;
        RECT 1024.120 677.125 1024.260 723.870 ;
        RECT 1024.050 676.755 1024.330 677.125 ;
        RECT 1024.510 676.075 1024.790 676.445 ;
        RECT 1024.580 651.850 1024.720 676.075 ;
        RECT 1024.580 651.710 1025.180 651.850 ;
        RECT 1025.040 628.050 1025.180 651.710 ;
        RECT 1025.040 627.910 1025.640 628.050 ;
        RECT 1025.500 580.030 1025.640 627.910 ;
        RECT 1024.520 579.710 1024.780 580.030 ;
        RECT 1025.440 579.710 1025.700 580.030 ;
        RECT 1024.580 531.750 1024.720 579.710 ;
        RECT 1023.600 531.430 1023.860 531.750 ;
        RECT 1024.520 531.430 1024.780 531.750 ;
        RECT 1023.660 483.470 1023.800 531.430 ;
        RECT 1023.600 483.150 1023.860 483.470 ;
        RECT 1024.520 483.150 1024.780 483.470 ;
        RECT 1024.580 435.190 1024.720 483.150 ;
        RECT 1023.600 434.870 1023.860 435.190 ;
        RECT 1024.520 434.870 1024.780 435.190 ;
        RECT 1023.660 427.710 1023.800 434.870 ;
        RECT 1023.600 427.390 1023.860 427.710 ;
        RECT 1024.520 379.450 1024.780 379.770 ;
        RECT 1024.580 331.150 1024.720 379.450 ;
        RECT 1024.520 330.830 1024.780 331.150 ;
        RECT 1024.520 282.890 1024.780 283.210 ;
        RECT 1024.580 234.590 1024.720 282.890 ;
        RECT 1024.520 234.270 1024.780 234.590 ;
        RECT 1024.520 186.330 1024.780 186.650 ;
        RECT 1024.580 138.030 1024.720 186.330 ;
        RECT 1024.520 137.710 1024.780 138.030 ;
        RECT 1024.520 89.770 1024.780 90.090 ;
        RECT 1024.580 48.690 1024.720 89.770 ;
        RECT 1024.120 48.550 1024.720 48.690 ;
        RECT 1024.120 35.350 1024.260 48.550 ;
        RECT 1024.060 35.030 1024.320 35.350 ;
        RECT 1287.180 22.790 1287.440 23.110 ;
        RECT 1159.300 21.770 1159.560 22.090 ;
        RECT 1159.360 21.490 1159.500 21.770 ;
        RECT 1159.360 21.410 1159.960 21.490 ;
        RECT 1159.360 21.350 1160.020 21.410 ;
        RECT 1159.760 21.090 1160.020 21.350 ;
        RECT 1287.240 2.400 1287.380 22.790 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
      LAYER via2 ;
        RECT 1024.050 773.360 1024.330 773.640 ;
        RECT 1024.510 772.680 1024.790 772.960 ;
        RECT 1024.050 676.800 1024.330 677.080 ;
        RECT 1024.510 676.120 1024.790 676.400 ;
      LAYER met3 ;
        RECT 1024.025 773.650 1024.355 773.665 ;
        RECT 1024.025 773.335 1024.570 773.650 ;
        RECT 1024.270 772.985 1024.570 773.335 ;
        RECT 1024.270 772.670 1024.815 772.985 ;
        RECT 1024.485 772.655 1024.815 772.670 ;
        RECT 1024.025 677.090 1024.355 677.105 ;
        RECT 1024.025 676.775 1024.570 677.090 ;
        RECT 1024.270 676.425 1024.570 676.775 ;
        RECT 1024.270 676.110 1024.815 676.425 ;
        RECT 1024.485 676.095 1024.815 676.110 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1287.225 23.885 1287.395 25.075 ;
        RECT 1058.605 22.525 1061.995 22.695 ;
        RECT 1058.605 22.185 1058.775 22.525 ;
        RECT 1129.445 21.165 1129.615 22.355 ;
        RECT 1159.805 21.335 1159.975 22.015 ;
        RECT 1163.025 21.845 1163.655 22.015 ;
        RECT 1159.345 21.165 1159.975 21.335 ;
      LAYER mcon ;
        RECT 1287.225 24.905 1287.395 25.075 ;
        RECT 1061.825 22.525 1061.995 22.695 ;
        RECT 1129.445 22.185 1129.615 22.355 ;
        RECT 1159.805 21.845 1159.975 22.015 ;
        RECT 1163.485 21.845 1163.655 22.015 ;
      LAYER met1 ;
        RECT 1045.190 1592.120 1045.510 1592.180 ;
        RECT 1003.880 1591.980 1045.510 1592.120 ;
        RECT 802.310 1591.780 802.630 1591.840 ;
        RECT 1003.880 1591.780 1004.020 1591.980 ;
        RECT 1045.190 1591.920 1045.510 1591.980 ;
        RECT 802.310 1591.640 1004.020 1591.780 ;
        RECT 802.310 1591.580 802.630 1591.640 ;
        RECT 1287.165 25.060 1287.455 25.105 ;
        RECT 1305.090 25.060 1305.410 25.120 ;
        RECT 1287.165 24.920 1305.410 25.060 ;
        RECT 1287.165 24.875 1287.455 24.920 ;
        RECT 1305.090 24.860 1305.410 24.920 ;
        RECT 1287.165 24.040 1287.455 24.085 ;
        RECT 1274.820 23.900 1287.455 24.040 ;
        RECT 1245.290 23.700 1245.610 23.760 ;
        RECT 1274.820 23.700 1274.960 23.900 ;
        RECT 1287.165 23.855 1287.455 23.900 ;
        RECT 1245.290 23.560 1274.960 23.700 ;
        RECT 1245.290 23.500 1245.610 23.560 ;
        RECT 1061.765 22.680 1062.055 22.725 ;
        RECT 1075.550 22.680 1075.870 22.740 ;
        RECT 1061.765 22.540 1075.870 22.680 ;
        RECT 1061.765 22.495 1062.055 22.540 ;
        RECT 1075.550 22.480 1075.870 22.540 ;
        RECT 1045.190 22.340 1045.510 22.400 ;
        RECT 1058.545 22.340 1058.835 22.385 ;
        RECT 1045.190 22.200 1058.835 22.340 ;
        RECT 1045.190 22.140 1045.510 22.200 ;
        RECT 1058.545 22.155 1058.835 22.200 ;
        RECT 1076.470 22.340 1076.790 22.400 ;
        RECT 1129.385 22.340 1129.675 22.385 ;
        RECT 1220.910 22.340 1221.230 22.400 ;
        RECT 1076.470 22.200 1129.675 22.340 ;
        RECT 1076.470 22.140 1076.790 22.200 ;
        RECT 1129.385 22.155 1129.675 22.200 ;
        RECT 1196.620 22.200 1221.230 22.340 ;
        RECT 1159.745 22.000 1160.035 22.045 ;
        RECT 1162.965 22.000 1163.255 22.045 ;
        RECT 1159.745 21.860 1163.255 22.000 ;
        RECT 1159.745 21.815 1160.035 21.860 ;
        RECT 1162.965 21.815 1163.255 21.860 ;
        RECT 1163.425 22.000 1163.715 22.045 ;
        RECT 1196.620 22.000 1196.760 22.200 ;
        RECT 1220.910 22.140 1221.230 22.200 ;
        RECT 1163.425 21.860 1196.760 22.000 ;
        RECT 1163.425 21.815 1163.715 21.860 ;
        RECT 1129.385 21.320 1129.675 21.365 ;
        RECT 1159.285 21.320 1159.575 21.365 ;
        RECT 1129.385 21.180 1159.575 21.320 ;
        RECT 1129.385 21.135 1129.675 21.180 ;
        RECT 1159.285 21.135 1159.575 21.180 ;
      LAYER via ;
        RECT 802.340 1591.580 802.600 1591.840 ;
        RECT 1045.220 1591.920 1045.480 1592.180 ;
        RECT 1305.120 24.860 1305.380 25.120 ;
        RECT 1245.320 23.500 1245.580 23.760 ;
        RECT 1075.580 22.480 1075.840 22.740 ;
        RECT 1045.220 22.140 1045.480 22.400 ;
        RECT 1076.500 22.140 1076.760 22.400 ;
        RECT 1220.940 22.140 1221.200 22.400 ;
      LAYER met2 ;
        RECT 802.200 1600.380 802.480 1604.000 ;
        RECT 802.200 1600.000 802.540 1600.380 ;
        RECT 802.400 1591.870 802.540 1600.000 ;
        RECT 1045.220 1591.890 1045.480 1592.210 ;
        RECT 802.340 1591.550 802.600 1591.870 ;
        RECT 1045.280 22.430 1045.420 1591.890 ;
        RECT 1305.120 24.830 1305.380 25.150 ;
        RECT 1245.320 23.470 1245.580 23.790 ;
        RECT 1245.380 22.965 1245.520 23.470 ;
        RECT 1075.580 22.450 1075.840 22.770 ;
        RECT 1220.930 22.595 1221.210 22.965 ;
        RECT 1245.310 22.595 1245.590 22.965 ;
        RECT 1045.220 22.110 1045.480 22.430 ;
        RECT 1075.640 22.285 1075.780 22.450 ;
        RECT 1221.000 22.430 1221.140 22.595 ;
        RECT 1076.500 22.285 1076.760 22.430 ;
        RECT 1075.570 21.915 1075.850 22.285 ;
        RECT 1076.490 21.915 1076.770 22.285 ;
        RECT 1220.940 22.110 1221.200 22.430 ;
        RECT 1305.180 2.400 1305.320 24.830 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
      LAYER via2 ;
        RECT 1220.930 22.640 1221.210 22.920 ;
        RECT 1245.310 22.640 1245.590 22.920 ;
        RECT 1075.570 21.960 1075.850 22.240 ;
        RECT 1076.490 21.960 1076.770 22.240 ;
      LAYER met3 ;
        RECT 1220.905 22.930 1221.235 22.945 ;
        RECT 1245.285 22.930 1245.615 22.945 ;
        RECT 1220.905 22.630 1245.615 22.930 ;
        RECT 1220.905 22.615 1221.235 22.630 ;
        RECT 1245.285 22.615 1245.615 22.630 ;
        RECT 1075.545 22.250 1075.875 22.265 ;
        RECT 1076.465 22.250 1076.795 22.265 ;
        RECT 1075.545 21.950 1076.795 22.250 ;
        RECT 1075.545 21.935 1075.875 21.950 ;
        RECT 1076.465 21.935 1076.795 21.950 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1003.405 1590.605 1003.575 1592.475 ;
        RECT 1059.525 786.505 1059.695 821.015 ;
        RECT 1059.525 689.605 1059.695 724.455 ;
        RECT 1059.525 593.045 1059.695 627.895 ;
        RECT 1059.525 496.485 1059.695 531.335 ;
        RECT 1059.525 386.325 1059.695 434.775 ;
        RECT 1059.525 351.645 1059.695 379.355 ;
        RECT 1059.525 253.385 1059.695 289.595 ;
        RECT 1059.525 144.925 1059.695 193.035 ;
        RECT 1076.085 22.185 1076.255 24.055 ;
        RECT 1077.005 23.885 1077.635 24.055 ;
        RECT 1274.345 23.885 1274.515 25.415 ;
        RECT 1077.465 23.545 1077.635 23.885 ;
        RECT 1095.865 22.525 1096.035 23.375 ;
        RECT 1148.305 20.825 1148.475 22.695 ;
        RECT 1197.065 20.825 1197.235 22.695 ;
      LAYER mcon ;
        RECT 1003.405 1592.305 1003.575 1592.475 ;
        RECT 1059.525 820.845 1059.695 821.015 ;
        RECT 1059.525 724.285 1059.695 724.455 ;
        RECT 1059.525 627.725 1059.695 627.895 ;
        RECT 1059.525 531.165 1059.695 531.335 ;
        RECT 1059.525 434.605 1059.695 434.775 ;
        RECT 1059.525 379.185 1059.695 379.355 ;
        RECT 1059.525 289.425 1059.695 289.595 ;
        RECT 1059.525 192.865 1059.695 193.035 ;
        RECT 1274.345 25.245 1274.515 25.415 ;
        RECT 1076.085 23.885 1076.255 24.055 ;
        RECT 1095.865 23.205 1096.035 23.375 ;
        RECT 1148.305 22.525 1148.475 22.695 ;
        RECT 1197.065 22.525 1197.235 22.695 ;
      LAYER met1 ;
        RECT 808.290 1592.460 808.610 1592.520 ;
        RECT 1003.345 1592.460 1003.635 1592.505 ;
        RECT 808.290 1592.320 1003.635 1592.460 ;
        RECT 808.290 1592.260 808.610 1592.320 ;
        RECT 1003.345 1592.275 1003.635 1592.320 ;
        RECT 1003.345 1590.760 1003.635 1590.805 ;
        RECT 1059.910 1590.760 1060.230 1590.820 ;
        RECT 1003.345 1590.620 1060.230 1590.760 ;
        RECT 1003.345 1590.575 1003.635 1590.620 ;
        RECT 1059.910 1590.560 1060.230 1590.620 ;
        RECT 1058.990 1511.200 1059.310 1511.260 ;
        RECT 1059.910 1511.200 1060.230 1511.260 ;
        RECT 1058.990 1511.060 1060.230 1511.200 ;
        RECT 1058.990 1511.000 1059.310 1511.060 ;
        RECT 1059.910 1511.000 1060.230 1511.060 ;
        RECT 1058.990 1414.640 1059.310 1414.700 ;
        RECT 1059.910 1414.640 1060.230 1414.700 ;
        RECT 1058.990 1414.500 1060.230 1414.640 ;
        RECT 1058.990 1414.440 1059.310 1414.500 ;
        RECT 1059.910 1414.440 1060.230 1414.500 ;
        RECT 1058.990 1318.080 1059.310 1318.140 ;
        RECT 1059.910 1318.080 1060.230 1318.140 ;
        RECT 1058.990 1317.940 1060.230 1318.080 ;
        RECT 1058.990 1317.880 1059.310 1317.940 ;
        RECT 1059.910 1317.880 1060.230 1317.940 ;
        RECT 1058.990 1221.520 1059.310 1221.580 ;
        RECT 1059.910 1221.520 1060.230 1221.580 ;
        RECT 1058.990 1221.380 1060.230 1221.520 ;
        RECT 1058.990 1221.320 1059.310 1221.380 ;
        RECT 1059.910 1221.320 1060.230 1221.380 ;
        RECT 1058.990 1124.960 1059.310 1125.020 ;
        RECT 1059.910 1124.960 1060.230 1125.020 ;
        RECT 1058.990 1124.820 1060.230 1124.960 ;
        RECT 1058.990 1124.760 1059.310 1124.820 ;
        RECT 1059.910 1124.760 1060.230 1124.820 ;
        RECT 1058.990 1028.400 1059.310 1028.460 ;
        RECT 1059.910 1028.400 1060.230 1028.460 ;
        RECT 1058.990 1028.260 1060.230 1028.400 ;
        RECT 1058.990 1028.200 1059.310 1028.260 ;
        RECT 1059.910 1028.200 1060.230 1028.260 ;
        RECT 1058.990 931.840 1059.310 931.900 ;
        RECT 1059.910 931.840 1060.230 931.900 ;
        RECT 1058.990 931.700 1060.230 931.840 ;
        RECT 1058.990 931.640 1059.310 931.700 ;
        RECT 1059.910 931.640 1060.230 931.700 ;
        RECT 1058.530 869.620 1058.850 869.680 ;
        RECT 1059.910 869.620 1060.230 869.680 ;
        RECT 1058.530 869.480 1060.230 869.620 ;
        RECT 1058.530 869.420 1058.850 869.480 ;
        RECT 1059.910 869.420 1060.230 869.480 ;
        RECT 1058.990 835.280 1059.310 835.340 ;
        RECT 1059.910 835.280 1060.230 835.340 ;
        RECT 1058.990 835.140 1060.230 835.280 ;
        RECT 1058.990 835.080 1059.310 835.140 ;
        RECT 1059.910 835.080 1060.230 835.140 ;
        RECT 1059.450 821.000 1059.770 821.060 ;
        RECT 1059.255 820.860 1059.770 821.000 ;
        RECT 1059.450 820.800 1059.770 820.860 ;
        RECT 1059.450 786.660 1059.770 786.720 ;
        RECT 1059.255 786.520 1059.770 786.660 ;
        RECT 1059.450 786.460 1059.770 786.520 ;
        RECT 1058.990 738.380 1059.310 738.440 ;
        RECT 1059.910 738.380 1060.230 738.440 ;
        RECT 1058.990 738.240 1060.230 738.380 ;
        RECT 1058.990 738.180 1059.310 738.240 ;
        RECT 1059.910 738.180 1060.230 738.240 ;
        RECT 1059.450 724.440 1059.770 724.500 ;
        RECT 1059.255 724.300 1059.770 724.440 ;
        RECT 1059.450 724.240 1059.770 724.300 ;
        RECT 1059.450 689.760 1059.770 689.820 ;
        RECT 1059.255 689.620 1059.770 689.760 ;
        RECT 1059.450 689.560 1059.770 689.620 ;
        RECT 1058.990 641.820 1059.310 641.880 ;
        RECT 1059.910 641.820 1060.230 641.880 ;
        RECT 1058.990 641.680 1060.230 641.820 ;
        RECT 1058.990 641.620 1059.310 641.680 ;
        RECT 1059.910 641.620 1060.230 641.680 ;
        RECT 1059.450 627.880 1059.770 627.940 ;
        RECT 1059.255 627.740 1059.770 627.880 ;
        RECT 1059.450 627.680 1059.770 627.740 ;
        RECT 1059.450 593.200 1059.770 593.260 ;
        RECT 1059.255 593.060 1059.770 593.200 ;
        RECT 1059.450 593.000 1059.770 593.060 ;
        RECT 1058.990 545.260 1059.310 545.320 ;
        RECT 1059.910 545.260 1060.230 545.320 ;
        RECT 1058.990 545.120 1060.230 545.260 ;
        RECT 1058.990 545.060 1059.310 545.120 ;
        RECT 1059.910 545.060 1060.230 545.120 ;
        RECT 1059.450 531.320 1059.770 531.380 ;
        RECT 1059.255 531.180 1059.770 531.320 ;
        RECT 1059.450 531.120 1059.770 531.180 ;
        RECT 1059.450 496.640 1059.770 496.700 ;
        RECT 1059.255 496.500 1059.770 496.640 ;
        RECT 1059.450 496.440 1059.770 496.500 ;
        RECT 1058.990 448.700 1059.310 448.760 ;
        RECT 1059.910 448.700 1060.230 448.760 ;
        RECT 1058.990 448.560 1060.230 448.700 ;
        RECT 1058.990 448.500 1059.310 448.560 ;
        RECT 1059.910 448.500 1060.230 448.560 ;
        RECT 1059.450 434.760 1059.770 434.820 ;
        RECT 1059.255 434.620 1059.770 434.760 ;
        RECT 1059.450 434.560 1059.770 434.620 ;
        RECT 1059.465 386.480 1059.755 386.525 ;
        RECT 1059.910 386.480 1060.230 386.540 ;
        RECT 1059.465 386.340 1060.230 386.480 ;
        RECT 1059.465 386.295 1059.755 386.340 ;
        RECT 1059.910 386.280 1060.230 386.340 ;
        RECT 1059.465 379.340 1059.755 379.385 ;
        RECT 1059.910 379.340 1060.230 379.400 ;
        RECT 1059.465 379.200 1060.230 379.340 ;
        RECT 1059.465 379.155 1059.755 379.200 ;
        RECT 1059.910 379.140 1060.230 379.200 ;
        RECT 1059.450 351.800 1059.770 351.860 ;
        RECT 1059.255 351.660 1059.770 351.800 ;
        RECT 1059.450 351.600 1059.770 351.660 ;
        RECT 1059.465 289.580 1059.755 289.625 ;
        RECT 1059.910 289.580 1060.230 289.640 ;
        RECT 1059.465 289.440 1060.230 289.580 ;
        RECT 1059.465 289.395 1059.755 289.440 ;
        RECT 1059.910 289.380 1060.230 289.440 ;
        RECT 1059.450 253.540 1059.770 253.600 ;
        RECT 1059.255 253.400 1059.770 253.540 ;
        RECT 1059.450 253.340 1059.770 253.400 ;
        RECT 1059.465 193.020 1059.755 193.065 ;
        RECT 1059.910 193.020 1060.230 193.080 ;
        RECT 1059.465 192.880 1060.230 193.020 ;
        RECT 1059.465 192.835 1059.755 192.880 ;
        RECT 1059.910 192.820 1060.230 192.880 ;
        RECT 1059.450 145.080 1059.770 145.140 ;
        RECT 1059.255 144.940 1059.770 145.080 ;
        RECT 1059.450 144.880 1059.770 144.940 ;
        RECT 1274.285 25.400 1274.575 25.445 ;
        RECT 1323.030 25.400 1323.350 25.460 ;
        RECT 1274.285 25.260 1323.350 25.400 ;
        RECT 1274.285 25.215 1274.575 25.260 ;
        RECT 1323.030 25.200 1323.350 25.260 ;
        RECT 1076.025 24.040 1076.315 24.085 ;
        RECT 1076.945 24.040 1077.235 24.085 ;
        RECT 1274.285 24.040 1274.575 24.085 ;
        RECT 1076.025 23.900 1077.235 24.040 ;
        RECT 1076.025 23.855 1076.315 23.900 ;
        RECT 1076.945 23.855 1077.235 23.900 ;
        RECT 1244.920 23.900 1274.575 24.040 ;
        RECT 1077.405 23.700 1077.695 23.745 ;
        RECT 1077.405 23.560 1096.020 23.700 ;
        RECT 1077.405 23.515 1077.695 23.560 ;
        RECT 1095.880 23.405 1096.020 23.560 ;
        RECT 1095.805 23.175 1096.095 23.405 ;
        RECT 1095.805 22.680 1096.095 22.725 ;
        RECT 1148.245 22.680 1148.535 22.725 ;
        RECT 1095.805 22.540 1148.535 22.680 ;
        RECT 1095.805 22.495 1096.095 22.540 ;
        RECT 1148.245 22.495 1148.535 22.540 ;
        RECT 1197.005 22.680 1197.295 22.725 ;
        RECT 1244.920 22.680 1245.060 23.900 ;
        RECT 1274.285 23.855 1274.575 23.900 ;
        RECT 1197.005 22.540 1245.060 22.680 ;
        RECT 1197.005 22.495 1197.295 22.540 ;
        RECT 1058.990 22.340 1059.310 22.400 ;
        RECT 1076.025 22.340 1076.315 22.385 ;
        RECT 1058.990 22.200 1076.315 22.340 ;
        RECT 1058.990 22.140 1059.310 22.200 ;
        RECT 1076.025 22.155 1076.315 22.200 ;
        RECT 1148.245 20.980 1148.535 21.025 ;
        RECT 1197.005 20.980 1197.295 21.025 ;
        RECT 1148.245 20.840 1197.295 20.980 ;
        RECT 1148.245 20.795 1148.535 20.840 ;
        RECT 1197.005 20.795 1197.295 20.840 ;
      LAYER via ;
        RECT 808.320 1592.260 808.580 1592.520 ;
        RECT 1059.940 1590.560 1060.200 1590.820 ;
        RECT 1059.020 1511.000 1059.280 1511.260 ;
        RECT 1059.940 1511.000 1060.200 1511.260 ;
        RECT 1059.020 1414.440 1059.280 1414.700 ;
        RECT 1059.940 1414.440 1060.200 1414.700 ;
        RECT 1059.020 1317.880 1059.280 1318.140 ;
        RECT 1059.940 1317.880 1060.200 1318.140 ;
        RECT 1059.020 1221.320 1059.280 1221.580 ;
        RECT 1059.940 1221.320 1060.200 1221.580 ;
        RECT 1059.020 1124.760 1059.280 1125.020 ;
        RECT 1059.940 1124.760 1060.200 1125.020 ;
        RECT 1059.020 1028.200 1059.280 1028.460 ;
        RECT 1059.940 1028.200 1060.200 1028.460 ;
        RECT 1059.020 931.640 1059.280 931.900 ;
        RECT 1059.940 931.640 1060.200 931.900 ;
        RECT 1058.560 869.420 1058.820 869.680 ;
        RECT 1059.940 869.420 1060.200 869.680 ;
        RECT 1059.020 835.080 1059.280 835.340 ;
        RECT 1059.940 835.080 1060.200 835.340 ;
        RECT 1059.480 820.800 1059.740 821.060 ;
        RECT 1059.480 786.460 1059.740 786.720 ;
        RECT 1059.020 738.180 1059.280 738.440 ;
        RECT 1059.940 738.180 1060.200 738.440 ;
        RECT 1059.480 724.240 1059.740 724.500 ;
        RECT 1059.480 689.560 1059.740 689.820 ;
        RECT 1059.020 641.620 1059.280 641.880 ;
        RECT 1059.940 641.620 1060.200 641.880 ;
        RECT 1059.480 627.680 1059.740 627.940 ;
        RECT 1059.480 593.000 1059.740 593.260 ;
        RECT 1059.020 545.060 1059.280 545.320 ;
        RECT 1059.940 545.060 1060.200 545.320 ;
        RECT 1059.480 531.120 1059.740 531.380 ;
        RECT 1059.480 496.440 1059.740 496.700 ;
        RECT 1059.020 448.500 1059.280 448.760 ;
        RECT 1059.940 448.500 1060.200 448.760 ;
        RECT 1059.480 434.560 1059.740 434.820 ;
        RECT 1059.940 386.280 1060.200 386.540 ;
        RECT 1059.940 379.140 1060.200 379.400 ;
        RECT 1059.480 351.600 1059.740 351.860 ;
        RECT 1059.940 289.380 1060.200 289.640 ;
        RECT 1059.480 253.340 1059.740 253.600 ;
        RECT 1059.940 192.820 1060.200 193.080 ;
        RECT 1059.480 144.880 1059.740 145.140 ;
        RECT 1323.060 25.200 1323.320 25.460 ;
        RECT 1059.020 22.140 1059.280 22.400 ;
      LAYER met2 ;
        RECT 808.180 1600.380 808.460 1604.000 ;
        RECT 808.180 1600.000 808.520 1600.380 ;
        RECT 808.380 1592.550 808.520 1600.000 ;
        RECT 808.320 1592.230 808.580 1592.550 ;
        RECT 1059.940 1590.530 1060.200 1590.850 ;
        RECT 1060.000 1511.290 1060.140 1590.530 ;
        RECT 1059.020 1510.970 1059.280 1511.290 ;
        RECT 1059.940 1510.970 1060.200 1511.290 ;
        RECT 1059.080 1510.690 1059.220 1510.970 ;
        RECT 1059.080 1510.550 1059.680 1510.690 ;
        RECT 1059.540 1463.090 1059.680 1510.550 ;
        RECT 1059.540 1462.950 1060.140 1463.090 ;
        RECT 1060.000 1414.730 1060.140 1462.950 ;
        RECT 1059.020 1414.410 1059.280 1414.730 ;
        RECT 1059.940 1414.410 1060.200 1414.730 ;
        RECT 1059.080 1414.130 1059.220 1414.410 ;
        RECT 1059.080 1413.990 1059.680 1414.130 ;
        RECT 1059.540 1366.530 1059.680 1413.990 ;
        RECT 1059.540 1366.390 1060.140 1366.530 ;
        RECT 1060.000 1318.170 1060.140 1366.390 ;
        RECT 1059.020 1317.850 1059.280 1318.170 ;
        RECT 1059.940 1317.850 1060.200 1318.170 ;
        RECT 1059.080 1317.570 1059.220 1317.850 ;
        RECT 1059.080 1317.430 1059.680 1317.570 ;
        RECT 1059.540 1269.970 1059.680 1317.430 ;
        RECT 1059.540 1269.830 1060.140 1269.970 ;
        RECT 1060.000 1221.610 1060.140 1269.830 ;
        RECT 1059.020 1221.290 1059.280 1221.610 ;
        RECT 1059.940 1221.290 1060.200 1221.610 ;
        RECT 1059.080 1221.010 1059.220 1221.290 ;
        RECT 1059.080 1220.870 1059.680 1221.010 ;
        RECT 1059.540 1173.410 1059.680 1220.870 ;
        RECT 1059.540 1173.270 1060.140 1173.410 ;
        RECT 1060.000 1125.050 1060.140 1173.270 ;
        RECT 1059.020 1124.730 1059.280 1125.050 ;
        RECT 1059.940 1124.730 1060.200 1125.050 ;
        RECT 1059.080 1124.450 1059.220 1124.730 ;
        RECT 1059.080 1124.310 1059.680 1124.450 ;
        RECT 1059.540 1076.850 1059.680 1124.310 ;
        RECT 1059.540 1076.710 1060.140 1076.850 ;
        RECT 1060.000 1028.490 1060.140 1076.710 ;
        RECT 1059.020 1028.170 1059.280 1028.490 ;
        RECT 1059.940 1028.170 1060.200 1028.490 ;
        RECT 1059.080 1027.890 1059.220 1028.170 ;
        RECT 1059.080 1027.750 1059.680 1027.890 ;
        RECT 1059.540 980.290 1059.680 1027.750 ;
        RECT 1059.540 980.150 1060.140 980.290 ;
        RECT 1060.000 931.930 1060.140 980.150 ;
        RECT 1059.020 931.610 1059.280 931.930 ;
        RECT 1059.940 931.610 1060.200 931.930 ;
        RECT 1059.080 931.330 1059.220 931.610 ;
        RECT 1059.080 931.190 1059.680 931.330 ;
        RECT 1059.540 917.845 1059.680 931.190 ;
        RECT 1058.550 917.475 1058.830 917.845 ;
        RECT 1059.470 917.475 1059.750 917.845 ;
        RECT 1058.620 869.710 1058.760 917.475 ;
        RECT 1058.560 869.390 1058.820 869.710 ;
        RECT 1059.940 869.390 1060.200 869.710 ;
        RECT 1060.000 835.370 1060.140 869.390 ;
        RECT 1059.020 835.050 1059.280 835.370 ;
        RECT 1059.940 835.050 1060.200 835.370 ;
        RECT 1059.080 834.770 1059.220 835.050 ;
        RECT 1059.080 834.630 1059.680 834.770 ;
        RECT 1059.540 821.090 1059.680 834.630 ;
        RECT 1059.480 820.770 1059.740 821.090 ;
        RECT 1059.480 786.430 1059.740 786.750 ;
        RECT 1059.540 772.890 1059.680 786.430 ;
        RECT 1059.540 772.750 1060.140 772.890 ;
        RECT 1060.000 738.470 1060.140 772.750 ;
        RECT 1059.020 738.210 1059.280 738.470 ;
        RECT 1059.020 738.150 1059.680 738.210 ;
        RECT 1059.940 738.150 1060.200 738.470 ;
        RECT 1059.080 738.070 1059.680 738.150 ;
        RECT 1059.540 724.530 1059.680 738.070 ;
        RECT 1059.480 724.210 1059.740 724.530 ;
        RECT 1059.480 689.530 1059.740 689.850 ;
        RECT 1059.540 676.330 1059.680 689.530 ;
        RECT 1059.540 676.190 1060.140 676.330 ;
        RECT 1060.000 641.910 1060.140 676.190 ;
        RECT 1059.020 641.650 1059.280 641.910 ;
        RECT 1059.020 641.590 1059.680 641.650 ;
        RECT 1059.940 641.590 1060.200 641.910 ;
        RECT 1059.080 641.510 1059.680 641.590 ;
        RECT 1059.540 627.970 1059.680 641.510 ;
        RECT 1059.480 627.650 1059.740 627.970 ;
        RECT 1059.480 592.970 1059.740 593.290 ;
        RECT 1059.540 579.770 1059.680 592.970 ;
        RECT 1059.540 579.630 1060.140 579.770 ;
        RECT 1060.000 545.350 1060.140 579.630 ;
        RECT 1059.020 545.090 1059.280 545.350 ;
        RECT 1059.020 545.030 1059.680 545.090 ;
        RECT 1059.940 545.030 1060.200 545.350 ;
        RECT 1059.080 544.950 1059.680 545.030 ;
        RECT 1059.540 531.410 1059.680 544.950 ;
        RECT 1059.480 531.090 1059.740 531.410 ;
        RECT 1059.480 496.410 1059.740 496.730 ;
        RECT 1059.540 483.210 1059.680 496.410 ;
        RECT 1059.540 483.070 1060.140 483.210 ;
        RECT 1060.000 448.790 1060.140 483.070 ;
        RECT 1059.020 448.530 1059.280 448.790 ;
        RECT 1059.020 448.470 1059.680 448.530 ;
        RECT 1059.940 448.470 1060.200 448.790 ;
        RECT 1059.080 448.390 1059.680 448.470 ;
        RECT 1059.540 434.850 1059.680 448.390 ;
        RECT 1059.480 434.530 1059.740 434.850 ;
        RECT 1059.940 386.250 1060.200 386.570 ;
        RECT 1060.000 379.430 1060.140 386.250 ;
        RECT 1059.940 379.110 1060.200 379.430 ;
        RECT 1059.480 351.570 1059.740 351.890 ;
        RECT 1059.540 303.690 1059.680 351.570 ;
        RECT 1059.540 303.550 1060.140 303.690 ;
        RECT 1060.000 289.670 1060.140 303.550 ;
        RECT 1059.940 289.350 1060.200 289.670 ;
        RECT 1059.480 253.310 1059.740 253.630 ;
        RECT 1059.540 207.130 1059.680 253.310 ;
        RECT 1059.540 206.990 1060.140 207.130 ;
        RECT 1060.000 193.110 1060.140 206.990 ;
        RECT 1059.940 192.790 1060.200 193.110 ;
        RECT 1059.480 144.850 1059.740 145.170 ;
        RECT 1059.540 110.570 1059.680 144.850 ;
        RECT 1059.540 110.430 1060.140 110.570 ;
        RECT 1060.000 62.290 1060.140 110.430 ;
        RECT 1059.080 62.150 1060.140 62.290 ;
        RECT 1059.080 22.430 1059.220 62.150 ;
        RECT 1323.060 25.170 1323.320 25.490 ;
        RECT 1059.020 22.110 1059.280 22.430 ;
        RECT 1323.120 2.400 1323.260 25.170 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
      LAYER via2 ;
        RECT 1058.550 917.520 1058.830 917.800 ;
        RECT 1059.470 917.520 1059.750 917.800 ;
      LAYER met3 ;
        RECT 1058.525 917.810 1058.855 917.825 ;
        RECT 1059.445 917.810 1059.775 917.825 ;
        RECT 1058.525 917.510 1059.775 917.810 ;
        RECT 1058.525 917.495 1058.855 917.510 ;
        RECT 1059.445 917.495 1059.775 917.510 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1290.445 24.565 1291.535 24.735 ;
        RECT 1290.445 24.225 1290.615 24.565 ;
        RECT 1095.405 23.545 1096.955 23.715 ;
        RECT 1095.405 22.525 1095.575 23.545 ;
        RECT 1115.185 22.865 1115.355 23.715 ;
        RECT 1148.765 22.865 1148.935 24.055 ;
      LAYER mcon ;
        RECT 1291.365 24.565 1291.535 24.735 ;
        RECT 1148.765 23.885 1148.935 24.055 ;
        RECT 1096.785 23.545 1096.955 23.715 ;
        RECT 1115.185 23.545 1115.355 23.715 ;
      LAYER met1 ;
        RECT 821.170 1593.620 821.490 1593.880 ;
        RECT 834.970 1593.820 835.290 1593.880 ;
        RECT 834.970 1593.680 956.180 1593.820 ;
        RECT 834.970 1593.620 835.290 1593.680 ;
        RECT 820.710 1593.480 821.030 1593.540 ;
        RECT 821.260 1593.480 821.400 1593.620 ;
        RECT 820.710 1593.340 821.400 1593.480 ;
        RECT 820.710 1593.280 821.030 1593.340 ;
        RECT 814.730 1593.140 815.050 1593.200 ;
        RECT 820.250 1593.140 820.570 1593.200 ;
        RECT 814.730 1593.000 820.570 1593.140 ;
        RECT 814.730 1592.940 815.050 1593.000 ;
        RECT 820.250 1592.940 820.570 1593.000 ;
        RECT 956.040 1592.800 956.180 1593.680 ;
        RECT 956.040 1592.660 1004.020 1592.800 ;
        RECT 1003.880 1592.460 1004.020 1592.660 ;
        RECT 1079.690 1592.460 1080.010 1592.520 ;
        RECT 1003.880 1592.320 1080.010 1592.460 ;
        RECT 1079.690 1592.260 1080.010 1592.320 ;
        RECT 1291.305 24.720 1291.595 24.765 ;
        RECT 1340.510 24.720 1340.830 24.780 ;
        RECT 1291.305 24.580 1340.830 24.720 ;
        RECT 1291.305 24.535 1291.595 24.580 ;
        RECT 1340.510 24.520 1340.830 24.580 ;
        RECT 1290.385 24.380 1290.675 24.425 ;
        RECT 1244.460 24.240 1290.675 24.380 ;
        RECT 1148.705 24.040 1148.995 24.085 ;
        RECT 1148.705 23.900 1195.380 24.040 ;
        RECT 1148.705 23.855 1148.995 23.900 ;
        RECT 1096.725 23.700 1097.015 23.745 ;
        RECT 1115.125 23.700 1115.415 23.745 ;
        RECT 1096.725 23.560 1115.415 23.700 ;
        RECT 1096.725 23.515 1097.015 23.560 ;
        RECT 1115.125 23.515 1115.415 23.560 ;
        RECT 1115.125 23.020 1115.415 23.065 ;
        RECT 1148.705 23.020 1148.995 23.065 ;
        RECT 1115.125 22.880 1148.995 23.020 ;
        RECT 1195.240 23.020 1195.380 23.900 ;
        RECT 1244.460 23.020 1244.600 24.240 ;
        RECT 1290.385 24.195 1290.675 24.240 ;
        RECT 1195.240 22.880 1244.600 23.020 ;
        RECT 1115.125 22.835 1115.415 22.880 ;
        RECT 1148.705 22.835 1148.995 22.880 ;
        RECT 1080.150 22.680 1080.470 22.740 ;
        RECT 1095.345 22.680 1095.635 22.725 ;
        RECT 1080.150 22.540 1095.635 22.680 ;
        RECT 1080.150 22.480 1080.470 22.540 ;
        RECT 1095.345 22.495 1095.635 22.540 ;
      LAYER via ;
        RECT 821.200 1593.620 821.460 1593.880 ;
        RECT 835.000 1593.620 835.260 1593.880 ;
        RECT 820.740 1593.280 821.000 1593.540 ;
        RECT 814.760 1592.940 815.020 1593.200 ;
        RECT 820.280 1592.940 820.540 1593.200 ;
        RECT 1079.720 1592.260 1079.980 1592.520 ;
        RECT 1340.540 24.520 1340.800 24.780 ;
        RECT 1080.180 22.480 1080.440 22.740 ;
      LAYER met2 ;
        RECT 814.620 1600.380 814.900 1604.000 ;
        RECT 814.620 1600.000 814.960 1600.380 ;
        RECT 814.820 1593.230 814.960 1600.000 ;
        RECT 821.200 1593.765 821.460 1593.910 ;
        RECT 835.000 1593.765 835.260 1593.910 ;
        RECT 820.740 1593.250 821.000 1593.570 ;
        RECT 821.190 1593.395 821.470 1593.765 ;
        RECT 834.990 1593.395 835.270 1593.765 ;
        RECT 814.760 1592.910 815.020 1593.230 ;
        RECT 820.280 1592.970 820.540 1593.230 ;
        RECT 820.800 1592.970 820.940 1593.250 ;
        RECT 820.280 1592.910 820.940 1592.970 ;
        RECT 820.340 1592.830 820.940 1592.910 ;
        RECT 1079.720 1592.230 1079.980 1592.550 ;
        RECT 1079.780 22.680 1079.920 1592.230 ;
        RECT 1340.540 24.490 1340.800 24.810 ;
        RECT 1080.180 22.680 1080.440 22.770 ;
        RECT 1079.780 22.540 1080.440 22.680 ;
        RECT 1080.180 22.450 1080.440 22.540 ;
        RECT 1340.600 2.400 1340.740 24.490 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
      LAYER via2 ;
        RECT 821.190 1593.440 821.470 1593.720 ;
        RECT 834.990 1593.440 835.270 1593.720 ;
      LAYER met3 ;
        RECT 821.165 1593.730 821.495 1593.745 ;
        RECT 834.965 1593.730 835.295 1593.745 ;
        RECT 821.165 1593.430 835.295 1593.730 ;
        RECT 821.165 1593.415 821.495 1593.430 ;
        RECT 834.965 1593.415 835.295 1593.430 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 592.090 1593.820 592.410 1593.880 ;
        RECT 665.690 1593.820 666.010 1593.880 ;
        RECT 592.090 1593.680 666.010 1593.820 ;
        RECT 592.090 1593.620 592.410 1593.680 ;
        RECT 665.690 1593.620 666.010 1593.680 ;
        RECT 665.690 17.240 666.010 17.300 ;
        RECT 698.350 17.240 698.670 17.300 ;
        RECT 665.690 17.100 698.670 17.240 ;
        RECT 665.690 17.040 666.010 17.100 ;
        RECT 698.350 17.040 698.670 17.100 ;
      LAYER via ;
        RECT 592.120 1593.620 592.380 1593.880 ;
        RECT 665.720 1593.620 665.980 1593.880 ;
        RECT 665.720 17.040 665.980 17.300 ;
        RECT 698.380 17.040 698.640 17.300 ;
      LAYER met2 ;
        RECT 591.980 1600.380 592.260 1604.000 ;
        RECT 591.980 1600.000 592.320 1600.380 ;
        RECT 592.180 1593.910 592.320 1600.000 ;
        RECT 592.120 1593.590 592.380 1593.910 ;
        RECT 665.720 1593.590 665.980 1593.910 ;
        RECT 665.780 17.330 665.920 1593.590 ;
        RECT 665.720 17.010 665.980 17.330 ;
        RECT 698.380 17.010 698.640 17.330 ;
        RECT 698.440 2.400 698.580 17.010 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1287.685 23.885 1287.855 24.735 ;
        RECT 1196.145 22.185 1196.315 23.375 ;
      LAYER mcon ;
        RECT 1287.685 24.565 1287.855 24.735 ;
        RECT 1196.145 23.205 1196.315 23.375 ;
      LAYER met1 ;
        RECT 819.790 1591.100 820.110 1591.160 ;
        RECT 1093.490 1591.100 1093.810 1591.160 ;
        RECT 819.790 1590.960 1093.810 1591.100 ;
        RECT 819.790 1590.900 820.110 1590.960 ;
        RECT 1093.490 1590.900 1093.810 1590.960 ;
        RECT 1093.490 39.680 1093.810 39.740 ;
        RECT 1096.250 39.680 1096.570 39.740 ;
        RECT 1093.490 39.540 1096.570 39.680 ;
        RECT 1093.490 39.480 1093.810 39.540 ;
        RECT 1096.250 39.480 1096.570 39.540 ;
        RECT 1287.625 24.720 1287.915 24.765 ;
        RECT 1244.000 24.580 1287.915 24.720 ;
        RECT 1125.320 23.560 1149.380 23.700 ;
        RECT 1096.250 23.360 1096.570 23.420 ;
        RECT 1125.320 23.360 1125.460 23.560 ;
        RECT 1096.250 23.220 1125.460 23.360 ;
        RECT 1096.250 23.160 1096.570 23.220 ;
        RECT 1149.240 22.680 1149.380 23.560 ;
        RECT 1196.085 23.360 1196.375 23.405 ;
        RECT 1244.000 23.360 1244.140 24.580 ;
        RECT 1287.625 24.535 1287.915 24.580 ;
        RECT 1287.625 24.040 1287.915 24.085 ;
        RECT 1358.450 24.040 1358.770 24.100 ;
        RECT 1287.625 23.900 1358.770 24.040 ;
        RECT 1287.625 23.855 1287.915 23.900 ;
        RECT 1358.450 23.840 1358.770 23.900 ;
        RECT 1196.085 23.220 1244.140 23.360 ;
        RECT 1196.085 23.175 1196.375 23.220 ;
        RECT 1149.240 22.540 1172.840 22.680 ;
        RECT 1172.700 22.340 1172.840 22.540 ;
        RECT 1196.085 22.340 1196.375 22.385 ;
        RECT 1172.700 22.200 1196.375 22.340 ;
        RECT 1196.085 22.155 1196.375 22.200 ;
      LAYER via ;
        RECT 819.820 1590.900 820.080 1591.160 ;
        RECT 1093.520 1590.900 1093.780 1591.160 ;
        RECT 1093.520 39.480 1093.780 39.740 ;
        RECT 1096.280 39.480 1096.540 39.740 ;
        RECT 1096.280 23.160 1096.540 23.420 ;
        RECT 1358.480 23.840 1358.740 24.100 ;
      LAYER met2 ;
        RECT 820.600 1601.130 820.880 1604.000 ;
        RECT 819.880 1600.990 820.880 1601.130 ;
        RECT 819.880 1597.050 820.020 1600.990 ;
        RECT 820.600 1600.000 820.880 1600.990 ;
        RECT 819.880 1596.910 820.480 1597.050 ;
        RECT 820.340 1593.650 820.480 1596.910 ;
        RECT 819.880 1593.510 820.480 1593.650 ;
        RECT 819.880 1591.190 820.020 1593.510 ;
        RECT 819.820 1590.870 820.080 1591.190 ;
        RECT 1093.520 1590.870 1093.780 1591.190 ;
        RECT 1093.580 39.770 1093.720 1590.870 ;
        RECT 1093.520 39.450 1093.780 39.770 ;
        RECT 1096.280 39.450 1096.540 39.770 ;
        RECT 1096.340 23.450 1096.480 39.450 ;
        RECT 1358.480 23.810 1358.740 24.130 ;
        RECT 1096.280 23.130 1096.540 23.450 ;
        RECT 1358.540 2.400 1358.680 23.810 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 827.150 55.660 827.470 55.720 ;
        RECT 1373.170 55.660 1373.490 55.720 ;
        RECT 827.150 55.520 1373.490 55.660 ;
        RECT 827.150 55.460 827.470 55.520 ;
        RECT 1373.170 55.460 1373.490 55.520 ;
        RECT 1373.170 2.960 1373.490 3.020 ;
        RECT 1376.390 2.960 1376.710 3.020 ;
        RECT 1373.170 2.820 1376.710 2.960 ;
        RECT 1373.170 2.760 1373.490 2.820 ;
        RECT 1376.390 2.760 1376.710 2.820 ;
      LAYER via ;
        RECT 827.180 55.460 827.440 55.720 ;
        RECT 1373.200 55.460 1373.460 55.720 ;
        RECT 1373.200 2.760 1373.460 3.020 ;
        RECT 1376.420 2.760 1376.680 3.020 ;
      LAYER met2 ;
        RECT 827.040 1600.380 827.320 1604.000 ;
        RECT 827.040 1600.000 827.380 1600.380 ;
        RECT 827.240 55.750 827.380 1600.000 ;
        RECT 827.180 55.430 827.440 55.750 ;
        RECT 1373.200 55.430 1373.460 55.750 ;
        RECT 1373.260 3.050 1373.400 55.430 ;
        RECT 1373.200 2.730 1373.460 3.050 ;
        RECT 1376.420 2.730 1376.680 3.050 ;
        RECT 1376.480 2.400 1376.620 2.730 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 833.590 70.280 833.910 70.340 ;
        RECT 1394.330 70.280 1394.650 70.340 ;
        RECT 833.590 70.140 1394.650 70.280 ;
        RECT 833.590 70.080 833.910 70.140 ;
        RECT 1394.330 70.080 1394.650 70.140 ;
      LAYER via ;
        RECT 833.620 70.080 833.880 70.340 ;
        RECT 1394.360 70.080 1394.620 70.340 ;
      LAYER met2 ;
        RECT 833.020 1600.450 833.300 1604.000 ;
        RECT 833.020 1600.310 833.820 1600.450 ;
        RECT 833.020 1600.000 833.300 1600.310 ;
        RECT 833.680 70.370 833.820 1600.310 ;
        RECT 833.620 70.050 833.880 70.370 ;
        RECT 1394.360 70.050 1394.620 70.370 ;
        RECT 1394.420 2.400 1394.560 70.050 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.030 70.620 840.350 70.680 ;
        RECT 1407.670 70.620 1407.990 70.680 ;
        RECT 840.030 70.480 1407.990 70.620 ;
        RECT 840.030 70.420 840.350 70.480 ;
        RECT 1407.670 70.420 1407.990 70.480 ;
        RECT 1407.670 2.960 1407.990 3.020 ;
        RECT 1412.270 2.960 1412.590 3.020 ;
        RECT 1407.670 2.820 1412.590 2.960 ;
        RECT 1407.670 2.760 1407.990 2.820 ;
        RECT 1412.270 2.760 1412.590 2.820 ;
      LAYER via ;
        RECT 840.060 70.420 840.320 70.680 ;
        RECT 1407.700 70.420 1407.960 70.680 ;
        RECT 1407.700 2.760 1407.960 3.020 ;
        RECT 1412.300 2.760 1412.560 3.020 ;
      LAYER met2 ;
        RECT 839.460 1600.450 839.740 1604.000 ;
        RECT 839.460 1600.310 840.260 1600.450 ;
        RECT 839.460 1600.000 839.740 1600.310 ;
        RECT 840.120 70.710 840.260 1600.310 ;
        RECT 840.060 70.390 840.320 70.710 ;
        RECT 1407.700 70.390 1407.960 70.710 ;
        RECT 1407.760 3.050 1407.900 70.390 ;
        RECT 1407.700 2.730 1407.960 3.050 ;
        RECT 1412.300 2.730 1412.560 3.050 ;
        RECT 1412.360 2.400 1412.500 2.730 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 847.390 82.180 847.710 82.240 ;
        RECT 1428.370 82.180 1428.690 82.240 ;
        RECT 847.390 82.040 1428.690 82.180 ;
        RECT 847.390 81.980 847.710 82.040 ;
        RECT 1428.370 81.980 1428.690 82.040 ;
        RECT 1428.370 2.960 1428.690 3.020 ;
        RECT 1429.750 2.960 1430.070 3.020 ;
        RECT 1428.370 2.820 1430.070 2.960 ;
        RECT 1428.370 2.760 1428.690 2.820 ;
        RECT 1429.750 2.760 1430.070 2.820 ;
      LAYER via ;
        RECT 847.420 81.980 847.680 82.240 ;
        RECT 1428.400 81.980 1428.660 82.240 ;
        RECT 1428.400 2.760 1428.660 3.020 ;
        RECT 1429.780 2.760 1430.040 3.020 ;
      LAYER met2 ;
        RECT 845.440 1600.450 845.720 1604.000 ;
        RECT 845.440 1600.310 846.700 1600.450 ;
        RECT 845.440 1600.000 845.720 1600.310 ;
        RECT 846.560 1580.050 846.700 1600.310 ;
        RECT 846.560 1579.910 847.620 1580.050 ;
        RECT 847.480 82.270 847.620 1579.910 ;
        RECT 847.420 81.950 847.680 82.270 ;
        RECT 1428.400 81.950 1428.660 82.270 ;
        RECT 1428.460 3.050 1428.600 81.950 ;
        RECT 1428.400 2.730 1428.660 3.050 ;
        RECT 1429.780 2.730 1430.040 3.050 ;
        RECT 1429.840 2.400 1429.980 2.730 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 854.290 81.840 854.610 81.900 ;
        RECT 1442.170 81.840 1442.490 81.900 ;
        RECT 854.290 81.700 1442.490 81.840 ;
        RECT 854.290 81.640 854.610 81.700 ;
        RECT 1442.170 81.640 1442.490 81.700 ;
        RECT 1442.170 2.960 1442.490 3.020 ;
        RECT 1447.690 2.960 1448.010 3.020 ;
        RECT 1442.170 2.820 1448.010 2.960 ;
        RECT 1442.170 2.760 1442.490 2.820 ;
        RECT 1447.690 2.760 1448.010 2.820 ;
      LAYER via ;
        RECT 854.320 81.640 854.580 81.900 ;
        RECT 1442.200 81.640 1442.460 81.900 ;
        RECT 1442.200 2.760 1442.460 3.020 ;
        RECT 1447.720 2.760 1447.980 3.020 ;
      LAYER met2 ;
        RECT 851.880 1600.450 852.160 1604.000 ;
        RECT 851.880 1600.310 852.680 1600.450 ;
        RECT 851.880 1600.000 852.160 1600.310 ;
        RECT 852.540 1580.050 852.680 1600.310 ;
        RECT 852.540 1579.910 854.520 1580.050 ;
        RECT 854.380 81.930 854.520 1579.910 ;
        RECT 854.320 81.610 854.580 81.930 ;
        RECT 1442.200 81.610 1442.460 81.930 ;
        RECT 1442.260 3.050 1442.400 81.610 ;
        RECT 1442.200 2.730 1442.460 3.050 ;
        RECT 1447.720 2.730 1447.980 3.050 ;
        RECT 1447.780 2.400 1447.920 2.730 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 857.970 1588.040 858.290 1588.100 ;
        RECT 860.730 1588.040 861.050 1588.100 ;
        RECT 857.970 1587.900 861.050 1588.040 ;
        RECT 857.970 1587.840 858.290 1587.900 ;
        RECT 860.730 1587.840 861.050 1587.900 ;
        RECT 860.730 81.500 861.050 81.560 ;
        RECT 1462.870 81.500 1463.190 81.560 ;
        RECT 860.730 81.360 1463.190 81.500 ;
        RECT 860.730 81.300 861.050 81.360 ;
        RECT 1462.870 81.300 1463.190 81.360 ;
        RECT 1462.870 2.960 1463.190 3.020 ;
        RECT 1465.630 2.960 1465.950 3.020 ;
        RECT 1462.870 2.820 1465.950 2.960 ;
        RECT 1462.870 2.760 1463.190 2.820 ;
        RECT 1465.630 2.760 1465.950 2.820 ;
      LAYER via ;
        RECT 858.000 1587.840 858.260 1588.100 ;
        RECT 860.760 1587.840 861.020 1588.100 ;
        RECT 860.760 81.300 861.020 81.560 ;
        RECT 1462.900 81.300 1463.160 81.560 ;
        RECT 1462.900 2.760 1463.160 3.020 ;
        RECT 1465.660 2.760 1465.920 3.020 ;
      LAYER met2 ;
        RECT 857.860 1600.380 858.140 1604.000 ;
        RECT 857.860 1600.000 858.200 1600.380 ;
        RECT 858.060 1588.130 858.200 1600.000 ;
        RECT 858.000 1587.810 858.260 1588.130 ;
        RECT 860.760 1587.810 861.020 1588.130 ;
        RECT 860.820 81.590 860.960 1587.810 ;
        RECT 860.760 81.270 861.020 81.590 ;
        RECT 1462.900 81.270 1463.160 81.590 ;
        RECT 1462.960 3.050 1463.100 81.270 ;
        RECT 1462.900 2.730 1463.160 3.050 ;
        RECT 1465.660 2.730 1465.920 3.050 ;
        RECT 1465.720 2.400 1465.860 2.730 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 863.950 1587.360 864.270 1587.420 ;
        RECT 868.090 1587.360 868.410 1587.420 ;
        RECT 863.950 1587.220 868.410 1587.360 ;
        RECT 863.950 1587.160 864.270 1587.220 ;
        RECT 868.090 1587.160 868.410 1587.220 ;
        RECT 868.090 81.160 868.410 81.220 ;
        RECT 1483.570 81.160 1483.890 81.220 ;
        RECT 868.090 81.020 1483.890 81.160 ;
        RECT 868.090 80.960 868.410 81.020 ;
        RECT 1483.570 80.960 1483.890 81.020 ;
      LAYER via ;
        RECT 863.980 1587.160 864.240 1587.420 ;
        RECT 868.120 1587.160 868.380 1587.420 ;
        RECT 868.120 80.960 868.380 81.220 ;
        RECT 1483.600 80.960 1483.860 81.220 ;
      LAYER met2 ;
        RECT 863.840 1600.380 864.120 1604.000 ;
        RECT 863.840 1600.000 864.180 1600.380 ;
        RECT 864.040 1587.450 864.180 1600.000 ;
        RECT 863.980 1587.130 864.240 1587.450 ;
        RECT 868.120 1587.130 868.380 1587.450 ;
        RECT 868.180 81.250 868.320 1587.130 ;
        RECT 868.120 80.930 868.380 81.250 ;
        RECT 1483.600 80.930 1483.860 81.250 ;
        RECT 1483.660 2.400 1483.800 80.930 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 870.390 1587.700 870.710 1587.760 ;
        RECT 875.910 1587.700 876.230 1587.760 ;
        RECT 870.390 1587.560 876.230 1587.700 ;
        RECT 870.390 1587.500 870.710 1587.560 ;
        RECT 875.910 1587.500 876.230 1587.560 ;
        RECT 875.910 16.560 876.230 16.620 ;
        RECT 1501.510 16.560 1501.830 16.620 ;
        RECT 875.910 16.420 1501.830 16.560 ;
        RECT 875.910 16.360 876.230 16.420 ;
        RECT 1501.510 16.360 1501.830 16.420 ;
      LAYER via ;
        RECT 870.420 1587.500 870.680 1587.760 ;
        RECT 875.940 1587.500 876.200 1587.760 ;
        RECT 875.940 16.360 876.200 16.620 ;
        RECT 1501.540 16.360 1501.800 16.620 ;
      LAYER met2 ;
        RECT 870.280 1600.380 870.560 1604.000 ;
        RECT 870.280 1600.000 870.620 1600.380 ;
        RECT 870.480 1587.790 870.620 1600.000 ;
        RECT 870.420 1587.470 870.680 1587.790 ;
        RECT 875.940 1587.470 876.200 1587.790 ;
        RECT 876.000 16.650 876.140 1587.470 ;
        RECT 875.940 16.330 876.200 16.650 ;
        RECT 1501.540 16.330 1501.800 16.650 ;
        RECT 1501.600 2.400 1501.740 16.330 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 876.370 1587.360 876.690 1587.420 ;
        RECT 881.430 1587.360 881.750 1587.420 ;
        RECT 876.370 1587.220 881.750 1587.360 ;
        RECT 876.370 1587.160 876.690 1587.220 ;
        RECT 881.430 1587.160 881.750 1587.220 ;
        RECT 881.430 80.820 881.750 80.880 ;
        RECT 1518.070 80.820 1518.390 80.880 ;
        RECT 881.430 80.680 1518.390 80.820 ;
        RECT 881.430 80.620 881.750 80.680 ;
        RECT 1518.070 80.620 1518.390 80.680 ;
        RECT 1518.070 2.960 1518.390 3.020 ;
        RECT 1518.990 2.960 1519.310 3.020 ;
        RECT 1518.070 2.820 1519.310 2.960 ;
        RECT 1518.070 2.760 1518.390 2.820 ;
        RECT 1518.990 2.760 1519.310 2.820 ;
      LAYER via ;
        RECT 876.400 1587.160 876.660 1587.420 ;
        RECT 881.460 1587.160 881.720 1587.420 ;
        RECT 881.460 80.620 881.720 80.880 ;
        RECT 1518.100 80.620 1518.360 80.880 ;
        RECT 1518.100 2.760 1518.360 3.020 ;
        RECT 1519.020 2.760 1519.280 3.020 ;
      LAYER met2 ;
        RECT 876.260 1600.380 876.540 1604.000 ;
        RECT 876.260 1600.000 876.600 1600.380 ;
        RECT 876.460 1587.450 876.600 1600.000 ;
        RECT 876.400 1587.130 876.660 1587.450 ;
        RECT 881.460 1587.130 881.720 1587.450 ;
        RECT 881.520 80.910 881.660 1587.130 ;
        RECT 881.460 80.590 881.720 80.910 ;
        RECT 1518.100 80.590 1518.360 80.910 ;
        RECT 1518.160 3.050 1518.300 80.590 ;
        RECT 1518.100 2.730 1518.360 3.050 ;
        RECT 1519.020 2.730 1519.280 3.050 ;
        RECT 1519.080 2.400 1519.220 2.730 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 680.945 17.425 681.115 20.995 ;
        RECT 693.365 15.045 693.535 17.595 ;
      LAYER mcon ;
        RECT 680.945 20.825 681.115 20.995 ;
        RECT 693.365 17.425 693.535 17.595 ;
      LAYER met1 ;
        RECT 613.800 1589.940 664.080 1590.080 ;
        RECT 613.800 1589.740 613.940 1589.940 ;
        RECT 613.340 1589.600 613.940 1589.740 ;
        RECT 663.940 1589.740 664.080 1589.940 ;
        RECT 672.590 1589.740 672.910 1589.800 ;
        RECT 663.940 1589.600 672.910 1589.740 ;
        RECT 598.070 1589.400 598.390 1589.460 ;
        RECT 613.340 1589.400 613.480 1589.600 ;
        RECT 672.590 1589.540 672.910 1589.600 ;
        RECT 598.070 1589.260 613.480 1589.400 ;
        RECT 598.070 1589.200 598.390 1589.260 ;
        RECT 672.590 20.980 672.910 21.040 ;
        RECT 680.885 20.980 681.175 21.025 ;
        RECT 672.590 20.840 681.175 20.980 ;
        RECT 672.590 20.780 672.910 20.840 ;
        RECT 680.885 20.795 681.175 20.840 ;
        RECT 680.885 17.580 681.175 17.625 ;
        RECT 693.305 17.580 693.595 17.625 ;
        RECT 680.885 17.440 693.595 17.580 ;
        RECT 680.885 17.395 681.175 17.440 ;
        RECT 693.305 17.395 693.595 17.440 ;
        RECT 693.305 15.200 693.595 15.245 ;
        RECT 716.290 15.200 716.610 15.260 ;
        RECT 693.305 15.060 716.610 15.200 ;
        RECT 693.305 15.015 693.595 15.060 ;
        RECT 716.290 15.000 716.610 15.060 ;
      LAYER via ;
        RECT 598.100 1589.200 598.360 1589.460 ;
        RECT 672.620 1589.540 672.880 1589.800 ;
        RECT 672.620 20.780 672.880 21.040 ;
        RECT 716.320 15.000 716.580 15.260 ;
      LAYER met2 ;
        RECT 597.960 1600.380 598.240 1604.000 ;
        RECT 597.960 1600.000 598.300 1600.380 ;
        RECT 598.160 1589.490 598.300 1600.000 ;
        RECT 672.620 1589.510 672.880 1589.830 ;
        RECT 598.100 1589.170 598.360 1589.490 ;
        RECT 672.680 21.070 672.820 1589.510 ;
        RECT 672.620 20.750 672.880 21.070 ;
        RECT 716.320 14.970 716.580 15.290 ;
        RECT 716.380 2.400 716.520 14.970 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 966.145 41.225 966.315 43.095 ;
        RECT 980.405 41.225 980.575 42.415 ;
        RECT 1075.625 39.865 1075.795 42.415 ;
        RECT 1077.005 39.865 1077.175 42.415 ;
      LAYER mcon ;
        RECT 966.145 42.925 966.315 43.095 ;
        RECT 980.405 42.245 980.575 42.415 ;
        RECT 1075.625 42.245 1075.795 42.415 ;
        RECT 1077.005 42.245 1077.175 42.415 ;
      LAYER met1 ;
        RECT 966.085 43.080 966.375 43.125 ;
        RECT 907.280 42.940 966.375 43.080 ;
        RECT 882.350 42.400 882.670 42.460 ;
        RECT 907.280 42.400 907.420 42.940 ;
        RECT 966.085 42.895 966.375 42.940 ;
        RECT 1214.470 42.740 1214.790 42.800 ;
        RECT 1198.460 42.600 1214.790 42.740 ;
        RECT 882.350 42.260 907.420 42.400 ;
        RECT 980.345 42.400 980.635 42.445 ;
        RECT 1075.565 42.400 1075.855 42.445 ;
        RECT 980.345 42.260 1075.855 42.400 ;
        RECT 882.350 42.200 882.670 42.260 ;
        RECT 980.345 42.215 980.635 42.260 ;
        RECT 1075.565 42.215 1075.855 42.260 ;
        RECT 1076.945 42.400 1077.235 42.445 ;
        RECT 1076.945 42.260 1172.840 42.400 ;
        RECT 1076.945 42.215 1077.235 42.260 ;
        RECT 1172.700 42.060 1172.840 42.260 ;
        RECT 1198.460 42.060 1198.600 42.600 ;
        RECT 1214.470 42.540 1214.790 42.600 ;
        RECT 1172.700 41.920 1198.600 42.060 ;
        RECT 966.085 41.380 966.375 41.425 ;
        RECT 980.345 41.380 980.635 41.425 ;
        RECT 966.085 41.240 980.635 41.380 ;
        RECT 966.085 41.195 966.375 41.240 ;
        RECT 980.345 41.195 980.635 41.240 ;
        RECT 1075.565 40.020 1075.855 40.065 ;
        RECT 1076.945 40.020 1077.235 40.065 ;
        RECT 1075.565 39.880 1077.235 40.020 ;
        RECT 1075.565 39.835 1075.855 39.880 ;
        RECT 1076.945 39.835 1077.235 39.880 ;
        RECT 1214.470 14.860 1214.790 14.920 ;
        RECT 1536.930 14.860 1537.250 14.920 ;
        RECT 1214.470 14.720 1537.250 14.860 ;
        RECT 1214.470 14.660 1214.790 14.720 ;
        RECT 1536.930 14.660 1537.250 14.720 ;
      LAYER via ;
        RECT 882.380 42.200 882.640 42.460 ;
        RECT 1214.500 42.540 1214.760 42.800 ;
        RECT 1214.500 14.660 1214.760 14.920 ;
        RECT 1536.960 14.660 1537.220 14.920 ;
      LAYER met2 ;
        RECT 882.700 1600.380 882.980 1604.000 ;
        RECT 882.700 1600.000 883.040 1600.380 ;
        RECT 882.900 1588.210 883.040 1600.000 ;
        RECT 882.440 1588.070 883.040 1588.210 ;
        RECT 882.440 42.490 882.580 1588.070 ;
        RECT 1214.500 42.510 1214.760 42.830 ;
        RECT 882.380 42.170 882.640 42.490 ;
        RECT 1214.560 14.950 1214.700 42.510 ;
        RECT 1214.500 14.630 1214.760 14.950 ;
        RECT 1536.960 14.630 1537.220 14.950 ;
        RECT 1537.020 2.400 1537.160 14.630 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 924.745 1587.545 924.915 1588.735 ;
      LAYER mcon ;
        RECT 924.745 1588.565 924.915 1588.735 ;
      LAYER met1 ;
        RECT 888.790 1588.720 889.110 1588.780 ;
        RECT 924.685 1588.720 924.975 1588.765 ;
        RECT 888.790 1588.580 924.975 1588.720 ;
        RECT 888.790 1588.520 889.110 1588.580 ;
        RECT 924.685 1588.535 924.975 1588.580 ;
        RECT 924.685 1587.700 924.975 1587.745 ;
        RECT 1500.590 1587.700 1500.910 1587.760 ;
        RECT 924.685 1587.560 1500.910 1587.700 ;
        RECT 924.685 1587.515 924.975 1587.560 ;
        RECT 1500.590 1587.500 1500.910 1587.560 ;
        RECT 1500.590 16.900 1500.910 16.960 ;
        RECT 1500.590 16.760 1502.200 16.900 ;
        RECT 1500.590 16.700 1500.910 16.760 ;
        RECT 1502.060 16.560 1502.200 16.760 ;
        RECT 1554.870 16.560 1555.190 16.620 ;
        RECT 1502.060 16.420 1555.190 16.560 ;
        RECT 1554.870 16.360 1555.190 16.420 ;
      LAYER via ;
        RECT 888.820 1588.520 889.080 1588.780 ;
        RECT 1500.620 1587.500 1500.880 1587.760 ;
        RECT 1500.620 16.700 1500.880 16.960 ;
        RECT 1554.900 16.360 1555.160 16.620 ;
      LAYER met2 ;
        RECT 888.680 1600.380 888.960 1604.000 ;
        RECT 888.680 1600.000 889.020 1600.380 ;
        RECT 888.880 1588.810 889.020 1600.000 ;
        RECT 888.820 1588.490 889.080 1588.810 ;
        RECT 1500.620 1587.470 1500.880 1587.790 ;
        RECT 1500.680 16.990 1500.820 1587.470 ;
        RECT 1500.620 16.670 1500.880 16.990 ;
        RECT 1554.900 16.330 1555.160 16.650 ;
        RECT 1554.960 2.400 1555.100 16.330 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 901.285 14.365 901.455 18.615 ;
      LAYER mcon ;
        RECT 901.285 18.445 901.455 18.615 ;
      LAYER met1 ;
        RECT 896.610 18.600 896.930 18.660 ;
        RECT 901.225 18.600 901.515 18.645 ;
        RECT 896.610 18.460 901.515 18.600 ;
        RECT 896.610 18.400 896.930 18.460 ;
        RECT 901.225 18.415 901.515 18.460 ;
        RECT 901.225 14.520 901.515 14.565 ;
        RECT 1572.810 14.520 1573.130 14.580 ;
        RECT 901.225 14.380 1573.130 14.520 ;
        RECT 901.225 14.335 901.515 14.380 ;
        RECT 1572.810 14.320 1573.130 14.380 ;
      LAYER via ;
        RECT 896.640 18.400 896.900 18.660 ;
        RECT 1572.840 14.320 1573.100 14.580 ;
      LAYER met2 ;
        RECT 895.120 1600.450 895.400 1604.000 ;
        RECT 895.120 1600.310 896.380 1600.450 ;
        RECT 895.120 1600.000 895.400 1600.310 ;
        RECT 896.240 1580.050 896.380 1600.310 ;
        RECT 896.240 1579.910 896.840 1580.050 ;
        RECT 896.700 18.690 896.840 1579.910 ;
        RECT 896.640 18.370 896.900 18.690 ;
        RECT 1572.840 14.290 1573.100 14.610 ;
        RECT 1572.900 2.400 1573.040 14.290 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1573.805 14.705 1573.975 16.915 ;
      LAYER mcon ;
        RECT 1573.805 16.745 1573.975 16.915 ;
      LAYER met1 ;
        RECT 901.210 1588.380 901.530 1588.440 ;
        RECT 901.210 1588.240 924.900 1588.380 ;
        RECT 901.210 1588.180 901.530 1588.240 ;
        RECT 924.760 1588.040 924.900 1588.240 ;
        RECT 1535.090 1588.040 1535.410 1588.100 ;
        RECT 924.760 1587.900 1535.410 1588.040 ;
        RECT 1535.090 1587.840 1535.410 1587.900 ;
        RECT 1535.090 16.900 1535.410 16.960 ;
        RECT 1573.745 16.900 1574.035 16.945 ;
        RECT 1535.090 16.760 1574.035 16.900 ;
        RECT 1535.090 16.700 1535.410 16.760 ;
        RECT 1573.745 16.715 1574.035 16.760 ;
        RECT 1573.745 14.860 1574.035 14.905 ;
        RECT 1590.290 14.860 1590.610 14.920 ;
        RECT 1573.745 14.720 1590.610 14.860 ;
        RECT 1573.745 14.675 1574.035 14.720 ;
        RECT 1590.290 14.660 1590.610 14.720 ;
      LAYER via ;
        RECT 901.240 1588.180 901.500 1588.440 ;
        RECT 1535.120 1587.840 1535.380 1588.100 ;
        RECT 1535.120 16.700 1535.380 16.960 ;
        RECT 1590.320 14.660 1590.580 14.920 ;
      LAYER met2 ;
        RECT 901.100 1600.380 901.380 1604.000 ;
        RECT 901.100 1600.000 901.440 1600.380 ;
        RECT 901.300 1588.470 901.440 1600.000 ;
        RECT 901.240 1588.150 901.500 1588.470 ;
        RECT 1535.120 1587.810 1535.380 1588.130 ;
        RECT 1535.180 16.990 1535.320 1587.810 ;
        RECT 1535.120 16.670 1535.380 16.990 ;
        RECT 1590.320 14.630 1590.580 14.950 ;
        RECT 1590.380 2.400 1590.520 14.630 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1197.525 42.585 1197.695 47.515 ;
        RECT 1224.205 43.605 1224.375 47.515 ;
      LAYER mcon ;
        RECT 1197.525 47.345 1197.695 47.515 ;
        RECT 1224.205 47.345 1224.375 47.515 ;
      LAYER met1 ;
        RECT 1197.465 47.500 1197.755 47.545 ;
        RECT 1224.145 47.500 1224.435 47.545 ;
        RECT 1197.465 47.360 1224.435 47.500 ;
        RECT 1197.465 47.315 1197.755 47.360 ;
        RECT 1224.145 47.315 1224.435 47.360 ;
        RECT 1224.145 43.760 1224.435 43.805 ;
        RECT 1240.690 43.760 1241.010 43.820 ;
        RECT 1224.145 43.620 1241.010 43.760 ;
        RECT 1224.145 43.575 1224.435 43.620 ;
        RECT 1240.690 43.560 1241.010 43.620 ;
        RECT 909.950 42.740 910.270 42.800 ;
        RECT 1197.465 42.740 1197.755 42.785 ;
        RECT 909.950 42.600 1197.755 42.740 ;
        RECT 909.950 42.540 910.270 42.600 ;
        RECT 1197.465 42.555 1197.755 42.600 ;
        RECT 1248.970 15.200 1249.290 15.260 ;
        RECT 1608.230 15.200 1608.550 15.260 ;
        RECT 1248.970 15.060 1608.550 15.200 ;
        RECT 1248.970 15.000 1249.290 15.060 ;
        RECT 1608.230 15.000 1608.550 15.060 ;
      LAYER via ;
        RECT 1240.720 43.560 1240.980 43.820 ;
        RECT 909.980 42.540 910.240 42.800 ;
        RECT 1249.000 15.000 1249.260 15.260 ;
        RECT 1608.260 15.000 1608.520 15.260 ;
      LAYER met2 ;
        RECT 907.540 1600.450 907.820 1604.000 ;
        RECT 907.540 1600.310 908.800 1600.450 ;
        RECT 907.540 1600.000 907.820 1600.310 ;
        RECT 908.660 1580.050 908.800 1600.310 ;
        RECT 908.660 1579.910 910.180 1580.050 ;
        RECT 910.040 42.830 910.180 1579.910 ;
        RECT 1240.720 43.530 1240.980 43.850 ;
        RECT 1240.780 43.365 1240.920 43.530 ;
        RECT 1240.710 42.995 1240.990 43.365 ;
        RECT 1248.990 42.995 1249.270 43.365 ;
        RECT 909.980 42.510 910.240 42.830 ;
        RECT 1249.060 15.290 1249.200 42.995 ;
        RECT 1249.000 14.970 1249.260 15.290 ;
        RECT 1608.260 14.970 1608.520 15.290 ;
        RECT 1608.320 2.400 1608.460 14.970 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
      LAYER via2 ;
        RECT 1240.710 43.040 1240.990 43.320 ;
        RECT 1248.990 43.040 1249.270 43.320 ;
      LAYER met3 ;
        RECT 1240.685 43.330 1241.015 43.345 ;
        RECT 1248.965 43.330 1249.295 43.345 ;
        RECT 1240.685 43.030 1249.295 43.330 ;
        RECT 1240.685 43.015 1241.015 43.030 ;
        RECT 1248.965 43.015 1249.295 43.030 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 950.045 1588.905 950.215 1590.435 ;
        RECT 994.665 1590.265 995.755 1590.435 ;
        RECT 1020.885 1588.565 1021.055 1590.435 ;
        RECT 1062.745 1586.865 1062.915 1588.735 ;
        RECT 1124.385 1586.865 1124.555 1588.735 ;
        RECT 1352.545 1586.865 1352.715 1588.735 ;
        RECT 1400.385 1586.865 1400.555 1588.735 ;
        RECT 1449.145 1587.205 1449.315 1588.735 ;
        RECT 1496.985 1587.205 1497.155 1588.735 ;
        RECT 1545.745 1587.885 1545.915 1588.735 ;
      LAYER mcon ;
        RECT 950.045 1590.265 950.215 1590.435 ;
        RECT 995.585 1590.265 995.755 1590.435 ;
        RECT 1020.885 1590.265 1021.055 1590.435 ;
        RECT 1062.745 1588.565 1062.915 1588.735 ;
        RECT 1124.385 1588.565 1124.555 1588.735 ;
        RECT 1352.545 1588.565 1352.715 1588.735 ;
        RECT 1400.385 1588.565 1400.555 1588.735 ;
        RECT 1449.145 1588.565 1449.315 1588.735 ;
        RECT 1496.985 1588.565 1497.155 1588.735 ;
        RECT 1545.745 1588.565 1545.915 1588.735 ;
      LAYER met1 ;
        RECT 949.985 1590.420 950.275 1590.465 ;
        RECT 994.605 1590.420 994.895 1590.465 ;
        RECT 949.985 1590.280 994.895 1590.420 ;
        RECT 949.985 1590.235 950.275 1590.280 ;
        RECT 994.605 1590.235 994.895 1590.280 ;
        RECT 995.525 1590.420 995.815 1590.465 ;
        RECT 1020.825 1590.420 1021.115 1590.465 ;
        RECT 995.525 1590.280 1021.115 1590.420 ;
        RECT 995.525 1590.235 995.815 1590.280 ;
        RECT 1020.825 1590.235 1021.115 1590.280 ;
        RECT 913.630 1589.060 913.950 1589.120 ;
        RECT 949.985 1589.060 950.275 1589.105 ;
        RECT 913.630 1588.920 950.275 1589.060 ;
        RECT 913.630 1588.860 913.950 1588.920 ;
        RECT 949.985 1588.875 950.275 1588.920 ;
        RECT 1020.825 1588.720 1021.115 1588.765 ;
        RECT 1062.685 1588.720 1062.975 1588.765 ;
        RECT 1020.825 1588.580 1062.975 1588.720 ;
        RECT 1020.825 1588.535 1021.115 1588.580 ;
        RECT 1062.685 1588.535 1062.975 1588.580 ;
        RECT 1124.325 1588.720 1124.615 1588.765 ;
        RECT 1352.485 1588.720 1352.775 1588.765 ;
        RECT 1124.325 1588.580 1352.775 1588.720 ;
        RECT 1124.325 1588.535 1124.615 1588.580 ;
        RECT 1352.485 1588.535 1352.775 1588.580 ;
        RECT 1400.325 1588.720 1400.615 1588.765 ;
        RECT 1449.085 1588.720 1449.375 1588.765 ;
        RECT 1400.325 1588.580 1449.375 1588.720 ;
        RECT 1400.325 1588.535 1400.615 1588.580 ;
        RECT 1449.085 1588.535 1449.375 1588.580 ;
        RECT 1496.925 1588.720 1497.215 1588.765 ;
        RECT 1545.685 1588.720 1545.975 1588.765 ;
        RECT 1496.925 1588.580 1545.975 1588.720 ;
        RECT 1496.925 1588.535 1497.215 1588.580 ;
        RECT 1545.685 1588.535 1545.975 1588.580 ;
        RECT 1545.685 1588.040 1545.975 1588.085 ;
        RECT 1555.790 1588.040 1556.110 1588.100 ;
        RECT 1545.685 1587.900 1556.110 1588.040 ;
        RECT 1545.685 1587.855 1545.975 1587.900 ;
        RECT 1555.790 1587.840 1556.110 1587.900 ;
        RECT 1449.085 1587.360 1449.375 1587.405 ;
        RECT 1496.925 1587.360 1497.215 1587.405 ;
        RECT 1449.085 1587.220 1497.215 1587.360 ;
        RECT 1449.085 1587.175 1449.375 1587.220 ;
        RECT 1496.925 1587.175 1497.215 1587.220 ;
        RECT 1062.685 1587.020 1062.975 1587.065 ;
        RECT 1124.325 1587.020 1124.615 1587.065 ;
        RECT 1062.685 1586.880 1124.615 1587.020 ;
        RECT 1062.685 1586.835 1062.975 1586.880 ;
        RECT 1124.325 1586.835 1124.615 1586.880 ;
        RECT 1352.485 1587.020 1352.775 1587.065 ;
        RECT 1400.325 1587.020 1400.615 1587.065 ;
        RECT 1352.485 1586.880 1400.615 1587.020 ;
        RECT 1352.485 1586.835 1352.775 1586.880 ;
        RECT 1400.325 1586.835 1400.615 1586.880 ;
        RECT 1555.790 16.560 1556.110 16.620 ;
        RECT 1626.170 16.560 1626.490 16.620 ;
        RECT 1555.790 16.420 1626.490 16.560 ;
        RECT 1555.790 16.360 1556.110 16.420 ;
        RECT 1626.170 16.360 1626.490 16.420 ;
      LAYER via ;
        RECT 913.660 1588.860 913.920 1589.120 ;
        RECT 1555.820 1587.840 1556.080 1588.100 ;
        RECT 1555.820 16.360 1556.080 16.620 ;
        RECT 1626.200 16.360 1626.460 16.620 ;
      LAYER met2 ;
        RECT 913.520 1600.380 913.800 1604.000 ;
        RECT 913.520 1600.000 913.860 1600.380 ;
        RECT 913.720 1589.150 913.860 1600.000 ;
        RECT 913.660 1588.830 913.920 1589.150 ;
        RECT 1555.820 1587.810 1556.080 1588.130 ;
        RECT 1555.880 16.650 1556.020 1587.810 ;
        RECT 1555.820 16.330 1556.080 16.650 ;
        RECT 1626.200 16.330 1626.460 16.650 ;
        RECT 1626.260 2.400 1626.400 16.330 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 919.610 1588.040 919.930 1588.100 ;
        RECT 924.210 1588.040 924.530 1588.100 ;
        RECT 919.610 1587.900 924.530 1588.040 ;
        RECT 919.610 1587.840 919.930 1587.900 ;
        RECT 924.210 1587.840 924.530 1587.900 ;
        RECT 923.750 20.640 924.070 20.700 ;
        RECT 1644.110 20.640 1644.430 20.700 ;
        RECT 923.750 20.500 1644.430 20.640 ;
        RECT 923.750 20.440 924.070 20.500 ;
        RECT 1644.110 20.440 1644.430 20.500 ;
      LAYER via ;
        RECT 919.640 1587.840 919.900 1588.100 ;
        RECT 924.240 1587.840 924.500 1588.100 ;
        RECT 923.780 20.440 924.040 20.700 ;
        RECT 1644.140 20.440 1644.400 20.700 ;
      LAYER met2 ;
        RECT 919.500 1600.380 919.780 1604.000 ;
        RECT 919.500 1600.000 919.840 1600.380 ;
        RECT 919.700 1588.130 919.840 1600.000 ;
        RECT 919.640 1587.810 919.900 1588.130 ;
        RECT 924.240 1587.810 924.500 1588.130 ;
        RECT 924.300 32.370 924.440 1587.810 ;
        RECT 923.840 32.230 924.440 32.370 ;
        RECT 923.840 20.730 923.980 32.230 ;
        RECT 923.780 20.410 924.040 20.730 ;
        RECT 1644.140 20.410 1644.400 20.730 ;
        RECT 1644.200 2.400 1644.340 20.410 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 955.105 1591.285 955.275 1592.815 ;
        RECT 979.485 1588.225 979.655 1591.455 ;
      LAYER mcon ;
        RECT 955.105 1592.645 955.275 1592.815 ;
        RECT 979.485 1591.285 979.655 1591.455 ;
      LAYER met1 ;
        RECT 926.050 1592.800 926.370 1592.860 ;
        RECT 955.045 1592.800 955.335 1592.845 ;
        RECT 926.050 1592.660 955.335 1592.800 ;
        RECT 926.050 1592.600 926.370 1592.660 ;
        RECT 955.045 1592.615 955.335 1592.660 ;
        RECT 955.045 1591.440 955.335 1591.485 ;
        RECT 979.425 1591.440 979.715 1591.485 ;
        RECT 955.045 1591.300 979.715 1591.440 ;
        RECT 955.045 1591.255 955.335 1591.300 ;
        RECT 979.425 1591.255 979.715 1591.300 ;
        RECT 979.425 1588.380 979.715 1588.425 ;
        RECT 1569.590 1588.380 1569.910 1588.440 ;
        RECT 979.425 1588.240 1569.910 1588.380 ;
        RECT 979.425 1588.195 979.715 1588.240 ;
        RECT 1569.590 1588.180 1569.910 1588.240 ;
        RECT 1569.590 14.860 1569.910 14.920 ;
        RECT 1569.590 14.720 1573.500 14.860 ;
        RECT 1569.590 14.660 1569.910 14.720 ;
        RECT 1573.360 14.520 1573.500 14.720 ;
        RECT 1662.050 14.520 1662.370 14.580 ;
        RECT 1573.360 14.380 1662.370 14.520 ;
        RECT 1662.050 14.320 1662.370 14.380 ;
      LAYER via ;
        RECT 926.080 1592.600 926.340 1592.860 ;
        RECT 1569.620 1588.180 1569.880 1588.440 ;
        RECT 1569.620 14.660 1569.880 14.920 ;
        RECT 1662.080 14.320 1662.340 14.580 ;
      LAYER met2 ;
        RECT 925.940 1600.380 926.220 1604.000 ;
        RECT 925.940 1600.000 926.280 1600.380 ;
        RECT 926.140 1592.890 926.280 1600.000 ;
        RECT 926.080 1592.570 926.340 1592.890 ;
        RECT 1569.620 1588.150 1569.880 1588.470 ;
        RECT 1569.680 14.950 1569.820 1588.150 ;
        RECT 1569.620 14.630 1569.880 14.950 ;
        RECT 1662.080 14.290 1662.340 14.610 ;
        RECT 1662.140 2.400 1662.280 14.290 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 932.030 1588.380 932.350 1588.440 ;
        RECT 938.010 1588.380 938.330 1588.440 ;
        RECT 932.030 1588.240 938.330 1588.380 ;
        RECT 932.030 1588.180 932.350 1588.240 ;
        RECT 938.010 1588.180 938.330 1588.240 ;
        RECT 938.010 20.300 938.330 20.360 ;
        RECT 1679.530 20.300 1679.850 20.360 ;
        RECT 938.010 20.160 1679.850 20.300 ;
        RECT 938.010 20.100 938.330 20.160 ;
        RECT 1679.530 20.100 1679.850 20.160 ;
      LAYER via ;
        RECT 932.060 1588.180 932.320 1588.440 ;
        RECT 938.040 1588.180 938.300 1588.440 ;
        RECT 938.040 20.100 938.300 20.360 ;
        RECT 1679.560 20.100 1679.820 20.360 ;
      LAYER met2 ;
        RECT 931.920 1600.380 932.200 1604.000 ;
        RECT 931.920 1600.000 932.260 1600.380 ;
        RECT 932.120 1588.470 932.260 1600.000 ;
        RECT 932.060 1588.150 932.320 1588.470 ;
        RECT 938.040 1588.150 938.300 1588.470 ;
        RECT 938.100 20.390 938.240 1588.150 ;
        RECT 938.040 20.070 938.300 20.390 ;
        RECT 1679.560 20.070 1679.820 20.390 ;
        RECT 1679.620 2.400 1679.760 20.070 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1590.290 1589.060 1590.610 1589.120 ;
        RECT 969.380 1588.920 1590.610 1589.060 ;
        RECT 938.470 1588.720 938.790 1588.780 ;
        RECT 969.380 1588.720 969.520 1588.920 ;
        RECT 1590.290 1588.860 1590.610 1588.920 ;
        RECT 938.470 1588.580 969.520 1588.720 ;
        RECT 938.470 1588.520 938.790 1588.580 ;
        RECT 1590.750 14.860 1591.070 14.920 ;
        RECT 1697.470 14.860 1697.790 14.920 ;
        RECT 1590.750 14.720 1697.790 14.860 ;
        RECT 1590.750 14.660 1591.070 14.720 ;
        RECT 1697.470 14.660 1697.790 14.720 ;
      LAYER via ;
        RECT 938.500 1588.520 938.760 1588.780 ;
        RECT 1590.320 1588.860 1590.580 1589.120 ;
        RECT 1590.780 14.660 1591.040 14.920 ;
        RECT 1697.500 14.660 1697.760 14.920 ;
      LAYER met2 ;
        RECT 938.360 1600.380 938.640 1604.000 ;
        RECT 938.360 1600.000 938.700 1600.380 ;
        RECT 938.560 1588.810 938.700 1600.000 ;
        RECT 1590.320 1588.830 1590.580 1589.150 ;
        RECT 938.500 1588.490 938.760 1588.810 ;
        RECT 1590.380 24.890 1590.520 1588.830 ;
        RECT 1590.380 24.750 1590.980 24.890 ;
        RECT 1590.840 14.950 1590.980 24.750 ;
        RECT 1590.780 14.630 1591.040 14.950 ;
        RECT 1697.500 14.630 1697.760 14.950 ;
        RECT 1697.560 2.400 1697.700 14.630 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 613.340 1590.280 691.220 1590.420 ;
        RECT 604.510 1590.080 604.830 1590.140 ;
        RECT 613.340 1590.080 613.480 1590.280 ;
        RECT 604.510 1589.940 613.480 1590.080 ;
        RECT 691.080 1590.080 691.220 1590.280 ;
        RECT 732.850 1590.080 733.170 1590.140 ;
        RECT 691.080 1589.940 733.170 1590.080 ;
        RECT 604.510 1589.880 604.830 1589.940 ;
        RECT 732.850 1589.880 733.170 1589.940 ;
        RECT 732.850 2.960 733.170 3.020 ;
        RECT 734.230 2.960 734.550 3.020 ;
        RECT 732.850 2.820 734.550 2.960 ;
        RECT 732.850 2.760 733.170 2.820 ;
        RECT 734.230 2.760 734.550 2.820 ;
      LAYER via ;
        RECT 604.540 1589.880 604.800 1590.140 ;
        RECT 732.880 1589.880 733.140 1590.140 ;
        RECT 732.880 2.760 733.140 3.020 ;
        RECT 734.260 2.760 734.520 3.020 ;
      LAYER met2 ;
        RECT 604.400 1600.380 604.680 1604.000 ;
        RECT 604.400 1600.000 604.740 1600.380 ;
        RECT 604.600 1590.170 604.740 1600.000 ;
        RECT 604.540 1589.850 604.800 1590.170 ;
        RECT 732.880 1589.850 733.140 1590.170 ;
        RECT 732.940 3.050 733.080 1589.850 ;
        RECT 732.880 2.730 733.140 3.050 ;
        RECT 734.260 2.730 734.520 3.050 ;
        RECT 734.320 2.400 734.460 2.730 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 948.665 14.025 948.835 15.215 ;
      LAYER mcon ;
        RECT 948.665 15.045 948.835 15.215 ;
      LAYER met1 ;
        RECT 944.910 15.200 945.230 15.260 ;
        RECT 948.605 15.200 948.895 15.245 ;
        RECT 944.910 15.060 948.895 15.200 ;
        RECT 944.910 15.000 945.230 15.060 ;
        RECT 948.605 15.015 948.895 15.060 ;
        RECT 948.605 14.180 948.895 14.225 ;
        RECT 1715.410 14.180 1715.730 14.240 ;
        RECT 948.605 14.040 1715.730 14.180 ;
        RECT 948.605 13.995 948.895 14.040 ;
        RECT 1715.410 13.980 1715.730 14.040 ;
      LAYER via ;
        RECT 944.940 15.000 945.200 15.260 ;
        RECT 1715.440 13.980 1715.700 14.240 ;
      LAYER met2 ;
        RECT 944.340 1600.450 944.620 1604.000 ;
        RECT 944.340 1600.310 945.140 1600.450 ;
        RECT 944.340 1600.000 944.620 1600.310 ;
        RECT 945.000 15.290 945.140 1600.310 ;
        RECT 944.940 14.970 945.200 15.290 ;
        RECT 1715.440 13.950 1715.700 14.270 ;
        RECT 1715.500 2.400 1715.640 13.950 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 950.890 1589.740 951.210 1589.800 ;
        RECT 1610.990 1589.740 1611.310 1589.800 ;
        RECT 950.890 1589.600 1611.310 1589.740 ;
        RECT 950.890 1589.540 951.210 1589.600 ;
        RECT 1610.990 1589.540 1611.310 1589.600 ;
        RECT 1610.990 15.200 1611.310 15.260 ;
        RECT 1733.350 15.200 1733.670 15.260 ;
        RECT 1610.990 15.060 1733.670 15.200 ;
        RECT 1610.990 15.000 1611.310 15.060 ;
        RECT 1733.350 15.000 1733.670 15.060 ;
      LAYER via ;
        RECT 950.920 1589.540 951.180 1589.800 ;
        RECT 1611.020 1589.540 1611.280 1589.800 ;
        RECT 1611.020 15.000 1611.280 15.260 ;
        RECT 1733.380 15.000 1733.640 15.260 ;
      LAYER met2 ;
        RECT 950.780 1600.380 951.060 1604.000 ;
        RECT 950.780 1600.000 951.120 1600.380 ;
        RECT 950.980 1589.830 951.120 1600.000 ;
        RECT 950.920 1589.510 951.180 1589.830 ;
        RECT 1611.020 1589.510 1611.280 1589.830 ;
        RECT 1611.080 15.290 1611.220 1589.510 ;
        RECT 1611.020 14.970 1611.280 15.290 ;
        RECT 1733.380 14.970 1733.640 15.290 ;
        RECT 1733.440 2.400 1733.580 14.970 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1244.905 42.245 1245.075 44.455 ;
        RECT 1274.805 44.285 1274.975 46.495 ;
        RECT 985.925 40.885 986.095 42.075 ;
        RECT 1014.445 40.885 1014.615 42.075 ;
        RECT 1027.785 41.905 1028.415 42.075 ;
        RECT 1076.085 40.205 1076.255 42.075 ;
        RECT 1076.545 40.205 1076.715 42.075 ;
      LAYER mcon ;
        RECT 1274.805 46.325 1274.975 46.495 ;
        RECT 1244.905 44.285 1245.075 44.455 ;
        RECT 985.925 41.905 986.095 42.075 ;
        RECT 1014.445 41.905 1014.615 42.075 ;
        RECT 1028.245 41.905 1028.415 42.075 ;
        RECT 1076.085 41.905 1076.255 42.075 ;
        RECT 1076.545 41.905 1076.715 42.075 ;
      LAYER met1 ;
        RECT 1274.745 46.480 1275.035 46.525 ;
        RECT 1274.745 46.340 1281.860 46.480 ;
        RECT 1274.745 46.295 1275.035 46.340 ;
        RECT 1281.720 46.140 1281.860 46.340 ;
        RECT 1288.990 46.140 1289.310 46.200 ;
        RECT 1281.720 46.000 1289.310 46.140 ;
        RECT 1288.990 45.940 1289.310 46.000 ;
        RECT 1244.845 44.440 1245.135 44.485 ;
        RECT 1274.745 44.440 1275.035 44.485 ;
        RECT 1244.845 44.300 1275.035 44.440 ;
        RECT 1244.845 44.255 1245.135 44.300 ;
        RECT 1274.745 44.255 1275.035 44.300 ;
        RECT 1198.830 42.400 1199.150 42.460 ;
        RECT 1244.845 42.400 1245.135 42.445 ;
        RECT 1198.830 42.260 1245.135 42.400 ;
        RECT 1198.830 42.200 1199.150 42.260 ;
        RECT 1244.845 42.215 1245.135 42.260 ;
        RECT 958.250 42.060 958.570 42.120 ;
        RECT 985.865 42.060 986.155 42.105 ;
        RECT 958.250 41.920 986.155 42.060 ;
        RECT 958.250 41.860 958.570 41.920 ;
        RECT 985.865 41.875 986.155 41.920 ;
        RECT 1014.385 42.060 1014.675 42.105 ;
        RECT 1027.725 42.060 1028.015 42.105 ;
        RECT 1014.385 41.920 1028.015 42.060 ;
        RECT 1014.385 41.875 1014.675 41.920 ;
        RECT 1027.725 41.875 1028.015 41.920 ;
        RECT 1028.185 42.060 1028.475 42.105 ;
        RECT 1076.025 42.060 1076.315 42.105 ;
        RECT 1028.185 41.920 1076.315 42.060 ;
        RECT 1028.185 41.875 1028.475 41.920 ;
        RECT 1076.025 41.875 1076.315 41.920 ;
        RECT 1076.485 42.060 1076.775 42.105 ;
        RECT 1172.150 42.060 1172.470 42.120 ;
        RECT 1076.485 41.920 1172.470 42.060 ;
        RECT 1076.485 41.875 1076.775 41.920 ;
        RECT 1172.150 41.860 1172.470 41.920 ;
        RECT 985.865 41.040 986.155 41.085 ;
        RECT 1014.385 41.040 1014.675 41.085 ;
        RECT 985.865 40.900 1014.675 41.040 ;
        RECT 985.865 40.855 986.155 40.900 ;
        RECT 1014.385 40.855 1014.675 40.900 ;
        RECT 1076.025 40.360 1076.315 40.405 ;
        RECT 1076.485 40.360 1076.775 40.405 ;
        RECT 1076.025 40.220 1076.775 40.360 ;
        RECT 1076.025 40.175 1076.315 40.220 ;
        RECT 1076.485 40.175 1076.775 40.220 ;
        RECT 1288.990 15.540 1289.310 15.600 ;
        RECT 1751.290 15.540 1751.610 15.600 ;
        RECT 1288.990 15.400 1751.610 15.540 ;
        RECT 1288.990 15.340 1289.310 15.400 ;
        RECT 1751.290 15.340 1751.610 15.400 ;
      LAYER via ;
        RECT 1289.020 45.940 1289.280 46.200 ;
        RECT 1198.860 42.200 1199.120 42.460 ;
        RECT 958.280 41.860 958.540 42.120 ;
        RECT 1172.180 41.860 1172.440 42.120 ;
        RECT 1289.020 15.340 1289.280 15.600 ;
        RECT 1751.320 15.340 1751.580 15.600 ;
      LAYER met2 ;
        RECT 956.760 1600.450 957.040 1604.000 ;
        RECT 956.760 1600.310 958.480 1600.450 ;
        RECT 956.760 1600.000 957.040 1600.310 ;
        RECT 958.340 42.150 958.480 1600.310 ;
        RECT 1289.020 45.910 1289.280 46.230 ;
        RECT 1198.860 42.170 1199.120 42.490 ;
        RECT 958.280 41.830 958.540 42.150 ;
        RECT 1172.180 42.005 1172.440 42.150 ;
        RECT 1198.920 42.005 1199.060 42.170 ;
        RECT 1172.170 41.635 1172.450 42.005 ;
        RECT 1198.850 41.635 1199.130 42.005 ;
        RECT 1289.080 15.630 1289.220 45.910 ;
        RECT 1289.020 15.310 1289.280 15.630 ;
        RECT 1751.320 15.310 1751.580 15.630 ;
        RECT 1751.380 2.400 1751.520 15.310 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
      LAYER via2 ;
        RECT 1172.170 41.680 1172.450 41.960 ;
        RECT 1198.850 41.680 1199.130 41.960 ;
      LAYER met3 ;
        RECT 1172.145 41.970 1172.475 41.985 ;
        RECT 1198.825 41.970 1199.155 41.985 ;
        RECT 1172.145 41.670 1199.155 41.970 ;
        RECT 1172.145 41.655 1172.475 41.670 ;
        RECT 1198.825 41.655 1199.155 41.670 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1003.865 1589.245 1004.035 1593.835 ;
        RECT 1624.865 1497.445 1625.035 1545.555 ;
        RECT 1624.865 1400.885 1625.035 1448.995 ;
        RECT 1624.865 1304.325 1625.035 1352.435 ;
        RECT 1623.945 1207.765 1624.115 1255.535 ;
        RECT 1624.405 1173.085 1624.575 1207.255 ;
        RECT 1624.865 338.045 1625.035 386.155 ;
        RECT 1624.405 192.525 1624.575 234.515 ;
        RECT 1738.485 15.045 1738.655 16.575 ;
      LAYER mcon ;
        RECT 1003.865 1593.665 1004.035 1593.835 ;
        RECT 1624.865 1545.385 1625.035 1545.555 ;
        RECT 1624.865 1448.825 1625.035 1448.995 ;
        RECT 1624.865 1352.265 1625.035 1352.435 ;
        RECT 1623.945 1255.365 1624.115 1255.535 ;
        RECT 1624.405 1207.085 1624.575 1207.255 ;
        RECT 1624.865 385.985 1625.035 386.155 ;
        RECT 1624.405 234.345 1624.575 234.515 ;
        RECT 1738.485 16.405 1738.655 16.575 ;
      LAYER met1 ;
        RECT 963.310 1593.820 963.630 1593.880 ;
        RECT 1003.805 1593.820 1004.095 1593.865 ;
        RECT 963.310 1593.680 1004.095 1593.820 ;
        RECT 963.310 1593.620 963.630 1593.680 ;
        RECT 1003.805 1593.635 1004.095 1593.680 ;
        RECT 1003.805 1589.400 1004.095 1589.445 ;
        RECT 1625.250 1589.400 1625.570 1589.460 ;
        RECT 1003.805 1589.260 1625.570 1589.400 ;
        RECT 1003.805 1589.215 1004.095 1589.260 ;
        RECT 1625.250 1589.200 1625.570 1589.260 ;
        RECT 1624.805 1545.540 1625.095 1545.585 ;
        RECT 1625.250 1545.540 1625.570 1545.600 ;
        RECT 1624.805 1545.400 1625.570 1545.540 ;
        RECT 1624.805 1545.355 1625.095 1545.400 ;
        RECT 1625.250 1545.340 1625.570 1545.400 ;
        RECT 1624.790 1497.600 1625.110 1497.660 ;
        RECT 1624.595 1497.460 1625.110 1497.600 ;
        RECT 1624.790 1497.400 1625.110 1497.460 ;
        RECT 1624.805 1448.980 1625.095 1449.025 ;
        RECT 1625.250 1448.980 1625.570 1449.040 ;
        RECT 1624.805 1448.840 1625.570 1448.980 ;
        RECT 1624.805 1448.795 1625.095 1448.840 ;
        RECT 1625.250 1448.780 1625.570 1448.840 ;
        RECT 1624.790 1401.040 1625.110 1401.100 ;
        RECT 1624.595 1400.900 1625.110 1401.040 ;
        RECT 1624.790 1400.840 1625.110 1400.900 ;
        RECT 1624.805 1352.420 1625.095 1352.465 ;
        RECT 1625.250 1352.420 1625.570 1352.480 ;
        RECT 1624.805 1352.280 1625.570 1352.420 ;
        RECT 1624.805 1352.235 1625.095 1352.280 ;
        RECT 1625.250 1352.220 1625.570 1352.280 ;
        RECT 1624.790 1304.480 1625.110 1304.540 ;
        RECT 1624.595 1304.340 1625.110 1304.480 ;
        RECT 1624.790 1304.280 1625.110 1304.340 ;
        RECT 1623.870 1256.200 1624.190 1256.260 ;
        RECT 1624.790 1256.200 1625.110 1256.260 ;
        RECT 1623.870 1256.060 1625.110 1256.200 ;
        RECT 1623.870 1256.000 1624.190 1256.060 ;
        RECT 1624.790 1256.000 1625.110 1256.060 ;
        RECT 1623.870 1255.520 1624.190 1255.580 ;
        RECT 1623.675 1255.380 1624.190 1255.520 ;
        RECT 1623.870 1255.320 1624.190 1255.380 ;
        RECT 1623.885 1207.920 1624.175 1207.965 ;
        RECT 1624.330 1207.920 1624.650 1207.980 ;
        RECT 1623.885 1207.780 1624.650 1207.920 ;
        RECT 1623.885 1207.735 1624.175 1207.780 ;
        RECT 1624.330 1207.720 1624.650 1207.780 ;
        RECT 1624.330 1207.240 1624.650 1207.300 ;
        RECT 1624.135 1207.100 1624.650 1207.240 ;
        RECT 1624.330 1207.040 1624.650 1207.100 ;
        RECT 1624.345 1173.240 1624.635 1173.285 ;
        RECT 1625.250 1173.240 1625.570 1173.300 ;
        RECT 1624.345 1173.100 1625.570 1173.240 ;
        RECT 1624.345 1173.055 1624.635 1173.100 ;
        RECT 1625.250 1173.040 1625.570 1173.100 ;
        RECT 1624.330 1111.020 1624.650 1111.080 ;
        RECT 1625.710 1111.020 1626.030 1111.080 ;
        RECT 1624.330 1110.880 1626.030 1111.020 ;
        RECT 1624.330 1110.820 1624.650 1110.880 ;
        RECT 1625.710 1110.820 1626.030 1110.880 ;
        RECT 1625.710 1077.020 1626.030 1077.080 ;
        RECT 1625.340 1076.880 1626.030 1077.020 ;
        RECT 1625.340 1076.400 1625.480 1076.880 ;
        RECT 1625.710 1076.820 1626.030 1076.880 ;
        RECT 1625.250 1076.140 1625.570 1076.400 ;
        RECT 1624.330 1014.460 1624.650 1014.520 ;
        RECT 1625.710 1014.460 1626.030 1014.520 ;
        RECT 1624.330 1014.320 1626.030 1014.460 ;
        RECT 1624.330 1014.260 1624.650 1014.320 ;
        RECT 1625.710 1014.260 1626.030 1014.320 ;
        RECT 1625.710 980.460 1626.030 980.520 ;
        RECT 1625.340 980.320 1626.030 980.460 ;
        RECT 1625.340 979.840 1625.480 980.320 ;
        RECT 1625.710 980.260 1626.030 980.320 ;
        RECT 1625.250 979.580 1625.570 979.840 ;
        RECT 1624.330 917.900 1624.650 917.960 ;
        RECT 1625.710 917.900 1626.030 917.960 ;
        RECT 1624.330 917.760 1626.030 917.900 ;
        RECT 1624.330 917.700 1624.650 917.760 ;
        RECT 1625.710 917.700 1626.030 917.760 ;
        RECT 1625.710 883.900 1626.030 883.960 ;
        RECT 1625.340 883.760 1626.030 883.900 ;
        RECT 1625.340 883.280 1625.480 883.760 ;
        RECT 1625.710 883.700 1626.030 883.760 ;
        RECT 1625.250 883.020 1625.570 883.280 ;
        RECT 1624.330 834.940 1624.650 835.000 ;
        RECT 1625.250 834.940 1625.570 835.000 ;
        RECT 1624.330 834.800 1625.570 834.940 ;
        RECT 1624.330 834.740 1624.650 834.800 ;
        RECT 1625.250 834.740 1625.570 834.800 ;
        RECT 1625.710 787.340 1626.030 787.400 ;
        RECT 1625.340 787.200 1626.030 787.340 ;
        RECT 1625.340 786.380 1625.480 787.200 ;
        RECT 1625.710 787.140 1626.030 787.200 ;
        RECT 1625.250 786.120 1625.570 786.380 ;
        RECT 1625.250 772.720 1625.570 772.780 ;
        RECT 1626.170 772.720 1626.490 772.780 ;
        RECT 1625.250 772.580 1626.490 772.720 ;
        RECT 1625.250 772.520 1625.570 772.580 ;
        RECT 1626.170 772.520 1626.490 772.580 ;
        RECT 1624.790 689.900 1625.110 690.160 ;
        RECT 1624.880 689.760 1625.020 689.900 ;
        RECT 1625.250 689.760 1625.570 689.820 ;
        RECT 1624.880 689.620 1625.570 689.760 ;
        RECT 1625.250 689.560 1625.570 689.620 ;
        RECT 1625.250 676.160 1625.570 676.220 ;
        RECT 1626.170 676.160 1626.490 676.220 ;
        RECT 1625.250 676.020 1626.490 676.160 ;
        RECT 1625.250 675.960 1625.570 676.020 ;
        RECT 1626.170 675.960 1626.490 676.020 ;
        RECT 1624.790 593.340 1625.110 593.600 ;
        RECT 1624.880 593.200 1625.020 593.340 ;
        RECT 1625.250 593.200 1625.570 593.260 ;
        RECT 1624.880 593.060 1625.570 593.200 ;
        RECT 1625.250 593.000 1625.570 593.060 ;
        RECT 1625.250 579.600 1625.570 579.660 ;
        RECT 1626.170 579.600 1626.490 579.660 ;
        RECT 1625.250 579.460 1626.490 579.600 ;
        RECT 1625.250 579.400 1625.570 579.460 ;
        RECT 1626.170 579.400 1626.490 579.460 ;
        RECT 1623.870 507.180 1624.190 507.240 ;
        RECT 1624.790 507.180 1625.110 507.240 ;
        RECT 1623.870 507.040 1625.110 507.180 ;
        RECT 1623.870 506.980 1624.190 507.040 ;
        RECT 1624.790 506.980 1625.110 507.040 ;
        RECT 1624.790 400.220 1625.110 400.480 ;
        RECT 1624.880 399.740 1625.020 400.220 ;
        RECT 1625.250 399.740 1625.570 399.800 ;
        RECT 1624.880 399.600 1625.570 399.740 ;
        RECT 1625.250 399.540 1625.570 399.600 ;
        RECT 1624.805 386.140 1625.095 386.185 ;
        RECT 1625.250 386.140 1625.570 386.200 ;
        RECT 1624.805 386.000 1625.570 386.140 ;
        RECT 1624.805 385.955 1625.095 386.000 ;
        RECT 1625.250 385.940 1625.570 386.000 ;
        RECT 1624.790 338.200 1625.110 338.260 ;
        RECT 1624.595 338.060 1625.110 338.200 ;
        RECT 1624.790 338.000 1625.110 338.060 ;
        RECT 1622.950 241.300 1623.270 241.360 ;
        RECT 1623.870 241.300 1624.190 241.360 ;
        RECT 1622.950 241.160 1624.190 241.300 ;
        RECT 1622.950 241.100 1623.270 241.160 ;
        RECT 1623.870 241.100 1624.190 241.160 ;
        RECT 1622.950 234.500 1623.270 234.560 ;
        RECT 1624.345 234.500 1624.635 234.545 ;
        RECT 1622.950 234.360 1624.635 234.500 ;
        RECT 1622.950 234.300 1623.270 234.360 ;
        RECT 1624.345 234.315 1624.635 234.360 ;
        RECT 1624.330 192.680 1624.650 192.740 ;
        RECT 1624.135 192.540 1624.650 192.680 ;
        RECT 1624.330 192.480 1624.650 192.540 ;
        RECT 1624.330 158.820 1624.650 159.080 ;
        RECT 1624.420 158.400 1624.560 158.820 ;
        RECT 1624.330 158.140 1624.650 158.400 ;
        RECT 1626.630 16.560 1626.950 16.620 ;
        RECT 1738.425 16.560 1738.715 16.605 ;
        RECT 1626.630 16.420 1738.715 16.560 ;
        RECT 1626.630 16.360 1626.950 16.420 ;
        RECT 1738.425 16.375 1738.715 16.420 ;
        RECT 1738.425 15.200 1738.715 15.245 ;
        RECT 1768.770 15.200 1769.090 15.260 ;
        RECT 1738.425 15.060 1769.090 15.200 ;
        RECT 1738.425 15.015 1738.715 15.060 ;
        RECT 1768.770 15.000 1769.090 15.060 ;
      LAYER via ;
        RECT 963.340 1593.620 963.600 1593.880 ;
        RECT 1625.280 1589.200 1625.540 1589.460 ;
        RECT 1625.280 1545.340 1625.540 1545.600 ;
        RECT 1624.820 1497.400 1625.080 1497.660 ;
        RECT 1625.280 1448.780 1625.540 1449.040 ;
        RECT 1624.820 1400.840 1625.080 1401.100 ;
        RECT 1625.280 1352.220 1625.540 1352.480 ;
        RECT 1624.820 1304.280 1625.080 1304.540 ;
        RECT 1623.900 1256.000 1624.160 1256.260 ;
        RECT 1624.820 1256.000 1625.080 1256.260 ;
        RECT 1623.900 1255.320 1624.160 1255.580 ;
        RECT 1624.360 1207.720 1624.620 1207.980 ;
        RECT 1624.360 1207.040 1624.620 1207.300 ;
        RECT 1625.280 1173.040 1625.540 1173.300 ;
        RECT 1624.360 1110.820 1624.620 1111.080 ;
        RECT 1625.740 1110.820 1626.000 1111.080 ;
        RECT 1625.740 1076.820 1626.000 1077.080 ;
        RECT 1625.280 1076.140 1625.540 1076.400 ;
        RECT 1624.360 1014.260 1624.620 1014.520 ;
        RECT 1625.740 1014.260 1626.000 1014.520 ;
        RECT 1625.740 980.260 1626.000 980.520 ;
        RECT 1625.280 979.580 1625.540 979.840 ;
        RECT 1624.360 917.700 1624.620 917.960 ;
        RECT 1625.740 917.700 1626.000 917.960 ;
        RECT 1625.740 883.700 1626.000 883.960 ;
        RECT 1625.280 883.020 1625.540 883.280 ;
        RECT 1624.360 834.740 1624.620 835.000 ;
        RECT 1625.280 834.740 1625.540 835.000 ;
        RECT 1625.740 787.140 1626.000 787.400 ;
        RECT 1625.280 786.120 1625.540 786.380 ;
        RECT 1625.280 772.520 1625.540 772.780 ;
        RECT 1626.200 772.520 1626.460 772.780 ;
        RECT 1624.820 689.900 1625.080 690.160 ;
        RECT 1625.280 689.560 1625.540 689.820 ;
        RECT 1625.280 675.960 1625.540 676.220 ;
        RECT 1626.200 675.960 1626.460 676.220 ;
        RECT 1624.820 593.340 1625.080 593.600 ;
        RECT 1625.280 593.000 1625.540 593.260 ;
        RECT 1625.280 579.400 1625.540 579.660 ;
        RECT 1626.200 579.400 1626.460 579.660 ;
        RECT 1623.900 506.980 1624.160 507.240 ;
        RECT 1624.820 506.980 1625.080 507.240 ;
        RECT 1624.820 400.220 1625.080 400.480 ;
        RECT 1625.280 399.540 1625.540 399.800 ;
        RECT 1625.280 385.940 1625.540 386.200 ;
        RECT 1624.820 338.000 1625.080 338.260 ;
        RECT 1622.980 241.100 1623.240 241.360 ;
        RECT 1623.900 241.100 1624.160 241.360 ;
        RECT 1622.980 234.300 1623.240 234.560 ;
        RECT 1624.360 192.480 1624.620 192.740 ;
        RECT 1624.360 158.820 1624.620 159.080 ;
        RECT 1624.360 158.140 1624.620 158.400 ;
        RECT 1626.660 16.360 1626.920 16.620 ;
        RECT 1768.800 15.000 1769.060 15.260 ;
      LAYER met2 ;
        RECT 963.200 1600.380 963.480 1604.000 ;
        RECT 963.200 1600.000 963.540 1600.380 ;
        RECT 963.400 1593.910 963.540 1600.000 ;
        RECT 963.340 1593.590 963.600 1593.910 ;
        RECT 1625.280 1589.170 1625.540 1589.490 ;
        RECT 1625.340 1545.630 1625.480 1589.170 ;
        RECT 1625.280 1545.310 1625.540 1545.630 ;
        RECT 1624.820 1497.370 1625.080 1497.690 ;
        RECT 1624.880 1463.090 1625.020 1497.370 ;
        RECT 1624.880 1462.950 1625.480 1463.090 ;
        RECT 1625.340 1449.070 1625.480 1462.950 ;
        RECT 1625.280 1448.750 1625.540 1449.070 ;
        RECT 1624.820 1400.810 1625.080 1401.130 ;
        RECT 1624.880 1366.530 1625.020 1400.810 ;
        RECT 1624.880 1366.390 1625.480 1366.530 ;
        RECT 1625.340 1352.510 1625.480 1366.390 ;
        RECT 1625.280 1352.190 1625.540 1352.510 ;
        RECT 1624.820 1304.250 1625.080 1304.570 ;
        RECT 1624.880 1256.290 1625.020 1304.250 ;
        RECT 1623.900 1255.970 1624.160 1256.290 ;
        RECT 1624.820 1255.970 1625.080 1256.290 ;
        RECT 1623.960 1255.610 1624.100 1255.970 ;
        RECT 1623.900 1255.290 1624.160 1255.610 ;
        RECT 1624.360 1207.690 1624.620 1208.010 ;
        RECT 1624.420 1207.330 1624.560 1207.690 ;
        RECT 1624.360 1207.010 1624.620 1207.330 ;
        RECT 1625.280 1173.010 1625.540 1173.330 ;
        RECT 1625.340 1159.245 1625.480 1173.010 ;
        RECT 1624.350 1158.875 1624.630 1159.245 ;
        RECT 1625.270 1158.875 1625.550 1159.245 ;
        RECT 1624.420 1111.110 1624.560 1158.875 ;
        RECT 1624.360 1110.790 1624.620 1111.110 ;
        RECT 1625.740 1110.790 1626.000 1111.110 ;
        RECT 1625.800 1077.110 1625.940 1110.790 ;
        RECT 1625.740 1076.790 1626.000 1077.110 ;
        RECT 1625.280 1076.110 1625.540 1076.430 ;
        RECT 1625.340 1062.685 1625.480 1076.110 ;
        RECT 1624.350 1062.315 1624.630 1062.685 ;
        RECT 1625.270 1062.315 1625.550 1062.685 ;
        RECT 1624.420 1014.550 1624.560 1062.315 ;
        RECT 1624.360 1014.230 1624.620 1014.550 ;
        RECT 1625.740 1014.230 1626.000 1014.550 ;
        RECT 1625.800 980.550 1625.940 1014.230 ;
        RECT 1625.740 980.230 1626.000 980.550 ;
        RECT 1625.280 979.550 1625.540 979.870 ;
        RECT 1625.340 966.125 1625.480 979.550 ;
        RECT 1624.350 965.755 1624.630 966.125 ;
        RECT 1625.270 965.755 1625.550 966.125 ;
        RECT 1624.420 917.990 1624.560 965.755 ;
        RECT 1624.360 917.670 1624.620 917.990 ;
        RECT 1625.740 917.670 1626.000 917.990 ;
        RECT 1625.800 883.990 1625.940 917.670 ;
        RECT 1625.740 883.670 1626.000 883.990 ;
        RECT 1625.280 882.990 1625.540 883.310 ;
        RECT 1625.340 869.565 1625.480 882.990 ;
        RECT 1624.350 869.195 1624.630 869.565 ;
        RECT 1625.270 869.195 1625.550 869.565 ;
        RECT 1624.420 835.030 1624.560 869.195 ;
        RECT 1624.360 834.710 1624.620 835.030 ;
        RECT 1625.280 834.710 1625.540 835.030 ;
        RECT 1625.340 821.170 1625.480 834.710 ;
        RECT 1625.340 821.030 1625.940 821.170 ;
        RECT 1625.800 787.430 1625.940 821.030 ;
        RECT 1625.740 787.110 1626.000 787.430 ;
        RECT 1625.280 786.090 1625.540 786.410 ;
        RECT 1625.340 772.810 1625.480 786.090 ;
        RECT 1625.280 772.490 1625.540 772.810 ;
        RECT 1626.200 772.490 1626.460 772.810 ;
        RECT 1626.260 724.725 1626.400 772.490 ;
        RECT 1624.810 724.355 1625.090 724.725 ;
        RECT 1626.190 724.355 1626.470 724.725 ;
        RECT 1624.880 690.190 1625.020 724.355 ;
        RECT 1624.820 689.870 1625.080 690.190 ;
        RECT 1625.280 689.530 1625.540 689.850 ;
        RECT 1625.340 676.250 1625.480 689.530 ;
        RECT 1625.280 675.930 1625.540 676.250 ;
        RECT 1626.200 675.930 1626.460 676.250 ;
        RECT 1626.260 628.165 1626.400 675.930 ;
        RECT 1624.810 627.795 1625.090 628.165 ;
        RECT 1626.190 627.795 1626.470 628.165 ;
        RECT 1624.880 593.630 1625.020 627.795 ;
        RECT 1624.820 593.310 1625.080 593.630 ;
        RECT 1625.280 592.970 1625.540 593.290 ;
        RECT 1625.340 579.690 1625.480 592.970 ;
        RECT 1625.280 579.370 1625.540 579.690 ;
        RECT 1626.200 579.370 1626.460 579.690 ;
        RECT 1626.260 531.605 1626.400 579.370 ;
        RECT 1624.810 531.235 1625.090 531.605 ;
        RECT 1626.190 531.235 1626.470 531.605 ;
        RECT 1624.880 507.270 1625.020 531.235 ;
        RECT 1623.900 506.950 1624.160 507.270 ;
        RECT 1624.820 506.950 1625.080 507.270 ;
        RECT 1623.960 448.530 1624.100 506.950 ;
        RECT 1623.960 448.390 1625.020 448.530 ;
        RECT 1624.880 400.510 1625.020 448.390 ;
        RECT 1624.820 400.190 1625.080 400.510 ;
        RECT 1625.280 399.510 1625.540 399.830 ;
        RECT 1625.340 386.230 1625.480 399.510 ;
        RECT 1625.280 385.910 1625.540 386.230 ;
        RECT 1624.820 337.970 1625.080 338.290 ;
        RECT 1624.880 303.690 1625.020 337.970 ;
        RECT 1623.960 303.550 1625.020 303.690 ;
        RECT 1623.960 241.390 1624.100 303.550 ;
        RECT 1622.980 241.070 1623.240 241.390 ;
        RECT 1623.900 241.070 1624.160 241.390 ;
        RECT 1623.040 234.590 1623.180 241.070 ;
        RECT 1622.980 234.270 1623.240 234.590 ;
        RECT 1624.360 192.450 1624.620 192.770 ;
        RECT 1624.420 159.110 1624.560 192.450 ;
        RECT 1624.360 158.790 1624.620 159.110 ;
        RECT 1624.360 158.110 1624.620 158.430 ;
        RECT 1624.420 110.570 1624.560 158.110 ;
        RECT 1624.420 110.430 1625.940 110.570 ;
        RECT 1625.800 109.890 1625.940 110.430 ;
        RECT 1625.800 109.750 1626.860 109.890 ;
        RECT 1626.720 16.650 1626.860 109.750 ;
        RECT 1626.660 16.330 1626.920 16.650 ;
        RECT 1768.800 14.970 1769.060 15.290 ;
        RECT 1768.860 2.400 1769.000 14.970 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
      LAYER via2 ;
        RECT 1624.350 1158.920 1624.630 1159.200 ;
        RECT 1625.270 1158.920 1625.550 1159.200 ;
        RECT 1624.350 1062.360 1624.630 1062.640 ;
        RECT 1625.270 1062.360 1625.550 1062.640 ;
        RECT 1624.350 965.800 1624.630 966.080 ;
        RECT 1625.270 965.800 1625.550 966.080 ;
        RECT 1624.350 869.240 1624.630 869.520 ;
        RECT 1625.270 869.240 1625.550 869.520 ;
        RECT 1624.810 724.400 1625.090 724.680 ;
        RECT 1626.190 724.400 1626.470 724.680 ;
        RECT 1624.810 627.840 1625.090 628.120 ;
        RECT 1626.190 627.840 1626.470 628.120 ;
        RECT 1624.810 531.280 1625.090 531.560 ;
        RECT 1626.190 531.280 1626.470 531.560 ;
      LAYER met3 ;
        RECT 1624.325 1159.210 1624.655 1159.225 ;
        RECT 1625.245 1159.210 1625.575 1159.225 ;
        RECT 1624.325 1158.910 1625.575 1159.210 ;
        RECT 1624.325 1158.895 1624.655 1158.910 ;
        RECT 1625.245 1158.895 1625.575 1158.910 ;
        RECT 1624.325 1062.650 1624.655 1062.665 ;
        RECT 1625.245 1062.650 1625.575 1062.665 ;
        RECT 1624.325 1062.350 1625.575 1062.650 ;
        RECT 1624.325 1062.335 1624.655 1062.350 ;
        RECT 1625.245 1062.335 1625.575 1062.350 ;
        RECT 1624.325 966.090 1624.655 966.105 ;
        RECT 1625.245 966.090 1625.575 966.105 ;
        RECT 1624.325 965.790 1625.575 966.090 ;
        RECT 1624.325 965.775 1624.655 965.790 ;
        RECT 1625.245 965.775 1625.575 965.790 ;
        RECT 1624.325 869.530 1624.655 869.545 ;
        RECT 1625.245 869.530 1625.575 869.545 ;
        RECT 1624.325 869.230 1625.575 869.530 ;
        RECT 1624.325 869.215 1624.655 869.230 ;
        RECT 1625.245 869.215 1625.575 869.230 ;
        RECT 1624.785 724.690 1625.115 724.705 ;
        RECT 1626.165 724.690 1626.495 724.705 ;
        RECT 1624.785 724.390 1626.495 724.690 ;
        RECT 1624.785 724.375 1625.115 724.390 ;
        RECT 1626.165 724.375 1626.495 724.390 ;
        RECT 1624.785 628.130 1625.115 628.145 ;
        RECT 1626.165 628.130 1626.495 628.145 ;
        RECT 1624.785 627.830 1626.495 628.130 ;
        RECT 1624.785 627.815 1625.115 627.830 ;
        RECT 1626.165 627.815 1626.495 627.830 ;
        RECT 1624.785 531.570 1625.115 531.585 ;
        RECT 1626.165 531.570 1626.495 531.585 ;
        RECT 1624.785 531.270 1626.495 531.570 ;
        RECT 1624.785 531.255 1625.115 531.270 ;
        RECT 1626.165 531.255 1626.495 531.270 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 969.290 1588.380 969.610 1588.440 ;
        RECT 972.510 1588.380 972.830 1588.440 ;
        RECT 969.290 1588.240 972.830 1588.380 ;
        RECT 969.290 1588.180 969.610 1588.240 ;
        RECT 972.510 1588.180 972.830 1588.240 ;
        RECT 972.510 19.620 972.830 19.680 ;
        RECT 1786.710 19.620 1787.030 19.680 ;
        RECT 972.510 19.480 1787.030 19.620 ;
        RECT 972.510 19.420 972.830 19.480 ;
        RECT 1786.710 19.420 1787.030 19.480 ;
      LAYER via ;
        RECT 969.320 1588.180 969.580 1588.440 ;
        RECT 972.540 1588.180 972.800 1588.440 ;
        RECT 972.540 19.420 972.800 19.680 ;
        RECT 1786.740 19.420 1787.000 19.680 ;
      LAYER met2 ;
        RECT 969.180 1600.380 969.460 1604.000 ;
        RECT 969.180 1600.000 969.520 1600.380 ;
        RECT 969.380 1588.470 969.520 1600.000 ;
        RECT 969.320 1588.150 969.580 1588.470 ;
        RECT 972.540 1588.150 972.800 1588.470 ;
        RECT 972.600 19.710 972.740 1588.150 ;
        RECT 972.540 19.390 972.800 19.710 ;
        RECT 1786.740 19.390 1787.000 19.710 ;
        RECT 1786.800 2.400 1786.940 19.390 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1789.085 16.745 1789.255 19.635 ;
      LAYER mcon ;
        RECT 1789.085 19.465 1789.255 19.635 ;
      LAYER met1 ;
        RECT 975.270 1593.140 975.590 1593.200 ;
        RECT 1645.490 1593.140 1645.810 1593.200 ;
        RECT 975.270 1593.000 1645.810 1593.140 ;
        RECT 975.270 1592.940 975.590 1593.000 ;
        RECT 1645.490 1592.940 1645.810 1593.000 ;
        RECT 1789.025 19.620 1789.315 19.665 ;
        RECT 1804.650 19.620 1804.970 19.680 ;
        RECT 1789.025 19.480 1804.970 19.620 ;
        RECT 1789.025 19.435 1789.315 19.480 ;
        RECT 1804.650 19.420 1804.970 19.480 ;
        RECT 1645.490 16.900 1645.810 16.960 ;
        RECT 1789.025 16.900 1789.315 16.945 ;
        RECT 1645.490 16.760 1789.315 16.900 ;
        RECT 1645.490 16.700 1645.810 16.760 ;
        RECT 1789.025 16.715 1789.315 16.760 ;
      LAYER via ;
        RECT 975.300 1592.940 975.560 1593.200 ;
        RECT 1645.520 1592.940 1645.780 1593.200 ;
        RECT 1804.680 19.420 1804.940 19.680 ;
        RECT 1645.520 16.700 1645.780 16.960 ;
      LAYER met2 ;
        RECT 975.160 1600.380 975.440 1604.000 ;
        RECT 975.160 1600.000 975.500 1600.380 ;
        RECT 975.360 1593.230 975.500 1600.000 ;
        RECT 975.300 1592.910 975.560 1593.230 ;
        RECT 1645.520 1592.910 1645.780 1593.230 ;
        RECT 1645.580 16.990 1645.720 1592.910 ;
        RECT 1804.680 19.390 1804.940 19.710 ;
        RECT 1645.520 16.670 1645.780 16.990 ;
        RECT 1804.740 2.400 1804.880 19.390 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1246.285 43.265 1246.455 45.475 ;
      LAYER mcon ;
        RECT 1246.285 45.305 1246.455 45.475 ;
      LAYER met1 ;
        RECT 981.710 1588.720 982.030 1588.780 ;
        RECT 985.850 1588.720 986.170 1588.780 ;
        RECT 981.710 1588.580 986.170 1588.720 ;
        RECT 981.710 1588.520 982.030 1588.580 ;
        RECT 985.850 1588.520 986.170 1588.580 ;
        RECT 1246.225 45.460 1246.515 45.505 ;
        RECT 1336.830 45.460 1337.150 45.520 ;
        RECT 1246.225 45.320 1337.150 45.460 ;
        RECT 1246.225 45.275 1246.515 45.320 ;
        RECT 1336.830 45.260 1337.150 45.320 ;
        RECT 1246.225 43.420 1246.515 43.465 ;
        RECT 1231.580 43.280 1246.515 43.420 ;
        RECT 985.850 43.080 986.170 43.140 ;
        RECT 1231.580 43.080 1231.720 43.280 ;
        RECT 1246.225 43.235 1246.515 43.280 ;
        RECT 985.850 42.940 1231.720 43.080 ;
        RECT 985.850 42.880 986.170 42.940 ;
        RECT 1336.830 15.880 1337.150 15.940 ;
        RECT 1822.590 15.880 1822.910 15.940 ;
        RECT 1336.830 15.740 1822.910 15.880 ;
        RECT 1336.830 15.680 1337.150 15.740 ;
        RECT 1822.590 15.680 1822.910 15.740 ;
      LAYER via ;
        RECT 981.740 1588.520 982.000 1588.780 ;
        RECT 985.880 1588.520 986.140 1588.780 ;
        RECT 1336.860 45.260 1337.120 45.520 ;
        RECT 985.880 42.880 986.140 43.140 ;
        RECT 1336.860 15.680 1337.120 15.940 ;
        RECT 1822.620 15.680 1822.880 15.940 ;
      LAYER met2 ;
        RECT 981.600 1600.380 981.880 1604.000 ;
        RECT 981.600 1600.000 981.940 1600.380 ;
        RECT 981.800 1588.810 981.940 1600.000 ;
        RECT 981.740 1588.490 982.000 1588.810 ;
        RECT 985.880 1588.490 986.140 1588.810 ;
        RECT 985.940 43.170 986.080 1588.490 ;
        RECT 1336.860 45.230 1337.120 45.550 ;
        RECT 985.880 42.850 986.140 43.170 ;
        RECT 1336.920 15.970 1337.060 45.230 ;
        RECT 1336.860 15.650 1337.120 15.970 ;
        RECT 1822.620 15.650 1822.880 15.970 ;
        RECT 1822.680 2.400 1822.820 15.650 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1008.005 1592.645 1008.175 1593.495 ;
        RECT 1700.765 19.805 1700.935 20.655 ;
      LAYER mcon ;
        RECT 1008.005 1593.325 1008.175 1593.495 ;
        RECT 1700.765 20.485 1700.935 20.655 ;
      LAYER met1 ;
        RECT 987.690 1593.480 988.010 1593.540 ;
        RECT 1007.945 1593.480 1008.235 1593.525 ;
        RECT 987.690 1593.340 1008.235 1593.480 ;
        RECT 987.690 1593.280 988.010 1593.340 ;
        RECT 1007.945 1593.295 1008.235 1593.340 ;
        RECT 1007.945 1592.800 1008.235 1592.845 ;
        RECT 1659.290 1592.800 1659.610 1592.860 ;
        RECT 1007.945 1592.660 1659.610 1592.800 ;
        RECT 1007.945 1592.615 1008.235 1592.660 ;
        RECT 1659.290 1592.600 1659.610 1592.660 ;
        RECT 1700.705 20.640 1700.995 20.685 ;
        RECT 1725.070 20.640 1725.390 20.700 ;
        RECT 1700.705 20.500 1725.390 20.640 ;
        RECT 1700.705 20.455 1700.995 20.500 ;
        RECT 1725.070 20.440 1725.390 20.500 ;
        RECT 1772.910 20.640 1773.230 20.700 ;
        RECT 1840.070 20.640 1840.390 20.700 ;
        RECT 1772.910 20.500 1840.390 20.640 ;
        RECT 1772.910 20.440 1773.230 20.500 ;
        RECT 1840.070 20.440 1840.390 20.500 ;
        RECT 1659.290 19.960 1659.610 20.020 ;
        RECT 1700.705 19.960 1700.995 20.005 ;
        RECT 1659.290 19.820 1700.995 19.960 ;
        RECT 1659.290 19.760 1659.610 19.820 ;
        RECT 1700.705 19.775 1700.995 19.820 ;
      LAYER via ;
        RECT 987.720 1593.280 987.980 1593.540 ;
        RECT 1659.320 1592.600 1659.580 1592.860 ;
        RECT 1725.100 20.440 1725.360 20.700 ;
        RECT 1772.940 20.440 1773.200 20.700 ;
        RECT 1840.100 20.440 1840.360 20.700 ;
        RECT 1659.320 19.760 1659.580 20.020 ;
      LAYER met2 ;
        RECT 987.580 1600.380 987.860 1604.000 ;
        RECT 987.580 1600.000 987.920 1600.380 ;
        RECT 987.780 1593.570 987.920 1600.000 ;
        RECT 987.720 1593.250 987.980 1593.570 ;
        RECT 1659.320 1592.570 1659.580 1592.890 ;
        RECT 1659.380 20.050 1659.520 1592.570 ;
        RECT 1725.090 20.555 1725.370 20.925 ;
        RECT 1772.930 20.555 1773.210 20.925 ;
        RECT 1725.100 20.410 1725.360 20.555 ;
        RECT 1772.940 20.410 1773.200 20.555 ;
        RECT 1840.100 20.410 1840.360 20.730 ;
        RECT 1659.320 19.730 1659.580 20.050 ;
        RECT 1840.160 2.400 1840.300 20.410 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
      LAYER via2 ;
        RECT 1725.090 20.600 1725.370 20.880 ;
        RECT 1772.930 20.600 1773.210 20.880 ;
      LAYER met3 ;
        RECT 1725.065 20.890 1725.395 20.905 ;
        RECT 1772.905 20.890 1773.235 20.905 ;
        RECT 1725.065 20.590 1773.235 20.890 ;
        RECT 1725.065 20.575 1725.395 20.590 ;
        RECT 1772.905 20.575 1773.235 20.590 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 994.130 1588.720 994.450 1588.780 ;
        RECT 1000.110 1588.720 1000.430 1588.780 ;
        RECT 994.130 1588.580 1000.430 1588.720 ;
        RECT 994.130 1588.520 994.450 1588.580 ;
        RECT 1000.110 1588.520 1000.430 1588.580 ;
        RECT 1000.110 19.280 1000.430 19.340 ;
        RECT 1858.010 19.280 1858.330 19.340 ;
        RECT 1000.110 19.140 1858.330 19.280 ;
        RECT 1000.110 19.080 1000.430 19.140 ;
        RECT 1858.010 19.080 1858.330 19.140 ;
      LAYER via ;
        RECT 994.160 1588.520 994.420 1588.780 ;
        RECT 1000.140 1588.520 1000.400 1588.780 ;
        RECT 1000.140 19.080 1000.400 19.340 ;
        RECT 1858.040 19.080 1858.300 19.340 ;
      LAYER met2 ;
        RECT 994.020 1600.380 994.300 1604.000 ;
        RECT 994.020 1600.000 994.360 1600.380 ;
        RECT 994.220 1588.810 994.360 1600.000 ;
        RECT 994.160 1588.490 994.420 1588.810 ;
        RECT 1000.140 1588.490 1000.400 1588.810 ;
        RECT 1000.200 19.370 1000.340 1588.490 ;
        RECT 1000.140 19.050 1000.400 19.370 ;
        RECT 1858.040 19.050 1858.300 19.370 ;
        RECT 1858.100 2.400 1858.240 19.050 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1000.110 1591.440 1000.430 1591.500 ;
        RECT 1679.990 1591.440 1680.310 1591.500 ;
        RECT 1000.110 1591.300 1680.310 1591.440 ;
        RECT 1000.110 1591.240 1000.430 1591.300 ;
        RECT 1679.990 1591.240 1680.310 1591.300 ;
        RECT 1679.990 20.300 1680.310 20.360 ;
        RECT 1824.430 20.300 1824.750 20.360 ;
        RECT 1679.990 20.160 1824.750 20.300 ;
        RECT 1679.990 20.100 1680.310 20.160 ;
        RECT 1824.430 20.100 1824.750 20.160 ;
        RECT 1835.010 15.880 1835.330 15.940 ;
        RECT 1875.950 15.880 1876.270 15.940 ;
        RECT 1835.010 15.740 1876.270 15.880 ;
        RECT 1835.010 15.680 1835.330 15.740 ;
        RECT 1875.950 15.680 1876.270 15.740 ;
      LAYER via ;
        RECT 1000.140 1591.240 1000.400 1591.500 ;
        RECT 1680.020 1591.240 1680.280 1591.500 ;
        RECT 1680.020 20.100 1680.280 20.360 ;
        RECT 1824.460 20.100 1824.720 20.360 ;
        RECT 1835.040 15.680 1835.300 15.940 ;
        RECT 1875.980 15.680 1876.240 15.940 ;
      LAYER met2 ;
        RECT 1000.000 1600.380 1000.280 1604.000 ;
        RECT 1000.000 1600.000 1000.340 1600.380 ;
        RECT 1000.200 1591.530 1000.340 1600.000 ;
        RECT 1000.140 1591.210 1000.400 1591.530 ;
        RECT 1680.020 1591.210 1680.280 1591.530 ;
        RECT 1680.080 20.390 1680.220 1591.210 ;
        RECT 1680.020 20.070 1680.280 20.390 ;
        RECT 1824.460 20.245 1824.720 20.390 ;
        RECT 1824.450 19.875 1824.730 20.245 ;
        RECT 1835.030 19.875 1835.310 20.245 ;
        RECT 1835.100 15.970 1835.240 19.875 ;
        RECT 1835.040 15.650 1835.300 15.970 ;
        RECT 1875.980 15.650 1876.240 15.970 ;
        RECT 1876.040 2.400 1876.180 15.650 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
      LAYER via2 ;
        RECT 1824.450 19.920 1824.730 20.200 ;
        RECT 1835.030 19.920 1835.310 20.200 ;
      LAYER met3 ;
        RECT 1824.425 20.210 1824.755 20.225 ;
        RECT 1835.005 20.210 1835.335 20.225 ;
        RECT 1824.425 19.910 1835.335 20.210 ;
        RECT 1824.425 19.895 1824.755 19.910 ;
        RECT 1835.005 19.895 1835.335 19.910 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 610.490 1589.060 610.810 1589.120 ;
        RECT 613.710 1589.060 614.030 1589.120 ;
        RECT 610.490 1588.920 614.030 1589.060 ;
        RECT 610.490 1588.860 610.810 1588.920 ;
        RECT 613.710 1588.860 614.030 1588.920 ;
        RECT 613.710 15.880 614.030 15.940 ;
        RECT 752.170 15.880 752.490 15.940 ;
        RECT 613.710 15.740 752.490 15.880 ;
        RECT 613.710 15.680 614.030 15.740 ;
        RECT 752.170 15.680 752.490 15.740 ;
      LAYER via ;
        RECT 610.520 1588.860 610.780 1589.120 ;
        RECT 613.740 1588.860 614.000 1589.120 ;
        RECT 613.740 15.680 614.000 15.940 ;
        RECT 752.200 15.680 752.460 15.940 ;
      LAYER met2 ;
        RECT 610.380 1600.380 610.660 1604.000 ;
        RECT 610.380 1600.000 610.720 1600.380 ;
        RECT 610.580 1589.150 610.720 1600.000 ;
        RECT 610.520 1588.830 610.780 1589.150 ;
        RECT 613.740 1588.830 614.000 1589.150 ;
        RECT 613.800 15.970 613.940 1588.830 ;
        RECT 613.740 15.650 614.000 15.970 ;
        RECT 752.200 15.650 752.460 15.970 ;
        RECT 752.260 2.400 752.400 15.650 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 18.940 1007.330 19.000 ;
        RECT 1893.890 18.940 1894.210 19.000 ;
        RECT 1007.010 18.800 1894.210 18.940 ;
        RECT 1007.010 18.740 1007.330 18.800 ;
        RECT 1893.890 18.740 1894.210 18.800 ;
      LAYER via ;
        RECT 1007.040 18.740 1007.300 19.000 ;
        RECT 1893.920 18.740 1894.180 19.000 ;
      LAYER met2 ;
        RECT 1006.440 1600.450 1006.720 1604.000 ;
        RECT 1006.440 1600.310 1007.240 1600.450 ;
        RECT 1006.440 1600.000 1006.720 1600.310 ;
        RECT 1007.100 19.030 1007.240 1600.310 ;
        RECT 1007.040 18.710 1007.300 19.030 ;
        RECT 1893.920 18.710 1894.180 19.030 ;
        RECT 1893.980 2.400 1894.120 18.710 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1052.165 1590.265 1052.335 1591.795 ;
      LAYER mcon ;
        RECT 1052.165 1591.625 1052.335 1591.795 ;
      LAYER met1 ;
        RECT 1012.530 1591.780 1012.850 1591.840 ;
        RECT 1052.105 1591.780 1052.395 1591.825 ;
        RECT 1012.530 1591.640 1052.395 1591.780 ;
        RECT 1012.530 1591.580 1012.850 1591.640 ;
        RECT 1052.105 1591.595 1052.395 1591.640 ;
        RECT 1052.105 1590.420 1052.395 1590.465 ;
        RECT 1700.690 1590.420 1701.010 1590.480 ;
        RECT 1052.105 1590.280 1701.010 1590.420 ;
        RECT 1052.105 1590.235 1052.395 1590.280 ;
        RECT 1700.690 1590.220 1701.010 1590.280 ;
        RECT 1701.150 19.960 1701.470 20.020 ;
        RECT 1911.370 19.960 1911.690 20.020 ;
        RECT 1701.150 19.820 1911.690 19.960 ;
        RECT 1701.150 19.760 1701.470 19.820 ;
        RECT 1911.370 19.760 1911.690 19.820 ;
      LAYER via ;
        RECT 1012.560 1591.580 1012.820 1591.840 ;
        RECT 1700.720 1590.220 1700.980 1590.480 ;
        RECT 1701.180 19.760 1701.440 20.020 ;
        RECT 1911.400 19.760 1911.660 20.020 ;
      LAYER met2 ;
        RECT 1012.420 1600.380 1012.700 1604.000 ;
        RECT 1012.420 1600.000 1012.760 1600.380 ;
        RECT 1012.620 1591.870 1012.760 1600.000 ;
        RECT 1012.560 1591.550 1012.820 1591.870 ;
        RECT 1700.720 1590.190 1700.980 1590.510 ;
        RECT 1700.780 26.930 1700.920 1590.190 ;
        RECT 1700.780 26.790 1701.380 26.930 ;
        RECT 1701.240 20.050 1701.380 26.790 ;
        RECT 1701.180 19.730 1701.440 20.050 ;
        RECT 1911.400 19.730 1911.660 20.050 ;
        RECT 1911.460 18.090 1911.600 19.730 ;
        RECT 1911.460 17.950 1912.060 18.090 ;
        RECT 1911.920 2.400 1912.060 17.950 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1018.970 1587.360 1019.290 1587.420 ;
        RECT 1020.810 1587.360 1021.130 1587.420 ;
        RECT 1018.970 1587.220 1021.130 1587.360 ;
        RECT 1018.970 1587.160 1019.290 1587.220 ;
        RECT 1020.810 1587.160 1021.130 1587.220 ;
        RECT 1020.810 18.600 1021.130 18.660 ;
        RECT 1929.310 18.600 1929.630 18.660 ;
        RECT 1020.810 18.460 1929.630 18.600 ;
        RECT 1020.810 18.400 1021.130 18.460 ;
        RECT 1929.310 18.400 1929.630 18.460 ;
      LAYER via ;
        RECT 1019.000 1587.160 1019.260 1587.420 ;
        RECT 1020.840 1587.160 1021.100 1587.420 ;
        RECT 1020.840 18.400 1021.100 18.660 ;
        RECT 1929.340 18.400 1929.600 18.660 ;
      LAYER met2 ;
        RECT 1018.860 1600.380 1019.140 1604.000 ;
        RECT 1018.860 1600.000 1019.200 1600.380 ;
        RECT 1019.060 1587.450 1019.200 1600.000 ;
        RECT 1019.000 1587.130 1019.260 1587.450 ;
        RECT 1020.840 1587.130 1021.100 1587.450 ;
        RECT 1020.900 18.690 1021.040 1587.130 ;
        RECT 1020.840 18.370 1021.100 18.690 ;
        RECT 1929.340 18.370 1929.600 18.690 ;
        RECT 1929.400 2.400 1929.540 18.370 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1042.965 1589.925 1043.135 1593.835 ;
        RECT 1052.625 1589.925 1052.795 1591.795 ;
        RECT 1060.445 1590.605 1060.615 1591.795 ;
        RECT 1076.085 1590.605 1076.255 1593.495 ;
        RECT 1111.045 1590.605 1111.215 1593.495 ;
      LAYER mcon ;
        RECT 1042.965 1593.665 1043.135 1593.835 ;
        RECT 1076.085 1593.325 1076.255 1593.495 ;
        RECT 1052.625 1591.625 1052.795 1591.795 ;
        RECT 1060.445 1591.625 1060.615 1591.795 ;
        RECT 1111.045 1593.325 1111.215 1593.495 ;
      LAYER met1 ;
        RECT 1024.950 1593.820 1025.270 1593.880 ;
        RECT 1042.905 1593.820 1043.195 1593.865 ;
        RECT 1024.950 1593.680 1043.195 1593.820 ;
        RECT 1024.950 1593.620 1025.270 1593.680 ;
        RECT 1042.905 1593.635 1043.195 1593.680 ;
        RECT 1076.025 1593.480 1076.315 1593.525 ;
        RECT 1110.985 1593.480 1111.275 1593.525 ;
        RECT 1076.025 1593.340 1111.275 1593.480 ;
        RECT 1076.025 1593.295 1076.315 1593.340 ;
        RECT 1110.985 1593.295 1111.275 1593.340 ;
        RECT 1052.565 1591.780 1052.855 1591.825 ;
        RECT 1060.385 1591.780 1060.675 1591.825 ;
        RECT 1052.565 1591.640 1060.675 1591.780 ;
        RECT 1052.565 1591.595 1052.855 1591.640 ;
        RECT 1060.385 1591.595 1060.675 1591.640 ;
        RECT 1060.385 1590.760 1060.675 1590.805 ;
        RECT 1076.025 1590.760 1076.315 1590.805 ;
        RECT 1060.385 1590.620 1076.315 1590.760 ;
        RECT 1060.385 1590.575 1060.675 1590.620 ;
        RECT 1076.025 1590.575 1076.315 1590.620 ;
        RECT 1110.985 1590.760 1111.275 1590.805 ;
        RECT 1714.490 1590.760 1714.810 1590.820 ;
        RECT 1110.985 1590.620 1714.810 1590.760 ;
        RECT 1110.985 1590.575 1111.275 1590.620 ;
        RECT 1714.490 1590.560 1714.810 1590.620 ;
        RECT 1042.905 1590.080 1043.195 1590.125 ;
        RECT 1052.565 1590.080 1052.855 1590.125 ;
        RECT 1042.905 1589.940 1052.855 1590.080 ;
        RECT 1042.905 1589.895 1043.195 1589.940 ;
        RECT 1052.565 1589.895 1052.855 1589.940 ;
        RECT 1714.490 14.520 1714.810 14.580 ;
        RECT 1714.490 14.380 1716.100 14.520 ;
        RECT 1714.490 14.320 1714.810 14.380 ;
        RECT 1715.960 14.180 1716.100 14.380 ;
        RECT 1947.250 14.180 1947.570 14.240 ;
        RECT 1715.960 14.040 1947.570 14.180 ;
        RECT 1947.250 13.980 1947.570 14.040 ;
      LAYER via ;
        RECT 1024.980 1593.620 1025.240 1593.880 ;
        RECT 1714.520 1590.560 1714.780 1590.820 ;
        RECT 1714.520 14.320 1714.780 14.580 ;
        RECT 1947.280 13.980 1947.540 14.240 ;
      LAYER met2 ;
        RECT 1024.840 1600.380 1025.120 1604.000 ;
        RECT 1024.840 1600.000 1025.180 1600.380 ;
        RECT 1025.040 1593.910 1025.180 1600.000 ;
        RECT 1024.980 1593.590 1025.240 1593.910 ;
        RECT 1714.520 1590.530 1714.780 1590.850 ;
        RECT 1714.580 14.610 1714.720 1590.530 ;
        RECT 1714.520 14.290 1714.780 14.610 ;
        RECT 1947.280 13.950 1947.540 14.270 ;
        RECT 1947.340 2.400 1947.480 13.950 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1030.930 1590.080 1031.250 1590.140 ;
        RECT 1033.230 1590.080 1033.550 1590.140 ;
        RECT 1030.930 1589.940 1033.550 1590.080 ;
        RECT 1030.930 1589.880 1031.250 1589.940 ;
        RECT 1033.230 1589.880 1033.550 1589.940 ;
        RECT 1033.690 80.480 1034.010 80.540 ;
        RECT 1959.670 80.480 1959.990 80.540 ;
        RECT 1033.690 80.340 1959.990 80.480 ;
        RECT 1033.690 80.280 1034.010 80.340 ;
        RECT 1959.670 80.280 1959.990 80.340 ;
      LAYER via ;
        RECT 1030.960 1589.880 1031.220 1590.140 ;
        RECT 1033.260 1589.880 1033.520 1590.140 ;
        RECT 1033.720 80.280 1033.980 80.540 ;
        RECT 1959.700 80.280 1959.960 80.540 ;
      LAYER met2 ;
        RECT 1030.820 1600.380 1031.100 1604.000 ;
        RECT 1030.820 1600.000 1031.160 1600.380 ;
        RECT 1031.020 1590.170 1031.160 1600.000 ;
        RECT 1030.960 1589.850 1031.220 1590.170 ;
        RECT 1033.260 1589.850 1033.520 1590.170 ;
        RECT 1033.320 1578.690 1033.460 1589.850 ;
        RECT 1033.320 1578.550 1033.920 1578.690 ;
        RECT 1033.780 80.570 1033.920 1578.550 ;
        RECT 1033.720 80.250 1033.980 80.570 ;
        RECT 1959.700 80.250 1959.960 80.570 ;
        RECT 1959.760 16.730 1959.900 80.250 ;
        RECT 1959.760 16.590 1965.420 16.730 ;
        RECT 1965.280 2.400 1965.420 16.590 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1037.370 1590.080 1037.690 1590.140 ;
        RECT 1041.050 1590.080 1041.370 1590.140 ;
        RECT 1037.370 1589.940 1041.370 1590.080 ;
        RECT 1037.370 1589.880 1037.690 1589.940 ;
        RECT 1041.050 1589.880 1041.370 1589.940 ;
        RECT 1041.510 18.260 1041.830 18.320 ;
        RECT 1983.130 18.260 1983.450 18.320 ;
        RECT 1041.510 18.120 1983.450 18.260 ;
        RECT 1041.510 18.060 1041.830 18.120 ;
        RECT 1983.130 18.060 1983.450 18.120 ;
      LAYER via ;
        RECT 1037.400 1589.880 1037.660 1590.140 ;
        RECT 1041.080 1589.880 1041.340 1590.140 ;
        RECT 1041.540 18.060 1041.800 18.320 ;
        RECT 1983.160 18.060 1983.420 18.320 ;
      LAYER met2 ;
        RECT 1037.260 1600.380 1037.540 1604.000 ;
        RECT 1037.260 1600.000 1037.600 1600.380 ;
        RECT 1037.460 1590.170 1037.600 1600.000 ;
        RECT 1037.400 1589.850 1037.660 1590.170 ;
        RECT 1041.080 1589.850 1041.340 1590.170 ;
        RECT 1041.140 1580.730 1041.280 1589.850 ;
        RECT 1041.140 1580.590 1041.740 1580.730 ;
        RECT 1041.600 18.350 1041.740 1580.590 ;
        RECT 1041.540 18.030 1041.800 18.350 ;
        RECT 1983.160 18.030 1983.420 18.350 ;
        RECT 1983.220 2.400 1983.360 18.030 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1069.185 1587.205 1069.355 1593.835 ;
      LAYER mcon ;
        RECT 1069.185 1593.665 1069.355 1593.835 ;
      LAYER met1 ;
        RECT 1043.350 1593.820 1043.670 1593.880 ;
        RECT 1069.125 1593.820 1069.415 1593.865 ;
        RECT 1043.350 1593.680 1069.415 1593.820 ;
        RECT 1043.350 1593.620 1043.670 1593.680 ;
        RECT 1069.125 1593.635 1069.415 1593.680 ;
        RECT 1069.125 1587.360 1069.415 1587.405 ;
        RECT 1383.290 1587.360 1383.610 1587.420 ;
        RECT 1069.125 1587.220 1383.610 1587.360 ;
        RECT 1069.125 1587.175 1069.415 1587.220 ;
        RECT 1383.290 1587.160 1383.610 1587.220 ;
        RECT 1383.290 16.220 1383.610 16.280 ;
        RECT 2001.070 16.220 2001.390 16.280 ;
        RECT 1383.290 16.080 2001.390 16.220 ;
        RECT 1383.290 16.020 1383.610 16.080 ;
        RECT 2001.070 16.020 2001.390 16.080 ;
      LAYER via ;
        RECT 1043.380 1593.620 1043.640 1593.880 ;
        RECT 1383.320 1587.160 1383.580 1587.420 ;
        RECT 1383.320 16.020 1383.580 16.280 ;
        RECT 2001.100 16.020 2001.360 16.280 ;
      LAYER met2 ;
        RECT 1043.240 1600.380 1043.520 1604.000 ;
        RECT 1043.240 1600.000 1043.580 1600.380 ;
        RECT 1043.440 1593.910 1043.580 1600.000 ;
        RECT 1043.380 1593.590 1043.640 1593.910 ;
        RECT 1383.320 1587.130 1383.580 1587.450 ;
        RECT 1383.380 16.310 1383.520 1587.130 ;
        RECT 1383.320 15.990 1383.580 16.310 ;
        RECT 2001.100 15.990 2001.360 16.310 ;
        RECT 2001.160 2.400 2001.300 15.990 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1741.705 13.685 1741.875 14.875 ;
        RECT 1751.825 13.685 1751.995 15.555 ;
        RECT 1769.305 14.535 1769.475 15.555 ;
        RECT 1769.305 14.365 1770.395 14.535 ;
      LAYER mcon ;
        RECT 1751.825 15.385 1751.995 15.555 ;
        RECT 1741.705 14.705 1741.875 14.875 ;
        RECT 1769.305 15.385 1769.475 15.555 ;
        RECT 1770.225 14.365 1770.395 14.535 ;
      LAYER met1 ;
        RECT 1049.790 1592.120 1050.110 1592.180 ;
        RECT 1049.790 1591.980 1061.980 1592.120 ;
        RECT 1049.790 1591.920 1050.110 1591.980 ;
        RECT 1061.840 1591.780 1061.980 1591.980 ;
        RECT 1728.290 1591.780 1728.610 1591.840 ;
        RECT 1061.840 1591.640 1728.610 1591.780 ;
        RECT 1728.290 1591.580 1728.610 1591.640 ;
        RECT 1751.765 15.540 1752.055 15.585 ;
        RECT 1769.245 15.540 1769.535 15.585 ;
        RECT 1751.765 15.400 1769.535 15.540 ;
        RECT 1751.765 15.355 1752.055 15.400 ;
        RECT 1769.245 15.355 1769.535 15.400 ;
        RECT 1728.290 14.860 1728.610 14.920 ;
        RECT 1741.645 14.860 1741.935 14.905 ;
        RECT 1728.290 14.720 1741.935 14.860 ;
        RECT 1728.290 14.660 1728.610 14.720 ;
        RECT 1741.645 14.675 1741.935 14.720 ;
        RECT 1770.165 14.520 1770.455 14.565 ;
        RECT 2018.550 14.520 2018.870 14.580 ;
        RECT 1770.165 14.380 2018.870 14.520 ;
        RECT 1770.165 14.335 1770.455 14.380 ;
        RECT 2018.550 14.320 2018.870 14.380 ;
        RECT 1741.645 13.840 1741.935 13.885 ;
        RECT 1751.765 13.840 1752.055 13.885 ;
        RECT 1741.645 13.700 1752.055 13.840 ;
        RECT 1741.645 13.655 1741.935 13.700 ;
        RECT 1751.765 13.655 1752.055 13.700 ;
      LAYER via ;
        RECT 1049.820 1591.920 1050.080 1592.180 ;
        RECT 1728.320 1591.580 1728.580 1591.840 ;
        RECT 1728.320 14.660 1728.580 14.920 ;
        RECT 2018.580 14.320 2018.840 14.580 ;
      LAYER met2 ;
        RECT 1049.680 1600.380 1049.960 1604.000 ;
        RECT 1049.680 1600.000 1050.020 1600.380 ;
        RECT 1049.880 1592.210 1050.020 1600.000 ;
        RECT 1049.820 1591.890 1050.080 1592.210 ;
        RECT 1728.320 1591.550 1728.580 1591.870 ;
        RECT 1728.380 14.950 1728.520 1591.550 ;
        RECT 1728.320 14.630 1728.580 14.950 ;
        RECT 2018.580 14.290 2018.840 14.610 ;
        RECT 2018.640 2.400 2018.780 14.290 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1055.770 1587.360 1056.090 1587.420 ;
        RECT 1060.370 1587.360 1060.690 1587.420 ;
        RECT 1055.770 1587.220 1060.690 1587.360 ;
        RECT 1055.770 1587.160 1056.090 1587.220 ;
        RECT 1060.370 1587.160 1060.690 1587.220 ;
        RECT 1061.290 80.140 1061.610 80.200 ;
        RECT 2035.570 80.140 2035.890 80.200 ;
        RECT 1061.290 80.000 2035.890 80.140 ;
        RECT 1061.290 79.940 1061.610 80.000 ;
        RECT 2035.570 79.940 2035.890 80.000 ;
      LAYER via ;
        RECT 1055.800 1587.160 1056.060 1587.420 ;
        RECT 1060.400 1587.160 1060.660 1587.420 ;
        RECT 1061.320 79.940 1061.580 80.200 ;
        RECT 2035.600 79.940 2035.860 80.200 ;
      LAYER met2 ;
        RECT 1055.660 1600.380 1055.940 1604.000 ;
        RECT 1055.660 1600.000 1056.000 1600.380 ;
        RECT 1055.860 1587.450 1056.000 1600.000 ;
        RECT 1055.800 1587.130 1056.060 1587.450 ;
        RECT 1060.400 1587.130 1060.660 1587.450 ;
        RECT 1060.460 1579.370 1060.600 1587.130 ;
        RECT 1060.460 1579.230 1061.520 1579.370 ;
        RECT 1061.380 80.230 1061.520 1579.230 ;
        RECT 1061.320 79.910 1061.580 80.230 ;
        RECT 2035.600 79.910 2035.860 80.230 ;
        RECT 2035.660 17.410 2035.800 79.910 ;
        RECT 2035.660 17.270 2036.720 17.410 ;
        RECT 2036.580 2.400 2036.720 17.270 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1062.210 1592.120 1062.530 1592.180 ;
        RECT 1735.190 1592.120 1735.510 1592.180 ;
        RECT 1062.210 1591.980 1735.510 1592.120 ;
        RECT 1062.210 1591.920 1062.530 1591.980 ;
        RECT 1735.190 1591.920 1735.510 1591.980 ;
        RECT 2054.430 14.860 2054.750 14.920 ;
        RECT 1769.780 14.720 2054.750 14.860 ;
        RECT 1735.190 14.520 1735.510 14.580 ;
        RECT 1769.780 14.520 1769.920 14.720 ;
        RECT 2054.430 14.660 2054.750 14.720 ;
        RECT 1735.190 14.380 1769.920 14.520 ;
        RECT 1735.190 14.320 1735.510 14.380 ;
      LAYER via ;
        RECT 1062.240 1591.920 1062.500 1592.180 ;
        RECT 1735.220 1591.920 1735.480 1592.180 ;
        RECT 1735.220 14.320 1735.480 14.580 ;
        RECT 2054.460 14.660 2054.720 14.920 ;
      LAYER met2 ;
        RECT 1062.100 1600.380 1062.380 1604.000 ;
        RECT 1062.100 1600.000 1062.440 1600.380 ;
        RECT 1062.300 1592.210 1062.440 1600.000 ;
        RECT 1062.240 1591.890 1062.500 1592.210 ;
        RECT 1735.220 1591.890 1735.480 1592.210 ;
        RECT 1735.280 14.610 1735.420 1591.890 ;
        RECT 2054.460 14.630 2054.720 14.950 ;
        RECT 1735.220 14.290 1735.480 14.610 ;
        RECT 2054.520 2.400 2054.660 14.630 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 639.085 16.065 639.255 18.275 ;
      LAYER mcon ;
        RECT 639.085 18.105 639.255 18.275 ;
      LAYER met1 ;
        RECT 616.930 1588.720 617.250 1588.780 ;
        RECT 620.150 1588.720 620.470 1588.780 ;
        RECT 616.930 1588.580 620.470 1588.720 ;
        RECT 616.930 1588.520 617.250 1588.580 ;
        RECT 620.150 1588.520 620.470 1588.580 ;
        RECT 639.025 18.260 639.315 18.305 ;
        RECT 769.650 18.260 769.970 18.320 ;
        RECT 639.025 18.120 769.970 18.260 ;
        RECT 639.025 18.075 639.315 18.120 ;
        RECT 769.650 18.060 769.970 18.120 ;
        RECT 620.150 16.220 620.470 16.280 ;
        RECT 639.025 16.220 639.315 16.265 ;
        RECT 620.150 16.080 639.315 16.220 ;
        RECT 620.150 16.020 620.470 16.080 ;
        RECT 639.025 16.035 639.315 16.080 ;
      LAYER via ;
        RECT 616.960 1588.520 617.220 1588.780 ;
        RECT 620.180 1588.520 620.440 1588.780 ;
        RECT 769.680 18.060 769.940 18.320 ;
        RECT 620.180 16.020 620.440 16.280 ;
      LAYER met2 ;
        RECT 616.820 1600.380 617.100 1604.000 ;
        RECT 616.820 1600.000 617.160 1600.380 ;
        RECT 617.020 1588.810 617.160 1600.000 ;
        RECT 616.960 1588.490 617.220 1588.810 ;
        RECT 620.180 1588.490 620.440 1588.810 ;
        RECT 620.240 16.310 620.380 1588.490 ;
        RECT 769.680 18.030 769.940 18.350 ;
        RECT 620.180 15.990 620.440 16.310 ;
        RECT 769.740 2.400 769.880 18.030 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1069.110 17.920 1069.430 17.980 ;
        RECT 2072.370 17.920 2072.690 17.980 ;
        RECT 1069.110 17.780 2072.690 17.920 ;
        RECT 1069.110 17.720 1069.430 17.780 ;
        RECT 2072.370 17.720 2072.690 17.780 ;
      LAYER via ;
        RECT 1069.140 17.720 1069.400 17.980 ;
        RECT 2072.400 17.720 2072.660 17.980 ;
      LAYER met2 ;
        RECT 1068.080 1600.450 1068.360 1604.000 ;
        RECT 1068.080 1600.310 1069.340 1600.450 ;
        RECT 1068.080 1600.000 1068.360 1600.310 ;
        RECT 1069.200 18.010 1069.340 1600.310 ;
        RECT 1069.140 17.690 1069.400 18.010 ;
        RECT 2072.400 17.690 2072.660 18.010 ;
        RECT 2072.460 2.400 2072.600 17.690 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1100.465 1592.305 1100.635 1593.835 ;
        RECT 1745.845 14.705 1746.015 16.575 ;
        RECT 1797.825 15.045 1797.995 16.915 ;
      LAYER mcon ;
        RECT 1100.465 1593.665 1100.635 1593.835 ;
        RECT 1797.825 16.745 1797.995 16.915 ;
        RECT 1745.845 16.405 1746.015 16.575 ;
      LAYER met1 ;
        RECT 1074.630 1593.820 1074.950 1593.880 ;
        RECT 1100.405 1593.820 1100.695 1593.865 ;
        RECT 1074.630 1593.680 1100.695 1593.820 ;
        RECT 1074.630 1593.620 1074.950 1593.680 ;
        RECT 1100.405 1593.635 1100.695 1593.680 ;
        RECT 1100.405 1592.460 1100.695 1592.505 ;
        RECT 1742.090 1592.460 1742.410 1592.520 ;
        RECT 1100.405 1592.320 1742.410 1592.460 ;
        RECT 1100.405 1592.275 1100.695 1592.320 ;
        RECT 1742.090 1592.260 1742.410 1592.320 ;
        RECT 1797.765 16.900 1798.055 16.945 ;
        RECT 1796.460 16.760 1798.055 16.900 ;
        RECT 1745.785 16.560 1746.075 16.605 ;
        RECT 1796.460 16.560 1796.600 16.760 ;
        RECT 1797.765 16.715 1798.055 16.760 ;
        RECT 1745.785 16.420 1796.600 16.560 ;
        RECT 1745.785 16.375 1746.075 16.420 ;
        RECT 1797.765 15.200 1798.055 15.245 ;
        RECT 2089.850 15.200 2090.170 15.260 ;
        RECT 1797.765 15.060 2090.170 15.200 ;
        RECT 1797.765 15.015 1798.055 15.060 ;
        RECT 2089.850 15.000 2090.170 15.060 ;
        RECT 1742.090 14.860 1742.410 14.920 ;
        RECT 1745.785 14.860 1746.075 14.905 ;
        RECT 1742.090 14.720 1746.075 14.860 ;
        RECT 1742.090 14.660 1742.410 14.720 ;
        RECT 1745.785 14.675 1746.075 14.720 ;
      LAYER via ;
        RECT 1074.660 1593.620 1074.920 1593.880 ;
        RECT 1742.120 1592.260 1742.380 1592.520 ;
        RECT 2089.880 15.000 2090.140 15.260 ;
        RECT 1742.120 14.660 1742.380 14.920 ;
      LAYER met2 ;
        RECT 1074.520 1600.380 1074.800 1604.000 ;
        RECT 1074.520 1600.000 1074.860 1600.380 ;
        RECT 1074.720 1593.910 1074.860 1600.000 ;
        RECT 1074.660 1593.590 1074.920 1593.910 ;
        RECT 1742.120 1592.230 1742.380 1592.550 ;
        RECT 1742.180 14.950 1742.320 1592.230 ;
        RECT 2089.880 14.970 2090.140 15.290 ;
        RECT 1742.120 14.630 1742.380 14.950 ;
        RECT 2089.940 2.400 2090.080 14.970 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1081.530 79.800 1081.850 79.860 ;
        RECT 2104.570 79.800 2104.890 79.860 ;
        RECT 1081.530 79.660 2104.890 79.800 ;
        RECT 1081.530 79.600 1081.850 79.660 ;
        RECT 2104.570 79.600 2104.890 79.660 ;
        RECT 2104.570 2.960 2104.890 3.020 ;
        RECT 2107.790 2.960 2108.110 3.020 ;
        RECT 2104.570 2.820 2108.110 2.960 ;
        RECT 2104.570 2.760 2104.890 2.820 ;
        RECT 2107.790 2.760 2108.110 2.820 ;
      LAYER via ;
        RECT 1081.560 79.600 1081.820 79.860 ;
        RECT 2104.600 79.600 2104.860 79.860 ;
        RECT 2104.600 2.760 2104.860 3.020 ;
        RECT 2107.820 2.760 2108.080 3.020 ;
      LAYER met2 ;
        RECT 1080.500 1600.450 1080.780 1604.000 ;
        RECT 1080.500 1600.310 1081.760 1600.450 ;
        RECT 1080.500 1600.000 1080.780 1600.310 ;
        RECT 1081.620 79.890 1081.760 1600.310 ;
        RECT 1081.560 79.570 1081.820 79.890 ;
        RECT 2104.600 79.570 2104.860 79.890 ;
        RECT 2104.660 3.050 2104.800 79.570 ;
        RECT 2104.600 2.730 2104.860 3.050 ;
        RECT 2107.820 2.730 2108.080 3.050 ;
        RECT 2107.880 2.400 2108.020 2.730 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1100.005 1590.945 1100.175 1592.475 ;
        RECT 1124.385 1591.115 1124.555 1593.835 ;
        RECT 1124.845 1593.665 1125.015 1594.515 ;
        RECT 1123.465 1590.945 1124.555 1591.115 ;
        RECT 1171.765 1589.925 1171.935 1594.515 ;
      LAYER mcon ;
        RECT 1124.845 1594.345 1125.015 1594.515 ;
        RECT 1124.385 1593.665 1124.555 1593.835 ;
        RECT 1171.765 1594.345 1171.935 1594.515 ;
        RECT 1100.005 1592.305 1100.175 1592.475 ;
      LAYER met1 ;
        RECT 1124.785 1594.500 1125.075 1594.545 ;
        RECT 1171.705 1594.500 1171.995 1594.545 ;
        RECT 1124.785 1594.360 1171.995 1594.500 ;
        RECT 1124.785 1594.315 1125.075 1594.360 ;
        RECT 1171.705 1594.315 1171.995 1594.360 ;
        RECT 1124.325 1593.820 1124.615 1593.865 ;
        RECT 1124.785 1593.820 1125.075 1593.865 ;
        RECT 1124.325 1593.680 1125.075 1593.820 ;
        RECT 1124.325 1593.635 1124.615 1593.680 ;
        RECT 1124.785 1593.635 1125.075 1593.680 ;
        RECT 1086.590 1592.460 1086.910 1592.520 ;
        RECT 1099.945 1592.460 1100.235 1592.505 ;
        RECT 1086.590 1592.320 1100.235 1592.460 ;
        RECT 1086.590 1592.260 1086.910 1592.320 ;
        RECT 1099.945 1592.275 1100.235 1592.320 ;
        RECT 1099.945 1591.100 1100.235 1591.145 ;
        RECT 1123.405 1591.100 1123.695 1591.145 ;
        RECT 1099.945 1590.960 1123.695 1591.100 ;
        RECT 1099.945 1590.915 1100.235 1590.960 ;
        RECT 1123.405 1590.915 1123.695 1590.960 ;
        RECT 1171.705 1590.080 1171.995 1590.125 ;
        RECT 1748.990 1590.080 1749.310 1590.140 ;
        RECT 1171.705 1589.940 1749.310 1590.080 ;
        RECT 1171.705 1589.895 1171.995 1589.940 ;
        RECT 1748.990 1589.880 1749.310 1589.940 ;
        RECT 2125.730 15.540 2126.050 15.600 ;
        RECT 1797.380 15.400 2126.050 15.540 ;
        RECT 1797.380 15.200 1797.520 15.400 ;
        RECT 2125.730 15.340 2126.050 15.400 ;
        RECT 1769.320 15.060 1797.520 15.200 ;
        RECT 1748.990 14.860 1749.310 14.920 ;
        RECT 1769.320 14.860 1769.460 15.060 ;
        RECT 1748.990 14.720 1769.460 14.860 ;
        RECT 1748.990 14.660 1749.310 14.720 ;
      LAYER via ;
        RECT 1086.620 1592.260 1086.880 1592.520 ;
        RECT 1749.020 1589.880 1749.280 1590.140 ;
        RECT 2125.760 15.340 2126.020 15.600 ;
        RECT 1749.020 14.660 1749.280 14.920 ;
      LAYER met2 ;
        RECT 1086.480 1600.380 1086.760 1604.000 ;
        RECT 1086.480 1600.000 1086.820 1600.380 ;
        RECT 1086.680 1592.550 1086.820 1600.000 ;
        RECT 1086.620 1592.230 1086.880 1592.550 ;
        RECT 1749.020 1589.850 1749.280 1590.170 ;
        RECT 1749.080 14.950 1749.220 1589.850 ;
        RECT 2125.760 15.310 2126.020 15.630 ;
        RECT 1749.020 14.630 1749.280 14.950 ;
        RECT 2125.820 2.400 2125.960 15.310 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1093.030 1590.760 1093.350 1590.820 ;
        RECT 1096.710 1590.760 1097.030 1590.820 ;
        RECT 1093.030 1590.620 1097.030 1590.760 ;
        RECT 1093.030 1590.560 1093.350 1590.620 ;
        RECT 1096.710 1590.560 1097.030 1590.620 ;
        RECT 1095.330 82.860 1095.650 82.920 ;
        RECT 1096.710 82.860 1097.030 82.920 ;
        RECT 1095.330 82.720 1097.030 82.860 ;
        RECT 1095.330 82.660 1095.650 82.720 ;
        RECT 1096.710 82.660 1097.030 82.720 ;
        RECT 1095.790 17.580 1096.110 17.640 ;
        RECT 2143.670 17.580 2143.990 17.640 ;
        RECT 1095.790 17.440 2143.990 17.580 ;
        RECT 1095.790 17.380 1096.110 17.440 ;
        RECT 2143.670 17.380 2143.990 17.440 ;
      LAYER via ;
        RECT 1093.060 1590.560 1093.320 1590.820 ;
        RECT 1096.740 1590.560 1097.000 1590.820 ;
        RECT 1095.360 82.660 1095.620 82.920 ;
        RECT 1096.740 82.660 1097.000 82.920 ;
        RECT 1095.820 17.380 1096.080 17.640 ;
        RECT 2143.700 17.380 2143.960 17.640 ;
      LAYER met2 ;
        RECT 1092.920 1600.380 1093.200 1604.000 ;
        RECT 1092.920 1600.000 1093.260 1600.380 ;
        RECT 1093.120 1590.850 1093.260 1600.000 ;
        RECT 1093.060 1590.530 1093.320 1590.850 ;
        RECT 1096.740 1590.530 1097.000 1590.850 ;
        RECT 1096.800 82.950 1096.940 1590.530 ;
        RECT 1095.360 82.630 1095.620 82.950 ;
        RECT 1096.740 82.630 1097.000 82.950 ;
        RECT 1095.420 39.170 1095.560 82.630 ;
        RECT 1095.420 39.030 1096.020 39.170 ;
        RECT 1095.880 17.670 1096.020 39.030 ;
        RECT 1095.820 17.350 1096.080 17.670 ;
        RECT 2143.700 17.350 2143.960 17.670 ;
        RECT 2143.760 2.400 2143.900 17.350 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1796.905 15.385 1797.075 16.575 ;
      LAYER mcon ;
        RECT 1796.905 16.405 1797.075 16.575 ;
      LAYER met1 ;
        RECT 1123.940 1594.020 1125.460 1594.160 ;
        RECT 1100.850 1593.820 1101.170 1593.880 ;
        RECT 1123.940 1593.820 1124.080 1594.020 ;
        RECT 1100.850 1593.680 1124.080 1593.820 ;
        RECT 1125.320 1593.820 1125.460 1594.020 ;
        RECT 1769.690 1593.820 1770.010 1593.880 ;
        RECT 1125.320 1593.680 1770.010 1593.820 ;
        RECT 1100.850 1593.620 1101.170 1593.680 ;
        RECT 1769.690 1593.620 1770.010 1593.680 ;
        RECT 1796.845 16.560 1797.135 16.605 ;
        RECT 2161.610 16.560 2161.930 16.620 ;
        RECT 1796.845 16.420 2161.930 16.560 ;
        RECT 1796.845 16.375 1797.135 16.420 ;
        RECT 2161.610 16.360 2161.930 16.420 ;
        RECT 1769.690 15.540 1770.010 15.600 ;
        RECT 1796.845 15.540 1797.135 15.585 ;
        RECT 1769.690 15.400 1797.135 15.540 ;
        RECT 1769.690 15.340 1770.010 15.400 ;
        RECT 1796.845 15.355 1797.135 15.400 ;
      LAYER via ;
        RECT 1100.880 1593.620 1101.140 1593.880 ;
        RECT 1769.720 1593.620 1769.980 1593.880 ;
        RECT 2161.640 16.360 2161.900 16.620 ;
        RECT 1769.720 15.340 1769.980 15.600 ;
      LAYER met2 ;
        RECT 1098.900 1600.450 1099.180 1604.000 ;
        RECT 1098.900 1600.310 1100.620 1600.450 ;
        RECT 1098.900 1600.000 1099.180 1600.310 ;
        RECT 1100.480 1593.820 1100.620 1600.310 ;
        RECT 1100.880 1593.820 1101.140 1593.910 ;
        RECT 1100.480 1593.680 1101.140 1593.820 ;
        RECT 1100.880 1593.590 1101.140 1593.680 ;
        RECT 1769.720 1593.590 1769.980 1593.910 ;
        RECT 1769.780 15.630 1769.920 1593.590 ;
        RECT 2161.640 16.330 2161.900 16.650 ;
        RECT 1769.720 15.310 1769.980 15.630 ;
        RECT 2161.700 2.400 2161.840 16.330 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1105.450 1590.760 1105.770 1590.820 ;
        RECT 1110.510 1590.760 1110.830 1590.820 ;
        RECT 1105.450 1590.620 1110.830 1590.760 ;
        RECT 1105.450 1590.560 1105.770 1590.620 ;
        RECT 1110.510 1590.560 1110.830 1590.620 ;
        RECT 1110.510 17.240 1110.830 17.300 ;
        RECT 2179.090 17.240 2179.410 17.300 ;
        RECT 1110.510 17.100 2179.410 17.240 ;
        RECT 1110.510 17.040 1110.830 17.100 ;
        RECT 2179.090 17.040 2179.410 17.100 ;
      LAYER via ;
        RECT 1105.480 1590.560 1105.740 1590.820 ;
        RECT 1110.540 1590.560 1110.800 1590.820 ;
        RECT 1110.540 17.040 1110.800 17.300 ;
        RECT 2179.120 17.040 2179.380 17.300 ;
      LAYER met2 ;
        RECT 1105.340 1600.380 1105.620 1604.000 ;
        RECT 1105.340 1600.000 1105.680 1600.380 ;
        RECT 1105.540 1590.850 1105.680 1600.000 ;
        RECT 1105.480 1590.530 1105.740 1590.850 ;
        RECT 1110.540 1590.530 1110.800 1590.850 ;
        RECT 1110.600 17.330 1110.740 1590.530 ;
        RECT 1110.540 17.010 1110.800 17.330 ;
        RECT 2179.120 17.010 2179.380 17.330 ;
        RECT 2179.180 2.400 2179.320 17.010 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1111.430 1593.480 1111.750 1593.540 ;
        RECT 1783.490 1593.480 1783.810 1593.540 ;
        RECT 1111.430 1593.340 1783.810 1593.480 ;
        RECT 1111.430 1593.280 1111.750 1593.340 ;
        RECT 1783.490 1593.280 1783.810 1593.340 ;
        RECT 1798.210 16.900 1798.530 16.960 ;
        RECT 2197.030 16.900 2197.350 16.960 ;
        RECT 1798.210 16.760 2197.350 16.900 ;
        RECT 1798.210 16.700 1798.530 16.760 ;
        RECT 2197.030 16.700 2197.350 16.760 ;
      LAYER via ;
        RECT 1111.460 1593.280 1111.720 1593.540 ;
        RECT 1783.520 1593.280 1783.780 1593.540 ;
        RECT 1798.240 16.700 1798.500 16.960 ;
        RECT 2197.060 16.700 2197.320 16.960 ;
      LAYER met2 ;
        RECT 1111.320 1600.380 1111.600 1604.000 ;
        RECT 1111.320 1600.000 1111.660 1600.380 ;
        RECT 1111.520 1593.570 1111.660 1600.000 ;
        RECT 1111.460 1593.250 1111.720 1593.570 ;
        RECT 1783.520 1593.250 1783.780 1593.570 ;
        RECT 1783.580 16.165 1783.720 1593.250 ;
        RECT 1798.240 16.670 1798.500 16.990 ;
        RECT 2197.060 16.670 2197.320 16.990 ;
        RECT 1798.300 16.165 1798.440 16.670 ;
        RECT 1783.510 15.795 1783.790 16.165 ;
        RECT 1798.230 15.795 1798.510 16.165 ;
        RECT 2197.120 2.400 2197.260 16.670 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
      LAYER via2 ;
        RECT 1783.510 15.840 1783.790 16.120 ;
        RECT 1798.230 15.840 1798.510 16.120 ;
      LAYER met3 ;
        RECT 1783.485 16.130 1783.815 16.145 ;
        RECT 1798.205 16.130 1798.535 16.145 ;
        RECT 1783.485 15.830 1798.535 16.130 ;
        RECT 1783.485 15.815 1783.815 15.830 ;
        RECT 1798.205 15.815 1798.535 15.830 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1118.330 1556.080 1118.650 1556.140 ;
        RECT 1124.310 1556.080 1124.630 1556.140 ;
        RECT 1118.330 1555.940 1124.630 1556.080 ;
        RECT 1118.330 1555.880 1118.650 1555.940 ;
        RECT 1124.310 1555.880 1124.630 1555.940 ;
      LAYER via ;
        RECT 1118.360 1555.880 1118.620 1556.140 ;
        RECT 1124.340 1555.880 1124.600 1556.140 ;
      LAYER met2 ;
        RECT 1117.760 1600.450 1118.040 1604.000 ;
        RECT 1117.760 1600.310 1118.560 1600.450 ;
        RECT 1117.760 1600.000 1118.040 1600.310 ;
        RECT 1118.420 1556.170 1118.560 1600.310 ;
        RECT 1118.360 1555.850 1118.620 1556.170 ;
        RECT 1124.340 1555.850 1124.600 1556.170 ;
        RECT 1124.400 19.565 1124.540 1555.850 ;
        RECT 1124.330 19.195 1124.610 19.565 ;
        RECT 2214.990 19.195 2215.270 19.565 ;
        RECT 2215.060 2.400 2215.200 19.195 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
      LAYER via2 ;
        RECT 1124.330 19.240 1124.610 19.520 ;
        RECT 2214.990 19.240 2215.270 19.520 ;
      LAYER met3 ;
        RECT 1124.305 19.530 1124.635 19.545 ;
        RECT 2214.965 19.530 2215.295 19.545 ;
        RECT 1124.305 19.230 2215.295 19.530 ;
        RECT 1124.305 19.215 1124.635 19.230 ;
        RECT 2214.965 19.215 2215.295 19.230 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1123.850 1591.100 1124.170 1591.160 ;
        RECT 1804.190 1591.100 1804.510 1591.160 ;
        RECT 1123.850 1590.960 1804.510 1591.100 ;
        RECT 1123.850 1590.900 1124.170 1590.960 ;
        RECT 1804.190 1590.900 1804.510 1590.960 ;
        RECT 1845.590 20.640 1845.910 20.700 ;
        RECT 2232.910 20.640 2233.230 20.700 ;
        RECT 1845.590 20.500 2233.230 20.640 ;
        RECT 1845.590 20.440 1845.910 20.500 ;
        RECT 2232.910 20.440 2233.230 20.500 ;
        RECT 1805.110 19.620 1805.430 19.680 ;
        RECT 1845.590 19.620 1845.910 19.680 ;
        RECT 1805.110 19.480 1845.910 19.620 ;
        RECT 1805.110 19.420 1805.430 19.480 ;
        RECT 1845.590 19.420 1845.910 19.480 ;
      LAYER via ;
        RECT 1123.880 1590.900 1124.140 1591.160 ;
        RECT 1804.220 1590.900 1804.480 1591.160 ;
        RECT 1845.620 20.440 1845.880 20.700 ;
        RECT 2232.940 20.440 2233.200 20.700 ;
        RECT 1805.140 19.420 1805.400 19.680 ;
        RECT 1845.620 19.420 1845.880 19.680 ;
      LAYER met2 ;
        RECT 1123.740 1600.380 1124.020 1604.000 ;
        RECT 1123.740 1600.000 1124.080 1600.380 ;
        RECT 1123.940 1591.190 1124.080 1600.000 ;
        RECT 1123.880 1590.870 1124.140 1591.190 ;
        RECT 1804.220 1590.870 1804.480 1591.190 ;
        RECT 1804.280 26.930 1804.420 1590.870 ;
        RECT 1804.280 26.790 1805.340 26.930 ;
        RECT 1805.200 19.710 1805.340 26.790 ;
        RECT 1845.620 20.410 1845.880 20.730 ;
        RECT 2232.940 20.410 2233.200 20.730 ;
        RECT 1845.680 19.710 1845.820 20.410 ;
        RECT 1805.140 19.390 1805.400 19.710 ;
        RECT 1845.620 19.390 1845.880 19.710 ;
        RECT 2233.000 2.400 2233.140 20.410 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 622.910 1589.740 623.230 1589.800 ;
        RECT 627.510 1589.740 627.830 1589.800 ;
        RECT 622.910 1589.600 627.830 1589.740 ;
        RECT 622.910 1589.540 623.230 1589.600 ;
        RECT 627.510 1589.540 627.830 1589.600 ;
        RECT 627.510 16.900 627.830 16.960 ;
        RECT 627.510 16.760 638.780 16.900 ;
        RECT 627.510 16.700 627.830 16.760 ;
        RECT 638.640 16.560 638.780 16.760 ;
        RECT 787.590 16.560 787.910 16.620 ;
        RECT 638.640 16.420 787.910 16.560 ;
        RECT 787.590 16.360 787.910 16.420 ;
      LAYER via ;
        RECT 622.940 1589.540 623.200 1589.800 ;
        RECT 627.540 1589.540 627.800 1589.800 ;
        RECT 627.540 16.700 627.800 16.960 ;
        RECT 787.620 16.360 787.880 16.620 ;
      LAYER met2 ;
        RECT 622.800 1600.380 623.080 1604.000 ;
        RECT 622.800 1600.000 623.140 1600.380 ;
        RECT 623.000 1589.830 623.140 1600.000 ;
        RECT 622.940 1589.510 623.200 1589.830 ;
        RECT 627.540 1589.510 627.800 1589.830 ;
        RECT 627.600 16.990 627.740 1589.510 ;
        RECT 627.540 16.670 627.800 16.990 ;
        RECT 787.620 16.330 787.880 16.650 ;
        RECT 787.680 2.400 787.820 16.330 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1130.180 1600.450 1130.460 1604.000 ;
        RECT 1130.180 1600.310 1131.440 1600.450 ;
        RECT 1130.180 1600.000 1130.460 1600.310 ;
        RECT 1131.300 18.885 1131.440 1600.310 ;
        RECT 1131.230 18.515 1131.510 18.885 ;
        RECT 2250.870 18.515 2251.150 18.885 ;
        RECT 2250.940 2.400 2251.080 18.515 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
      LAYER via2 ;
        RECT 1131.230 18.560 1131.510 18.840 ;
        RECT 2250.870 18.560 2251.150 18.840 ;
      LAYER met3 ;
        RECT 1131.205 18.850 1131.535 18.865 ;
        RECT 2250.845 18.850 2251.175 18.865 ;
        RECT 1131.205 18.550 2251.175 18.850 ;
        RECT 1131.205 18.535 1131.535 18.550 ;
        RECT 2250.845 18.535 2251.175 18.550 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.890 20.300 1825.210 20.360 ;
        RECT 2268.330 20.300 2268.650 20.360 ;
        RECT 1824.890 20.160 2268.650 20.300 ;
        RECT 1824.890 20.100 1825.210 20.160 ;
        RECT 2268.330 20.100 2268.650 20.160 ;
      LAYER via ;
        RECT 1824.920 20.100 1825.180 20.360 ;
        RECT 2268.360 20.100 2268.620 20.360 ;
      LAYER met2 ;
        RECT 1136.160 1600.380 1136.440 1604.000 ;
        RECT 1136.160 1600.000 1136.500 1600.380 ;
        RECT 1136.360 1591.045 1136.500 1600.000 ;
        RECT 1136.290 1590.675 1136.570 1591.045 ;
        RECT 1824.910 1590.675 1825.190 1591.045 ;
        RECT 1824.980 20.390 1825.120 1590.675 ;
        RECT 1824.920 20.070 1825.180 20.390 ;
        RECT 2268.360 20.070 2268.620 20.390 ;
        RECT 2268.420 2.400 2268.560 20.070 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
      LAYER via2 ;
        RECT 1136.290 1590.720 1136.570 1591.000 ;
        RECT 1824.910 1590.720 1825.190 1591.000 ;
      LAYER met3 ;
        RECT 1136.265 1591.010 1136.595 1591.025 ;
        RECT 1824.885 1591.010 1825.215 1591.025 ;
        RECT 1136.265 1590.710 1825.215 1591.010 ;
        RECT 1136.265 1590.695 1136.595 1590.710 ;
        RECT 1824.885 1590.695 1825.215 1590.710 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1143.630 1579.880 1143.950 1579.940 ;
        RECT 1145.010 1579.880 1145.330 1579.940 ;
        RECT 1143.630 1579.740 1145.330 1579.880 ;
        RECT 1143.630 1579.680 1143.950 1579.740 ;
        RECT 1145.010 1579.680 1145.330 1579.740 ;
      LAYER via ;
        RECT 1143.660 1579.680 1143.920 1579.940 ;
        RECT 1145.040 1579.680 1145.300 1579.940 ;
      LAYER met2 ;
        RECT 1142.140 1600.450 1142.420 1604.000 ;
        RECT 1142.140 1600.310 1143.860 1600.450 ;
        RECT 1142.140 1600.000 1142.420 1600.310 ;
        RECT 1143.720 1579.970 1143.860 1600.310 ;
        RECT 1143.660 1579.650 1143.920 1579.970 ;
        RECT 1145.040 1579.650 1145.300 1579.970 ;
        RECT 1145.100 18.205 1145.240 1579.650 ;
        RECT 1145.030 17.835 1145.310 18.205 ;
        RECT 2286.290 17.835 2286.570 18.205 ;
        RECT 2286.360 2.400 2286.500 17.835 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
      LAYER via2 ;
        RECT 1145.030 17.880 1145.310 18.160 ;
        RECT 2286.290 17.880 2286.570 18.160 ;
      LAYER met3 ;
        RECT 1145.005 18.170 1145.335 18.185 ;
        RECT 2286.265 18.170 2286.595 18.185 ;
        RECT 1145.005 17.870 2286.595 18.170 ;
        RECT 1145.005 17.855 1145.335 17.870 ;
        RECT 2286.265 17.855 2286.595 17.870 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1845.205 19.635 1845.375 20.655 ;
        RECT 1845.205 19.465 1846.295 19.635 ;
        RECT 1893.505 15.725 1893.675 19.295 ;
      LAYER mcon ;
        RECT 1845.205 20.485 1845.375 20.655 ;
        RECT 1846.125 19.465 1846.295 19.635 ;
        RECT 1893.505 19.125 1893.675 19.295 ;
      LAYER met1 ;
        RECT 1838.690 27.780 1839.010 27.840 ;
        RECT 1840.990 27.780 1841.310 27.840 ;
        RECT 1838.690 27.640 1841.310 27.780 ;
        RECT 1838.690 27.580 1839.010 27.640 ;
        RECT 1840.990 27.580 1841.310 27.640 ;
        RECT 1840.990 20.640 1841.310 20.700 ;
        RECT 1845.145 20.640 1845.435 20.685 ;
        RECT 1840.990 20.500 1845.435 20.640 ;
        RECT 1840.990 20.440 1841.310 20.500 ;
        RECT 1845.145 20.455 1845.435 20.500 ;
        RECT 1846.065 19.620 1846.355 19.665 ;
        RECT 1846.065 19.480 1858.700 19.620 ;
        RECT 1846.065 19.435 1846.355 19.480 ;
        RECT 1858.560 19.280 1858.700 19.480 ;
        RECT 1893.445 19.280 1893.735 19.325 ;
        RECT 1858.560 19.140 1893.735 19.280 ;
        RECT 1893.445 19.095 1893.735 19.140 ;
        RECT 1893.445 15.880 1893.735 15.925 ;
        RECT 2304.210 15.880 2304.530 15.940 ;
        RECT 1893.445 15.740 2304.530 15.880 ;
        RECT 1893.445 15.695 1893.735 15.740 ;
        RECT 2304.210 15.680 2304.530 15.740 ;
      LAYER via ;
        RECT 1838.720 27.580 1838.980 27.840 ;
        RECT 1841.020 27.580 1841.280 27.840 ;
        RECT 1841.020 20.440 1841.280 20.700 ;
        RECT 2304.240 15.680 2304.500 15.940 ;
      LAYER met2 ;
        RECT 1148.580 1600.380 1148.860 1604.000 ;
        RECT 1148.580 1600.000 1148.920 1600.380 ;
        RECT 1148.780 1593.085 1148.920 1600.000 ;
        RECT 1148.710 1592.715 1148.990 1593.085 ;
        RECT 1838.710 1592.035 1838.990 1592.405 ;
        RECT 1838.780 27.870 1838.920 1592.035 ;
        RECT 1838.720 27.550 1838.980 27.870 ;
        RECT 1841.020 27.550 1841.280 27.870 ;
        RECT 1841.080 20.730 1841.220 27.550 ;
        RECT 1841.020 20.410 1841.280 20.730 ;
        RECT 2304.240 15.650 2304.500 15.970 ;
        RECT 2304.300 2.400 2304.440 15.650 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
      LAYER via2 ;
        RECT 1148.710 1592.760 1148.990 1593.040 ;
        RECT 1838.710 1592.080 1838.990 1592.360 ;
      LAYER met3 ;
        RECT 1148.685 1593.050 1149.015 1593.065 ;
        RECT 1148.685 1592.750 1185.570 1593.050 ;
        RECT 1148.685 1592.735 1149.015 1592.750 ;
        RECT 1185.270 1592.370 1185.570 1592.750 ;
        RECT 1838.685 1592.370 1839.015 1592.385 ;
        RECT 1185.270 1592.070 1839.015 1592.370 ;
        RECT 1838.685 1592.055 1839.015 1592.070 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1153.750 1535.000 1154.070 1535.060 ;
        RECT 1158.810 1535.000 1159.130 1535.060 ;
        RECT 1153.750 1534.860 1159.130 1535.000 ;
        RECT 1153.750 1534.800 1154.070 1534.860 ;
        RECT 1158.810 1534.800 1159.130 1534.860 ;
      LAYER via ;
        RECT 1153.780 1534.800 1154.040 1535.060 ;
        RECT 1158.840 1534.800 1159.100 1535.060 ;
      LAYER met2 ;
        RECT 1154.560 1600.450 1154.840 1604.000 ;
        RECT 1153.840 1600.310 1154.840 1600.450 ;
        RECT 1153.840 1535.090 1153.980 1600.310 ;
        RECT 1154.560 1600.000 1154.840 1600.310 ;
        RECT 1153.780 1534.770 1154.040 1535.090 ;
        RECT 1158.840 1534.770 1159.100 1535.090 ;
        RECT 1158.900 17.525 1159.040 1534.770 ;
        RECT 1158.830 17.155 1159.110 17.525 ;
        RECT 2322.170 17.155 2322.450 17.525 ;
        RECT 2322.240 2.400 2322.380 17.155 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
      LAYER via2 ;
        RECT 1158.830 17.200 1159.110 17.480 ;
        RECT 2322.170 17.200 2322.450 17.480 ;
      LAYER met3 ;
        RECT 1158.805 17.490 1159.135 17.505 ;
        RECT 2322.145 17.490 2322.475 17.505 ;
        RECT 1158.805 17.190 2322.475 17.490 ;
        RECT 1158.805 17.175 1159.135 17.190 ;
        RECT 2322.145 17.175 2322.475 17.190 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1859.390 19.620 1859.710 19.680 ;
        RECT 2339.630 19.620 2339.950 19.680 ;
        RECT 1859.390 19.480 2339.950 19.620 ;
        RECT 1859.390 19.420 1859.710 19.480 ;
        RECT 2339.630 19.420 2339.950 19.480 ;
      LAYER via ;
        RECT 1859.420 19.420 1859.680 19.680 ;
        RECT 2339.660 19.420 2339.920 19.680 ;
      LAYER met2 ;
        RECT 1161.000 1600.380 1161.280 1604.000 ;
        RECT 1161.000 1600.000 1161.340 1600.380 ;
        RECT 1161.200 1590.365 1161.340 1600.000 ;
        RECT 1161.130 1589.995 1161.410 1590.365 ;
        RECT 1859.410 1589.995 1859.690 1590.365 ;
        RECT 1859.480 19.710 1859.620 1589.995 ;
        RECT 1859.420 19.390 1859.680 19.710 ;
        RECT 2339.660 19.390 2339.920 19.710 ;
        RECT 2339.720 2.400 2339.860 19.390 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
      LAYER via2 ;
        RECT 1161.130 1590.040 1161.410 1590.320 ;
        RECT 1859.410 1590.040 1859.690 1590.320 ;
      LAYER met3 ;
        RECT 1161.105 1590.330 1161.435 1590.345 ;
        RECT 1859.385 1590.330 1859.715 1590.345 ;
        RECT 1161.105 1590.030 1859.715 1590.330 ;
        RECT 1161.105 1590.015 1161.435 1590.030 ;
        RECT 1859.385 1590.015 1859.715 1590.030 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1166.170 1535.340 1166.490 1535.400 ;
        RECT 1172.610 1535.340 1172.930 1535.400 ;
        RECT 1166.170 1535.200 1172.930 1535.340 ;
        RECT 1166.170 1535.140 1166.490 1535.200 ;
        RECT 1172.610 1535.140 1172.930 1535.200 ;
      LAYER via ;
        RECT 1166.200 1535.140 1166.460 1535.400 ;
        RECT 1172.640 1535.140 1172.900 1535.400 ;
      LAYER met2 ;
        RECT 1166.980 1600.450 1167.260 1604.000 ;
        RECT 1166.260 1600.310 1167.260 1600.450 ;
        RECT 1166.260 1535.430 1166.400 1600.310 ;
        RECT 1166.980 1600.000 1167.260 1600.310 ;
        RECT 1166.200 1535.110 1166.460 1535.430 ;
        RECT 1172.640 1535.110 1172.900 1535.430 ;
        RECT 1172.700 16.845 1172.840 1535.110 ;
        RECT 1172.630 16.475 1172.910 16.845 ;
        RECT 2357.590 16.475 2357.870 16.845 ;
        RECT 2357.660 2.400 2357.800 16.475 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
      LAYER via2 ;
        RECT 1172.630 16.520 1172.910 16.800 ;
        RECT 2357.590 16.520 2357.870 16.800 ;
      LAYER met3 ;
        RECT 1172.605 16.810 1172.935 16.825 ;
        RECT 2357.565 16.810 2357.895 16.825 ;
        RECT 1172.605 16.510 2357.895 16.810 ;
        RECT 1172.605 16.495 1172.935 16.510 ;
        RECT 2357.565 16.495 2357.895 16.510 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1173.420 1600.380 1173.700 1604.000 ;
        RECT 1173.420 1600.000 1173.760 1600.380 ;
        RECT 1173.620 1591.725 1173.760 1600.000 ;
        RECT 1173.550 1591.355 1173.830 1591.725 ;
        RECT 1866.310 1591.355 1866.590 1591.725 ;
        RECT 1866.380 20.245 1866.520 1591.355 ;
        RECT 1866.310 19.875 1866.590 20.245 ;
        RECT 2375.530 19.875 2375.810 20.245 ;
        RECT 2375.600 2.400 2375.740 19.875 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
      LAYER via2 ;
        RECT 1173.550 1591.400 1173.830 1591.680 ;
        RECT 1866.310 1591.400 1866.590 1591.680 ;
        RECT 1866.310 19.920 1866.590 20.200 ;
        RECT 2375.530 19.920 2375.810 20.200 ;
      LAYER met3 ;
        RECT 1173.525 1591.690 1173.855 1591.705 ;
        RECT 1866.285 1591.690 1866.615 1591.705 ;
        RECT 1173.525 1591.390 1866.615 1591.690 ;
        RECT 1173.525 1591.375 1173.855 1591.390 ;
        RECT 1866.285 1591.375 1866.615 1591.390 ;
        RECT 1866.285 20.210 1866.615 20.225 ;
        RECT 2375.505 20.210 2375.835 20.225 ;
        RECT 1866.285 19.910 2375.835 20.210 ;
        RECT 1866.285 19.895 1866.615 19.910 ;
        RECT 2375.505 19.895 2375.835 19.910 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1178.665 1435.565 1178.835 1483.335 ;
        RECT 1177.745 1000.705 1177.915 1048.815 ;
        RECT 1178.205 855.525 1178.375 903.975 ;
        RECT 1178.665 434.945 1178.835 483.055 ;
        RECT 1178.665 338.045 1178.835 386.155 ;
        RECT 1178.665 241.485 1178.835 289.595 ;
        RECT 1178.665 144.925 1178.835 193.035 ;
        RECT 1178.665 79.305 1178.835 96.475 ;
      LAYER mcon ;
        RECT 1178.665 1483.165 1178.835 1483.335 ;
        RECT 1177.745 1048.645 1177.915 1048.815 ;
        RECT 1178.205 903.805 1178.375 903.975 ;
        RECT 1178.665 482.885 1178.835 483.055 ;
        RECT 1178.665 385.985 1178.835 386.155 ;
        RECT 1178.665 289.425 1178.835 289.595 ;
        RECT 1178.665 192.865 1178.835 193.035 ;
        RECT 1178.665 96.305 1178.835 96.475 ;
      LAYER met1 ;
        RECT 1174.450 1580.220 1174.770 1580.280 ;
        RECT 1178.130 1580.220 1178.450 1580.280 ;
        RECT 1174.450 1580.080 1178.450 1580.220 ;
        RECT 1174.450 1580.020 1174.770 1580.080 ;
        RECT 1178.130 1580.020 1178.450 1580.080 ;
        RECT 1174.450 1484.000 1174.770 1484.060 ;
        RECT 1178.590 1484.000 1178.910 1484.060 ;
        RECT 1174.450 1483.860 1178.910 1484.000 ;
        RECT 1174.450 1483.800 1174.770 1483.860 ;
        RECT 1178.590 1483.800 1178.910 1483.860 ;
        RECT 1178.590 1483.320 1178.910 1483.380 ;
        RECT 1178.395 1483.180 1178.910 1483.320 ;
        RECT 1178.590 1483.120 1178.910 1483.180 ;
        RECT 1178.590 1435.720 1178.910 1435.780 ;
        RECT 1178.395 1435.580 1178.910 1435.720 ;
        RECT 1178.590 1435.520 1178.910 1435.580 ;
        RECT 1177.685 1048.800 1177.975 1048.845 ;
        RECT 1178.590 1048.800 1178.910 1048.860 ;
        RECT 1177.685 1048.660 1178.910 1048.800 ;
        RECT 1177.685 1048.615 1177.975 1048.660 ;
        RECT 1178.590 1048.600 1178.910 1048.660 ;
        RECT 1177.670 1000.860 1177.990 1000.920 ;
        RECT 1177.475 1000.720 1177.990 1000.860 ;
        RECT 1177.670 1000.660 1177.990 1000.720 ;
        RECT 1178.145 903.960 1178.435 904.005 ;
        RECT 1178.590 903.960 1178.910 904.020 ;
        RECT 1178.145 903.820 1178.910 903.960 ;
        RECT 1178.145 903.775 1178.435 903.820 ;
        RECT 1178.590 903.760 1178.910 903.820 ;
        RECT 1178.130 855.680 1178.450 855.740 ;
        RECT 1177.935 855.540 1178.450 855.680 ;
        RECT 1178.130 855.480 1178.450 855.540 ;
        RECT 1178.590 483.040 1178.910 483.100 ;
        RECT 1178.395 482.900 1178.910 483.040 ;
        RECT 1178.590 482.840 1178.910 482.900 ;
        RECT 1178.590 435.100 1178.910 435.160 ;
        RECT 1178.395 434.960 1178.910 435.100 ;
        RECT 1178.590 434.900 1178.910 434.960 ;
        RECT 1178.590 386.140 1178.910 386.200 ;
        RECT 1178.395 386.000 1178.910 386.140 ;
        RECT 1178.590 385.940 1178.910 386.000 ;
        RECT 1178.590 338.200 1178.910 338.260 ;
        RECT 1178.395 338.060 1178.910 338.200 ;
        RECT 1178.590 338.000 1178.910 338.060 ;
        RECT 1178.590 289.580 1178.910 289.640 ;
        RECT 1178.395 289.440 1178.910 289.580 ;
        RECT 1178.590 289.380 1178.910 289.440 ;
        RECT 1178.590 241.640 1178.910 241.700 ;
        RECT 1178.395 241.500 1178.910 241.640 ;
        RECT 1178.590 241.440 1178.910 241.500 ;
        RECT 1178.590 193.020 1178.910 193.080 ;
        RECT 1178.395 192.880 1178.910 193.020 ;
        RECT 1178.590 192.820 1178.910 192.880 ;
        RECT 1178.590 145.080 1178.910 145.140 ;
        RECT 1178.395 144.940 1178.910 145.080 ;
        RECT 1178.590 144.880 1178.910 144.940 ;
        RECT 1178.590 96.460 1178.910 96.520 ;
        RECT 1178.395 96.320 1178.910 96.460 ;
        RECT 1178.590 96.260 1178.910 96.320 ;
        RECT 1178.605 79.460 1178.895 79.505 ;
        RECT 2387.470 79.460 2387.790 79.520 ;
        RECT 1178.605 79.320 2387.790 79.460 ;
        RECT 1178.605 79.275 1178.895 79.320 ;
        RECT 2387.470 79.260 2387.790 79.320 ;
        RECT 2387.470 17.920 2387.790 17.980 ;
        RECT 2393.450 17.920 2393.770 17.980 ;
        RECT 2387.470 17.780 2393.770 17.920 ;
        RECT 2387.470 17.720 2387.790 17.780 ;
        RECT 2393.450 17.720 2393.770 17.780 ;
      LAYER via ;
        RECT 1174.480 1580.020 1174.740 1580.280 ;
        RECT 1178.160 1580.020 1178.420 1580.280 ;
        RECT 1174.480 1483.800 1174.740 1484.060 ;
        RECT 1178.620 1483.800 1178.880 1484.060 ;
        RECT 1178.620 1483.120 1178.880 1483.380 ;
        RECT 1178.620 1435.520 1178.880 1435.780 ;
        RECT 1178.620 1048.600 1178.880 1048.860 ;
        RECT 1177.700 1000.660 1177.960 1000.920 ;
        RECT 1178.620 903.760 1178.880 904.020 ;
        RECT 1178.160 855.480 1178.420 855.740 ;
        RECT 1178.620 482.840 1178.880 483.100 ;
        RECT 1178.620 434.900 1178.880 435.160 ;
        RECT 1178.620 385.940 1178.880 386.200 ;
        RECT 1178.620 338.000 1178.880 338.260 ;
        RECT 1178.620 289.380 1178.880 289.640 ;
        RECT 1178.620 241.440 1178.880 241.700 ;
        RECT 1178.620 192.820 1178.880 193.080 ;
        RECT 1178.620 144.880 1178.880 145.140 ;
        RECT 1178.620 96.260 1178.880 96.520 ;
        RECT 2387.500 79.260 2387.760 79.520 ;
        RECT 2387.500 17.720 2387.760 17.980 ;
        RECT 2393.480 17.720 2393.740 17.980 ;
      LAYER met2 ;
        RECT 1179.400 1600.450 1179.680 1604.000 ;
        RECT 1178.220 1600.310 1179.680 1600.450 ;
        RECT 1178.220 1580.310 1178.360 1600.310 ;
        RECT 1179.400 1600.000 1179.680 1600.310 ;
        RECT 1174.480 1579.990 1174.740 1580.310 ;
        RECT 1178.160 1579.990 1178.420 1580.310 ;
        RECT 1174.540 1484.090 1174.680 1579.990 ;
        RECT 1174.480 1483.770 1174.740 1484.090 ;
        RECT 1178.620 1483.770 1178.880 1484.090 ;
        RECT 1178.680 1483.410 1178.820 1483.770 ;
        RECT 1178.620 1483.090 1178.880 1483.410 ;
        RECT 1178.620 1435.490 1178.880 1435.810 ;
        RECT 1178.680 1048.890 1178.820 1435.490 ;
        RECT 1178.620 1048.570 1178.880 1048.890 ;
        RECT 1177.700 1000.630 1177.960 1000.950 ;
        RECT 1177.760 904.245 1177.900 1000.630 ;
        RECT 1177.690 903.875 1177.970 904.245 ;
        RECT 1178.610 903.875 1178.890 904.245 ;
        RECT 1178.620 903.730 1178.880 903.875 ;
        RECT 1178.160 855.450 1178.420 855.770 ;
        RECT 1178.220 846.330 1178.360 855.450 ;
        RECT 1177.760 846.190 1178.360 846.330 ;
        RECT 1177.760 773.005 1177.900 846.190 ;
        RECT 1177.690 772.635 1177.970 773.005 ;
        RECT 1178.610 772.635 1178.890 773.005 ;
        RECT 1178.680 483.130 1178.820 772.635 ;
        RECT 1178.620 482.810 1178.880 483.130 ;
        RECT 1178.620 434.870 1178.880 435.190 ;
        RECT 1178.680 386.230 1178.820 434.870 ;
        RECT 1178.620 385.910 1178.880 386.230 ;
        RECT 1178.620 337.970 1178.880 338.290 ;
        RECT 1178.680 289.670 1178.820 337.970 ;
        RECT 1178.620 289.350 1178.880 289.670 ;
        RECT 1178.620 241.410 1178.880 241.730 ;
        RECT 1178.680 193.110 1178.820 241.410 ;
        RECT 1178.620 192.790 1178.880 193.110 ;
        RECT 1178.620 144.850 1178.880 145.170 ;
        RECT 1178.680 96.550 1178.820 144.850 ;
        RECT 1178.620 96.230 1178.880 96.550 ;
        RECT 2387.500 79.230 2387.760 79.550 ;
        RECT 2387.560 18.010 2387.700 79.230 ;
        RECT 2387.500 17.690 2387.760 18.010 ;
        RECT 2393.480 17.690 2393.740 18.010 ;
        RECT 2393.540 2.400 2393.680 17.690 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
      LAYER via2 ;
        RECT 1177.690 903.920 1177.970 904.200 ;
        RECT 1178.610 903.920 1178.890 904.200 ;
        RECT 1177.690 772.680 1177.970 772.960 ;
        RECT 1178.610 772.680 1178.890 772.960 ;
      LAYER met3 ;
        RECT 1177.665 904.210 1177.995 904.225 ;
        RECT 1178.585 904.210 1178.915 904.225 ;
        RECT 1177.665 903.910 1178.915 904.210 ;
        RECT 1177.665 903.895 1177.995 903.910 ;
        RECT 1178.585 903.895 1178.915 903.910 ;
        RECT 1177.665 772.970 1177.995 772.985 ;
        RECT 1178.585 772.970 1178.915 772.985 ;
        RECT 1177.665 772.670 1178.915 772.970 ;
        RECT 1177.665 772.655 1177.995 772.670 ;
        RECT 1178.585 772.655 1178.915 772.670 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1893.045 19.465 1894.135 19.635 ;
        RECT 1893.045 15.725 1893.215 19.465 ;
        RECT 1893.965 19.295 1894.135 19.465 ;
        RECT 1893.965 19.125 1894.595 19.295 ;
      LAYER mcon ;
        RECT 1894.425 19.125 1894.595 19.295 ;
      LAYER met1 ;
        RECT 1894.365 19.280 1894.655 19.325 ;
        RECT 2411.390 19.280 2411.710 19.340 ;
        RECT 1894.365 19.140 2411.710 19.280 ;
        RECT 1894.365 19.095 1894.655 19.140 ;
        RECT 2411.390 19.080 2411.710 19.140 ;
        RECT 1876.410 15.880 1876.730 15.940 ;
        RECT 1892.985 15.880 1893.275 15.925 ;
        RECT 1876.410 15.740 1893.275 15.880 ;
        RECT 1876.410 15.680 1876.730 15.740 ;
        RECT 1892.985 15.695 1893.275 15.740 ;
      LAYER via ;
        RECT 2411.420 19.080 2411.680 19.340 ;
        RECT 1876.440 15.680 1876.700 15.940 ;
      LAYER met2 ;
        RECT 1185.840 1600.380 1186.120 1604.000 ;
        RECT 1185.840 1600.000 1186.180 1600.380 ;
        RECT 1186.040 1593.085 1186.180 1600.000 ;
        RECT 1185.970 1592.715 1186.250 1593.085 ;
        RECT 1873.210 1592.715 1873.490 1593.085 ;
        RECT 1873.280 26.930 1873.420 1592.715 ;
        RECT 1873.280 26.790 1876.640 26.930 ;
        RECT 1876.500 15.970 1876.640 26.790 ;
        RECT 2411.420 19.050 2411.680 19.370 ;
        RECT 1876.440 15.650 1876.700 15.970 ;
        RECT 2411.480 2.400 2411.620 19.050 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
      LAYER via2 ;
        RECT 1185.970 1592.760 1186.250 1593.040 ;
        RECT 1873.210 1592.760 1873.490 1593.040 ;
      LAYER met3 ;
        RECT 1185.945 1593.050 1186.275 1593.065 ;
        RECT 1873.185 1593.050 1873.515 1593.065 ;
        RECT 1185.945 1592.750 1873.515 1593.050 ;
        RECT 1185.945 1592.735 1186.275 1592.750 ;
        RECT 1873.185 1592.735 1873.515 1592.750 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 686.925 14.025 687.095 15.215 ;
        RECT 793.185 14.705 793.355 15.895 ;
      LAYER mcon ;
        RECT 793.185 15.725 793.355 15.895 ;
        RECT 686.925 15.045 687.095 15.215 ;
      LAYER met1 ;
        RECT 655.660 1589.600 663.620 1589.740 ;
        RECT 629.350 1589.400 629.670 1589.460 ;
        RECT 655.660 1589.400 655.800 1589.600 ;
        RECT 629.350 1589.260 655.800 1589.400 ;
        RECT 629.350 1589.200 629.670 1589.260 ;
        RECT 663.480 1588.380 663.620 1589.600 ;
        RECT 679.490 1588.380 679.810 1588.440 ;
        RECT 663.480 1588.240 679.810 1588.380 ;
        RECT 679.490 1588.180 679.810 1588.240 ;
        RECT 793.125 15.880 793.415 15.925 ;
        RECT 805.530 15.880 805.850 15.940 ;
        RECT 793.125 15.740 805.850 15.880 ;
        RECT 793.125 15.695 793.415 15.740 ;
        RECT 805.530 15.680 805.850 15.740 ;
        RECT 679.490 15.200 679.810 15.260 ;
        RECT 686.865 15.200 687.155 15.245 ;
        RECT 679.490 15.060 687.155 15.200 ;
        RECT 679.490 15.000 679.810 15.060 ;
        RECT 686.865 15.015 687.155 15.060 ;
        RECT 786.210 14.860 786.530 14.920 ;
        RECT 793.125 14.860 793.415 14.905 ;
        RECT 786.210 14.720 793.415 14.860 ;
        RECT 786.210 14.660 786.530 14.720 ;
        RECT 793.125 14.675 793.415 14.720 ;
        RECT 758.610 14.520 758.930 14.580 ;
        RECT 748.120 14.380 758.930 14.520 ;
        RECT 686.865 14.180 687.155 14.225 ;
        RECT 748.120 14.180 748.260 14.380 ;
        RECT 758.610 14.320 758.930 14.380 ;
        RECT 686.865 14.040 748.260 14.180 ;
        RECT 686.865 13.995 687.155 14.040 ;
      LAYER via ;
        RECT 629.380 1589.200 629.640 1589.460 ;
        RECT 679.520 1588.180 679.780 1588.440 ;
        RECT 805.560 15.680 805.820 15.940 ;
        RECT 679.520 15.000 679.780 15.260 ;
        RECT 786.240 14.660 786.500 14.920 ;
        RECT 758.640 14.320 758.900 14.580 ;
      LAYER met2 ;
        RECT 629.240 1600.380 629.520 1604.000 ;
        RECT 629.240 1600.000 629.580 1600.380 ;
        RECT 629.440 1589.490 629.580 1600.000 ;
        RECT 629.380 1589.170 629.640 1589.490 ;
        RECT 679.520 1588.150 679.780 1588.470 ;
        RECT 679.580 15.290 679.720 1588.150 ;
        RECT 805.560 15.650 805.820 15.970 ;
        RECT 679.520 14.970 679.780 15.290 ;
        RECT 786.240 14.805 786.500 14.950 ;
        RECT 758.630 14.435 758.910 14.805 ;
        RECT 786.230 14.435 786.510 14.805 ;
        RECT 758.640 14.290 758.900 14.435 ;
        RECT 805.620 2.400 805.760 15.650 ;
        RECT 805.410 -4.800 805.970 2.400 ;
      LAYER via2 ;
        RECT 758.630 14.480 758.910 14.760 ;
        RECT 786.230 14.480 786.510 14.760 ;
      LAYER met3 ;
        RECT 758.605 14.770 758.935 14.785 ;
        RECT 786.205 14.770 786.535 14.785 ;
        RECT 758.605 14.470 786.535 14.770 ;
        RECT 758.605 14.455 758.935 14.470 ;
        RECT 786.205 14.455 786.535 14.470 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.050 2837.880 972.370 2837.940 ;
        RECT 1260.930 2837.880 1261.250 2837.940 ;
        RECT 972.050 2837.740 1261.250 2837.880 ;
        RECT 972.050 2837.680 972.370 2837.740 ;
        RECT 1260.930 2837.680 1261.250 2837.740 ;
        RECT 1262.770 2787.900 1263.090 2787.960 ;
        RECT 1262.770 2787.760 1269.900 2787.900 ;
        RECT 1262.770 2787.700 1263.090 2787.760 ;
        RECT 1269.760 2787.560 1269.900 2787.760 ;
        RECT 1289.910 2787.560 1290.230 2787.620 ;
        RECT 1269.760 2787.420 1290.230 2787.560 ;
        RECT 1289.910 2787.360 1290.230 2787.420 ;
        RECT 1290.370 2758.320 1290.690 2758.380 ;
        RECT 1298.650 2758.320 1298.970 2758.380 ;
        RECT 1290.370 2758.180 1298.970 2758.320 ;
        RECT 1290.370 2758.120 1290.690 2758.180 ;
        RECT 1298.650 2758.120 1298.970 2758.180 ;
        RECT 1298.650 2746.080 1298.970 2746.140 ;
        RECT 1307.390 2746.080 1307.710 2746.140 ;
        RECT 1298.650 2745.940 1307.710 2746.080 ;
        RECT 1298.650 2745.880 1298.970 2745.940 ;
        RECT 1307.390 2745.880 1307.710 2745.940 ;
        RECT 1307.390 2704.940 1307.710 2705.000 ;
        RECT 1307.390 2704.800 1311.300 2704.940 ;
        RECT 1307.390 2704.740 1307.710 2704.800 ;
        RECT 1311.160 2704.600 1311.300 2704.800 ;
        RECT 1317.970 2704.600 1318.290 2704.660 ;
        RECT 1311.160 2704.460 1318.290 2704.600 ;
        RECT 1317.970 2704.400 1318.290 2704.460 ;
        RECT 1317.970 2694.400 1318.290 2694.460 ;
        RECT 1360.290 2694.400 1360.610 2694.460 ;
        RECT 1317.970 2694.260 1360.610 2694.400 ;
        RECT 1317.970 2694.200 1318.290 2694.260 ;
        RECT 1360.290 2694.200 1360.610 2694.260 ;
        RECT 1360.290 2672.980 1360.610 2673.040 ;
        RECT 1369.490 2672.980 1369.810 2673.040 ;
        RECT 1360.290 2672.840 1369.810 2672.980 ;
        RECT 1360.290 2672.780 1360.610 2672.840 ;
        RECT 1369.490 2672.780 1369.810 2672.840 ;
        RECT 599.910 2628.440 600.230 2628.500 ;
        RECT 973.890 2628.440 974.210 2628.500 ;
        RECT 599.910 2628.300 974.210 2628.440 ;
        RECT 599.910 2628.240 600.230 2628.300 ;
        RECT 973.890 2628.240 974.210 2628.300 ;
        RECT 1369.490 2618.920 1369.810 2618.980 ;
        RECT 1376.850 2618.920 1377.170 2618.980 ;
        RECT 1369.490 2618.780 1377.170 2618.920 ;
        RECT 1369.490 2618.720 1369.810 2618.780 ;
        RECT 1376.850 2618.720 1377.170 2618.780 ;
        RECT 1376.850 2595.120 1377.170 2595.180 ;
        RECT 1393.870 2595.120 1394.190 2595.180 ;
        RECT 1376.850 2594.980 1394.190 2595.120 ;
        RECT 1376.850 2594.920 1377.170 2594.980 ;
        RECT 1393.870 2594.920 1394.190 2594.980 ;
        RECT 1393.870 2585.260 1394.190 2585.320 ;
        RECT 1400.310 2585.260 1400.630 2585.320 ;
        RECT 1393.870 2585.120 1400.630 2585.260 ;
        RECT 1393.870 2585.060 1394.190 2585.120 ;
        RECT 1400.310 2585.060 1400.630 2585.120 ;
        RECT 1400.310 2584.240 1400.630 2584.300 ;
        RECT 1600.870 2584.240 1601.190 2584.300 ;
        RECT 1400.310 2584.100 1601.190 2584.240 ;
        RECT 1400.310 2584.040 1400.630 2584.100 ;
        RECT 1600.870 2584.040 1601.190 2584.100 ;
        RECT 2.830 24.380 3.150 24.440 ;
        RECT 345.070 24.380 345.390 24.440 ;
        RECT 2.830 24.240 345.390 24.380 ;
        RECT 2.830 24.180 3.150 24.240 ;
        RECT 345.070 24.180 345.390 24.240 ;
      LAYER via ;
        RECT 972.080 2837.680 972.340 2837.940 ;
        RECT 1260.960 2837.680 1261.220 2837.940 ;
        RECT 1262.800 2787.700 1263.060 2787.960 ;
        RECT 1289.940 2787.360 1290.200 2787.620 ;
        RECT 1290.400 2758.120 1290.660 2758.380 ;
        RECT 1298.680 2758.120 1298.940 2758.380 ;
        RECT 1298.680 2745.880 1298.940 2746.140 ;
        RECT 1307.420 2745.880 1307.680 2746.140 ;
        RECT 1307.420 2704.740 1307.680 2705.000 ;
        RECT 1318.000 2704.400 1318.260 2704.660 ;
        RECT 1318.000 2694.200 1318.260 2694.460 ;
        RECT 1360.320 2694.200 1360.580 2694.460 ;
        RECT 1360.320 2672.780 1360.580 2673.040 ;
        RECT 1369.520 2672.780 1369.780 2673.040 ;
        RECT 599.940 2628.240 600.200 2628.500 ;
        RECT 973.920 2628.240 974.180 2628.500 ;
        RECT 1369.520 2618.720 1369.780 2618.980 ;
        RECT 1376.880 2618.720 1377.140 2618.980 ;
        RECT 1376.880 2594.920 1377.140 2595.180 ;
        RECT 1393.900 2594.920 1394.160 2595.180 ;
        RECT 1393.900 2585.060 1394.160 2585.320 ;
        RECT 1400.340 2585.060 1400.600 2585.320 ;
        RECT 1400.340 2584.040 1400.600 2584.300 ;
        RECT 1600.900 2584.040 1601.160 2584.300 ;
        RECT 2.860 24.180 3.120 24.440 ;
        RECT 345.100 24.180 345.360 24.440 ;
      LAYER met2 ;
        RECT 599.930 2850.715 600.210 2851.085 ;
        RECT 600.000 2628.530 600.140 2850.715 ;
        RECT 972.070 2841.875 972.350 2842.245 ;
        RECT 972.140 2838.165 972.280 2841.875 ;
        RECT 972.070 2837.795 972.350 2838.165 ;
        RECT 972.080 2837.650 972.340 2837.795 ;
        RECT 1260.960 2837.650 1261.220 2837.970 ;
        RECT 972.140 2837.495 972.280 2837.650 ;
        RECT 1261.020 2808.130 1261.160 2837.650 ;
        RECT 1261.020 2807.990 1263.000 2808.130 ;
        RECT 1262.860 2787.990 1263.000 2807.990 ;
        RECT 1262.800 2787.670 1263.060 2787.990 ;
        RECT 1289.940 2787.330 1290.200 2787.650 ;
        RECT 1290.000 2777.530 1290.140 2787.330 ;
        RECT 1290.000 2777.390 1290.600 2777.530 ;
        RECT 1290.460 2758.410 1290.600 2777.390 ;
        RECT 1290.400 2758.090 1290.660 2758.410 ;
        RECT 1298.680 2758.090 1298.940 2758.410 ;
        RECT 1298.740 2746.170 1298.880 2758.090 ;
        RECT 1298.680 2745.850 1298.940 2746.170 ;
        RECT 1307.420 2745.850 1307.680 2746.170 ;
        RECT 1307.480 2705.030 1307.620 2745.850 ;
        RECT 1307.420 2704.710 1307.680 2705.030 ;
        RECT 1318.000 2704.370 1318.260 2704.690 ;
        RECT 1318.060 2694.490 1318.200 2704.370 ;
        RECT 1318.000 2694.170 1318.260 2694.490 ;
        RECT 1360.320 2694.170 1360.580 2694.490 ;
        RECT 1360.380 2673.070 1360.520 2694.170 ;
        RECT 1360.320 2672.750 1360.580 2673.070 ;
        RECT 1369.520 2672.750 1369.780 2673.070 ;
        RECT 599.940 2628.210 600.200 2628.530 ;
        RECT 973.920 2628.210 974.180 2628.530 ;
        RECT 973.980 2610.000 974.120 2628.210 ;
        RECT 1369.580 2619.010 1369.720 2672.750 ;
        RECT 1369.520 2618.690 1369.780 2619.010 ;
        RECT 1376.880 2618.690 1377.140 2619.010 ;
        RECT 973.780 2609.500 974.120 2610.000 ;
        RECT 973.780 2606.000 974.060 2609.500 ;
        RECT 1376.940 2595.210 1377.080 2618.690 ;
        RECT 1376.880 2594.890 1377.140 2595.210 ;
        RECT 1393.900 2594.890 1394.160 2595.210 ;
        RECT 1393.960 2585.350 1394.100 2594.890 ;
        RECT 1393.900 2585.030 1394.160 2585.350 ;
        RECT 1400.340 2585.030 1400.600 2585.350 ;
        RECT 1400.400 2584.330 1400.540 2585.030 ;
        RECT 1400.340 2584.010 1400.600 2584.330 ;
        RECT 1600.900 2584.010 1601.160 2584.330 ;
        RECT 1400.400 1980.685 1400.540 2584.010 ;
        RECT 1600.960 2583.845 1601.100 2584.010 ;
        RECT 1600.890 2583.475 1601.170 2583.845 ;
        RECT 1400.330 1980.315 1400.610 1980.685 ;
        RECT 350.940 1603.170 351.220 1604.000 ;
        RECT 351.530 1603.170 351.810 1603.285 ;
        RECT 350.940 1603.030 351.810 1603.170 ;
        RECT 350.940 1600.000 351.280 1603.030 ;
        RECT 351.530 1602.915 351.810 1603.030 ;
        RECT 351.140 1593.765 351.280 1600.000 ;
        RECT 345.090 1593.395 345.370 1593.765 ;
        RECT 351.070 1593.395 351.350 1593.765 ;
        RECT 345.160 24.470 345.300 1593.395 ;
        RECT 2.860 24.150 3.120 24.470 ;
        RECT 345.100 24.150 345.360 24.470 ;
        RECT 2.920 2.400 3.060 24.150 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 599.930 2850.760 600.210 2851.040 ;
        RECT 972.070 2841.920 972.350 2842.200 ;
        RECT 972.070 2837.840 972.350 2838.120 ;
        RECT 1600.890 2583.520 1601.170 2583.800 ;
        RECT 1400.330 1980.360 1400.610 1980.640 ;
        RECT 351.530 1602.960 351.810 1603.240 ;
        RECT 345.090 1593.440 345.370 1593.720 ;
        RECT 351.070 1593.440 351.350 1593.720 ;
      LAYER met3 ;
        RECT 599.190 2851.050 599.570 2851.060 ;
        RECT 599.905 2851.050 600.235 2851.065 ;
        RECT 599.190 2850.750 600.235 2851.050 ;
        RECT 599.190 2850.740 599.570 2850.750 ;
        RECT 599.905 2850.735 600.235 2850.750 ;
        RECT 972.045 2842.220 972.375 2842.225 ;
        RECT 971.790 2842.210 972.375 2842.220 ;
        RECT 971.590 2841.910 972.375 2842.210 ;
        RECT 971.790 2841.900 972.375 2841.910 ;
        RECT 972.045 2841.895 972.375 2841.900 ;
        RECT 417.030 2838.130 417.410 2838.140 ;
        RECT 972.045 2838.130 972.375 2838.145 ;
        RECT 417.030 2837.830 972.375 2838.130 ;
        RECT 417.030 2837.820 417.410 2837.830 ;
        RECT 972.045 2837.815 972.375 2837.830 ;
        RECT 1600.865 2583.820 1601.195 2583.825 ;
        RECT 1600.865 2583.810 1601.450 2583.820 ;
        RECT 1600.640 2583.510 1601.450 2583.810 ;
        RECT 1600.865 2583.500 1601.450 2583.510 ;
        RECT 1600.865 2583.495 1601.195 2583.500 ;
        RECT 1399.590 1980.650 1399.970 1980.660 ;
        RECT 1400.305 1980.650 1400.635 1980.665 ;
        RECT 1399.590 1980.350 1400.635 1980.650 ;
        RECT 1399.590 1980.340 1399.970 1980.350 ;
        RECT 1400.305 1980.335 1400.635 1980.350 ;
        RECT 350.790 1603.250 351.170 1603.260 ;
        RECT 351.505 1603.250 351.835 1603.265 ;
        RECT 350.790 1602.950 351.835 1603.250 ;
        RECT 350.790 1602.940 351.170 1602.950 ;
        RECT 351.505 1602.935 351.835 1602.950 ;
        RECT 345.065 1593.730 345.395 1593.745 ;
        RECT 351.045 1593.730 351.375 1593.745 ;
        RECT 345.065 1593.430 351.375 1593.730 ;
        RECT 345.065 1593.415 345.395 1593.430 ;
        RECT 351.045 1593.415 351.375 1593.430 ;
      LAYER via3 ;
        RECT 599.220 2850.740 599.540 2851.060 ;
        RECT 971.820 2841.900 972.140 2842.220 ;
        RECT 417.060 2837.820 417.380 2838.140 ;
        RECT 1601.100 2583.500 1601.420 2583.820 ;
        RECT 1399.620 1980.340 1399.940 1980.660 ;
        RECT 350.820 1602.940 351.140 1603.260 ;
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 418.020 3306.235 421.020 3557.200 ;
        RECT 598.020 3306.235 601.020 3557.200 ;
        RECT 778.020 3306.235 781.020 3557.200 ;
        RECT 958.020 3306.235 961.020 3557.200 ;
        RECT 1138.020 3306.235 1141.020 3557.200 ;
        RECT 1318.020 3306.235 1321.020 3557.200 ;
        RECT 600.105 3301.635 600.405 3306.235 ;
        RECT 1317.865 3301.635 1318.165 3306.235 ;
        RECT 419.015 2851.050 419.315 2854.600 ;
        RECT 417.070 2850.750 419.315 2851.050 ;
        RECT 417.070 2838.145 417.370 2850.750 ;
        RECT 419.015 2850.000 419.315 2850.750 ;
        RECT 598.150 2851.050 598.450 2854.600 ;
        RECT 599.215 2851.050 599.545 2851.065 ;
        RECT 598.150 2850.750 599.545 2851.050 ;
        RECT 598.150 2850.000 598.450 2850.750 ;
        RECT 599.215 2850.735 599.545 2850.750 ;
        RECT 969.015 2851.050 969.315 2854.600 ;
        RECT 969.015 2850.750 972.130 2851.050 ;
        RECT 969.015 2850.000 969.315 2850.750 ;
        RECT 417.055 2837.815 417.385 2838.145 ;
        RECT 350.390 1979.910 351.570 1981.090 ;
        RECT 350.830 1603.265 351.130 1979.910 ;
        RECT 350.815 1602.935 351.145 1603.265 ;
        RECT 418.020 -37.520 421.020 2850.000 ;
        RECT 598.020 -37.520 601.020 2850.000 ;
        RECT 778.020 -37.520 781.020 2850.000 ;
        RECT 958.020 -37.520 961.020 2850.000 ;
        RECT 971.830 2842.225 972.130 2850.750 ;
        RECT 971.815 2841.895 972.145 2842.225 ;
        RECT 1138.020 -37.520 1141.020 2850.000 ;
        RECT 1318.020 -37.520 1321.020 2850.000 ;
        RECT 1399.190 1979.910 1400.370 1981.090 ;
        RECT 1498.020 -37.520 1501.020 3557.200 ;
        RECT 1678.020 2586.480 1681.020 3557.200 ;
        RECT 1858.020 2586.480 1861.020 3557.200 ;
        RECT 2038.020 2586.480 2041.020 3557.200 ;
        RECT 1601.095 2583.495 1601.425 2583.825 ;
        RECT 1601.110 2567.465 1601.410 2583.495 ;
        RECT 1600.000 2567.165 1604.600 2567.465 ;
        RECT 1678.020 1986.480 1681.020 2200.000 ;
        RECT 1858.020 1986.480 1861.020 2200.000 ;
        RECT 2038.020 1986.480 2041.020 2200.000 ;
        RECT 1600.670 1979.910 1601.850 1981.090 ;
        RECT 1601.110 1967.465 1601.410 1979.910 ;
        RECT 1600.000 1967.165 1604.600 1967.465 ;
        RECT 1678.020 -37.520 1681.020 1600.000 ;
        RECT 1858.020 -37.520 1861.020 1600.000 ;
        RECT 2038.020 -37.520 2041.020 1600.000 ;
        RECT 2218.020 -37.520 2221.020 3557.200 ;
        RECT 2398.020 -37.520 2401.020 3557.200 ;
        RECT 2578.020 -37.520 2581.020 3557.200 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT 350.180 1979.700 1602.060 1981.300 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 352.505 1449.165 352.675 1497.275 ;
      LAYER mcon ;
        RECT 352.505 1497.105 352.675 1497.275 ;
      LAYER met1 ;
        RECT 352.890 1511.540 353.210 1511.600 ;
        RECT 352.520 1511.400 353.210 1511.540 ;
        RECT 352.520 1510.920 352.660 1511.400 ;
        RECT 352.890 1511.340 353.210 1511.400 ;
        RECT 352.430 1510.660 352.750 1510.920 ;
        RECT 352.430 1497.260 352.750 1497.320 ;
        RECT 352.235 1497.120 352.750 1497.260 ;
        RECT 352.430 1497.060 352.750 1497.120 ;
        RECT 352.445 1449.320 352.735 1449.365 ;
        RECT 352.890 1449.320 353.210 1449.380 ;
        RECT 352.445 1449.180 353.210 1449.320 ;
        RECT 352.445 1449.135 352.735 1449.180 ;
        RECT 352.890 1449.120 353.210 1449.180 ;
        RECT 352.430 1320.460 352.750 1320.520 ;
        RECT 353.350 1320.460 353.670 1320.520 ;
        RECT 352.430 1320.320 353.670 1320.460 ;
        RECT 352.430 1320.260 352.750 1320.320 ;
        RECT 353.350 1320.260 353.670 1320.320 ;
        RECT 352.430 1269.460 352.750 1269.520 ;
        RECT 353.350 1269.460 353.670 1269.520 ;
        RECT 352.430 1269.320 353.670 1269.460 ;
        RECT 352.430 1269.260 352.750 1269.320 ;
        RECT 353.350 1269.260 353.670 1269.320 ;
        RECT 353.350 1221.860 353.670 1221.920 ;
        RECT 352.520 1221.720 353.670 1221.860 ;
        RECT 352.520 1221.580 352.660 1221.720 ;
        RECT 353.350 1221.660 353.670 1221.720 ;
        RECT 352.430 1221.320 352.750 1221.580 ;
        RECT 352.430 1172.900 352.750 1172.960 ;
        RECT 353.350 1172.900 353.670 1172.960 ;
        RECT 352.430 1172.760 353.670 1172.900 ;
        RECT 352.430 1172.700 352.750 1172.760 ;
        RECT 353.350 1172.700 353.670 1172.760 ;
        RECT 353.350 1125.300 353.670 1125.360 ;
        RECT 352.520 1125.160 353.670 1125.300 ;
        RECT 352.520 1125.020 352.660 1125.160 ;
        RECT 353.350 1125.100 353.670 1125.160 ;
        RECT 352.430 1124.760 352.750 1125.020 ;
        RECT 352.430 1076.340 352.750 1076.400 ;
        RECT 353.350 1076.340 353.670 1076.400 ;
        RECT 352.430 1076.200 353.670 1076.340 ;
        RECT 352.430 1076.140 352.750 1076.200 ;
        RECT 353.350 1076.140 353.670 1076.200 ;
        RECT 353.350 1028.740 353.670 1028.800 ;
        RECT 352.520 1028.600 353.670 1028.740 ;
        RECT 352.520 1028.460 352.660 1028.600 ;
        RECT 353.350 1028.540 353.670 1028.600 ;
        RECT 352.430 1028.200 352.750 1028.460 ;
        RECT 352.430 979.780 352.750 979.840 ;
        RECT 353.350 979.780 353.670 979.840 ;
        RECT 352.430 979.640 353.670 979.780 ;
        RECT 352.430 979.580 352.750 979.640 ;
        RECT 353.350 979.580 353.670 979.640 ;
        RECT 353.350 932.180 353.670 932.240 ;
        RECT 352.520 932.040 353.670 932.180 ;
        RECT 352.520 931.900 352.660 932.040 ;
        RECT 353.350 931.980 353.670 932.040 ;
        RECT 352.430 931.640 352.750 931.900 ;
        RECT 352.430 883.220 352.750 883.280 ;
        RECT 353.350 883.220 353.670 883.280 ;
        RECT 352.430 883.080 353.670 883.220 ;
        RECT 352.430 883.020 352.750 883.080 ;
        RECT 353.350 883.020 353.670 883.080 ;
        RECT 353.350 835.620 353.670 835.680 ;
        RECT 352.520 835.480 353.670 835.620 ;
        RECT 352.520 835.340 352.660 835.480 ;
        RECT 353.350 835.420 353.670 835.480 ;
        RECT 352.430 835.080 352.750 835.340 ;
        RECT 352.430 786.660 352.750 786.720 ;
        RECT 353.810 786.660 354.130 786.720 ;
        RECT 352.430 786.520 354.130 786.660 ;
        RECT 352.430 786.460 352.750 786.520 ;
        RECT 353.810 786.460 354.130 786.520 ;
        RECT 352.430 738.380 352.750 738.440 ;
        RECT 353.810 738.380 354.130 738.440 ;
        RECT 352.430 738.240 354.130 738.380 ;
        RECT 352.430 738.180 352.750 738.240 ;
        RECT 353.810 738.180 354.130 738.240 ;
        RECT 353.350 642.160 353.670 642.220 ;
        RECT 352.520 642.020 353.670 642.160 ;
        RECT 352.520 641.880 352.660 642.020 ;
        RECT 353.350 641.960 353.670 642.020 ;
        RECT 352.430 641.620 352.750 641.880 ;
        RECT 352.430 627.880 352.750 627.940 ;
        RECT 353.350 627.880 353.670 627.940 ;
        RECT 352.430 627.740 353.670 627.880 ;
        RECT 352.430 627.680 352.750 627.740 ;
        RECT 353.350 627.680 353.670 627.740 ;
        RECT 353.350 545.600 353.670 545.660 ;
        RECT 352.520 545.460 353.670 545.600 ;
        RECT 352.520 545.320 352.660 545.460 ;
        RECT 353.350 545.400 353.670 545.460 ;
        RECT 352.430 545.060 352.750 545.320 ;
        RECT 352.430 476.240 352.750 476.300 ;
        RECT 353.350 476.240 353.670 476.300 ;
        RECT 352.430 476.100 353.670 476.240 ;
        RECT 352.430 476.040 352.750 476.100 ;
        RECT 353.350 476.040 353.670 476.100 ;
        RECT 353.350 449.040 353.670 449.100 ;
        RECT 352.520 448.900 353.670 449.040 ;
        RECT 352.520 448.760 352.660 448.900 ;
        RECT 353.350 448.840 353.670 448.900 ;
        RECT 352.430 448.500 352.750 448.760 ;
        RECT 352.430 357.240 352.750 357.300 ;
        RECT 353.350 357.240 353.670 357.300 ;
        RECT 352.430 357.100 353.670 357.240 ;
        RECT 352.430 357.040 352.750 357.100 ;
        RECT 353.350 357.040 353.670 357.100 ;
        RECT 352.430 335.820 352.750 335.880 ;
        RECT 353.350 335.820 353.670 335.880 ;
        RECT 352.430 335.680 353.670 335.820 ;
        RECT 352.430 335.620 352.750 335.680 ;
        RECT 353.350 335.620 353.670 335.680 ;
        RECT 352.430 265.780 352.750 265.840 ;
        RECT 353.350 265.780 353.670 265.840 ;
        RECT 352.430 265.640 353.670 265.780 ;
        RECT 352.430 265.580 352.750 265.640 ;
        RECT 353.350 265.580 353.670 265.640 ;
        RECT 352.430 206.960 352.750 207.020 ;
        RECT 353.350 206.960 353.670 207.020 ;
        RECT 352.430 206.820 353.670 206.960 ;
        RECT 352.430 206.760 352.750 206.820 ;
        RECT 353.350 206.760 353.670 206.820 ;
        RECT 352.430 169.220 352.750 169.280 ;
        RECT 353.350 169.220 353.670 169.280 ;
        RECT 352.430 169.080 353.670 169.220 ;
        RECT 352.430 169.020 352.750 169.080 ;
        RECT 353.350 169.020 353.670 169.080 ;
        RECT 352.430 113.460 352.750 113.520 ;
        RECT 353.350 113.460 353.670 113.520 ;
        RECT 352.430 113.320 353.670 113.460 ;
        RECT 352.430 113.260 352.750 113.320 ;
        RECT 353.350 113.260 353.670 113.320 ;
        RECT 353.350 62.800 353.670 62.860 ;
        RECT 352.520 62.660 353.670 62.800 ;
        RECT 352.520 62.520 352.660 62.660 ;
        RECT 353.350 62.600 353.670 62.660 ;
        RECT 352.430 62.260 352.750 62.520 ;
        RECT 8.350 24.040 8.670 24.100 ;
        RECT 352.430 24.040 352.750 24.100 ;
        RECT 8.350 23.900 352.750 24.040 ;
        RECT 8.350 23.840 8.670 23.900 ;
        RECT 352.430 23.840 352.750 23.900 ;
      LAYER via ;
        RECT 352.920 1511.340 353.180 1511.600 ;
        RECT 352.460 1510.660 352.720 1510.920 ;
        RECT 352.460 1497.060 352.720 1497.320 ;
        RECT 352.920 1449.120 353.180 1449.380 ;
        RECT 352.460 1320.260 352.720 1320.520 ;
        RECT 353.380 1320.260 353.640 1320.520 ;
        RECT 352.460 1269.260 352.720 1269.520 ;
        RECT 353.380 1269.260 353.640 1269.520 ;
        RECT 353.380 1221.660 353.640 1221.920 ;
        RECT 352.460 1221.320 352.720 1221.580 ;
        RECT 352.460 1172.700 352.720 1172.960 ;
        RECT 353.380 1172.700 353.640 1172.960 ;
        RECT 353.380 1125.100 353.640 1125.360 ;
        RECT 352.460 1124.760 352.720 1125.020 ;
        RECT 352.460 1076.140 352.720 1076.400 ;
        RECT 353.380 1076.140 353.640 1076.400 ;
        RECT 353.380 1028.540 353.640 1028.800 ;
        RECT 352.460 1028.200 352.720 1028.460 ;
        RECT 352.460 979.580 352.720 979.840 ;
        RECT 353.380 979.580 353.640 979.840 ;
        RECT 353.380 931.980 353.640 932.240 ;
        RECT 352.460 931.640 352.720 931.900 ;
        RECT 352.460 883.020 352.720 883.280 ;
        RECT 353.380 883.020 353.640 883.280 ;
        RECT 353.380 835.420 353.640 835.680 ;
        RECT 352.460 835.080 352.720 835.340 ;
        RECT 352.460 786.460 352.720 786.720 ;
        RECT 353.840 786.460 354.100 786.720 ;
        RECT 352.460 738.180 352.720 738.440 ;
        RECT 353.840 738.180 354.100 738.440 ;
        RECT 353.380 641.960 353.640 642.220 ;
        RECT 352.460 641.620 352.720 641.880 ;
        RECT 352.460 627.680 352.720 627.940 ;
        RECT 353.380 627.680 353.640 627.940 ;
        RECT 353.380 545.400 353.640 545.660 ;
        RECT 352.460 545.060 352.720 545.320 ;
        RECT 352.460 476.040 352.720 476.300 ;
        RECT 353.380 476.040 353.640 476.300 ;
        RECT 353.380 448.840 353.640 449.100 ;
        RECT 352.460 448.500 352.720 448.760 ;
        RECT 352.460 357.040 352.720 357.300 ;
        RECT 353.380 357.040 353.640 357.300 ;
        RECT 352.460 335.620 352.720 335.880 ;
        RECT 353.380 335.620 353.640 335.880 ;
        RECT 352.460 265.580 352.720 265.840 ;
        RECT 353.380 265.580 353.640 265.840 ;
        RECT 352.460 206.760 352.720 207.020 ;
        RECT 353.380 206.760 353.640 207.020 ;
        RECT 352.460 169.020 352.720 169.280 ;
        RECT 353.380 169.020 353.640 169.280 ;
        RECT 352.460 113.260 352.720 113.520 ;
        RECT 353.380 113.260 353.640 113.520 ;
        RECT 353.380 62.600 353.640 62.860 ;
        RECT 352.460 62.260 352.720 62.520 ;
        RECT 8.380 23.840 8.640 24.100 ;
        RECT 352.460 23.840 352.720 24.100 ;
      LAYER met2 ;
        RECT 352.780 1601.130 353.060 1604.000 ;
        RECT 352.060 1600.990 353.060 1601.130 ;
        RECT 352.060 1597.050 352.200 1600.990 ;
        RECT 352.780 1600.000 353.060 1600.990 ;
        RECT 352.060 1596.910 352.660 1597.050 ;
        RECT 352.520 1569.850 352.660 1596.910 ;
        RECT 352.520 1569.710 353.120 1569.850 ;
        RECT 352.980 1511.630 353.120 1569.710 ;
        RECT 352.920 1511.310 353.180 1511.630 ;
        RECT 352.460 1510.630 352.720 1510.950 ;
        RECT 352.520 1497.350 352.660 1510.630 ;
        RECT 352.460 1497.030 352.720 1497.350 ;
        RECT 352.920 1449.090 353.180 1449.410 ;
        RECT 352.980 1400.530 353.120 1449.090 ;
        RECT 352.980 1400.390 353.580 1400.530 ;
        RECT 353.440 1320.550 353.580 1400.390 ;
        RECT 352.460 1320.230 352.720 1320.550 ;
        RECT 353.380 1320.230 353.640 1320.550 ;
        RECT 352.520 1269.550 352.660 1320.230 ;
        RECT 352.460 1269.230 352.720 1269.550 ;
        RECT 353.380 1269.230 353.640 1269.550 ;
        RECT 353.440 1221.950 353.580 1269.230 ;
        RECT 353.380 1221.630 353.640 1221.950 ;
        RECT 352.460 1221.290 352.720 1221.610 ;
        RECT 352.520 1172.990 352.660 1221.290 ;
        RECT 352.460 1172.670 352.720 1172.990 ;
        RECT 353.380 1172.670 353.640 1172.990 ;
        RECT 353.440 1125.390 353.580 1172.670 ;
        RECT 353.380 1125.070 353.640 1125.390 ;
        RECT 352.460 1124.730 352.720 1125.050 ;
        RECT 352.520 1076.430 352.660 1124.730 ;
        RECT 352.460 1076.110 352.720 1076.430 ;
        RECT 353.380 1076.110 353.640 1076.430 ;
        RECT 353.440 1028.830 353.580 1076.110 ;
        RECT 353.380 1028.510 353.640 1028.830 ;
        RECT 352.460 1028.170 352.720 1028.490 ;
        RECT 352.520 979.870 352.660 1028.170 ;
        RECT 352.460 979.550 352.720 979.870 ;
        RECT 353.380 979.550 353.640 979.870 ;
        RECT 353.440 932.270 353.580 979.550 ;
        RECT 353.380 931.950 353.640 932.270 ;
        RECT 352.460 931.610 352.720 931.930 ;
        RECT 352.520 883.310 352.660 931.610 ;
        RECT 352.460 882.990 352.720 883.310 ;
        RECT 353.380 882.990 353.640 883.310 ;
        RECT 353.440 835.710 353.580 882.990 ;
        RECT 353.380 835.390 353.640 835.710 ;
        RECT 352.460 835.050 352.720 835.370 ;
        RECT 352.520 786.750 352.660 835.050 ;
        RECT 352.460 786.430 352.720 786.750 ;
        RECT 353.840 786.430 354.100 786.750 ;
        RECT 353.900 738.470 354.040 786.430 ;
        RECT 352.460 738.150 352.720 738.470 ;
        RECT 353.840 738.150 354.100 738.470 ;
        RECT 352.520 700.130 352.660 738.150 ;
        RECT 352.520 699.990 353.580 700.130 ;
        RECT 353.440 642.250 353.580 699.990 ;
        RECT 353.380 641.930 353.640 642.250 ;
        RECT 352.460 641.590 352.720 641.910 ;
        RECT 352.520 627.970 352.660 641.590 ;
        RECT 352.460 627.650 352.720 627.970 ;
        RECT 353.380 627.650 353.640 627.970 ;
        RECT 353.440 545.690 353.580 627.650 ;
        RECT 353.380 545.370 353.640 545.690 ;
        RECT 352.460 545.030 352.720 545.350 ;
        RECT 352.520 476.330 352.660 545.030 ;
        RECT 352.460 476.010 352.720 476.330 ;
        RECT 353.380 476.010 353.640 476.330 ;
        RECT 353.440 449.130 353.580 476.010 ;
        RECT 353.380 448.810 353.640 449.130 ;
        RECT 352.460 448.470 352.720 448.790 ;
        RECT 352.520 419.290 352.660 448.470 ;
        RECT 352.520 419.150 353.580 419.290 ;
        RECT 353.440 357.330 353.580 419.150 ;
        RECT 352.460 357.010 352.720 357.330 ;
        RECT 353.380 357.010 353.640 357.330 ;
        RECT 352.520 335.910 352.660 357.010 ;
        RECT 352.460 335.590 352.720 335.910 ;
        RECT 353.380 335.590 353.640 335.910 ;
        RECT 353.440 265.870 353.580 335.590 ;
        RECT 352.460 265.550 352.720 265.870 ;
        RECT 353.380 265.550 353.640 265.870 ;
        RECT 352.520 207.050 352.660 265.550 ;
        RECT 352.460 206.730 352.720 207.050 ;
        RECT 353.380 206.730 353.640 207.050 ;
        RECT 353.440 169.310 353.580 206.730 ;
        RECT 352.460 168.990 352.720 169.310 ;
        RECT 353.380 168.990 353.640 169.310 ;
        RECT 352.520 113.550 352.660 168.990 ;
        RECT 352.460 113.230 352.720 113.550 ;
        RECT 353.380 113.230 353.640 113.550 ;
        RECT 353.440 62.890 353.580 113.230 ;
        RECT 353.380 62.570 353.640 62.890 ;
        RECT 352.460 62.230 352.720 62.550 ;
        RECT 352.520 24.130 352.660 62.230 ;
        RECT 8.380 23.810 8.640 24.130 ;
        RECT 352.460 23.810 352.720 24.130 ;
        RECT 8.440 2.400 8.580 23.810 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 354.345 1538.925 354.515 1545.895 ;
        RECT 353.885 1442.025 354.055 1490.475 ;
        RECT 353.885 1207.425 354.055 1297.015 ;
        RECT 353.885 1159.145 354.055 1172.915 ;
        RECT 353.885 1062.585 354.055 1076.355 ;
        RECT 353.885 966.025 354.055 979.795 ;
        RECT 353.885 869.465 354.055 883.235 ;
        RECT 353.425 772.905 353.595 787.355 ;
        RECT 353.885 476.425 354.055 524.195 ;
        RECT 353.425 289.765 353.595 337.875 ;
      LAYER mcon ;
        RECT 354.345 1545.725 354.515 1545.895 ;
        RECT 353.885 1490.305 354.055 1490.475 ;
        RECT 353.885 1296.845 354.055 1297.015 ;
        RECT 353.885 1172.745 354.055 1172.915 ;
        RECT 353.885 1076.185 354.055 1076.355 ;
        RECT 353.885 979.625 354.055 979.795 ;
        RECT 353.885 883.065 354.055 883.235 ;
        RECT 353.425 787.185 353.595 787.355 ;
        RECT 353.885 524.025 354.055 524.195 ;
        RECT 353.425 337.705 353.595 337.875 ;
      LAYER met1 ;
        RECT 354.270 1545.880 354.590 1545.940 ;
        RECT 354.075 1545.740 354.590 1545.880 ;
        RECT 354.270 1545.680 354.590 1545.740 ;
        RECT 354.270 1539.080 354.590 1539.140 ;
        RECT 354.075 1538.940 354.590 1539.080 ;
        RECT 354.270 1538.880 354.590 1538.940 ;
        RECT 353.350 1497.600 353.670 1497.660 ;
        RECT 354.270 1497.600 354.590 1497.660 ;
        RECT 353.350 1497.460 354.590 1497.600 ;
        RECT 353.350 1497.400 353.670 1497.460 ;
        RECT 354.270 1497.400 354.590 1497.460 ;
        RECT 353.810 1490.460 354.130 1490.520 ;
        RECT 353.615 1490.320 354.130 1490.460 ;
        RECT 353.810 1490.260 354.130 1490.320 ;
        RECT 353.810 1442.180 354.130 1442.240 ;
        RECT 353.615 1442.040 354.130 1442.180 ;
        RECT 353.810 1441.980 354.130 1442.040 ;
        RECT 353.810 1414.440 354.130 1414.700 ;
        RECT 353.900 1414.300 354.040 1414.440 ;
        RECT 354.270 1414.300 354.590 1414.360 ;
        RECT 353.900 1414.160 354.590 1414.300 ;
        RECT 354.270 1414.100 354.590 1414.160 ;
        RECT 353.810 1352.760 354.130 1352.820 ;
        RECT 354.270 1352.760 354.590 1352.820 ;
        RECT 353.810 1352.620 354.590 1352.760 ;
        RECT 353.810 1352.560 354.130 1352.620 ;
        RECT 354.270 1352.560 354.590 1352.620 ;
        RECT 353.810 1318.080 354.130 1318.140 ;
        RECT 353.440 1317.940 354.130 1318.080 ;
        RECT 353.440 1317.800 353.580 1317.940 ;
        RECT 353.810 1317.880 354.130 1317.940 ;
        RECT 353.350 1317.540 353.670 1317.800 ;
        RECT 353.350 1297.000 353.670 1297.060 ;
        RECT 353.825 1297.000 354.115 1297.045 ;
        RECT 353.350 1296.860 354.115 1297.000 ;
        RECT 353.350 1296.800 353.670 1296.860 ;
        RECT 353.825 1296.815 354.115 1296.860 ;
        RECT 353.810 1207.580 354.130 1207.640 ;
        RECT 353.615 1207.440 354.130 1207.580 ;
        RECT 353.810 1207.380 354.130 1207.440 ;
        RECT 353.810 1172.900 354.130 1172.960 ;
        RECT 353.810 1172.760 354.325 1172.900 ;
        RECT 353.810 1172.700 354.130 1172.760 ;
        RECT 353.810 1159.300 354.130 1159.360 ;
        RECT 353.615 1159.160 354.130 1159.300 ;
        RECT 353.810 1159.100 354.130 1159.160 ;
        RECT 353.810 1076.340 354.130 1076.400 ;
        RECT 353.810 1076.200 354.325 1076.340 ;
        RECT 353.810 1076.140 354.130 1076.200 ;
        RECT 353.810 1062.740 354.130 1062.800 ;
        RECT 353.615 1062.600 354.130 1062.740 ;
        RECT 353.810 1062.540 354.130 1062.600 ;
        RECT 353.810 979.780 354.130 979.840 ;
        RECT 353.810 979.640 354.325 979.780 ;
        RECT 353.810 979.580 354.130 979.640 ;
        RECT 353.810 966.180 354.130 966.240 ;
        RECT 353.615 966.040 354.130 966.180 ;
        RECT 353.810 965.980 354.130 966.040 ;
        RECT 353.810 883.220 354.130 883.280 ;
        RECT 353.810 883.080 354.325 883.220 ;
        RECT 353.810 883.020 354.130 883.080 ;
        RECT 353.810 869.620 354.130 869.680 ;
        RECT 353.615 869.480 354.130 869.620 ;
        RECT 353.810 869.420 354.130 869.480 ;
        RECT 353.365 787.340 353.655 787.385 ;
        RECT 353.810 787.340 354.130 787.400 ;
        RECT 353.365 787.200 354.130 787.340 ;
        RECT 353.365 787.155 353.655 787.200 ;
        RECT 353.810 787.140 354.130 787.200 ;
        RECT 353.350 773.060 353.670 773.120 ;
        RECT 353.155 772.920 353.670 773.060 ;
        RECT 353.350 772.860 353.670 772.920 ;
        RECT 353.810 641.960 354.130 642.220 ;
        RECT 352.890 641.480 353.210 641.540 ;
        RECT 353.900 641.480 354.040 641.960 ;
        RECT 352.890 641.340 354.040 641.480 ;
        RECT 352.890 641.280 353.210 641.340 ;
        RECT 352.890 627.540 353.210 627.600 ;
        RECT 353.810 627.540 354.130 627.600 ;
        RECT 352.890 627.400 354.130 627.540 ;
        RECT 352.890 627.340 353.210 627.400 ;
        RECT 353.810 627.340 354.130 627.400 ;
        RECT 353.810 620.740 354.130 620.800 ;
        RECT 354.270 620.740 354.590 620.800 ;
        RECT 353.810 620.600 354.590 620.740 ;
        RECT 353.810 620.540 354.130 620.600 ;
        RECT 354.270 620.540 354.590 620.600 ;
        RECT 353.825 524.180 354.115 524.225 ;
        RECT 354.270 524.180 354.590 524.240 ;
        RECT 353.825 524.040 354.590 524.180 ;
        RECT 353.825 523.995 354.115 524.040 ;
        RECT 354.270 523.980 354.590 524.040 ;
        RECT 353.810 476.580 354.130 476.640 ;
        RECT 353.615 476.440 354.130 476.580 ;
        RECT 353.810 476.380 354.130 476.440 ;
        RECT 353.810 475.900 354.130 475.960 ;
        RECT 354.730 475.900 355.050 475.960 ;
        RECT 353.810 475.760 355.050 475.900 ;
        RECT 353.810 475.700 354.130 475.760 ;
        RECT 354.730 475.700 355.050 475.760 ;
        RECT 353.810 352.480 354.130 352.540 ;
        RECT 353.440 352.340 354.130 352.480 ;
        RECT 353.440 351.860 353.580 352.340 ;
        RECT 353.810 352.280 354.130 352.340 ;
        RECT 353.350 351.600 353.670 351.860 ;
        RECT 353.350 337.860 353.670 337.920 ;
        RECT 353.155 337.720 353.670 337.860 ;
        RECT 353.350 337.660 353.670 337.720 ;
        RECT 353.365 289.920 353.655 289.965 ;
        RECT 353.810 289.920 354.130 289.980 ;
        RECT 353.365 289.780 354.130 289.920 ;
        RECT 353.365 289.735 353.655 289.780 ;
        RECT 353.810 289.720 354.130 289.780 ;
        RECT 353.810 255.580 354.130 255.640 ;
        RECT 353.440 255.440 354.130 255.580 ;
        RECT 353.440 255.300 353.580 255.440 ;
        RECT 353.810 255.380 354.130 255.440 ;
        RECT 353.350 255.040 353.670 255.300 ;
        RECT 352.890 206.620 353.210 206.680 ;
        RECT 353.810 206.620 354.130 206.680 ;
        RECT 352.890 206.480 354.130 206.620 ;
        RECT 352.890 206.420 353.210 206.480 ;
        RECT 353.810 206.420 354.130 206.480 ;
        RECT 353.810 159.020 354.130 159.080 ;
        RECT 353.440 158.880 354.130 159.020 ;
        RECT 353.440 158.740 353.580 158.880 ;
        RECT 353.810 158.820 354.130 158.880 ;
        RECT 353.350 158.480 353.670 158.740 ;
        RECT 14.330 24.720 14.650 24.780 ;
        RECT 353.810 24.720 354.130 24.780 ;
        RECT 14.330 24.580 354.130 24.720 ;
        RECT 14.330 24.520 14.650 24.580 ;
        RECT 353.810 24.520 354.130 24.580 ;
      LAYER via ;
        RECT 354.300 1545.680 354.560 1545.940 ;
        RECT 354.300 1538.880 354.560 1539.140 ;
        RECT 353.380 1497.400 353.640 1497.660 ;
        RECT 354.300 1497.400 354.560 1497.660 ;
        RECT 353.840 1490.260 354.100 1490.520 ;
        RECT 353.840 1441.980 354.100 1442.240 ;
        RECT 353.840 1414.440 354.100 1414.700 ;
        RECT 354.300 1414.100 354.560 1414.360 ;
        RECT 353.840 1352.560 354.100 1352.820 ;
        RECT 354.300 1352.560 354.560 1352.820 ;
        RECT 353.840 1317.880 354.100 1318.140 ;
        RECT 353.380 1317.540 353.640 1317.800 ;
        RECT 353.380 1296.800 353.640 1297.060 ;
        RECT 353.840 1207.380 354.100 1207.640 ;
        RECT 353.840 1172.700 354.100 1172.960 ;
        RECT 353.840 1159.100 354.100 1159.360 ;
        RECT 353.840 1076.140 354.100 1076.400 ;
        RECT 353.840 1062.540 354.100 1062.800 ;
        RECT 353.840 979.580 354.100 979.840 ;
        RECT 353.840 965.980 354.100 966.240 ;
        RECT 353.840 883.020 354.100 883.280 ;
        RECT 353.840 869.420 354.100 869.680 ;
        RECT 353.840 787.140 354.100 787.400 ;
        RECT 353.380 772.860 353.640 773.120 ;
        RECT 353.840 641.960 354.100 642.220 ;
        RECT 352.920 641.280 353.180 641.540 ;
        RECT 352.920 627.340 353.180 627.600 ;
        RECT 353.840 627.340 354.100 627.600 ;
        RECT 353.840 620.540 354.100 620.800 ;
        RECT 354.300 620.540 354.560 620.800 ;
        RECT 354.300 523.980 354.560 524.240 ;
        RECT 353.840 476.380 354.100 476.640 ;
        RECT 353.840 475.700 354.100 475.960 ;
        RECT 354.760 475.700 355.020 475.960 ;
        RECT 353.840 352.280 354.100 352.540 ;
        RECT 353.380 351.600 353.640 351.860 ;
        RECT 353.380 337.660 353.640 337.920 ;
        RECT 353.840 289.720 354.100 289.980 ;
        RECT 353.840 255.380 354.100 255.640 ;
        RECT 353.380 255.040 353.640 255.300 ;
        RECT 352.920 206.420 353.180 206.680 ;
        RECT 353.840 206.420 354.100 206.680 ;
        RECT 353.840 158.820 354.100 159.080 ;
        RECT 353.380 158.480 353.640 158.740 ;
        RECT 14.360 24.520 14.620 24.780 ;
        RECT 353.840 24.520 354.100 24.780 ;
      LAYER met2 ;
        RECT 354.620 1601.130 354.900 1604.000 ;
        RECT 353.900 1600.990 354.900 1601.130 ;
        RECT 353.900 1597.050 354.040 1600.990 ;
        RECT 354.620 1600.000 354.900 1600.990 ;
        RECT 353.900 1596.910 354.500 1597.050 ;
        RECT 354.360 1545.970 354.500 1596.910 ;
        RECT 354.300 1545.650 354.560 1545.970 ;
        RECT 354.300 1538.850 354.560 1539.170 ;
        RECT 354.360 1497.690 354.500 1538.850 ;
        RECT 353.380 1497.370 353.640 1497.690 ;
        RECT 354.300 1497.370 354.560 1497.690 ;
        RECT 353.440 1497.090 353.580 1497.370 ;
        RECT 353.440 1496.950 354.040 1497.090 ;
        RECT 353.900 1490.550 354.040 1496.950 ;
        RECT 353.840 1490.230 354.100 1490.550 ;
        RECT 353.840 1441.950 354.100 1442.270 ;
        RECT 353.900 1414.730 354.040 1441.950 ;
        RECT 353.840 1414.410 354.100 1414.730 ;
        RECT 354.300 1414.070 354.560 1414.390 ;
        RECT 354.360 1352.850 354.500 1414.070 ;
        RECT 353.840 1352.530 354.100 1352.850 ;
        RECT 354.300 1352.530 354.560 1352.850 ;
        RECT 353.900 1318.170 354.040 1352.530 ;
        RECT 353.840 1317.850 354.100 1318.170 ;
        RECT 353.380 1317.510 353.640 1317.830 ;
        RECT 353.440 1297.090 353.580 1317.510 ;
        RECT 353.380 1296.770 353.640 1297.090 ;
        RECT 353.840 1207.350 354.100 1207.670 ;
        RECT 353.900 1172.990 354.040 1207.350 ;
        RECT 353.840 1172.670 354.100 1172.990 ;
        RECT 353.840 1159.070 354.100 1159.390 ;
        RECT 353.900 1076.430 354.040 1159.070 ;
        RECT 353.840 1076.110 354.100 1076.430 ;
        RECT 353.840 1062.510 354.100 1062.830 ;
        RECT 353.900 979.870 354.040 1062.510 ;
        RECT 353.840 979.550 354.100 979.870 ;
        RECT 353.840 965.950 354.100 966.270 ;
        RECT 353.900 883.310 354.040 965.950 ;
        RECT 353.840 882.990 354.100 883.310 ;
        RECT 353.840 869.390 354.100 869.710 ;
        RECT 353.900 787.430 354.040 869.390 ;
        RECT 353.840 787.110 354.100 787.430 ;
        RECT 353.380 772.830 353.640 773.150 ;
        RECT 353.440 702.170 353.580 772.830 ;
        RECT 353.440 702.030 354.960 702.170 ;
        RECT 354.820 676.445 354.960 702.030 ;
        RECT 353.830 676.075 354.110 676.445 ;
        RECT 354.750 676.075 355.030 676.445 ;
        RECT 353.900 642.250 354.040 676.075 ;
        RECT 353.840 641.930 354.100 642.250 ;
        RECT 352.920 641.250 353.180 641.570 ;
        RECT 352.980 627.630 353.120 641.250 ;
        RECT 352.920 627.310 353.180 627.630 ;
        RECT 353.840 627.310 354.100 627.630 ;
        RECT 353.900 620.830 354.040 627.310 ;
        RECT 353.840 620.510 354.100 620.830 ;
        RECT 354.300 620.510 354.560 620.830 ;
        RECT 354.360 524.270 354.500 620.510 ;
        RECT 354.300 523.950 354.560 524.270 ;
        RECT 353.840 476.350 354.100 476.670 ;
        RECT 353.900 475.990 354.040 476.350 ;
        RECT 353.840 475.670 354.100 475.990 ;
        RECT 354.760 475.670 355.020 475.990 ;
        RECT 354.820 386.765 354.960 475.670 ;
        RECT 353.830 386.395 354.110 386.765 ;
        RECT 354.750 386.395 355.030 386.765 ;
        RECT 353.900 352.570 354.040 386.395 ;
        RECT 353.840 352.250 354.100 352.570 ;
        RECT 353.380 351.570 353.640 351.890 ;
        RECT 353.440 337.950 353.580 351.570 ;
        RECT 353.380 337.630 353.640 337.950 ;
        RECT 353.840 289.690 354.100 290.010 ;
        RECT 353.900 255.670 354.040 289.690 ;
        RECT 353.840 255.350 354.100 255.670 ;
        RECT 353.380 255.010 353.640 255.330 ;
        RECT 353.440 230.930 353.580 255.010 ;
        RECT 352.980 230.790 353.580 230.930 ;
        RECT 352.980 206.710 353.120 230.790 ;
        RECT 352.920 206.390 353.180 206.710 ;
        RECT 353.840 206.390 354.100 206.710 ;
        RECT 353.900 159.110 354.040 206.390 ;
        RECT 353.840 158.790 354.100 159.110 ;
        RECT 353.380 158.450 353.640 158.770 ;
        RECT 353.440 114.650 353.580 158.450 ;
        RECT 353.440 114.510 354.040 114.650 ;
        RECT 353.900 24.810 354.040 114.510 ;
        RECT 14.360 24.490 14.620 24.810 ;
        RECT 353.840 24.490 354.100 24.810 ;
        RECT 14.420 2.400 14.560 24.490 ;
        RECT 14.210 -4.800 14.770 2.400 ;
      LAYER via2 ;
        RECT 353.830 676.120 354.110 676.400 ;
        RECT 354.750 676.120 355.030 676.400 ;
        RECT 353.830 386.440 354.110 386.720 ;
        RECT 354.750 386.440 355.030 386.720 ;
      LAYER met3 ;
        RECT 353.805 676.410 354.135 676.425 ;
        RECT 354.725 676.410 355.055 676.425 ;
        RECT 353.805 676.110 355.055 676.410 ;
        RECT 353.805 676.095 354.135 676.110 ;
        RECT 354.725 676.095 355.055 676.110 ;
        RECT 353.805 386.730 354.135 386.745 ;
        RECT 354.725 386.730 355.055 386.745 ;
        RECT 353.805 386.430 355.055 386.730 ;
        RECT 353.805 386.415 354.135 386.430 ;
        RECT 354.725 386.415 355.055 386.430 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 360.785 1441.685 360.955 1483.335 ;
        RECT 361.705 855.525 361.875 870.315 ;
        RECT 361.705 620.925 361.875 669.375 ;
        RECT 361.245 483.565 361.415 531.335 ;
        RECT 360.785 379.525 360.955 427.635 ;
        RECT 360.785 338.385 360.955 362.355 ;
        RECT 360.325 282.965 360.495 331.075 ;
        RECT 360.325 186.405 360.495 234.515 ;
      LAYER mcon ;
        RECT 360.785 1483.165 360.955 1483.335 ;
        RECT 361.705 870.145 361.875 870.315 ;
        RECT 361.705 669.205 361.875 669.375 ;
        RECT 361.245 531.165 361.415 531.335 ;
        RECT 360.785 427.465 360.955 427.635 ;
        RECT 360.785 362.185 360.955 362.355 ;
        RECT 360.325 330.905 360.495 331.075 ;
        RECT 360.325 234.345 360.495 234.515 ;
      LAYER met1 ;
        RECT 360.710 1483.320 361.030 1483.380 ;
        RECT 360.515 1483.180 361.030 1483.320 ;
        RECT 360.710 1483.120 361.030 1483.180 ;
        RECT 360.725 1441.840 361.015 1441.885 ;
        RECT 361.630 1441.840 361.950 1441.900 ;
        RECT 360.725 1441.700 361.950 1441.840 ;
        RECT 360.725 1441.655 361.015 1441.700 ;
        RECT 361.630 1441.640 361.950 1441.700 ;
        RECT 361.630 1387.100 361.950 1387.160 ;
        RECT 362.550 1387.100 362.870 1387.160 ;
        RECT 361.630 1386.960 362.870 1387.100 ;
        RECT 361.630 1386.900 361.950 1386.960 ;
        RECT 362.550 1386.900 362.870 1386.960 ;
        RECT 362.090 1338.820 362.410 1338.880 ;
        RECT 363.010 1338.820 363.330 1338.880 ;
        RECT 362.090 1338.680 363.330 1338.820 ;
        RECT 362.090 1338.620 362.410 1338.680 ;
        RECT 363.010 1338.620 363.330 1338.680 ;
        RECT 360.710 1249.060 361.030 1249.120 ;
        RECT 362.090 1249.060 362.410 1249.120 ;
        RECT 360.710 1248.920 362.410 1249.060 ;
        RECT 360.710 1248.860 361.030 1248.920 ;
        RECT 362.090 1248.860 362.410 1248.920 ;
        RECT 361.170 1200.780 361.490 1200.840 ;
        RECT 362.090 1200.780 362.410 1200.840 ;
        RECT 361.170 1200.640 362.410 1200.780 ;
        RECT 361.170 1200.580 361.490 1200.640 ;
        RECT 362.090 1200.580 362.410 1200.640 ;
        RECT 360.710 1159.300 361.030 1159.360 ;
        RECT 362.090 1159.300 362.410 1159.360 ;
        RECT 360.710 1159.160 362.410 1159.300 ;
        RECT 360.710 1159.100 361.030 1159.160 ;
        RECT 362.090 1159.100 362.410 1159.160 ;
        RECT 360.710 1111.020 361.030 1111.080 ;
        RECT 362.090 1111.020 362.410 1111.080 ;
        RECT 360.710 1110.880 362.410 1111.020 ;
        RECT 360.710 1110.820 361.030 1110.880 ;
        RECT 362.090 1110.820 362.410 1110.880 ;
        RECT 360.710 1062.740 361.030 1062.800 ;
        RECT 362.090 1062.740 362.410 1062.800 ;
        RECT 360.710 1062.600 362.410 1062.740 ;
        RECT 360.710 1062.540 361.030 1062.600 ;
        RECT 362.090 1062.540 362.410 1062.600 ;
        RECT 360.710 1014.460 361.030 1014.520 ;
        RECT 362.090 1014.460 362.410 1014.520 ;
        RECT 360.710 1014.320 362.410 1014.460 ;
        RECT 360.710 1014.260 361.030 1014.320 ;
        RECT 362.090 1014.260 362.410 1014.320 ;
        RECT 360.710 966.180 361.030 966.240 ;
        RECT 362.090 966.180 362.410 966.240 ;
        RECT 360.710 966.040 362.410 966.180 ;
        RECT 360.710 965.980 361.030 966.040 ;
        RECT 362.090 965.980 362.410 966.040 ;
        RECT 360.250 959.040 360.570 959.100 ;
        RECT 360.710 959.040 361.030 959.100 ;
        RECT 360.250 958.900 361.030 959.040 ;
        RECT 360.250 958.840 360.570 958.900 ;
        RECT 360.710 958.840 361.030 958.900 ;
        RECT 361.630 870.300 361.950 870.360 ;
        RECT 361.435 870.160 361.950 870.300 ;
        RECT 361.630 870.100 361.950 870.160 ;
        RECT 361.630 855.680 361.950 855.740 ;
        RECT 361.435 855.540 361.950 855.680 ;
        RECT 361.630 855.480 361.950 855.540 ;
        RECT 360.710 759.120 361.030 759.180 ;
        RECT 361.630 759.120 361.950 759.180 ;
        RECT 360.710 758.980 361.950 759.120 ;
        RECT 360.710 758.920 361.030 758.980 ;
        RECT 361.630 758.920 361.950 758.980 ;
        RECT 360.710 717.640 361.030 717.700 ;
        RECT 361.630 717.640 361.950 717.700 ;
        RECT 360.710 717.500 361.950 717.640 ;
        RECT 360.710 717.440 361.030 717.500 ;
        RECT 361.630 717.440 361.950 717.500 ;
        RECT 361.630 669.360 361.950 669.420 ;
        RECT 361.435 669.220 361.950 669.360 ;
        RECT 361.630 669.160 361.950 669.220 ;
        RECT 361.630 621.080 361.950 621.140 ;
        RECT 361.435 620.940 361.950 621.080 ;
        RECT 361.630 620.880 361.950 620.940 ;
        RECT 360.710 572.800 361.030 572.860 ;
        RECT 361.170 572.800 361.490 572.860 ;
        RECT 360.710 572.660 361.490 572.800 ;
        RECT 360.710 572.600 361.030 572.660 ;
        RECT 361.170 572.600 361.490 572.660 ;
        RECT 361.170 531.320 361.490 531.380 ;
        RECT 360.975 531.180 361.490 531.320 ;
        RECT 361.170 531.120 361.490 531.180 ;
        RECT 361.170 483.720 361.490 483.780 ;
        RECT 360.975 483.580 361.490 483.720 ;
        RECT 361.170 483.520 361.490 483.580 ;
        RECT 360.710 427.620 361.030 427.680 ;
        RECT 360.515 427.480 361.030 427.620 ;
        RECT 360.710 427.420 361.030 427.480 ;
        RECT 360.710 379.680 361.030 379.740 ;
        RECT 360.515 379.540 361.030 379.680 ;
        RECT 360.710 379.480 361.030 379.540 ;
        RECT 360.710 362.340 361.030 362.400 ;
        RECT 360.515 362.200 361.030 362.340 ;
        RECT 360.710 362.140 361.030 362.200 ;
        RECT 360.710 338.540 361.030 338.600 ;
        RECT 360.515 338.400 361.030 338.540 ;
        RECT 360.710 338.340 361.030 338.400 ;
        RECT 360.265 331.060 360.555 331.105 ;
        RECT 360.710 331.060 361.030 331.120 ;
        RECT 360.265 330.920 361.030 331.060 ;
        RECT 360.265 330.875 360.555 330.920 ;
        RECT 360.710 330.860 361.030 330.920 ;
        RECT 360.250 283.120 360.570 283.180 ;
        RECT 360.055 282.980 360.570 283.120 ;
        RECT 360.250 282.920 360.570 282.980 ;
        RECT 360.250 241.640 360.570 241.700 ;
        RECT 361.170 241.640 361.490 241.700 ;
        RECT 360.250 241.500 361.490 241.640 ;
        RECT 360.250 241.440 360.570 241.500 ;
        RECT 361.170 241.440 361.490 241.500 ;
        RECT 360.265 234.500 360.555 234.545 ;
        RECT 361.170 234.500 361.490 234.560 ;
        RECT 360.265 234.360 361.490 234.500 ;
        RECT 360.265 234.315 360.555 234.360 ;
        RECT 361.170 234.300 361.490 234.360 ;
        RECT 360.250 186.560 360.570 186.620 ;
        RECT 360.055 186.420 360.570 186.560 ;
        RECT 360.250 186.360 360.570 186.420 ;
        RECT 360.250 145.080 360.570 145.140 ;
        RECT 361.170 145.080 361.490 145.140 ;
        RECT 360.250 144.940 361.490 145.080 ;
        RECT 360.250 144.880 360.570 144.940 ;
        RECT 361.170 144.880 361.490 144.940 ;
        RECT 361.170 110.740 361.490 110.800 ;
        RECT 360.800 110.600 361.490 110.740 ;
        RECT 360.800 110.460 360.940 110.600 ;
        RECT 361.170 110.540 361.490 110.600 ;
        RECT 360.710 110.200 361.030 110.460 ;
        RECT 38.250 25.060 38.570 25.120 ;
        RECT 360.710 25.060 361.030 25.120 ;
        RECT 38.250 24.920 361.030 25.060 ;
        RECT 38.250 24.860 38.570 24.920 ;
        RECT 360.710 24.860 361.030 24.920 ;
      LAYER via ;
        RECT 360.740 1483.120 361.000 1483.380 ;
        RECT 361.660 1441.640 361.920 1441.900 ;
        RECT 361.660 1386.900 361.920 1387.160 ;
        RECT 362.580 1386.900 362.840 1387.160 ;
        RECT 362.120 1338.620 362.380 1338.880 ;
        RECT 363.040 1338.620 363.300 1338.880 ;
        RECT 360.740 1248.860 361.000 1249.120 ;
        RECT 362.120 1248.860 362.380 1249.120 ;
        RECT 361.200 1200.580 361.460 1200.840 ;
        RECT 362.120 1200.580 362.380 1200.840 ;
        RECT 360.740 1159.100 361.000 1159.360 ;
        RECT 362.120 1159.100 362.380 1159.360 ;
        RECT 360.740 1110.820 361.000 1111.080 ;
        RECT 362.120 1110.820 362.380 1111.080 ;
        RECT 360.740 1062.540 361.000 1062.800 ;
        RECT 362.120 1062.540 362.380 1062.800 ;
        RECT 360.740 1014.260 361.000 1014.520 ;
        RECT 362.120 1014.260 362.380 1014.520 ;
        RECT 360.740 965.980 361.000 966.240 ;
        RECT 362.120 965.980 362.380 966.240 ;
        RECT 360.280 958.840 360.540 959.100 ;
        RECT 360.740 958.840 361.000 959.100 ;
        RECT 361.660 870.100 361.920 870.360 ;
        RECT 361.660 855.480 361.920 855.740 ;
        RECT 360.740 758.920 361.000 759.180 ;
        RECT 361.660 758.920 361.920 759.180 ;
        RECT 360.740 717.440 361.000 717.700 ;
        RECT 361.660 717.440 361.920 717.700 ;
        RECT 361.660 669.160 361.920 669.420 ;
        RECT 361.660 620.880 361.920 621.140 ;
        RECT 360.740 572.600 361.000 572.860 ;
        RECT 361.200 572.600 361.460 572.860 ;
        RECT 361.200 531.120 361.460 531.380 ;
        RECT 361.200 483.520 361.460 483.780 ;
        RECT 360.740 427.420 361.000 427.680 ;
        RECT 360.740 379.480 361.000 379.740 ;
        RECT 360.740 362.140 361.000 362.400 ;
        RECT 360.740 338.340 361.000 338.600 ;
        RECT 360.740 330.860 361.000 331.120 ;
        RECT 360.280 282.920 360.540 283.180 ;
        RECT 360.280 241.440 360.540 241.700 ;
        RECT 361.200 241.440 361.460 241.700 ;
        RECT 361.200 234.300 361.460 234.560 ;
        RECT 360.280 186.360 360.540 186.620 ;
        RECT 360.280 144.880 360.540 145.140 ;
        RECT 361.200 144.880 361.460 145.140 ;
        RECT 361.200 110.540 361.460 110.800 ;
        RECT 360.740 110.200 361.000 110.460 ;
        RECT 38.280 24.860 38.540 25.120 ;
        RECT 360.740 24.860 361.000 25.120 ;
      LAYER met2 ;
        RECT 362.900 1600.450 363.180 1604.000 ;
        RECT 362.180 1600.310 363.180 1600.450 ;
        RECT 362.180 1546.560 362.320 1600.310 ;
        RECT 362.900 1600.000 363.180 1600.310 ;
        RECT 361.720 1546.420 362.320 1546.560 ;
        RECT 361.720 1546.050 361.860 1546.420 ;
        RECT 361.260 1545.910 361.860 1546.050 ;
        RECT 361.260 1512.050 361.400 1545.910 ;
        RECT 361.260 1511.910 361.860 1512.050 ;
        RECT 361.720 1510.690 361.860 1511.910 ;
        RECT 360.800 1510.550 361.860 1510.690 ;
        RECT 360.800 1483.410 360.940 1510.550 ;
        RECT 360.740 1483.090 361.000 1483.410 ;
        RECT 361.660 1441.610 361.920 1441.930 ;
        RECT 361.720 1435.325 361.860 1441.610 ;
        RECT 361.650 1434.955 361.930 1435.325 ;
        RECT 362.570 1434.955 362.850 1435.325 ;
        RECT 362.640 1387.190 362.780 1434.955 ;
        RECT 361.660 1387.045 361.920 1387.190 ;
        RECT 361.650 1386.675 361.930 1387.045 ;
        RECT 362.580 1386.870 362.840 1387.190 ;
        RECT 363.030 1386.675 363.310 1387.045 ;
        RECT 363.100 1338.910 363.240 1386.675 ;
        RECT 362.120 1338.590 362.380 1338.910 ;
        RECT 363.040 1338.590 363.300 1338.910 ;
        RECT 362.180 1249.150 362.320 1338.590 ;
        RECT 360.740 1248.890 361.000 1249.150 ;
        RECT 360.740 1248.830 361.400 1248.890 ;
        RECT 362.120 1248.830 362.380 1249.150 ;
        RECT 360.800 1248.750 361.400 1248.830 ;
        RECT 361.260 1200.870 361.400 1248.750 ;
        RECT 361.200 1200.550 361.460 1200.870 ;
        RECT 362.120 1200.550 362.380 1200.870 ;
        RECT 362.180 1159.390 362.320 1200.550 ;
        RECT 360.740 1159.070 361.000 1159.390 ;
        RECT 362.120 1159.070 362.380 1159.390 ;
        RECT 360.800 1111.110 360.940 1159.070 ;
        RECT 360.740 1110.790 361.000 1111.110 ;
        RECT 362.120 1110.790 362.380 1111.110 ;
        RECT 362.180 1062.830 362.320 1110.790 ;
        RECT 360.740 1062.510 361.000 1062.830 ;
        RECT 362.120 1062.510 362.380 1062.830 ;
        RECT 360.800 1014.550 360.940 1062.510 ;
        RECT 360.740 1014.230 361.000 1014.550 ;
        RECT 362.120 1014.230 362.380 1014.550 ;
        RECT 362.180 966.270 362.320 1014.230 ;
        RECT 360.740 965.950 361.000 966.270 ;
        RECT 362.120 965.950 362.380 966.270 ;
        RECT 360.800 959.130 360.940 965.950 ;
        RECT 360.280 958.810 360.540 959.130 ;
        RECT 360.740 958.810 361.000 959.130 ;
        RECT 360.340 911.045 360.480 958.810 ;
        RECT 360.270 910.675 360.550 911.045 ;
        RECT 361.650 910.675 361.930 911.045 ;
        RECT 361.720 870.390 361.860 910.675 ;
        RECT 361.660 870.070 361.920 870.390 ;
        RECT 361.660 855.450 361.920 855.770 ;
        RECT 361.720 759.210 361.860 855.450 ;
        RECT 360.740 758.890 361.000 759.210 ;
        RECT 361.660 758.890 361.920 759.210 ;
        RECT 360.800 717.730 360.940 758.890 ;
        RECT 360.740 717.410 361.000 717.730 ;
        RECT 361.660 717.410 361.920 717.730 ;
        RECT 361.720 669.450 361.860 717.410 ;
        RECT 361.660 669.130 361.920 669.450 ;
        RECT 361.660 620.850 361.920 621.170 ;
        RECT 361.720 580.450 361.860 620.850 ;
        RECT 361.260 580.310 361.860 580.450 ;
        RECT 361.260 572.890 361.400 580.310 ;
        RECT 360.740 572.570 361.000 572.890 ;
        RECT 361.200 572.570 361.460 572.890 ;
        RECT 360.800 544.920 360.940 572.570 ;
        RECT 360.800 544.780 361.400 544.920 ;
        RECT 361.260 531.410 361.400 544.780 ;
        RECT 361.200 531.090 361.460 531.410 ;
        RECT 361.200 483.490 361.460 483.810 ;
        RECT 361.260 435.725 361.400 483.490 ;
        RECT 361.190 435.355 361.470 435.725 ;
        RECT 360.730 434.675 361.010 435.045 ;
        RECT 360.800 427.710 360.940 434.675 ;
        RECT 360.740 427.390 361.000 427.710 ;
        RECT 360.740 379.450 361.000 379.770 ;
        RECT 360.800 362.430 360.940 379.450 ;
        RECT 360.740 362.110 361.000 362.430 ;
        RECT 360.740 338.310 361.000 338.630 ;
        RECT 360.800 331.150 360.940 338.310 ;
        RECT 360.740 330.830 361.000 331.150 ;
        RECT 360.280 282.890 360.540 283.210 ;
        RECT 360.340 241.730 360.480 282.890 ;
        RECT 360.280 241.410 360.540 241.730 ;
        RECT 361.200 241.410 361.460 241.730 ;
        RECT 361.260 234.590 361.400 241.410 ;
        RECT 361.200 234.270 361.460 234.590 ;
        RECT 360.280 186.330 360.540 186.650 ;
        RECT 360.340 145.170 360.480 186.330 ;
        RECT 360.280 144.850 360.540 145.170 ;
        RECT 361.200 144.850 361.460 145.170 ;
        RECT 361.260 110.830 361.400 144.850 ;
        RECT 361.200 110.510 361.460 110.830 ;
        RECT 360.740 110.170 361.000 110.490 ;
        RECT 360.800 25.150 360.940 110.170 ;
        RECT 38.280 24.830 38.540 25.150 ;
        RECT 360.740 24.830 361.000 25.150 ;
        RECT 38.340 2.400 38.480 24.830 ;
        RECT 38.130 -4.800 38.690 2.400 ;
      LAYER via2 ;
        RECT 361.650 1435.000 361.930 1435.280 ;
        RECT 362.570 1435.000 362.850 1435.280 ;
        RECT 361.650 1386.720 361.930 1387.000 ;
        RECT 363.030 1386.720 363.310 1387.000 ;
        RECT 360.270 910.720 360.550 911.000 ;
        RECT 361.650 910.720 361.930 911.000 ;
        RECT 361.190 435.400 361.470 435.680 ;
        RECT 360.730 434.720 361.010 435.000 ;
      LAYER met3 ;
        RECT 361.625 1435.290 361.955 1435.305 ;
        RECT 362.545 1435.290 362.875 1435.305 ;
        RECT 361.625 1434.990 362.875 1435.290 ;
        RECT 361.625 1434.975 361.955 1434.990 ;
        RECT 362.545 1434.975 362.875 1434.990 ;
        RECT 361.625 1387.010 361.955 1387.025 ;
        RECT 363.005 1387.010 363.335 1387.025 ;
        RECT 361.625 1386.710 363.335 1387.010 ;
        RECT 361.625 1386.695 361.955 1386.710 ;
        RECT 363.005 1386.695 363.335 1386.710 ;
        RECT 360.245 911.010 360.575 911.025 ;
        RECT 361.625 911.010 361.955 911.025 ;
        RECT 360.245 910.710 361.955 911.010 ;
        RECT 360.245 910.695 360.575 910.710 ;
        RECT 361.625 910.695 361.955 910.710 ;
        RECT 361.165 435.690 361.495 435.705 ;
        RECT 360.950 435.375 361.495 435.690 ;
        RECT 360.950 435.025 361.250 435.375 ;
        RECT 360.705 434.710 361.250 435.025 ;
        RECT 360.705 434.695 361.035 434.710 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 241.110 25.400 241.430 25.460 ;
        RECT 428.330 25.400 428.650 25.460 ;
        RECT 241.110 25.260 428.650 25.400 ;
        RECT 241.110 25.200 241.430 25.260 ;
        RECT 428.330 25.200 428.650 25.260 ;
      LAYER via ;
        RECT 241.140 25.200 241.400 25.460 ;
        RECT 428.360 25.200 428.620 25.460 ;
      LAYER met2 ;
        RECT 433.280 1600.450 433.560 1604.000 ;
        RECT 432.100 1600.310 433.560 1600.450 ;
        RECT 432.100 1580.050 432.240 1600.310 ;
        RECT 433.280 1600.000 433.560 1600.310 ;
        RECT 428.420 1579.910 432.240 1580.050 ;
        RECT 428.420 25.490 428.560 1579.910 ;
        RECT 241.140 25.170 241.400 25.490 ;
        RECT 428.360 25.170 428.620 25.490 ;
        RECT 241.200 12.650 241.340 25.170 ;
        RECT 240.740 12.510 241.340 12.650 ;
        RECT 240.740 2.400 240.880 12.510 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 25.740 258.450 25.800 ;
        RECT 435.230 25.740 435.550 25.800 ;
        RECT 258.130 25.600 435.550 25.740 ;
        RECT 258.130 25.540 258.450 25.600 ;
        RECT 435.230 25.540 435.550 25.600 ;
      LAYER via ;
        RECT 258.160 25.540 258.420 25.800 ;
        RECT 435.260 25.540 435.520 25.800 ;
      LAYER met2 ;
        RECT 439.260 1600.450 439.540 1604.000 ;
        RECT 438.540 1600.310 439.540 1600.450 ;
        RECT 438.540 1580.050 438.680 1600.310 ;
        RECT 439.260 1600.000 439.540 1600.310 ;
        RECT 435.320 1579.910 438.680 1580.050 ;
        RECT 435.320 25.830 435.460 1579.910 ;
        RECT 258.160 25.510 258.420 25.830 ;
        RECT 435.260 25.510 435.520 25.830 ;
        RECT 258.220 2.400 258.360 25.510 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 442.130 1579.880 442.450 1579.940 ;
        RECT 444.430 1579.880 444.750 1579.940 ;
        RECT 442.130 1579.740 444.750 1579.880 ;
        RECT 442.130 1579.680 442.450 1579.740 ;
        RECT 444.430 1579.680 444.750 1579.740 ;
        RECT 276.070 26.080 276.390 26.140 ;
        RECT 442.130 26.080 442.450 26.140 ;
        RECT 276.070 25.940 442.450 26.080 ;
        RECT 276.070 25.880 276.390 25.940 ;
        RECT 442.130 25.880 442.450 25.940 ;
      LAYER via ;
        RECT 442.160 1579.680 442.420 1579.940 ;
        RECT 444.460 1579.680 444.720 1579.940 ;
        RECT 276.100 25.880 276.360 26.140 ;
        RECT 442.160 25.880 442.420 26.140 ;
      LAYER met2 ;
        RECT 445.700 1600.450 445.980 1604.000 ;
        RECT 444.520 1600.310 445.980 1600.450 ;
        RECT 444.520 1579.970 444.660 1600.310 ;
        RECT 445.700 1600.000 445.980 1600.310 ;
        RECT 442.160 1579.650 442.420 1579.970 ;
        RECT 444.460 1579.650 444.720 1579.970 ;
        RECT 442.220 26.170 442.360 1579.650 ;
        RECT 276.100 25.850 276.360 26.170 ;
        RECT 442.160 25.850 442.420 26.170 ;
        RECT 276.160 2.400 276.300 25.850 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 26.420 294.330 26.480 ;
        RECT 449.030 26.420 449.350 26.480 ;
        RECT 294.010 26.280 449.350 26.420 ;
        RECT 294.010 26.220 294.330 26.280 ;
        RECT 449.030 26.220 449.350 26.280 ;
      LAYER via ;
        RECT 294.040 26.220 294.300 26.480 ;
        RECT 449.060 26.220 449.320 26.480 ;
      LAYER met2 ;
        RECT 451.680 1600.450 451.960 1604.000 ;
        RECT 450.500 1600.310 451.960 1600.450 ;
        RECT 450.500 1580.050 450.640 1600.310 ;
        RECT 451.680 1600.000 451.960 1600.310 ;
        RECT 449.120 1579.910 450.640 1580.050 ;
        RECT 449.120 26.510 449.260 1579.910 ;
        RECT 294.040 26.190 294.300 26.510 ;
        RECT 449.060 26.190 449.320 26.510 ;
        RECT 294.100 2.400 294.240 26.190 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.010 1588.380 317.330 1588.440 ;
        RECT 458.230 1588.380 458.550 1588.440 ;
        RECT 317.010 1588.240 458.550 1588.380 ;
        RECT 317.010 1588.180 317.330 1588.240 ;
        RECT 458.230 1588.180 458.550 1588.240 ;
        RECT 311.950 15.540 312.270 15.600 ;
        RECT 317.010 15.540 317.330 15.600 ;
        RECT 311.950 15.400 317.330 15.540 ;
        RECT 311.950 15.340 312.270 15.400 ;
        RECT 317.010 15.340 317.330 15.400 ;
      LAYER via ;
        RECT 317.040 1588.180 317.300 1588.440 ;
        RECT 458.260 1588.180 458.520 1588.440 ;
        RECT 311.980 15.340 312.240 15.600 ;
        RECT 317.040 15.340 317.300 15.600 ;
      LAYER met2 ;
        RECT 458.120 1600.380 458.400 1604.000 ;
        RECT 458.120 1600.000 458.460 1600.380 ;
        RECT 458.320 1588.470 458.460 1600.000 ;
        RECT 317.040 1588.150 317.300 1588.470 ;
        RECT 458.260 1588.150 458.520 1588.470 ;
        RECT 317.100 15.630 317.240 1588.150 ;
        RECT 311.980 15.310 312.240 15.630 ;
        RECT 317.040 15.310 317.300 15.630 ;
        RECT 312.040 2.400 312.180 15.310 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 352.045 1586.525 352.215 1588.055 ;
        RECT 423.345 1587.885 423.515 1590.095 ;
      LAYER mcon ;
        RECT 423.345 1589.925 423.515 1590.095 ;
        RECT 352.045 1587.885 352.215 1588.055 ;
      LAYER met1 ;
        RECT 423.285 1590.080 423.575 1590.125 ;
        RECT 464.210 1590.080 464.530 1590.140 ;
        RECT 423.285 1589.940 464.530 1590.080 ;
        RECT 423.285 1589.895 423.575 1589.940 ;
        RECT 464.210 1589.880 464.530 1589.940 ;
        RECT 351.985 1588.040 352.275 1588.085 ;
        RECT 423.285 1588.040 423.575 1588.085 ;
        RECT 351.985 1587.900 423.575 1588.040 ;
        RECT 351.985 1587.855 352.275 1587.900 ;
        RECT 423.285 1587.855 423.575 1587.900 ;
        RECT 341.390 1587.360 341.710 1587.420 ;
        RECT 341.390 1587.220 348.060 1587.360 ;
        RECT 341.390 1587.160 341.710 1587.220 ;
        RECT 347.920 1586.680 348.060 1587.220 ;
        RECT 351.985 1586.680 352.275 1586.725 ;
        RECT 347.920 1586.540 352.275 1586.680 ;
        RECT 351.985 1586.495 352.275 1586.540 ;
        RECT 329.890 14.180 330.210 14.240 ;
        RECT 340.930 14.180 341.250 14.240 ;
        RECT 329.890 14.040 341.250 14.180 ;
        RECT 329.890 13.980 330.210 14.040 ;
        RECT 340.930 13.980 341.250 14.040 ;
      LAYER via ;
        RECT 464.240 1589.880 464.500 1590.140 ;
        RECT 341.420 1587.160 341.680 1587.420 ;
        RECT 329.920 13.980 330.180 14.240 ;
        RECT 340.960 13.980 341.220 14.240 ;
      LAYER met2 ;
        RECT 464.100 1600.380 464.380 1604.000 ;
        RECT 464.100 1600.000 464.440 1600.380 ;
        RECT 464.300 1590.170 464.440 1600.000 ;
        RECT 464.240 1589.850 464.500 1590.170 ;
        RECT 341.420 1587.130 341.680 1587.450 ;
        RECT 341.480 14.690 341.620 1587.130 ;
        RECT 341.020 14.550 341.620 14.690 ;
        RECT 341.020 14.270 341.160 14.550 ;
        RECT 329.920 13.950 330.180 14.270 ;
        RECT 340.960 13.950 341.220 14.270 ;
        RECT 329.980 2.400 330.120 13.950 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 470.265 1539.265 470.435 1587.035 ;
        RECT 470.265 1490.645 470.435 1538.755 ;
        RECT 470.265 1159.145 470.435 1224.935 ;
        RECT 470.265 966.025 470.435 1014.135 ;
        RECT 470.265 734.825 470.435 783.275 ;
        RECT 470.265 476.085 470.435 524.195 ;
        RECT 470.265 404.685 470.435 427.635 ;
        RECT 470.725 324.445 470.895 372.555 ;
        RECT 470.725 253.045 470.895 300.135 ;
        RECT 471.185 14.365 471.355 48.195 ;
      LAYER mcon ;
        RECT 470.265 1586.865 470.435 1587.035 ;
        RECT 470.265 1538.585 470.435 1538.755 ;
        RECT 470.265 1224.765 470.435 1224.935 ;
        RECT 470.265 1013.965 470.435 1014.135 ;
        RECT 470.265 783.105 470.435 783.275 ;
        RECT 470.265 524.025 470.435 524.195 ;
        RECT 470.265 427.465 470.435 427.635 ;
        RECT 470.725 372.385 470.895 372.555 ;
        RECT 470.725 299.965 470.895 300.135 ;
        RECT 471.185 48.025 471.355 48.195 ;
      LAYER met1 ;
        RECT 470.190 1587.020 470.510 1587.080 ;
        RECT 469.995 1586.880 470.510 1587.020 ;
        RECT 470.190 1586.820 470.510 1586.880 ;
        RECT 470.190 1539.420 470.510 1539.480 ;
        RECT 469.995 1539.280 470.510 1539.420 ;
        RECT 470.190 1539.220 470.510 1539.280 ;
        RECT 470.190 1538.740 470.510 1538.800 ;
        RECT 469.995 1538.600 470.510 1538.740 ;
        RECT 470.190 1538.540 470.510 1538.600 ;
        RECT 470.190 1490.800 470.510 1490.860 ;
        RECT 469.995 1490.660 470.510 1490.800 ;
        RECT 470.190 1490.600 470.510 1490.660 ;
        RECT 470.190 1442.180 470.510 1442.240 ;
        RECT 470.650 1442.180 470.970 1442.240 ;
        RECT 470.190 1442.040 470.970 1442.180 ;
        RECT 470.190 1441.980 470.510 1442.040 ;
        RECT 470.650 1441.980 470.970 1442.040 ;
        RECT 470.650 1387.100 470.970 1387.160 ;
        RECT 471.570 1387.100 471.890 1387.160 ;
        RECT 470.650 1386.960 471.890 1387.100 ;
        RECT 470.650 1386.900 470.970 1386.960 ;
        RECT 471.570 1386.900 471.890 1386.960 ;
        RECT 470.190 1256.200 470.510 1256.260 ;
        RECT 470.650 1256.200 470.970 1256.260 ;
        RECT 470.190 1256.060 470.970 1256.200 ;
        RECT 470.190 1256.000 470.510 1256.060 ;
        RECT 470.650 1256.000 470.970 1256.060 ;
        RECT 470.205 1224.920 470.495 1224.965 ;
        RECT 470.650 1224.920 470.970 1224.980 ;
        RECT 470.205 1224.780 470.970 1224.920 ;
        RECT 470.205 1224.735 470.495 1224.780 ;
        RECT 470.650 1224.720 470.970 1224.780 ;
        RECT 470.205 1159.300 470.495 1159.345 ;
        RECT 470.650 1159.300 470.970 1159.360 ;
        RECT 470.205 1159.160 470.970 1159.300 ;
        RECT 470.205 1159.115 470.495 1159.160 ;
        RECT 470.650 1159.100 470.970 1159.160 ;
        RECT 470.650 1125.300 470.970 1125.360 ;
        RECT 470.280 1125.160 470.970 1125.300 ;
        RECT 470.280 1124.680 470.420 1125.160 ;
        RECT 470.650 1125.100 470.970 1125.160 ;
        RECT 470.190 1124.420 470.510 1124.680 ;
        RECT 470.650 1062.740 470.970 1062.800 ;
        RECT 471.570 1062.740 471.890 1062.800 ;
        RECT 470.650 1062.600 471.890 1062.740 ;
        RECT 470.650 1062.540 470.970 1062.600 ;
        RECT 471.570 1062.540 471.890 1062.600 ;
        RECT 470.650 1028.740 470.970 1028.800 ;
        RECT 470.280 1028.600 470.970 1028.740 ;
        RECT 470.280 1028.120 470.420 1028.600 ;
        RECT 470.650 1028.540 470.970 1028.600 ;
        RECT 470.190 1027.860 470.510 1028.120 ;
        RECT 470.190 1014.120 470.510 1014.180 ;
        RECT 469.995 1013.980 470.510 1014.120 ;
        RECT 470.190 1013.920 470.510 1013.980 ;
        RECT 470.205 966.180 470.495 966.225 ;
        RECT 470.650 966.180 470.970 966.240 ;
        RECT 470.205 966.040 470.970 966.180 ;
        RECT 470.205 965.995 470.495 966.040 ;
        RECT 470.650 965.980 470.970 966.040 ;
        RECT 470.650 869.620 470.970 869.680 ;
        RECT 471.110 869.620 471.430 869.680 ;
        RECT 470.650 869.480 471.430 869.620 ;
        RECT 470.650 869.420 470.970 869.480 ;
        RECT 471.110 869.420 471.430 869.480 ;
        RECT 470.650 862.480 470.970 862.540 ;
        RECT 471.570 862.480 471.890 862.540 ;
        RECT 470.650 862.340 471.890 862.480 ;
        RECT 470.650 862.280 470.970 862.340 ;
        RECT 471.570 862.280 471.890 862.340 ;
        RECT 470.205 783.260 470.495 783.305 ;
        RECT 470.650 783.260 470.970 783.320 ;
        RECT 470.205 783.120 470.970 783.260 ;
        RECT 470.205 783.075 470.495 783.120 ;
        RECT 470.650 783.060 470.970 783.120 ;
        RECT 470.205 734.980 470.495 735.025 ;
        RECT 471.570 734.980 471.890 735.040 ;
        RECT 470.205 734.840 471.890 734.980 ;
        RECT 470.205 734.795 470.495 734.840 ;
        RECT 471.570 734.780 471.890 734.840 ;
        RECT 470.190 591.980 470.510 592.240 ;
        RECT 470.280 591.840 470.420 591.980 ;
        RECT 470.650 591.840 470.970 591.900 ;
        RECT 470.280 591.700 470.970 591.840 ;
        RECT 470.650 591.640 470.970 591.700 ;
        RECT 470.190 524.180 470.510 524.240 ;
        RECT 469.995 524.040 470.510 524.180 ;
        RECT 470.190 523.980 470.510 524.040 ;
        RECT 470.190 476.240 470.510 476.300 ;
        RECT 469.995 476.100 470.510 476.240 ;
        RECT 470.190 476.040 470.510 476.100 ;
        RECT 470.190 427.620 470.510 427.680 ;
        RECT 469.995 427.480 470.510 427.620 ;
        RECT 470.190 427.420 470.510 427.480 ;
        RECT 470.205 404.840 470.495 404.885 ;
        RECT 471.570 404.840 471.890 404.900 ;
        RECT 470.205 404.700 471.890 404.840 ;
        RECT 470.205 404.655 470.495 404.700 ;
        RECT 471.570 404.640 471.890 404.700 ;
        RECT 470.665 372.540 470.955 372.585 ;
        RECT 471.570 372.540 471.890 372.600 ;
        RECT 470.665 372.400 471.890 372.540 ;
        RECT 470.665 372.355 470.955 372.400 ;
        RECT 471.570 372.340 471.890 372.400 ;
        RECT 470.650 324.600 470.970 324.660 ;
        RECT 470.455 324.460 470.970 324.600 ;
        RECT 470.650 324.400 470.970 324.460 ;
        RECT 470.650 300.120 470.970 300.180 ;
        RECT 470.455 299.980 470.970 300.120 ;
        RECT 470.650 299.920 470.970 299.980 ;
        RECT 470.650 253.200 470.970 253.260 ;
        RECT 470.455 253.060 470.970 253.200 ;
        RECT 470.650 253.000 470.970 253.060 ;
        RECT 470.650 158.820 470.970 159.080 ;
        RECT 470.740 158.060 470.880 158.820 ;
        RECT 470.650 157.800 470.970 158.060 ;
        RECT 470.650 62.260 470.970 62.520 ;
        RECT 470.740 61.780 470.880 62.260 ;
        RECT 471.110 61.780 471.430 61.840 ;
        RECT 470.740 61.640 471.430 61.780 ;
        RECT 471.110 61.580 471.430 61.640 ;
        RECT 471.110 48.180 471.430 48.240 ;
        RECT 470.915 48.040 471.430 48.180 ;
        RECT 471.110 47.980 471.430 48.040 ;
        RECT 347.370 14.520 347.690 14.580 ;
        RECT 471.125 14.520 471.415 14.565 ;
        RECT 347.370 14.380 471.415 14.520 ;
        RECT 347.370 14.320 347.690 14.380 ;
        RECT 471.125 14.335 471.415 14.380 ;
      LAYER via ;
        RECT 470.220 1586.820 470.480 1587.080 ;
        RECT 470.220 1539.220 470.480 1539.480 ;
        RECT 470.220 1538.540 470.480 1538.800 ;
        RECT 470.220 1490.600 470.480 1490.860 ;
        RECT 470.220 1441.980 470.480 1442.240 ;
        RECT 470.680 1441.980 470.940 1442.240 ;
        RECT 470.680 1386.900 470.940 1387.160 ;
        RECT 471.600 1386.900 471.860 1387.160 ;
        RECT 470.220 1256.000 470.480 1256.260 ;
        RECT 470.680 1256.000 470.940 1256.260 ;
        RECT 470.680 1224.720 470.940 1224.980 ;
        RECT 470.680 1159.100 470.940 1159.360 ;
        RECT 470.680 1125.100 470.940 1125.360 ;
        RECT 470.220 1124.420 470.480 1124.680 ;
        RECT 470.680 1062.540 470.940 1062.800 ;
        RECT 471.600 1062.540 471.860 1062.800 ;
        RECT 470.680 1028.540 470.940 1028.800 ;
        RECT 470.220 1027.860 470.480 1028.120 ;
        RECT 470.220 1013.920 470.480 1014.180 ;
        RECT 470.680 965.980 470.940 966.240 ;
        RECT 470.680 869.420 470.940 869.680 ;
        RECT 471.140 869.420 471.400 869.680 ;
        RECT 470.680 862.280 470.940 862.540 ;
        RECT 471.600 862.280 471.860 862.540 ;
        RECT 470.680 783.060 470.940 783.320 ;
        RECT 471.600 734.780 471.860 735.040 ;
        RECT 470.220 591.980 470.480 592.240 ;
        RECT 470.680 591.640 470.940 591.900 ;
        RECT 470.220 523.980 470.480 524.240 ;
        RECT 470.220 476.040 470.480 476.300 ;
        RECT 470.220 427.420 470.480 427.680 ;
        RECT 471.600 404.640 471.860 404.900 ;
        RECT 471.600 372.340 471.860 372.600 ;
        RECT 470.680 324.400 470.940 324.660 ;
        RECT 470.680 299.920 470.940 300.180 ;
        RECT 470.680 253.000 470.940 253.260 ;
        RECT 470.680 158.820 470.940 159.080 ;
        RECT 470.680 157.800 470.940 158.060 ;
        RECT 470.680 62.260 470.940 62.520 ;
        RECT 471.140 61.580 471.400 61.840 ;
        RECT 471.140 47.980 471.400 48.240 ;
        RECT 347.400 14.320 347.660 14.580 ;
      LAYER met2 ;
        RECT 470.080 1600.380 470.360 1604.000 ;
        RECT 470.080 1600.000 470.420 1600.380 ;
        RECT 470.280 1587.110 470.420 1600.000 ;
        RECT 470.220 1586.790 470.480 1587.110 ;
        RECT 470.220 1539.190 470.480 1539.510 ;
        RECT 470.280 1538.830 470.420 1539.190 ;
        RECT 470.220 1538.510 470.480 1538.830 ;
        RECT 470.220 1490.570 470.480 1490.890 ;
        RECT 470.280 1442.270 470.420 1490.570 ;
        RECT 470.220 1441.950 470.480 1442.270 ;
        RECT 470.680 1441.950 470.940 1442.270 ;
        RECT 470.740 1435.325 470.880 1441.950 ;
        RECT 470.670 1434.955 470.950 1435.325 ;
        RECT 471.590 1434.955 471.870 1435.325 ;
        RECT 471.660 1387.190 471.800 1434.955 ;
        RECT 470.680 1386.870 470.940 1387.190 ;
        RECT 471.600 1386.870 471.860 1387.190 ;
        RECT 470.740 1328.450 470.880 1386.870 ;
        RECT 470.280 1328.310 470.880 1328.450 ;
        RECT 470.280 1256.290 470.420 1328.310 ;
        RECT 470.220 1255.970 470.480 1256.290 ;
        RECT 470.680 1255.970 470.940 1256.290 ;
        RECT 470.740 1225.010 470.880 1255.970 ;
        RECT 470.680 1224.690 470.940 1225.010 ;
        RECT 470.680 1159.070 470.940 1159.390 ;
        RECT 470.740 1125.390 470.880 1159.070 ;
        RECT 470.680 1125.070 470.940 1125.390 ;
        RECT 470.220 1124.390 470.480 1124.710 ;
        RECT 470.280 1110.965 470.420 1124.390 ;
        RECT 470.210 1110.595 470.490 1110.965 ;
        RECT 471.590 1110.595 471.870 1110.965 ;
        RECT 471.660 1062.830 471.800 1110.595 ;
        RECT 470.680 1062.510 470.940 1062.830 ;
        RECT 471.600 1062.510 471.860 1062.830 ;
        RECT 470.740 1028.830 470.880 1062.510 ;
        RECT 470.680 1028.510 470.940 1028.830 ;
        RECT 470.220 1027.830 470.480 1028.150 ;
        RECT 470.280 1014.210 470.420 1027.830 ;
        RECT 470.220 1013.890 470.480 1014.210 ;
        RECT 470.680 965.950 470.940 966.270 ;
        RECT 470.740 942.210 470.880 965.950 ;
        RECT 470.740 942.070 471.340 942.210 ;
        RECT 471.200 869.710 471.340 942.070 ;
        RECT 470.680 869.390 470.940 869.710 ;
        RECT 471.140 869.390 471.400 869.710 ;
        RECT 470.740 862.570 470.880 869.390 ;
        RECT 470.680 862.250 470.940 862.570 ;
        RECT 471.600 862.250 471.860 862.570 ;
        RECT 471.660 814.485 471.800 862.250 ;
        RECT 470.670 814.115 470.950 814.485 ;
        RECT 471.590 814.115 471.870 814.485 ;
        RECT 470.740 783.350 470.880 814.115 ;
        RECT 470.680 783.030 470.940 783.350 ;
        RECT 471.600 734.750 471.860 735.070 ;
        RECT 471.660 669.645 471.800 734.750 ;
        RECT 470.670 669.275 470.950 669.645 ;
        RECT 471.590 669.275 471.870 669.645 ;
        RECT 470.740 628.050 470.880 669.275 ;
        RECT 470.280 627.910 470.880 628.050 ;
        RECT 470.280 592.270 470.420 627.910 ;
        RECT 470.220 591.950 470.480 592.270 ;
        RECT 470.680 591.610 470.940 591.930 ;
        RECT 470.740 532.965 470.880 591.610 ;
        RECT 470.670 532.595 470.950 532.965 ;
        RECT 470.210 531.235 470.490 531.605 ;
        RECT 470.280 524.270 470.420 531.235 ;
        RECT 470.220 523.950 470.480 524.270 ;
        RECT 470.220 476.010 470.480 476.330 ;
        RECT 470.280 435.725 470.420 476.010 ;
        RECT 470.210 435.355 470.490 435.725 ;
        RECT 470.210 434.675 470.490 435.045 ;
        RECT 470.280 427.710 470.420 434.675 ;
        RECT 470.220 427.390 470.480 427.710 ;
        RECT 471.600 404.610 471.860 404.930 ;
        RECT 471.660 372.630 471.800 404.610 ;
        RECT 471.600 372.310 471.860 372.630 ;
        RECT 470.680 324.370 470.940 324.690 ;
        RECT 470.740 300.210 470.880 324.370 ;
        RECT 470.680 299.890 470.940 300.210 ;
        RECT 470.680 252.970 470.940 253.290 ;
        RECT 470.740 159.110 470.880 252.970 ;
        RECT 470.680 158.790 470.940 159.110 ;
        RECT 470.680 157.770 470.940 158.090 ;
        RECT 470.740 110.570 470.880 157.770 ;
        RECT 470.280 110.430 470.880 110.570 ;
        RECT 470.280 96.970 470.420 110.430 ;
        RECT 470.280 96.830 470.880 96.970 ;
        RECT 470.740 62.550 470.880 96.830 ;
        RECT 470.680 62.230 470.940 62.550 ;
        RECT 471.140 61.550 471.400 61.870 ;
        RECT 471.200 48.270 471.340 61.550 ;
        RECT 471.140 47.950 471.400 48.270 ;
        RECT 347.400 14.290 347.660 14.610 ;
        RECT 347.460 2.400 347.600 14.290 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 470.670 1435.000 470.950 1435.280 ;
        RECT 471.590 1435.000 471.870 1435.280 ;
        RECT 470.210 1110.640 470.490 1110.920 ;
        RECT 471.590 1110.640 471.870 1110.920 ;
        RECT 470.670 814.160 470.950 814.440 ;
        RECT 471.590 814.160 471.870 814.440 ;
        RECT 470.670 669.320 470.950 669.600 ;
        RECT 471.590 669.320 471.870 669.600 ;
        RECT 470.670 532.640 470.950 532.920 ;
        RECT 470.210 531.280 470.490 531.560 ;
        RECT 470.210 435.400 470.490 435.680 ;
        RECT 470.210 434.720 470.490 435.000 ;
      LAYER met3 ;
        RECT 470.645 1435.290 470.975 1435.305 ;
        RECT 471.565 1435.290 471.895 1435.305 ;
        RECT 470.645 1434.990 471.895 1435.290 ;
        RECT 470.645 1434.975 470.975 1434.990 ;
        RECT 471.565 1434.975 471.895 1434.990 ;
        RECT 470.185 1110.930 470.515 1110.945 ;
        RECT 471.565 1110.930 471.895 1110.945 ;
        RECT 470.185 1110.630 471.895 1110.930 ;
        RECT 470.185 1110.615 470.515 1110.630 ;
        RECT 471.565 1110.615 471.895 1110.630 ;
        RECT 470.645 814.450 470.975 814.465 ;
        RECT 471.565 814.450 471.895 814.465 ;
        RECT 470.645 814.150 471.895 814.450 ;
        RECT 470.645 814.135 470.975 814.150 ;
        RECT 471.565 814.135 471.895 814.150 ;
        RECT 470.645 669.610 470.975 669.625 ;
        RECT 471.565 669.610 471.895 669.625 ;
        RECT 470.645 669.310 471.895 669.610 ;
        RECT 470.645 669.295 470.975 669.310 ;
        RECT 471.565 669.295 471.895 669.310 ;
        RECT 470.645 532.930 470.975 532.945 ;
        RECT 469.510 532.630 470.975 532.930 ;
        RECT 469.510 531.570 469.810 532.630 ;
        RECT 470.645 532.615 470.975 532.630 ;
        RECT 470.185 531.570 470.515 531.585 ;
        RECT 469.510 531.270 470.515 531.570 ;
        RECT 470.185 531.255 470.515 531.270 ;
        RECT 470.185 435.690 470.515 435.705 ;
        RECT 470.185 435.375 470.730 435.690 ;
        RECT 470.430 435.025 470.730 435.375 ;
        RECT 470.185 434.710 470.730 435.025 ;
        RECT 470.185 434.695 470.515 434.710 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 17.580 365.630 17.640 ;
        RECT 476.630 17.580 476.950 17.640 ;
        RECT 365.310 17.440 476.950 17.580 ;
        RECT 365.310 17.380 365.630 17.440 ;
        RECT 476.630 17.380 476.950 17.440 ;
      LAYER via ;
        RECT 365.340 17.380 365.600 17.640 ;
        RECT 476.660 17.380 476.920 17.640 ;
      LAYER met2 ;
        RECT 476.520 1600.380 476.800 1604.000 ;
        RECT 476.520 1600.000 476.860 1600.380 ;
        RECT 476.720 17.670 476.860 1600.000 ;
        RECT 365.340 17.350 365.600 17.670 ;
        RECT 476.660 17.350 476.920 17.670 ;
        RECT 365.400 2.400 365.540 17.350 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 412.305 16.745 412.475 19.295 ;
      LAYER mcon ;
        RECT 412.305 19.125 412.475 19.295 ;
      LAYER met1 ;
        RECT 478.470 1173.240 478.790 1173.300 ;
        RECT 478.100 1173.100 478.790 1173.240 ;
        RECT 478.100 1172.960 478.240 1173.100 ;
        RECT 478.470 1173.040 478.790 1173.100 ;
        RECT 478.010 1172.700 478.330 1172.960 ;
        RECT 478.470 1076.680 478.790 1076.740 ;
        RECT 478.100 1076.540 478.790 1076.680 ;
        RECT 478.100 1076.400 478.240 1076.540 ;
        RECT 478.470 1076.480 478.790 1076.540 ;
        RECT 478.010 1076.140 478.330 1076.400 ;
        RECT 478.470 980.120 478.790 980.180 ;
        RECT 478.100 979.980 478.790 980.120 ;
        RECT 478.100 979.840 478.240 979.980 ;
        RECT 478.470 979.920 478.790 979.980 ;
        RECT 478.010 979.580 478.330 979.840 ;
        RECT 477.550 883.560 477.870 883.620 ;
        RECT 477.550 883.420 478.240 883.560 ;
        RECT 477.550 883.360 477.870 883.420 ;
        RECT 478.100 883.280 478.240 883.420 ;
        RECT 478.010 883.020 478.330 883.280 ;
        RECT 478.010 593.680 478.330 593.940 ;
        RECT 478.100 593.260 478.240 593.680 ;
        RECT 478.010 593.000 478.330 593.260 ;
        RECT 412.245 19.280 412.535 19.325 ;
        RECT 478.470 19.280 478.790 19.340 ;
        RECT 412.245 19.140 478.790 19.280 ;
        RECT 412.245 19.095 412.535 19.140 ;
        RECT 478.470 19.080 478.790 19.140 ;
        RECT 383.250 17.240 383.570 17.300 ;
        RECT 383.250 17.100 399.580 17.240 ;
        RECT 383.250 17.040 383.570 17.100 ;
        RECT 399.440 16.900 399.580 17.100 ;
        RECT 412.245 16.900 412.535 16.945 ;
        RECT 399.440 16.760 412.535 16.900 ;
        RECT 412.245 16.715 412.535 16.760 ;
      LAYER via ;
        RECT 478.500 1173.040 478.760 1173.300 ;
        RECT 478.040 1172.700 478.300 1172.960 ;
        RECT 478.500 1076.480 478.760 1076.740 ;
        RECT 478.040 1076.140 478.300 1076.400 ;
        RECT 478.500 979.920 478.760 980.180 ;
        RECT 478.040 979.580 478.300 979.840 ;
        RECT 477.580 883.360 477.840 883.620 ;
        RECT 478.040 883.020 478.300 883.280 ;
        RECT 478.040 593.680 478.300 593.940 ;
        RECT 478.040 593.000 478.300 593.260 ;
        RECT 478.500 19.080 478.760 19.340 ;
        RECT 383.280 17.040 383.540 17.300 ;
      LAYER met2 ;
        RECT 482.500 1600.450 482.780 1604.000 ;
        RECT 481.320 1600.310 482.780 1600.450 ;
        RECT 481.320 1580.050 481.460 1600.310 ;
        RECT 482.500 1600.000 482.780 1600.310 ;
        RECT 478.100 1579.910 481.460 1580.050 ;
        RECT 478.100 1511.370 478.240 1579.910 ;
        RECT 477.640 1511.230 478.240 1511.370 ;
        RECT 477.640 1510.690 477.780 1511.230 ;
        RECT 477.640 1510.550 478.700 1510.690 ;
        RECT 478.560 1366.530 478.700 1510.550 ;
        RECT 477.640 1366.390 478.700 1366.530 ;
        RECT 477.640 1365.850 477.780 1366.390 ;
        RECT 477.640 1365.710 478.240 1365.850 ;
        RECT 478.100 1207.410 478.240 1365.710 ;
        RECT 478.100 1207.270 478.700 1207.410 ;
        RECT 478.560 1173.330 478.700 1207.270 ;
        RECT 478.500 1173.010 478.760 1173.330 ;
        RECT 478.040 1172.670 478.300 1172.990 ;
        RECT 478.100 1110.850 478.240 1172.670 ;
        RECT 478.100 1110.710 478.700 1110.850 ;
        RECT 478.560 1076.770 478.700 1110.710 ;
        RECT 478.500 1076.450 478.760 1076.770 ;
        RECT 478.040 1076.110 478.300 1076.430 ;
        RECT 478.100 1014.290 478.240 1076.110 ;
        RECT 478.100 1014.150 478.700 1014.290 ;
        RECT 478.560 980.210 478.700 1014.150 ;
        RECT 478.500 979.890 478.760 980.210 ;
        RECT 478.040 979.550 478.300 979.870 ;
        RECT 478.100 917.730 478.240 979.550 ;
        RECT 477.640 917.590 478.240 917.730 ;
        RECT 477.640 883.650 477.780 917.590 ;
        RECT 477.580 883.330 477.840 883.650 ;
        RECT 478.040 882.990 478.300 883.310 ;
        RECT 478.100 787.170 478.240 882.990 ;
        RECT 477.640 787.030 478.240 787.170 ;
        RECT 477.640 786.490 477.780 787.030 ;
        RECT 477.640 786.350 478.240 786.490 ;
        RECT 478.100 690.610 478.240 786.350 ;
        RECT 477.640 690.470 478.240 690.610 ;
        RECT 477.640 689.250 477.780 690.470 ;
        RECT 477.640 689.110 478.240 689.250 ;
        RECT 478.100 593.970 478.240 689.110 ;
        RECT 478.040 593.650 478.300 593.970 ;
        RECT 478.040 592.970 478.300 593.290 ;
        RECT 478.100 314.570 478.240 592.970 ;
        RECT 477.640 314.430 478.240 314.570 ;
        RECT 477.640 313.210 477.780 314.430 ;
        RECT 477.640 313.070 478.240 313.210 ;
        RECT 478.100 207.130 478.240 313.070 ;
        RECT 477.640 206.990 478.240 207.130 ;
        RECT 477.640 206.450 477.780 206.990 ;
        RECT 477.640 206.310 478.240 206.450 ;
        RECT 478.100 109.890 478.240 206.310 ;
        RECT 478.100 109.750 478.700 109.890 ;
        RECT 478.560 19.370 478.700 109.750 ;
        RECT 478.500 19.050 478.760 19.370 ;
        RECT 383.280 17.010 383.540 17.330 ;
        RECT 383.340 2.400 383.480 17.010 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 446.345 15.725 446.515 19.975 ;
      LAYER mcon ;
        RECT 446.345 19.805 446.515 19.975 ;
      LAYER met1 ;
        RECT 483.070 1579.880 483.390 1579.940 ;
        RECT 487.670 1579.880 487.990 1579.940 ;
        RECT 483.070 1579.740 487.990 1579.880 ;
        RECT 483.070 1579.680 483.390 1579.740 ;
        RECT 487.670 1579.680 487.990 1579.740 ;
        RECT 446.285 19.960 446.575 20.005 ;
        RECT 483.070 19.960 483.390 20.020 ;
        RECT 446.285 19.820 483.390 19.960 ;
        RECT 446.285 19.775 446.575 19.820 ;
        RECT 483.070 19.760 483.390 19.820 ;
        RECT 401.190 15.880 401.510 15.940 ;
        RECT 446.285 15.880 446.575 15.925 ;
        RECT 401.190 15.740 446.575 15.880 ;
        RECT 401.190 15.680 401.510 15.740 ;
        RECT 446.285 15.695 446.575 15.740 ;
      LAYER via ;
        RECT 483.100 1579.680 483.360 1579.940 ;
        RECT 487.700 1579.680 487.960 1579.940 ;
        RECT 483.100 19.760 483.360 20.020 ;
        RECT 401.220 15.680 401.480 15.940 ;
      LAYER met2 ;
        RECT 488.940 1600.450 489.220 1604.000 ;
        RECT 487.760 1600.310 489.220 1600.450 ;
        RECT 487.760 1579.970 487.900 1600.310 ;
        RECT 488.940 1600.000 489.220 1600.310 ;
        RECT 483.100 1579.650 483.360 1579.970 ;
        RECT 487.700 1579.650 487.960 1579.970 ;
        RECT 483.160 20.050 483.300 1579.650 ;
        RECT 483.100 19.730 483.360 20.050 ;
        RECT 401.220 15.650 401.480 15.970 ;
        RECT 401.280 2.400 401.420 15.650 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.770 1579.880 366.090 1579.940 ;
        RECT 369.910 1579.880 370.230 1579.940 ;
        RECT 365.770 1579.740 370.230 1579.880 ;
        RECT 365.770 1579.680 366.090 1579.740 ;
        RECT 369.910 1579.680 370.230 1579.740 ;
        RECT 365.770 18.940 366.090 19.000 ;
        RECT 352.980 18.800 366.090 18.940 ;
        RECT 62.170 18.600 62.490 18.660 ;
        RECT 352.980 18.600 353.120 18.800 ;
        RECT 365.770 18.740 366.090 18.800 ;
        RECT 62.170 18.460 353.120 18.600 ;
        RECT 62.170 18.400 62.490 18.460 ;
      LAYER via ;
        RECT 365.800 1579.680 366.060 1579.940 ;
        RECT 369.940 1579.680 370.200 1579.940 ;
        RECT 62.200 18.400 62.460 18.660 ;
        RECT 365.800 18.740 366.060 19.000 ;
      LAYER met2 ;
        RECT 371.180 1600.450 371.460 1604.000 ;
        RECT 370.000 1600.310 371.460 1600.450 ;
        RECT 370.000 1579.970 370.140 1600.310 ;
        RECT 371.180 1600.000 371.460 1600.310 ;
        RECT 365.800 1579.650 366.060 1579.970 ;
        RECT 369.940 1579.650 370.200 1579.970 ;
        RECT 365.860 19.030 366.000 1579.650 ;
        RECT 365.800 18.710 366.060 19.030 ;
        RECT 62.200 18.370 62.460 18.690 ;
        RECT 62.260 2.400 62.400 18.370 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 445.885 16.065 446.055 20.315 ;
        RECT 457.845 16.745 458.015 20.315 ;
      LAYER mcon ;
        RECT 445.885 20.145 446.055 20.315 ;
        RECT 457.845 20.145 458.015 20.315 ;
      LAYER met1 ;
        RECT 445.825 20.300 446.115 20.345 ;
        RECT 457.785 20.300 458.075 20.345 ;
        RECT 445.825 20.160 458.075 20.300 ;
        RECT 445.825 20.115 446.115 20.160 ;
        RECT 457.785 20.115 458.075 20.160 ;
        RECT 457.785 16.900 458.075 16.945 ;
        RECT 491.350 16.900 491.670 16.960 ;
        RECT 457.785 16.760 491.670 16.900 ;
        RECT 457.785 16.715 458.075 16.760 ;
        RECT 491.350 16.700 491.670 16.760 ;
        RECT 419.130 16.220 419.450 16.280 ;
        RECT 445.825 16.220 446.115 16.265 ;
        RECT 419.130 16.080 446.115 16.220 ;
        RECT 419.130 16.020 419.450 16.080 ;
        RECT 445.825 16.035 446.115 16.080 ;
      LAYER via ;
        RECT 491.380 16.700 491.640 16.960 ;
        RECT 419.160 16.020 419.420 16.280 ;
      LAYER met2 ;
        RECT 494.920 1600.450 495.200 1604.000 ;
        RECT 494.200 1600.310 495.200 1600.450 ;
        RECT 494.200 1580.050 494.340 1600.310 ;
        RECT 494.920 1600.000 495.200 1600.310 ;
        RECT 490.520 1579.910 494.340 1580.050 ;
        RECT 490.520 19.450 490.660 1579.910 ;
        RECT 490.520 19.310 491.580 19.450 ;
        RECT 491.440 16.990 491.580 19.310 ;
        RECT 491.380 16.670 491.640 16.990 ;
        RECT 419.160 15.990 419.420 16.310 ;
        RECT 419.220 2.400 419.360 15.990 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 501.470 1591.100 501.790 1591.160 ;
        RECT 472.580 1590.960 501.790 1591.100 ;
        RECT 441.210 1590.760 441.530 1590.820 ;
        RECT 472.580 1590.760 472.720 1590.960 ;
        RECT 501.470 1590.900 501.790 1590.960 ;
        RECT 441.210 1590.620 472.720 1590.760 ;
        RECT 441.210 1590.560 441.530 1590.620 ;
        RECT 436.610 20.640 436.930 20.700 ;
        RECT 441.210 20.640 441.530 20.700 ;
        RECT 436.610 20.500 441.530 20.640 ;
        RECT 436.610 20.440 436.930 20.500 ;
        RECT 441.210 20.440 441.530 20.500 ;
      LAYER via ;
        RECT 441.240 1590.560 441.500 1590.820 ;
        RECT 501.500 1590.900 501.760 1591.160 ;
        RECT 436.640 20.440 436.900 20.700 ;
        RECT 441.240 20.440 441.500 20.700 ;
      LAYER met2 ;
        RECT 501.360 1600.380 501.640 1604.000 ;
        RECT 501.360 1600.000 501.700 1600.380 ;
        RECT 501.560 1591.190 501.700 1600.000 ;
        RECT 501.500 1590.870 501.760 1591.190 ;
        RECT 441.240 1590.530 441.500 1590.850 ;
        RECT 441.300 20.730 441.440 1590.530 ;
        RECT 436.640 20.410 436.900 20.730 ;
        RECT 441.240 20.410 441.500 20.730 ;
        RECT 436.700 2.400 436.840 20.410 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 455.085 1062.245 455.255 1103.555 ;
        RECT 455.085 1013.965 455.255 1055.615 ;
        RECT 455.085 904.145 455.255 917.915 ;
        RECT 455.085 855.525 455.255 893.435 ;
        RECT 454.625 524.365 454.795 572.475 ;
        RECT 454.625 276.165 454.795 283.475 ;
        RECT 455.545 89.845 455.715 137.955 ;
      LAYER mcon ;
        RECT 455.085 1103.385 455.255 1103.555 ;
        RECT 455.085 1055.445 455.255 1055.615 ;
        RECT 455.085 917.745 455.255 917.915 ;
        RECT 455.085 893.265 455.255 893.435 ;
        RECT 454.625 572.305 454.795 572.475 ;
        RECT 454.625 283.305 454.795 283.475 ;
        RECT 455.545 137.785 455.715 137.955 ;
      LAYER met1 ;
        RECT 455.010 1593.140 455.330 1593.200 ;
        RECT 507.450 1593.140 507.770 1593.200 ;
        RECT 455.010 1593.000 507.770 1593.140 ;
        RECT 455.010 1592.940 455.330 1593.000 ;
        RECT 507.450 1592.940 507.770 1593.000 ;
        RECT 454.090 1152.500 454.410 1152.560 ;
        RECT 454.550 1152.500 454.870 1152.560 ;
        RECT 454.090 1152.360 454.870 1152.500 ;
        RECT 454.090 1152.300 454.410 1152.360 ;
        RECT 454.550 1152.300 454.870 1152.360 ;
        RECT 453.170 1104.220 453.490 1104.280 ;
        RECT 455.010 1104.220 455.330 1104.280 ;
        RECT 453.170 1104.080 455.330 1104.220 ;
        RECT 453.170 1104.020 453.490 1104.080 ;
        RECT 455.010 1104.020 455.330 1104.080 ;
        RECT 455.010 1103.540 455.330 1103.600 ;
        RECT 454.815 1103.400 455.330 1103.540 ;
        RECT 455.010 1103.340 455.330 1103.400 ;
        RECT 455.025 1062.400 455.315 1062.445 ;
        RECT 455.470 1062.400 455.790 1062.460 ;
        RECT 455.025 1062.260 455.790 1062.400 ;
        RECT 455.025 1062.215 455.315 1062.260 ;
        RECT 455.470 1062.200 455.790 1062.260 ;
        RECT 455.025 1055.600 455.315 1055.645 ;
        RECT 455.930 1055.600 456.250 1055.660 ;
        RECT 455.025 1055.460 456.250 1055.600 ;
        RECT 455.025 1055.415 455.315 1055.460 ;
        RECT 455.930 1055.400 456.250 1055.460 ;
        RECT 455.010 1014.120 455.330 1014.180 ;
        RECT 454.815 1013.980 455.330 1014.120 ;
        RECT 455.010 1013.920 455.330 1013.980 ;
        RECT 455.010 917.900 455.330 917.960 ;
        RECT 454.815 917.760 455.330 917.900 ;
        RECT 455.010 917.700 455.330 917.760 ;
        RECT 455.010 904.300 455.330 904.360 ;
        RECT 454.815 904.160 455.330 904.300 ;
        RECT 455.010 904.100 455.330 904.160 ;
        RECT 455.010 893.420 455.330 893.480 ;
        RECT 454.815 893.280 455.330 893.420 ;
        RECT 455.010 893.220 455.330 893.280 ;
        RECT 455.025 855.680 455.315 855.725 ;
        RECT 455.930 855.680 456.250 855.740 ;
        RECT 455.025 855.540 456.250 855.680 ;
        RECT 455.025 855.495 455.315 855.540 ;
        RECT 455.930 855.480 456.250 855.540 ;
        RECT 455.010 669.700 455.330 669.760 ;
        RECT 455.930 669.700 456.250 669.760 ;
        RECT 455.010 669.560 456.250 669.700 ;
        RECT 455.010 669.500 455.330 669.560 ;
        RECT 455.930 669.500 456.250 669.560 ;
        RECT 455.010 620.740 455.330 620.800 ;
        RECT 455.930 620.740 456.250 620.800 ;
        RECT 455.010 620.600 456.250 620.740 ;
        RECT 455.010 620.540 455.330 620.600 ;
        RECT 455.930 620.540 456.250 620.600 ;
        RECT 454.550 572.460 454.870 572.520 ;
        RECT 454.355 572.320 454.870 572.460 ;
        RECT 454.550 572.260 454.870 572.320 ;
        RECT 454.565 524.520 454.855 524.565 ;
        RECT 455.010 524.520 455.330 524.580 ;
        RECT 454.565 524.380 455.330 524.520 ;
        RECT 454.565 524.335 454.855 524.380 ;
        RECT 455.010 524.320 455.330 524.380 ;
        RECT 455.010 476.240 455.330 476.300 ;
        RECT 455.470 476.240 455.790 476.300 ;
        RECT 455.010 476.100 455.790 476.240 ;
        RECT 455.010 476.040 455.330 476.100 ;
        RECT 455.470 476.040 455.790 476.100 ;
        RECT 455.470 331.740 455.790 331.800 ;
        RECT 455.100 331.600 455.790 331.740 ;
        RECT 455.100 331.460 455.240 331.600 ;
        RECT 455.470 331.540 455.790 331.600 ;
        RECT 455.010 331.200 455.330 331.460 ;
        RECT 454.565 283.460 454.855 283.505 ;
        RECT 455.010 283.460 455.330 283.520 ;
        RECT 454.565 283.320 455.330 283.460 ;
        RECT 454.565 283.275 454.855 283.320 ;
        RECT 455.010 283.260 455.330 283.320 ;
        RECT 454.550 276.320 454.870 276.380 ;
        RECT 454.355 276.180 454.870 276.320 ;
        RECT 454.550 276.120 454.870 276.180 ;
        RECT 454.550 234.840 454.870 234.900 ;
        RECT 455.010 234.840 455.330 234.900 ;
        RECT 454.550 234.700 455.330 234.840 ;
        RECT 454.550 234.640 454.870 234.700 ;
        RECT 455.010 234.640 455.330 234.700 ;
        RECT 455.010 234.160 455.330 234.220 ;
        RECT 455.930 234.160 456.250 234.220 ;
        RECT 455.010 234.020 456.250 234.160 ;
        RECT 455.010 233.960 455.330 234.020 ;
        RECT 455.930 233.960 456.250 234.020 ;
        RECT 455.010 145.080 455.330 145.140 ;
        RECT 455.930 145.080 456.250 145.140 ;
        RECT 455.010 144.940 456.250 145.080 ;
        RECT 455.010 144.880 455.330 144.940 ;
        RECT 455.930 144.880 456.250 144.940 ;
        RECT 455.010 137.940 455.330 138.000 ;
        RECT 455.485 137.940 455.775 137.985 ;
        RECT 455.010 137.800 455.775 137.940 ;
        RECT 455.010 137.740 455.330 137.800 ;
        RECT 455.485 137.755 455.775 137.800 ;
        RECT 455.010 90.000 455.330 90.060 ;
        RECT 455.485 90.000 455.775 90.045 ;
        RECT 455.010 89.860 455.775 90.000 ;
        RECT 455.010 89.800 455.330 89.860 ;
        RECT 455.485 89.815 455.775 89.860 ;
        RECT 455.010 62.460 455.330 62.520 ;
        RECT 454.640 62.320 455.330 62.460 ;
        RECT 454.640 62.180 454.780 62.320 ;
        RECT 455.010 62.260 455.330 62.320 ;
        RECT 454.550 61.920 454.870 62.180 ;
        RECT 454.550 47.980 454.870 48.240 ;
        RECT 454.640 47.560 454.780 47.980 ;
        RECT 454.550 47.300 454.870 47.560 ;
      LAYER via ;
        RECT 455.040 1592.940 455.300 1593.200 ;
        RECT 507.480 1592.940 507.740 1593.200 ;
        RECT 454.120 1152.300 454.380 1152.560 ;
        RECT 454.580 1152.300 454.840 1152.560 ;
        RECT 453.200 1104.020 453.460 1104.280 ;
        RECT 455.040 1104.020 455.300 1104.280 ;
        RECT 455.040 1103.340 455.300 1103.600 ;
        RECT 455.500 1062.200 455.760 1062.460 ;
        RECT 455.960 1055.400 456.220 1055.660 ;
        RECT 455.040 1013.920 455.300 1014.180 ;
        RECT 455.040 917.700 455.300 917.960 ;
        RECT 455.040 904.100 455.300 904.360 ;
        RECT 455.040 893.220 455.300 893.480 ;
        RECT 455.960 855.480 456.220 855.740 ;
        RECT 455.040 669.500 455.300 669.760 ;
        RECT 455.960 669.500 456.220 669.760 ;
        RECT 455.040 620.540 455.300 620.800 ;
        RECT 455.960 620.540 456.220 620.800 ;
        RECT 454.580 572.260 454.840 572.520 ;
        RECT 455.040 524.320 455.300 524.580 ;
        RECT 455.040 476.040 455.300 476.300 ;
        RECT 455.500 476.040 455.760 476.300 ;
        RECT 455.500 331.540 455.760 331.800 ;
        RECT 455.040 331.200 455.300 331.460 ;
        RECT 455.040 283.260 455.300 283.520 ;
        RECT 454.580 276.120 454.840 276.380 ;
        RECT 454.580 234.640 454.840 234.900 ;
        RECT 455.040 234.640 455.300 234.900 ;
        RECT 455.040 233.960 455.300 234.220 ;
        RECT 455.960 233.960 456.220 234.220 ;
        RECT 455.040 144.880 455.300 145.140 ;
        RECT 455.960 144.880 456.220 145.140 ;
        RECT 455.040 137.740 455.300 138.000 ;
        RECT 455.040 89.800 455.300 90.060 ;
        RECT 455.040 62.260 455.300 62.520 ;
        RECT 454.580 61.920 454.840 62.180 ;
        RECT 454.580 47.980 454.840 48.240 ;
        RECT 454.580 47.300 454.840 47.560 ;
      LAYER met2 ;
        RECT 507.340 1600.380 507.620 1604.000 ;
        RECT 507.340 1600.000 507.680 1600.380 ;
        RECT 507.540 1593.230 507.680 1600.000 ;
        RECT 455.040 1592.910 455.300 1593.230 ;
        RECT 507.480 1592.910 507.740 1593.230 ;
        RECT 455.100 1200.610 455.240 1592.910 ;
        RECT 454.640 1200.470 455.240 1200.610 ;
        RECT 454.640 1152.590 454.780 1200.470 ;
        RECT 454.120 1152.445 454.380 1152.590 ;
        RECT 453.190 1152.075 453.470 1152.445 ;
        RECT 454.110 1152.075 454.390 1152.445 ;
        RECT 454.580 1152.270 454.840 1152.590 ;
        RECT 453.260 1104.310 453.400 1152.075 ;
        RECT 453.200 1103.990 453.460 1104.310 ;
        RECT 455.040 1103.990 455.300 1104.310 ;
        RECT 455.100 1103.630 455.240 1103.990 ;
        RECT 455.040 1103.310 455.300 1103.630 ;
        RECT 455.500 1062.170 455.760 1062.490 ;
        RECT 455.560 1055.770 455.700 1062.170 ;
        RECT 455.560 1055.690 456.160 1055.770 ;
        RECT 455.560 1055.630 456.220 1055.690 ;
        RECT 455.960 1055.370 456.220 1055.630 ;
        RECT 456.020 1055.215 456.160 1055.370 ;
        RECT 455.040 1013.890 455.300 1014.210 ;
        RECT 455.100 917.990 455.240 1013.890 ;
        RECT 455.040 917.670 455.300 917.990 ;
        RECT 455.040 904.070 455.300 904.390 ;
        RECT 455.100 893.510 455.240 904.070 ;
        RECT 455.040 893.190 455.300 893.510 ;
        RECT 455.960 855.450 456.220 855.770 ;
        RECT 456.020 814.485 456.160 855.450 ;
        RECT 455.950 814.115 456.230 814.485 ;
        RECT 455.490 812.755 455.770 813.125 ;
        RECT 455.560 766.205 455.700 812.755 ;
        RECT 455.490 765.835 455.770 766.205 ;
        RECT 455.950 765.155 456.230 765.525 ;
        RECT 456.020 669.790 456.160 765.155 ;
        RECT 455.040 669.470 455.300 669.790 ;
        RECT 455.960 669.470 456.220 669.790 ;
        RECT 455.100 620.830 455.240 669.470 ;
        RECT 455.040 620.510 455.300 620.830 ;
        RECT 455.960 620.510 456.220 620.830 ;
        RECT 456.020 573.085 456.160 620.510 ;
        RECT 455.030 572.970 455.310 573.085 ;
        RECT 454.640 572.830 455.310 572.970 ;
        RECT 454.640 572.550 454.780 572.830 ;
        RECT 455.030 572.715 455.310 572.830 ;
        RECT 455.950 572.715 456.230 573.085 ;
        RECT 454.580 572.230 454.840 572.550 ;
        RECT 455.040 524.290 455.300 524.610 ;
        RECT 455.100 524.010 455.240 524.290 ;
        RECT 455.100 523.870 455.700 524.010 ;
        RECT 455.560 476.330 455.700 523.870 ;
        RECT 455.040 476.010 455.300 476.330 ;
        RECT 455.500 476.010 455.760 476.330 ;
        RECT 455.100 427.565 455.240 476.010 ;
        RECT 455.030 427.195 455.310 427.565 ;
        RECT 455.490 426.515 455.770 426.885 ;
        RECT 455.560 331.830 455.700 426.515 ;
        RECT 455.500 331.510 455.760 331.830 ;
        RECT 455.040 331.170 455.300 331.490 ;
        RECT 455.100 283.550 455.240 331.170 ;
        RECT 455.040 283.230 455.300 283.550 ;
        RECT 454.580 276.090 454.840 276.410 ;
        RECT 454.640 234.930 454.780 276.090 ;
        RECT 454.580 234.610 454.840 234.930 ;
        RECT 455.040 234.610 455.300 234.930 ;
        RECT 455.100 234.250 455.240 234.610 ;
        RECT 455.040 233.930 455.300 234.250 ;
        RECT 455.960 233.930 456.220 234.250 ;
        RECT 456.020 145.170 456.160 233.930 ;
        RECT 455.040 144.850 455.300 145.170 ;
        RECT 455.960 144.850 456.220 145.170 ;
        RECT 455.100 138.030 455.240 144.850 ;
        RECT 455.040 137.710 455.300 138.030 ;
        RECT 455.040 89.770 455.300 90.090 ;
        RECT 455.100 62.550 455.240 89.770 ;
        RECT 455.040 62.230 455.300 62.550 ;
        RECT 454.580 61.890 454.840 62.210 ;
        RECT 454.640 48.270 454.780 61.890 ;
        RECT 454.580 47.950 454.840 48.270 ;
        RECT 454.580 47.270 454.840 47.590 ;
        RECT 454.640 2.400 454.780 47.270 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 453.190 1152.120 453.470 1152.400 ;
        RECT 454.110 1152.120 454.390 1152.400 ;
        RECT 455.950 814.160 456.230 814.440 ;
        RECT 455.490 812.800 455.770 813.080 ;
        RECT 455.490 765.880 455.770 766.160 ;
        RECT 455.950 765.200 456.230 765.480 ;
        RECT 455.030 572.760 455.310 573.040 ;
        RECT 455.950 572.760 456.230 573.040 ;
        RECT 455.030 427.240 455.310 427.520 ;
        RECT 455.490 426.560 455.770 426.840 ;
      LAYER met3 ;
        RECT 453.165 1152.410 453.495 1152.425 ;
        RECT 454.085 1152.410 454.415 1152.425 ;
        RECT 453.165 1152.110 454.415 1152.410 ;
        RECT 453.165 1152.095 453.495 1152.110 ;
        RECT 454.085 1152.095 454.415 1152.110 ;
        RECT 455.925 814.450 456.255 814.465 ;
        RECT 455.710 814.135 456.255 814.450 ;
        RECT 455.710 813.105 456.010 814.135 ;
        RECT 455.465 812.790 456.010 813.105 ;
        RECT 455.465 812.775 455.795 812.790 ;
        RECT 455.465 766.170 455.795 766.185 ;
        RECT 454.790 765.870 455.795 766.170 ;
        RECT 454.790 765.490 455.090 765.870 ;
        RECT 455.465 765.855 455.795 765.870 ;
        RECT 455.925 765.490 456.255 765.505 ;
        RECT 454.790 765.190 456.255 765.490 ;
        RECT 455.925 765.175 456.255 765.190 ;
        RECT 455.005 573.050 455.335 573.065 ;
        RECT 455.925 573.050 456.255 573.065 ;
        RECT 455.005 572.750 456.255 573.050 ;
        RECT 455.005 572.735 455.335 572.750 ;
        RECT 455.925 572.735 456.255 572.750 ;
        RECT 455.005 427.530 455.335 427.545 ;
        RECT 455.005 427.230 456.010 427.530 ;
        RECT 455.005 427.215 455.335 427.230 ;
        RECT 455.710 426.865 456.010 427.230 ;
        RECT 455.465 426.550 456.010 426.865 ;
        RECT 455.465 426.535 455.795 426.550 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 481.690 1589.060 482.010 1589.120 ;
        RECT 513.890 1589.060 514.210 1589.120 ;
        RECT 481.690 1588.920 514.210 1589.060 ;
        RECT 481.690 1588.860 482.010 1588.920 ;
        RECT 513.890 1588.860 514.210 1588.920 ;
        RECT 472.490 20.640 472.810 20.700 ;
        RECT 479.390 20.640 479.710 20.700 ;
        RECT 472.490 20.500 479.710 20.640 ;
        RECT 472.490 20.440 472.810 20.500 ;
        RECT 479.390 20.440 479.710 20.500 ;
      LAYER via ;
        RECT 481.720 1588.860 481.980 1589.120 ;
        RECT 513.920 1588.860 514.180 1589.120 ;
        RECT 472.520 20.440 472.780 20.700 ;
        RECT 479.420 20.440 479.680 20.700 ;
      LAYER met2 ;
        RECT 513.780 1600.380 514.060 1604.000 ;
        RECT 513.780 1600.000 514.120 1600.380 ;
        RECT 513.980 1589.150 514.120 1600.000 ;
        RECT 481.720 1588.830 481.980 1589.150 ;
        RECT 513.920 1588.830 514.180 1589.150 ;
        RECT 481.780 1573.930 481.920 1588.830 ;
        RECT 479.480 1573.790 481.920 1573.930 ;
        RECT 479.480 20.730 479.620 1573.790 ;
        RECT 472.520 20.410 472.780 20.730 ;
        RECT 479.420 20.410 479.680 20.730 ;
        RECT 472.580 2.400 472.720 20.410 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 513.890 1587.360 514.210 1587.420 ;
        RECT 519.870 1587.360 520.190 1587.420 ;
        RECT 513.890 1587.220 520.190 1587.360 ;
        RECT 513.890 1587.160 514.210 1587.220 ;
        RECT 519.870 1587.160 520.190 1587.220 ;
        RECT 490.430 18.260 490.750 18.320 ;
        RECT 512.970 18.260 513.290 18.320 ;
        RECT 490.430 18.120 513.290 18.260 ;
        RECT 490.430 18.060 490.750 18.120 ;
        RECT 512.970 18.060 513.290 18.120 ;
      LAYER via ;
        RECT 513.920 1587.160 514.180 1587.420 ;
        RECT 519.900 1587.160 520.160 1587.420 ;
        RECT 490.460 18.060 490.720 18.320 ;
        RECT 513.000 18.060 513.260 18.320 ;
      LAYER met2 ;
        RECT 519.760 1600.380 520.040 1604.000 ;
        RECT 519.760 1600.000 520.100 1600.380 ;
        RECT 519.960 1587.450 520.100 1600.000 ;
        RECT 513.920 1587.130 514.180 1587.450 ;
        RECT 519.900 1587.130 520.160 1587.450 ;
        RECT 513.980 21.490 514.120 1587.130 ;
        RECT 513.060 21.350 514.120 21.490 ;
        RECT 513.060 18.350 513.200 21.350 ;
        RECT 490.460 18.030 490.720 18.350 ;
        RECT 513.000 18.030 513.260 18.350 ;
        RECT 490.520 2.400 490.660 18.030 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 525.465 1490.645 525.635 1511.215 ;
        RECT 525.925 1365.525 526.095 1400.715 ;
        RECT 525.925 1317.245 526.095 1352.435 ;
        RECT 525.925 1268.965 526.095 1304.155 ;
        RECT 525.465 1207.425 525.635 1255.875 ;
        RECT 525.465 1110.865 525.635 1124.975 ;
        RECT 525.465 1014.305 525.635 1028.415 ;
        RECT 525.465 917.745 525.635 931.855 ;
        RECT 525.465 689.605 525.635 717.655 ;
        RECT 525.465 572.645 525.635 620.755 ;
        RECT 525.465 476.085 525.635 524.195 ;
        RECT 525.465 420.665 525.635 427.635 ;
        RECT 525.005 331.245 525.175 372.895 ;
      LAYER mcon ;
        RECT 525.465 1511.045 525.635 1511.215 ;
        RECT 525.925 1400.545 526.095 1400.715 ;
        RECT 525.925 1352.265 526.095 1352.435 ;
        RECT 525.925 1303.985 526.095 1304.155 ;
        RECT 525.465 1255.705 525.635 1255.875 ;
        RECT 525.465 1124.805 525.635 1124.975 ;
        RECT 525.465 1028.245 525.635 1028.415 ;
        RECT 525.465 931.685 525.635 931.855 ;
        RECT 525.465 717.485 525.635 717.655 ;
        RECT 525.465 620.585 525.635 620.755 ;
        RECT 525.465 524.025 525.635 524.195 ;
        RECT 525.465 427.465 525.635 427.635 ;
        RECT 525.005 372.725 525.175 372.895 ;
      LAYER met1 ;
        RECT 525.390 1559.620 525.710 1559.880 ;
        RECT 525.480 1558.800 525.620 1559.620 ;
        RECT 525.850 1558.800 526.170 1558.860 ;
        RECT 525.480 1558.660 526.170 1558.800 ;
        RECT 525.850 1558.600 526.170 1558.660 ;
        RECT 525.405 1511.200 525.695 1511.245 ;
        RECT 525.850 1511.200 526.170 1511.260 ;
        RECT 525.405 1511.060 526.170 1511.200 ;
        RECT 525.405 1511.015 525.695 1511.060 ;
        RECT 525.850 1511.000 526.170 1511.060 ;
        RECT 525.390 1490.800 525.710 1490.860 ;
        RECT 525.195 1490.660 525.710 1490.800 ;
        RECT 525.390 1490.600 525.710 1490.660 ;
        RECT 525.850 1462.240 526.170 1462.300 ;
        RECT 526.770 1462.240 527.090 1462.300 ;
        RECT 525.850 1462.100 527.090 1462.240 ;
        RECT 525.850 1462.040 526.170 1462.100 ;
        RECT 526.770 1462.040 527.090 1462.100 ;
        RECT 525.850 1414.780 526.170 1415.040 ;
        RECT 525.940 1414.020 526.080 1414.780 ;
        RECT 525.850 1413.760 526.170 1414.020 ;
        RECT 525.850 1400.700 526.170 1400.760 ;
        RECT 525.655 1400.560 526.170 1400.700 ;
        RECT 525.850 1400.500 526.170 1400.560 ;
        RECT 525.850 1365.680 526.170 1365.740 ;
        RECT 525.655 1365.540 526.170 1365.680 ;
        RECT 525.850 1365.480 526.170 1365.540 ;
        RECT 525.850 1352.420 526.170 1352.480 ;
        RECT 525.655 1352.280 526.170 1352.420 ;
        RECT 525.850 1352.220 526.170 1352.280 ;
        RECT 525.850 1317.400 526.170 1317.460 ;
        RECT 525.655 1317.260 526.170 1317.400 ;
        RECT 525.850 1317.200 526.170 1317.260 ;
        RECT 525.850 1304.140 526.170 1304.200 ;
        RECT 525.655 1304.000 526.170 1304.140 ;
        RECT 525.850 1303.940 526.170 1304.000 ;
        RECT 525.850 1269.120 526.170 1269.180 ;
        RECT 525.655 1268.980 526.170 1269.120 ;
        RECT 525.850 1268.920 526.170 1268.980 ;
        RECT 525.405 1255.860 525.695 1255.905 ;
        RECT 525.850 1255.860 526.170 1255.920 ;
        RECT 525.405 1255.720 526.170 1255.860 ;
        RECT 525.405 1255.675 525.695 1255.720 ;
        RECT 525.850 1255.660 526.170 1255.720 ;
        RECT 525.390 1207.580 525.710 1207.640 ;
        RECT 525.195 1207.440 525.710 1207.580 ;
        RECT 525.390 1207.380 525.710 1207.440 ;
        RECT 525.390 1173.040 525.710 1173.300 ;
        RECT 525.480 1172.560 525.620 1173.040 ;
        RECT 525.850 1172.560 526.170 1172.620 ;
        RECT 525.480 1172.420 526.170 1172.560 ;
        RECT 525.850 1172.360 526.170 1172.420 ;
        RECT 525.390 1124.960 525.710 1125.020 ;
        RECT 525.195 1124.820 525.710 1124.960 ;
        RECT 525.390 1124.760 525.710 1124.820 ;
        RECT 525.390 1111.020 525.710 1111.080 ;
        RECT 525.195 1110.880 525.710 1111.020 ;
        RECT 525.390 1110.820 525.710 1110.880 ;
        RECT 525.390 1076.480 525.710 1076.740 ;
        RECT 525.480 1076.000 525.620 1076.480 ;
        RECT 525.850 1076.000 526.170 1076.060 ;
        RECT 525.480 1075.860 526.170 1076.000 ;
        RECT 525.850 1075.800 526.170 1075.860 ;
        RECT 525.390 1028.400 525.710 1028.460 ;
        RECT 525.195 1028.260 525.710 1028.400 ;
        RECT 525.390 1028.200 525.710 1028.260 ;
        RECT 525.390 1014.460 525.710 1014.520 ;
        RECT 525.195 1014.320 525.710 1014.460 ;
        RECT 525.390 1014.260 525.710 1014.320 ;
        RECT 525.390 979.920 525.710 980.180 ;
        RECT 525.480 979.440 525.620 979.920 ;
        RECT 525.850 979.440 526.170 979.500 ;
        RECT 525.480 979.300 526.170 979.440 ;
        RECT 525.850 979.240 526.170 979.300 ;
        RECT 525.390 931.840 525.710 931.900 ;
        RECT 525.195 931.700 525.710 931.840 ;
        RECT 525.390 931.640 525.710 931.700 ;
        RECT 525.390 917.900 525.710 917.960 ;
        RECT 525.195 917.760 525.710 917.900 ;
        RECT 525.390 917.700 525.710 917.760 ;
        RECT 525.390 883.360 525.710 883.620 ;
        RECT 525.480 882.880 525.620 883.360 ;
        RECT 525.850 882.880 526.170 882.940 ;
        RECT 525.480 882.740 526.170 882.880 ;
        RECT 525.850 882.680 526.170 882.740 ;
        RECT 524.470 845.480 524.790 845.540 ;
        RECT 525.390 845.480 525.710 845.540 ;
        RECT 524.470 845.340 525.710 845.480 ;
        RECT 524.470 845.280 524.790 845.340 ;
        RECT 525.390 845.280 525.710 845.340 ;
        RECT 525.390 786.800 525.710 787.060 ;
        RECT 525.480 786.320 525.620 786.800 ;
        RECT 525.850 786.320 526.170 786.380 ;
        RECT 525.480 786.180 526.170 786.320 ;
        RECT 525.850 786.120 526.170 786.180 ;
        RECT 525.850 738.720 526.170 738.780 ;
        RECT 525.480 738.580 526.170 738.720 ;
        RECT 525.480 738.100 525.620 738.580 ;
        RECT 525.850 738.520 526.170 738.580 ;
        RECT 525.390 737.840 525.710 738.100 ;
        RECT 525.390 717.640 525.710 717.700 ;
        RECT 525.195 717.500 525.710 717.640 ;
        RECT 525.390 717.440 525.710 717.500 ;
        RECT 525.390 689.760 525.710 689.820 ;
        RECT 525.195 689.620 525.710 689.760 ;
        RECT 525.390 689.560 525.710 689.620 ;
        RECT 525.850 642.160 526.170 642.220 ;
        RECT 525.480 642.020 526.170 642.160 ;
        RECT 525.480 641.540 525.620 642.020 ;
        RECT 525.850 641.960 526.170 642.020 ;
        RECT 525.390 641.280 525.710 641.540 ;
        RECT 525.390 620.740 525.710 620.800 ;
        RECT 525.195 620.600 525.710 620.740 ;
        RECT 525.390 620.540 525.710 620.600 ;
        RECT 525.405 572.800 525.695 572.845 ;
        RECT 525.850 572.800 526.170 572.860 ;
        RECT 525.405 572.660 526.170 572.800 ;
        RECT 525.405 572.615 525.695 572.660 ;
        RECT 525.850 572.600 526.170 572.660 ;
        RECT 525.850 545.600 526.170 545.660 ;
        RECT 525.480 545.460 526.170 545.600 ;
        RECT 525.480 544.980 525.620 545.460 ;
        RECT 525.850 545.400 526.170 545.460 ;
        RECT 525.390 544.720 525.710 544.980 ;
        RECT 525.390 524.180 525.710 524.240 ;
        RECT 525.195 524.040 525.710 524.180 ;
        RECT 525.390 523.980 525.710 524.040 ;
        RECT 525.405 476.240 525.695 476.285 ;
        RECT 525.850 476.240 526.170 476.300 ;
        RECT 525.405 476.100 526.170 476.240 ;
        RECT 525.405 476.055 525.695 476.100 ;
        RECT 525.850 476.040 526.170 476.100 ;
        RECT 525.850 449.040 526.170 449.100 ;
        RECT 525.480 448.900 526.170 449.040 ;
        RECT 525.480 448.420 525.620 448.900 ;
        RECT 525.850 448.840 526.170 448.900 ;
        RECT 525.390 448.160 525.710 448.420 ;
        RECT 525.390 427.620 525.710 427.680 ;
        RECT 525.195 427.480 525.710 427.620 ;
        RECT 525.390 427.420 525.710 427.480 ;
        RECT 525.405 420.635 525.695 420.865 ;
        RECT 524.930 420.480 525.250 420.540 ;
        RECT 525.480 420.480 525.620 420.635 ;
        RECT 524.930 420.340 525.620 420.480 ;
        RECT 524.930 420.280 525.250 420.340 ;
        RECT 524.930 372.880 525.250 372.940 ;
        RECT 524.735 372.740 525.250 372.880 ;
        RECT 524.930 372.680 525.250 372.740 ;
        RECT 524.930 331.400 525.250 331.460 ;
        RECT 524.735 331.260 525.250 331.400 ;
        RECT 524.930 331.200 525.250 331.260 ;
        RECT 524.930 324.260 525.250 324.320 ;
        RECT 526.310 324.260 526.630 324.320 ;
        RECT 524.930 324.120 526.630 324.260 ;
        RECT 524.930 324.060 525.250 324.120 ;
        RECT 526.310 324.060 526.630 324.120 ;
        RECT 524.470 234.840 524.790 234.900 ;
        RECT 526.310 234.840 526.630 234.900 ;
        RECT 524.470 234.700 526.630 234.840 ;
        RECT 524.470 234.640 524.790 234.700 ;
        RECT 526.310 234.640 526.630 234.700 ;
        RECT 524.470 206.620 524.790 206.680 ;
        RECT 525.850 206.620 526.170 206.680 ;
        RECT 524.470 206.480 526.170 206.620 ;
        RECT 524.470 206.420 524.790 206.480 ;
        RECT 525.850 206.420 526.170 206.480 ;
        RECT 525.850 159.020 526.170 159.080 ;
        RECT 525.480 158.880 526.170 159.020 ;
        RECT 525.480 158.740 525.620 158.880 ;
        RECT 525.850 158.820 526.170 158.880 ;
        RECT 525.390 158.480 525.710 158.740 ;
        RECT 507.910 20.300 508.230 20.360 ;
        RECT 524.930 20.300 525.250 20.360 ;
        RECT 507.910 20.160 525.250 20.300 ;
        RECT 507.910 20.100 508.230 20.160 ;
        RECT 524.930 20.100 525.250 20.160 ;
      LAYER via ;
        RECT 525.420 1559.620 525.680 1559.880 ;
        RECT 525.880 1558.600 526.140 1558.860 ;
        RECT 525.880 1511.000 526.140 1511.260 ;
        RECT 525.420 1490.600 525.680 1490.860 ;
        RECT 525.880 1462.040 526.140 1462.300 ;
        RECT 526.800 1462.040 527.060 1462.300 ;
        RECT 525.880 1414.780 526.140 1415.040 ;
        RECT 525.880 1413.760 526.140 1414.020 ;
        RECT 525.880 1400.500 526.140 1400.760 ;
        RECT 525.880 1365.480 526.140 1365.740 ;
        RECT 525.880 1352.220 526.140 1352.480 ;
        RECT 525.880 1317.200 526.140 1317.460 ;
        RECT 525.880 1303.940 526.140 1304.200 ;
        RECT 525.880 1268.920 526.140 1269.180 ;
        RECT 525.880 1255.660 526.140 1255.920 ;
        RECT 525.420 1207.380 525.680 1207.640 ;
        RECT 525.420 1173.040 525.680 1173.300 ;
        RECT 525.880 1172.360 526.140 1172.620 ;
        RECT 525.420 1124.760 525.680 1125.020 ;
        RECT 525.420 1110.820 525.680 1111.080 ;
        RECT 525.420 1076.480 525.680 1076.740 ;
        RECT 525.880 1075.800 526.140 1076.060 ;
        RECT 525.420 1028.200 525.680 1028.460 ;
        RECT 525.420 1014.260 525.680 1014.520 ;
        RECT 525.420 979.920 525.680 980.180 ;
        RECT 525.880 979.240 526.140 979.500 ;
        RECT 525.420 931.640 525.680 931.900 ;
        RECT 525.420 917.700 525.680 917.960 ;
        RECT 525.420 883.360 525.680 883.620 ;
        RECT 525.880 882.680 526.140 882.940 ;
        RECT 524.500 845.280 524.760 845.540 ;
        RECT 525.420 845.280 525.680 845.540 ;
        RECT 525.420 786.800 525.680 787.060 ;
        RECT 525.880 786.120 526.140 786.380 ;
        RECT 525.880 738.520 526.140 738.780 ;
        RECT 525.420 737.840 525.680 738.100 ;
        RECT 525.420 717.440 525.680 717.700 ;
        RECT 525.420 689.560 525.680 689.820 ;
        RECT 525.880 641.960 526.140 642.220 ;
        RECT 525.420 641.280 525.680 641.540 ;
        RECT 525.420 620.540 525.680 620.800 ;
        RECT 525.880 572.600 526.140 572.860 ;
        RECT 525.880 545.400 526.140 545.660 ;
        RECT 525.420 544.720 525.680 544.980 ;
        RECT 525.420 523.980 525.680 524.240 ;
        RECT 525.880 476.040 526.140 476.300 ;
        RECT 525.880 448.840 526.140 449.100 ;
        RECT 525.420 448.160 525.680 448.420 ;
        RECT 525.420 427.420 525.680 427.680 ;
        RECT 524.960 420.280 525.220 420.540 ;
        RECT 524.960 372.680 525.220 372.940 ;
        RECT 524.960 331.200 525.220 331.460 ;
        RECT 524.960 324.060 525.220 324.320 ;
        RECT 526.340 324.060 526.600 324.320 ;
        RECT 524.500 234.640 524.760 234.900 ;
        RECT 526.340 234.640 526.600 234.900 ;
        RECT 524.500 206.420 524.760 206.680 ;
        RECT 525.880 206.420 526.140 206.680 ;
        RECT 525.880 158.820 526.140 159.080 ;
        RECT 525.420 158.480 525.680 158.740 ;
        RECT 507.940 20.100 508.200 20.360 ;
        RECT 524.960 20.100 525.220 20.360 ;
      LAYER met2 ;
        RECT 525.740 1601.130 526.020 1604.000 ;
        RECT 525.020 1600.990 526.020 1601.130 ;
        RECT 525.020 1597.050 525.160 1600.990 ;
        RECT 525.740 1600.000 526.020 1600.990 ;
        RECT 525.020 1596.910 525.620 1597.050 ;
        RECT 525.480 1559.910 525.620 1596.910 ;
        RECT 525.420 1559.590 525.680 1559.910 ;
        RECT 525.880 1558.570 526.140 1558.890 ;
        RECT 525.940 1511.290 526.080 1558.570 ;
        RECT 525.880 1510.970 526.140 1511.290 ;
        RECT 525.420 1490.570 525.680 1490.890 ;
        RECT 525.480 1490.290 525.620 1490.570 ;
        RECT 525.870 1490.290 526.150 1490.405 ;
        RECT 525.480 1490.150 526.150 1490.290 ;
        RECT 525.870 1490.035 526.150 1490.150 ;
        RECT 526.790 1490.035 527.070 1490.405 ;
        RECT 526.860 1462.330 527.000 1490.035 ;
        RECT 525.880 1462.010 526.140 1462.330 ;
        RECT 526.800 1462.010 527.060 1462.330 ;
        RECT 525.940 1415.070 526.080 1462.010 ;
        RECT 525.880 1414.750 526.140 1415.070 ;
        RECT 525.880 1413.730 526.140 1414.050 ;
        RECT 525.940 1400.790 526.080 1413.730 ;
        RECT 525.880 1400.470 526.140 1400.790 ;
        RECT 525.880 1365.450 526.140 1365.770 ;
        RECT 525.940 1352.510 526.080 1365.450 ;
        RECT 525.880 1352.190 526.140 1352.510 ;
        RECT 525.880 1317.170 526.140 1317.490 ;
        RECT 525.940 1304.230 526.080 1317.170 ;
        RECT 525.880 1303.910 526.140 1304.230 ;
        RECT 525.880 1268.890 526.140 1269.210 ;
        RECT 525.940 1255.950 526.080 1268.890 ;
        RECT 525.880 1255.630 526.140 1255.950 ;
        RECT 525.420 1207.350 525.680 1207.670 ;
        RECT 525.480 1173.330 525.620 1207.350 ;
        RECT 525.420 1173.010 525.680 1173.330 ;
        RECT 525.880 1172.330 526.140 1172.650 ;
        RECT 525.940 1159.130 526.080 1172.330 ;
        RECT 525.480 1158.990 526.080 1159.130 ;
        RECT 525.480 1125.050 525.620 1158.990 ;
        RECT 525.420 1124.730 525.680 1125.050 ;
        RECT 525.420 1110.790 525.680 1111.110 ;
        RECT 525.480 1076.770 525.620 1110.790 ;
        RECT 525.420 1076.450 525.680 1076.770 ;
        RECT 525.880 1075.770 526.140 1076.090 ;
        RECT 525.940 1062.570 526.080 1075.770 ;
        RECT 525.480 1062.430 526.080 1062.570 ;
        RECT 525.480 1028.490 525.620 1062.430 ;
        RECT 525.420 1028.170 525.680 1028.490 ;
        RECT 525.420 1014.230 525.680 1014.550 ;
        RECT 525.480 980.210 525.620 1014.230 ;
        RECT 525.420 979.890 525.680 980.210 ;
        RECT 525.880 979.210 526.140 979.530 ;
        RECT 525.940 966.010 526.080 979.210 ;
        RECT 525.480 965.870 526.080 966.010 ;
        RECT 525.480 931.930 525.620 965.870 ;
        RECT 525.420 931.610 525.680 931.930 ;
        RECT 525.420 917.670 525.680 917.990 ;
        RECT 525.480 883.650 525.620 917.670 ;
        RECT 525.420 883.330 525.680 883.650 ;
        RECT 525.880 882.650 526.140 882.970 ;
        RECT 525.940 869.450 526.080 882.650 ;
        RECT 525.480 869.310 526.080 869.450 ;
        RECT 525.480 845.570 525.620 869.310 ;
        RECT 524.500 845.250 524.760 845.570 ;
        RECT 525.420 845.250 525.680 845.570 ;
        RECT 524.560 821.285 524.700 845.250 ;
        RECT 524.490 820.915 524.770 821.285 ;
        RECT 525.410 820.915 525.690 821.285 ;
        RECT 525.480 787.090 525.620 820.915 ;
        RECT 525.420 786.770 525.680 787.090 ;
        RECT 525.880 786.090 526.140 786.410 ;
        RECT 525.940 738.810 526.080 786.090 ;
        RECT 525.880 738.490 526.140 738.810 ;
        RECT 525.420 737.810 525.680 738.130 ;
        RECT 525.480 717.730 525.620 737.810 ;
        RECT 525.420 717.410 525.680 717.730 ;
        RECT 525.420 689.530 525.680 689.850 ;
        RECT 525.480 669.530 525.620 689.530 ;
        RECT 525.480 669.390 526.080 669.530 ;
        RECT 525.940 642.250 526.080 669.390 ;
        RECT 525.880 641.930 526.140 642.250 ;
        RECT 525.420 641.250 525.680 641.570 ;
        RECT 525.480 620.830 525.620 641.250 ;
        RECT 525.420 620.510 525.680 620.830 ;
        RECT 525.880 572.570 526.140 572.890 ;
        RECT 525.940 545.690 526.080 572.570 ;
        RECT 525.880 545.370 526.140 545.690 ;
        RECT 525.420 544.690 525.680 545.010 ;
        RECT 525.480 524.270 525.620 544.690 ;
        RECT 525.420 523.950 525.680 524.270 ;
        RECT 525.880 476.010 526.140 476.330 ;
        RECT 525.940 449.130 526.080 476.010 ;
        RECT 525.880 448.810 526.140 449.130 ;
        RECT 525.420 448.130 525.680 448.450 ;
        RECT 525.480 427.710 525.620 448.130 ;
        RECT 525.420 427.390 525.680 427.710 ;
        RECT 524.960 420.250 525.220 420.570 ;
        RECT 525.020 372.970 525.160 420.250 ;
        RECT 524.960 372.650 525.220 372.970 ;
        RECT 524.960 331.170 525.220 331.490 ;
        RECT 525.020 324.350 525.160 331.170 ;
        RECT 524.960 324.030 525.220 324.350 ;
        RECT 526.340 324.030 526.600 324.350 ;
        RECT 526.400 234.930 526.540 324.030 ;
        RECT 524.500 234.610 524.760 234.930 ;
        RECT 526.340 234.610 526.600 234.930 ;
        RECT 524.560 206.710 524.700 234.610 ;
        RECT 524.500 206.390 524.760 206.710 ;
        RECT 525.880 206.390 526.140 206.710 ;
        RECT 525.940 159.110 526.080 206.390 ;
        RECT 525.880 158.790 526.140 159.110 ;
        RECT 525.420 158.450 525.680 158.770 ;
        RECT 525.480 144.570 525.620 158.450 ;
        RECT 525.480 144.430 526.080 144.570 ;
        RECT 525.940 21.490 526.080 144.430 ;
        RECT 525.020 21.350 526.080 21.490 ;
        RECT 525.020 20.390 525.160 21.350 ;
        RECT 507.940 20.070 508.200 20.390 ;
        RECT 524.960 20.070 525.220 20.390 ;
        RECT 508.000 2.400 508.140 20.070 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 525.870 1490.080 526.150 1490.360 ;
        RECT 526.790 1490.080 527.070 1490.360 ;
        RECT 524.490 820.960 524.770 821.240 ;
        RECT 525.410 820.960 525.690 821.240 ;
      LAYER met3 ;
        RECT 525.845 1490.370 526.175 1490.385 ;
        RECT 526.765 1490.370 527.095 1490.385 ;
        RECT 525.845 1490.070 527.095 1490.370 ;
        RECT 525.845 1490.055 526.175 1490.070 ;
        RECT 526.765 1490.055 527.095 1490.070 ;
        RECT 524.465 821.250 524.795 821.265 ;
        RECT 525.385 821.250 525.715 821.265 ;
        RECT 524.465 820.950 525.715 821.250 ;
        RECT 524.465 820.935 524.795 820.950 ;
        RECT 525.385 820.935 525.715 820.950 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 20.640 526.170 20.700 ;
        RECT 531.370 20.640 531.690 20.700 ;
        RECT 525.850 20.500 531.690 20.640 ;
        RECT 525.850 20.440 526.170 20.500 ;
        RECT 531.370 20.440 531.690 20.500 ;
      LAYER via ;
        RECT 525.880 20.440 526.140 20.700 ;
        RECT 531.400 20.440 531.660 20.700 ;
      LAYER met2 ;
        RECT 532.180 1600.450 532.460 1604.000 ;
        RECT 531.460 1600.310 532.460 1600.450 ;
        RECT 531.460 20.730 531.600 1600.310 ;
        RECT 532.180 1600.000 532.460 1600.310 ;
        RECT 525.880 20.410 526.140 20.730 ;
        RECT 531.400 20.410 531.660 20.730 ;
        RECT 525.940 2.400 526.080 20.410 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 539.190 20.640 539.510 20.700 ;
        RECT 543.790 20.640 544.110 20.700 ;
        RECT 539.190 20.500 544.110 20.640 ;
        RECT 539.190 20.440 539.510 20.500 ;
        RECT 543.790 20.440 544.110 20.500 ;
      LAYER via ;
        RECT 539.220 20.440 539.480 20.700 ;
        RECT 543.820 20.440 544.080 20.700 ;
      LAYER met2 ;
        RECT 538.160 1600.450 538.440 1604.000 ;
        RECT 538.160 1600.310 539.420 1600.450 ;
        RECT 538.160 1600.000 538.440 1600.310 ;
        RECT 539.280 20.730 539.420 1600.310 ;
        RECT 539.220 20.410 539.480 20.730 ;
        RECT 543.820 20.410 544.080 20.730 ;
        RECT 543.880 2.400 544.020 20.410 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 544.710 1591.440 545.030 1591.500 ;
        RECT 555.290 1591.440 555.610 1591.500 ;
        RECT 544.710 1591.300 555.610 1591.440 ;
        RECT 544.710 1591.240 545.030 1591.300 ;
        RECT 555.290 1591.240 555.610 1591.300 ;
        RECT 555.290 17.580 555.610 17.640 ;
        RECT 561.730 17.580 562.050 17.640 ;
        RECT 555.290 17.440 562.050 17.580 ;
        RECT 555.290 17.380 555.610 17.440 ;
        RECT 561.730 17.380 562.050 17.440 ;
      LAYER via ;
        RECT 544.740 1591.240 545.000 1591.500 ;
        RECT 555.320 1591.240 555.580 1591.500 ;
        RECT 555.320 17.380 555.580 17.640 ;
        RECT 561.760 17.380 562.020 17.640 ;
      LAYER met2 ;
        RECT 544.600 1600.380 544.880 1604.000 ;
        RECT 544.600 1600.000 544.940 1600.380 ;
        RECT 544.800 1591.530 544.940 1600.000 ;
        RECT 544.740 1591.210 545.000 1591.530 ;
        RECT 555.320 1591.210 555.580 1591.530 ;
        RECT 555.380 17.670 555.520 1591.210 ;
        RECT 555.320 17.350 555.580 17.670 ;
        RECT 561.760 17.350 562.020 17.670 ;
        RECT 561.820 2.400 561.960 17.350 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 550.690 1590.760 551.010 1590.820 ;
        RECT 555.750 1590.760 556.070 1590.820 ;
        RECT 550.690 1590.620 556.070 1590.760 ;
        RECT 550.690 1590.560 551.010 1590.620 ;
        RECT 555.750 1590.560 556.070 1590.620 ;
        RECT 555.750 18.260 556.070 18.320 ;
        RECT 555.750 18.120 562.420 18.260 ;
        RECT 555.750 18.060 556.070 18.120 ;
        RECT 562.280 17.580 562.420 18.120 ;
        RECT 579.670 17.580 579.990 17.640 ;
        RECT 562.280 17.440 579.990 17.580 ;
        RECT 579.670 17.380 579.990 17.440 ;
      LAYER via ;
        RECT 550.720 1590.560 550.980 1590.820 ;
        RECT 555.780 1590.560 556.040 1590.820 ;
        RECT 555.780 18.060 556.040 18.320 ;
        RECT 579.700 17.380 579.960 17.640 ;
      LAYER met2 ;
        RECT 550.580 1600.380 550.860 1604.000 ;
        RECT 550.580 1600.000 550.920 1600.380 ;
        RECT 550.780 1590.850 550.920 1600.000 ;
        RECT 550.720 1590.530 550.980 1590.850 ;
        RECT 555.780 1590.530 556.040 1590.850 ;
        RECT 555.840 18.350 555.980 1590.530 ;
        RECT 555.780 18.030 556.040 18.350 ;
        RECT 579.700 17.350 579.960 17.670 ;
        RECT 579.760 2.400 579.900 17.350 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 16.900 86.410 16.960 ;
        RECT 89.310 16.900 89.630 16.960 ;
        RECT 86.090 16.760 89.630 16.900 ;
        RECT 86.090 16.700 86.410 16.760 ;
        RECT 89.310 16.700 89.630 16.760 ;
      LAYER via ;
        RECT 86.120 16.700 86.380 16.960 ;
        RECT 89.340 16.700 89.600 16.960 ;
      LAYER met2 ;
        RECT 379.460 1600.380 379.740 1604.000 ;
        RECT 379.460 1600.000 379.800 1600.380 ;
        RECT 379.660 1592.405 379.800 1600.000 ;
        RECT 89.330 1592.035 89.610 1592.405 ;
        RECT 379.590 1592.035 379.870 1592.405 ;
        RECT 89.400 16.990 89.540 1592.035 ;
        RECT 86.120 16.670 86.380 16.990 ;
        RECT 89.340 16.670 89.600 16.990 ;
        RECT 86.180 2.400 86.320 16.670 ;
        RECT 85.970 -4.800 86.530 2.400 ;
      LAYER via2 ;
        RECT 89.330 1592.080 89.610 1592.360 ;
        RECT 379.590 1592.080 379.870 1592.360 ;
      LAYER met3 ;
        RECT 89.305 1592.370 89.635 1592.385 ;
        RECT 379.565 1592.370 379.895 1592.385 ;
        RECT 89.305 1592.070 379.895 1592.370 ;
        RECT 89.305 1592.055 89.635 1592.070 ;
        RECT 379.565 1592.055 379.895 1592.070 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 558.050 19.280 558.370 19.340 ;
        RECT 597.150 19.280 597.470 19.340 ;
        RECT 558.050 19.140 597.470 19.280 ;
        RECT 558.050 19.080 558.370 19.140 ;
        RECT 597.150 19.080 597.470 19.140 ;
      LAYER via ;
        RECT 558.080 19.080 558.340 19.340 ;
        RECT 597.180 19.080 597.440 19.340 ;
      LAYER met2 ;
        RECT 557.020 1600.450 557.300 1604.000 ;
        RECT 557.020 1600.310 558.280 1600.450 ;
        RECT 557.020 1600.000 557.300 1600.310 ;
        RECT 558.140 19.370 558.280 1600.310 ;
        RECT 558.080 19.050 558.340 19.370 ;
        RECT 597.180 19.050 597.440 19.370 ;
        RECT 597.240 2.400 597.380 19.050 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 563.110 1590.080 563.430 1590.140 ;
        RECT 565.410 1590.080 565.730 1590.140 ;
        RECT 563.110 1589.940 565.730 1590.080 ;
        RECT 563.110 1589.880 563.430 1589.940 ;
        RECT 565.410 1589.880 565.730 1589.940 ;
        RECT 565.410 18.260 565.730 18.320 ;
        RECT 615.090 18.260 615.410 18.320 ;
        RECT 565.410 18.120 615.410 18.260 ;
        RECT 565.410 18.060 565.730 18.120 ;
        RECT 615.090 18.060 615.410 18.120 ;
      LAYER via ;
        RECT 563.140 1589.880 563.400 1590.140 ;
        RECT 565.440 1589.880 565.700 1590.140 ;
        RECT 565.440 18.060 565.700 18.320 ;
        RECT 615.120 18.060 615.380 18.320 ;
      LAYER met2 ;
        RECT 563.000 1600.380 563.280 1604.000 ;
        RECT 563.000 1600.000 563.340 1600.380 ;
        RECT 563.200 1590.170 563.340 1600.000 ;
        RECT 563.140 1589.850 563.400 1590.170 ;
        RECT 565.440 1589.850 565.700 1590.170 ;
        RECT 565.500 18.350 565.640 1589.850 ;
        RECT 565.440 18.030 565.700 18.350 ;
        RECT 615.120 18.030 615.380 18.350 ;
        RECT 615.180 2.400 615.320 18.030 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 387.465 1086.725 387.635 1128.375 ;
        RECT 387.465 1014.305 387.635 1028.415 ;
        RECT 387.465 869.465 387.635 917.575 ;
        RECT 387.465 379.525 387.635 427.635 ;
        RECT 387.465 89.845 387.635 137.955 ;
        RECT 352.505 17.085 352.675 18.955 ;
        RECT 375.505 17.425 376.595 17.595 ;
        RECT 357.565 16.235 357.735 17.255 ;
        RECT 357.565 16.065 359.575 16.235 ;
        RECT 375.505 16.065 375.675 17.425 ;
        RECT 376.425 17.085 376.595 17.425 ;
        RECT 381.025 17.085 381.195 18.955 ;
      LAYER mcon ;
        RECT 387.465 1128.205 387.635 1128.375 ;
        RECT 387.465 1028.245 387.635 1028.415 ;
        RECT 387.465 917.405 387.635 917.575 ;
        RECT 387.465 427.465 387.635 427.635 ;
        RECT 387.465 137.785 387.635 137.955 ;
        RECT 352.505 18.785 352.675 18.955 ;
        RECT 381.025 18.785 381.195 18.955 ;
        RECT 357.565 17.085 357.735 17.255 ;
        RECT 359.405 16.065 359.575 16.235 ;
      LAYER met1 ;
        RECT 387.850 1546.360 388.170 1546.620 ;
        RECT 387.940 1545.940 388.080 1546.360 ;
        RECT 387.850 1545.680 388.170 1545.940 ;
        RECT 387.850 1449.320 388.170 1449.380 ;
        RECT 388.310 1449.320 388.630 1449.380 ;
        RECT 387.850 1449.180 388.630 1449.320 ;
        RECT 387.850 1449.120 388.170 1449.180 ;
        RECT 388.310 1449.120 388.630 1449.180 ;
        RECT 387.850 1414.980 388.170 1415.040 ;
        RECT 387.480 1414.840 388.170 1414.980 ;
        RECT 387.480 1414.360 387.620 1414.840 ;
        RECT 387.850 1414.780 388.170 1414.840 ;
        RECT 387.390 1414.100 387.710 1414.360 ;
        RECT 387.390 1352.420 387.710 1352.480 ;
        RECT 387.850 1352.420 388.170 1352.480 ;
        RECT 387.390 1352.280 388.170 1352.420 ;
        RECT 387.390 1352.220 387.710 1352.280 ;
        RECT 387.850 1352.220 388.170 1352.280 ;
        RECT 388.310 1224.920 388.630 1224.980 ;
        RECT 389.230 1224.920 389.550 1224.980 ;
        RECT 388.310 1224.780 389.550 1224.920 ;
        RECT 388.310 1224.720 388.630 1224.780 ;
        RECT 389.230 1224.720 389.550 1224.780 ;
        RECT 387.405 1128.360 387.695 1128.405 ;
        RECT 388.770 1128.360 389.090 1128.420 ;
        RECT 387.405 1128.220 389.090 1128.360 ;
        RECT 387.405 1128.175 387.695 1128.220 ;
        RECT 388.770 1128.160 389.090 1128.220 ;
        RECT 387.405 1086.880 387.695 1086.925 ;
        RECT 387.850 1086.880 388.170 1086.940 ;
        RECT 387.405 1086.740 388.170 1086.880 ;
        RECT 387.405 1086.695 387.695 1086.740 ;
        RECT 387.850 1086.680 388.170 1086.740 ;
        RECT 387.390 1028.400 387.710 1028.460 ;
        RECT 387.195 1028.260 387.710 1028.400 ;
        RECT 387.390 1028.200 387.710 1028.260 ;
        RECT 387.390 1014.460 387.710 1014.520 ;
        RECT 387.195 1014.320 387.710 1014.460 ;
        RECT 387.390 1014.260 387.710 1014.320 ;
        RECT 387.850 932.180 388.170 932.240 ;
        RECT 387.480 932.040 388.170 932.180 ;
        RECT 387.480 931.560 387.620 932.040 ;
        RECT 387.850 931.980 388.170 932.040 ;
        RECT 387.390 931.300 387.710 931.560 ;
        RECT 387.390 917.560 387.710 917.620 ;
        RECT 387.195 917.420 387.710 917.560 ;
        RECT 387.390 917.360 387.710 917.420 ;
        RECT 387.405 869.620 387.695 869.665 ;
        RECT 387.850 869.620 388.170 869.680 ;
        RECT 387.405 869.480 388.170 869.620 ;
        RECT 387.405 869.435 387.695 869.480 ;
        RECT 387.850 869.420 388.170 869.480 ;
        RECT 386.930 838.340 387.250 838.400 ;
        RECT 387.850 838.340 388.170 838.400 ;
        RECT 386.930 838.200 388.170 838.340 ;
        RECT 386.930 838.140 387.250 838.200 ;
        RECT 387.850 838.140 388.170 838.200 ;
        RECT 387.390 765.720 387.710 765.980 ;
        RECT 387.480 765.240 387.620 765.720 ;
        RECT 388.310 765.240 388.630 765.300 ;
        RECT 387.480 765.100 388.630 765.240 ;
        RECT 388.310 765.040 388.630 765.100 ;
        RECT 387.850 545.600 388.170 545.660 ;
        RECT 387.480 545.460 388.170 545.600 ;
        RECT 387.480 544.980 387.620 545.460 ;
        RECT 387.850 545.400 388.170 545.460 ;
        RECT 387.390 544.720 387.710 544.980 ;
        RECT 387.390 427.620 387.710 427.680 ;
        RECT 387.195 427.480 387.710 427.620 ;
        RECT 387.390 427.420 387.710 427.480 ;
        RECT 387.405 379.680 387.695 379.725 ;
        RECT 387.850 379.680 388.170 379.740 ;
        RECT 387.405 379.540 388.170 379.680 ;
        RECT 387.405 379.495 387.695 379.540 ;
        RECT 387.850 379.480 388.170 379.540 ;
        RECT 387.850 352.480 388.170 352.540 ;
        RECT 387.480 352.340 388.170 352.480 ;
        RECT 387.480 351.860 387.620 352.340 ;
        RECT 387.850 352.280 388.170 352.340 ;
        RECT 387.390 351.600 387.710 351.860 ;
        RECT 386.930 331.060 387.250 331.120 ;
        RECT 387.390 331.060 387.710 331.120 ;
        RECT 386.930 330.920 387.710 331.060 ;
        RECT 386.930 330.860 387.250 330.920 ;
        RECT 387.390 330.860 387.710 330.920 ;
        RECT 386.930 193.500 387.250 193.760 ;
        RECT 387.020 193.080 387.160 193.500 ;
        RECT 386.930 192.820 387.250 193.080 ;
        RECT 387.390 137.940 387.710 138.000 ;
        RECT 387.195 137.800 387.710 137.940 ;
        RECT 387.390 137.740 387.710 137.800 ;
        RECT 387.390 90.000 387.710 90.060 ;
        RECT 387.195 89.860 387.710 90.000 ;
        RECT 387.390 89.800 387.710 89.860 ;
        RECT 109.550 18.940 109.870 19.000 ;
        RECT 352.445 18.940 352.735 18.985 ;
        RECT 109.550 18.800 352.735 18.940 ;
        RECT 109.550 18.740 109.870 18.800 ;
        RECT 352.445 18.755 352.735 18.800 ;
        RECT 380.965 18.940 381.255 18.985 ;
        RECT 387.390 18.940 387.710 19.000 ;
        RECT 380.965 18.800 387.710 18.940 ;
        RECT 380.965 18.755 381.255 18.800 ;
        RECT 387.390 18.740 387.710 18.800 ;
        RECT 352.445 17.240 352.735 17.285 ;
        RECT 357.505 17.240 357.795 17.285 ;
        RECT 352.445 17.100 357.795 17.240 ;
        RECT 352.445 17.055 352.735 17.100 ;
        RECT 357.505 17.055 357.795 17.100 ;
        RECT 376.365 17.240 376.655 17.285 ;
        RECT 380.965 17.240 381.255 17.285 ;
        RECT 376.365 17.100 381.255 17.240 ;
        RECT 376.365 17.055 376.655 17.100 ;
        RECT 380.965 17.055 381.255 17.100 ;
        RECT 359.345 16.220 359.635 16.265 ;
        RECT 375.445 16.220 375.735 16.265 ;
        RECT 359.345 16.080 375.735 16.220 ;
        RECT 359.345 16.035 359.635 16.080 ;
        RECT 375.445 16.035 375.735 16.080 ;
      LAYER via ;
        RECT 387.880 1546.360 388.140 1546.620 ;
        RECT 387.880 1545.680 388.140 1545.940 ;
        RECT 387.880 1449.120 388.140 1449.380 ;
        RECT 388.340 1449.120 388.600 1449.380 ;
        RECT 387.880 1414.780 388.140 1415.040 ;
        RECT 387.420 1414.100 387.680 1414.360 ;
        RECT 387.420 1352.220 387.680 1352.480 ;
        RECT 387.880 1352.220 388.140 1352.480 ;
        RECT 388.340 1224.720 388.600 1224.980 ;
        RECT 389.260 1224.720 389.520 1224.980 ;
        RECT 388.800 1128.160 389.060 1128.420 ;
        RECT 387.880 1086.680 388.140 1086.940 ;
        RECT 387.420 1028.200 387.680 1028.460 ;
        RECT 387.420 1014.260 387.680 1014.520 ;
        RECT 387.880 931.980 388.140 932.240 ;
        RECT 387.420 931.300 387.680 931.560 ;
        RECT 387.420 917.360 387.680 917.620 ;
        RECT 387.880 869.420 388.140 869.680 ;
        RECT 386.960 838.140 387.220 838.400 ;
        RECT 387.880 838.140 388.140 838.400 ;
        RECT 387.420 765.720 387.680 765.980 ;
        RECT 388.340 765.040 388.600 765.300 ;
        RECT 387.880 545.400 388.140 545.660 ;
        RECT 387.420 544.720 387.680 544.980 ;
        RECT 387.420 427.420 387.680 427.680 ;
        RECT 387.880 379.480 388.140 379.740 ;
        RECT 387.880 352.280 388.140 352.540 ;
        RECT 387.420 351.600 387.680 351.860 ;
        RECT 386.960 330.860 387.220 331.120 ;
        RECT 387.420 330.860 387.680 331.120 ;
        RECT 386.960 193.500 387.220 193.760 ;
        RECT 386.960 192.820 387.220 193.080 ;
        RECT 387.420 137.740 387.680 138.000 ;
        RECT 387.420 89.800 387.680 90.060 ;
        RECT 109.580 18.740 109.840 19.000 ;
        RECT 387.420 18.740 387.680 19.000 ;
      LAYER met2 ;
        RECT 387.740 1601.130 388.020 1604.000 ;
        RECT 387.020 1600.990 388.020 1601.130 ;
        RECT 387.020 1597.050 387.160 1600.990 ;
        RECT 387.740 1600.000 388.020 1600.990 ;
        RECT 387.020 1596.910 387.620 1597.050 ;
        RECT 387.480 1593.820 387.620 1596.910 ;
        RECT 387.480 1593.680 388.080 1593.820 ;
        RECT 387.940 1546.650 388.080 1593.680 ;
        RECT 387.880 1546.330 388.140 1546.650 ;
        RECT 387.880 1545.650 388.140 1545.970 ;
        RECT 387.940 1545.370 388.080 1545.650 ;
        RECT 387.940 1545.230 388.540 1545.370 ;
        RECT 388.400 1449.410 388.540 1545.230 ;
        RECT 387.880 1449.090 388.140 1449.410 ;
        RECT 388.340 1449.090 388.600 1449.410 ;
        RECT 387.940 1415.070 388.080 1449.090 ;
        RECT 387.880 1414.750 388.140 1415.070 ;
        RECT 387.420 1414.070 387.680 1414.390 ;
        RECT 387.480 1352.510 387.620 1414.070 ;
        RECT 387.420 1352.190 387.680 1352.510 ;
        RECT 387.880 1352.190 388.140 1352.510 ;
        RECT 387.940 1265.890 388.080 1352.190 ;
        RECT 387.480 1265.750 388.080 1265.890 ;
        RECT 387.480 1242.205 387.620 1265.750 ;
        RECT 387.410 1241.835 387.690 1242.205 ;
        RECT 389.250 1241.835 389.530 1242.205 ;
        RECT 389.320 1225.010 389.460 1241.835 ;
        RECT 388.340 1224.690 388.600 1225.010 ;
        RECT 389.260 1224.690 389.520 1225.010 ;
        RECT 388.400 1152.330 388.540 1224.690 ;
        RECT 388.400 1152.190 389.000 1152.330 ;
        RECT 388.860 1128.450 389.000 1152.190 ;
        RECT 388.800 1128.130 389.060 1128.450 ;
        RECT 387.880 1086.650 388.140 1086.970 ;
        RECT 387.940 1062.570 388.080 1086.650 ;
        RECT 387.480 1062.430 388.080 1062.570 ;
        RECT 387.480 1028.490 387.620 1062.430 ;
        RECT 387.420 1028.170 387.680 1028.490 ;
        RECT 387.420 1014.405 387.680 1014.550 ;
        RECT 387.410 1014.035 387.690 1014.405 ;
        RECT 387.870 978.675 388.150 979.045 ;
        RECT 387.940 932.270 388.080 978.675 ;
        RECT 387.880 931.950 388.140 932.270 ;
        RECT 387.420 931.270 387.680 931.590 ;
        RECT 387.480 917.650 387.620 931.270 ;
        RECT 387.420 917.330 387.680 917.650 ;
        RECT 387.880 869.390 388.140 869.710 ;
        RECT 387.940 838.430 388.080 869.390 ;
        RECT 386.960 838.110 387.220 838.430 ;
        RECT 387.880 838.110 388.140 838.430 ;
        RECT 387.020 814.370 387.160 838.110 ;
        RECT 387.020 814.230 387.620 814.370 ;
        RECT 387.480 766.010 387.620 814.230 ;
        RECT 387.420 765.690 387.680 766.010 ;
        RECT 388.340 765.010 388.600 765.330 ;
        RECT 388.400 628.165 388.540 765.010 ;
        RECT 387.410 627.795 387.690 628.165 ;
        RECT 388.330 627.795 388.610 628.165 ;
        RECT 387.480 603.570 387.620 627.795 ;
        RECT 387.480 603.430 388.080 603.570 ;
        RECT 387.940 545.690 388.080 603.430 ;
        RECT 387.880 545.370 388.140 545.690 ;
        RECT 387.420 544.690 387.680 545.010 ;
        RECT 387.480 483.210 387.620 544.690 ;
        RECT 387.480 483.070 388.080 483.210 ;
        RECT 387.940 435.725 388.080 483.070 ;
        RECT 387.870 435.355 388.150 435.725 ;
        RECT 387.410 434.675 387.690 435.045 ;
        RECT 387.480 427.710 387.620 434.675 ;
        RECT 387.420 427.390 387.680 427.710 ;
        RECT 387.880 379.450 388.140 379.770 ;
        RECT 387.940 352.570 388.080 379.450 ;
        RECT 387.880 352.250 388.140 352.570 ;
        RECT 387.420 351.570 387.680 351.890 ;
        RECT 387.480 331.150 387.620 351.570 ;
        RECT 386.960 330.830 387.220 331.150 ;
        RECT 387.420 330.830 387.680 331.150 ;
        RECT 387.020 193.790 387.160 330.830 ;
        RECT 386.960 193.470 387.220 193.790 ;
        RECT 386.960 192.790 387.220 193.110 ;
        RECT 387.020 145.250 387.160 192.790 ;
        RECT 387.020 145.110 387.620 145.250 ;
        RECT 387.480 138.030 387.620 145.110 ;
        RECT 387.420 137.710 387.680 138.030 ;
        RECT 387.420 89.770 387.680 90.090 ;
        RECT 387.480 19.030 387.620 89.770 ;
        RECT 109.580 18.710 109.840 19.030 ;
        RECT 387.420 18.710 387.680 19.030 ;
        RECT 109.640 2.400 109.780 18.710 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 387.410 1241.880 387.690 1242.160 ;
        RECT 389.250 1241.880 389.530 1242.160 ;
        RECT 387.410 1014.080 387.690 1014.360 ;
        RECT 387.870 978.720 388.150 979.000 ;
        RECT 387.410 627.840 387.690 628.120 ;
        RECT 388.330 627.840 388.610 628.120 ;
        RECT 387.870 435.400 388.150 435.680 ;
        RECT 387.410 434.720 387.690 435.000 ;
      LAYER met3 ;
        RECT 387.385 1242.170 387.715 1242.185 ;
        RECT 389.225 1242.170 389.555 1242.185 ;
        RECT 387.385 1241.870 389.555 1242.170 ;
        RECT 387.385 1241.855 387.715 1241.870 ;
        RECT 389.225 1241.855 389.555 1241.870 ;
        RECT 387.385 1014.380 387.715 1014.385 ;
        RECT 387.385 1014.370 387.970 1014.380 ;
        RECT 387.160 1014.070 387.970 1014.370 ;
        RECT 387.385 1014.060 387.970 1014.070 ;
        RECT 387.385 1014.055 387.715 1014.060 ;
        RECT 387.845 979.020 388.175 979.025 ;
        RECT 387.590 979.010 388.175 979.020 ;
        RECT 387.390 978.710 388.175 979.010 ;
        RECT 387.590 978.700 388.175 978.710 ;
        RECT 387.845 978.695 388.175 978.700 ;
        RECT 387.385 628.130 387.715 628.145 ;
        RECT 388.305 628.130 388.635 628.145 ;
        RECT 387.385 627.830 388.635 628.130 ;
        RECT 387.385 627.815 387.715 627.830 ;
        RECT 388.305 627.815 388.635 627.830 ;
        RECT 387.845 435.690 388.175 435.705 ;
        RECT 387.630 435.375 388.175 435.690 ;
        RECT 387.630 435.025 387.930 435.375 ;
        RECT 387.385 434.710 387.930 435.025 ;
        RECT 387.385 434.695 387.715 434.710 ;
      LAYER via3 ;
        RECT 387.620 1014.060 387.940 1014.380 ;
        RECT 387.620 978.700 387.940 979.020 ;
      LAYER met4 ;
        RECT 387.615 1014.055 387.945 1014.385 ;
        RECT 387.630 979.025 387.930 1014.055 ;
        RECT 387.615 978.695 387.945 979.025 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 137.610 1591.440 137.930 1591.500 ;
        RECT 396.130 1591.440 396.450 1591.500 ;
        RECT 137.610 1591.300 396.450 1591.440 ;
        RECT 137.610 1591.240 137.930 1591.300 ;
        RECT 396.130 1591.240 396.450 1591.300 ;
        RECT 133.470 16.900 133.790 16.960 ;
        RECT 137.610 16.900 137.930 16.960 ;
        RECT 133.470 16.760 137.930 16.900 ;
        RECT 133.470 16.700 133.790 16.760 ;
        RECT 137.610 16.700 137.930 16.760 ;
      LAYER via ;
        RECT 137.640 1591.240 137.900 1591.500 ;
        RECT 396.160 1591.240 396.420 1591.500 ;
        RECT 133.500 16.700 133.760 16.960 ;
        RECT 137.640 16.700 137.900 16.960 ;
      LAYER met2 ;
        RECT 396.020 1600.380 396.300 1604.000 ;
        RECT 396.020 1600.000 396.360 1600.380 ;
        RECT 396.220 1591.530 396.360 1600.000 ;
        RECT 137.640 1591.210 137.900 1591.530 ;
        RECT 396.160 1591.210 396.420 1591.530 ;
        RECT 137.700 16.990 137.840 1591.210 ;
        RECT 133.500 16.670 133.760 16.990 ;
        RECT 137.640 16.670 137.900 16.990 ;
        RECT 133.560 2.400 133.700 16.670 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 19.960 151.730 20.020 ;
        RECT 401.650 19.960 401.970 20.020 ;
        RECT 151.410 19.820 401.970 19.960 ;
        RECT 151.410 19.760 151.730 19.820 ;
        RECT 401.650 19.760 401.970 19.820 ;
      LAYER via ;
        RECT 151.440 19.760 151.700 20.020 ;
        RECT 401.680 19.760 401.940 20.020 ;
      LAYER met2 ;
        RECT 402.460 1600.450 402.740 1604.000 ;
        RECT 401.740 1600.310 402.740 1600.450 ;
        RECT 401.740 20.050 401.880 1600.310 ;
        RECT 402.460 1600.000 402.740 1600.310 ;
        RECT 151.440 19.730 151.700 20.050 ;
        RECT 401.680 19.730 401.940 20.050 ;
        RECT 151.500 2.400 151.640 19.730 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 408.550 1592.460 408.870 1592.520 ;
        RECT 375.980 1592.320 408.870 1592.460 ;
        RECT 172.110 1592.120 172.430 1592.180 ;
        RECT 375.980 1592.120 376.120 1592.320 ;
        RECT 408.550 1592.260 408.870 1592.320 ;
        RECT 172.110 1591.980 376.120 1592.120 ;
        RECT 172.110 1591.920 172.430 1591.980 ;
        RECT 169.350 16.900 169.670 16.960 ;
        RECT 172.110 16.900 172.430 16.960 ;
        RECT 169.350 16.760 172.430 16.900 ;
        RECT 169.350 16.700 169.670 16.760 ;
        RECT 172.110 16.700 172.430 16.760 ;
      LAYER via ;
        RECT 172.140 1591.920 172.400 1592.180 ;
        RECT 408.580 1592.260 408.840 1592.520 ;
        RECT 169.380 16.700 169.640 16.960 ;
        RECT 172.140 16.700 172.400 16.960 ;
      LAYER met2 ;
        RECT 408.440 1600.380 408.720 1604.000 ;
        RECT 408.440 1600.000 408.780 1600.380 ;
        RECT 408.640 1592.550 408.780 1600.000 ;
        RECT 408.580 1592.230 408.840 1592.550 ;
        RECT 172.140 1591.890 172.400 1592.210 ;
        RECT 172.200 16.990 172.340 1591.890 ;
        RECT 169.380 16.670 169.640 16.990 ;
        RECT 172.140 16.670 172.400 16.990 ;
        RECT 169.440 2.400 169.580 16.670 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 226.925 15.045 227.095 16.915 ;
        RECT 276.145 14.025 276.315 16.915 ;
        RECT 323.985 14.025 324.155 16.915 ;
        RECT 375.965 16.065 376.135 17.255 ;
      LAYER mcon ;
        RECT 375.965 17.085 376.135 17.255 ;
        RECT 226.925 16.745 227.095 16.915 ;
        RECT 276.145 16.745 276.315 16.915 ;
        RECT 323.985 16.745 324.155 16.915 ;
      LAYER met1 ;
        RECT 375.905 17.240 376.195 17.285 ;
        RECT 358.040 17.100 376.195 17.240 ;
        RECT 226.865 16.900 227.155 16.945 ;
        RECT 276.085 16.900 276.375 16.945 ;
        RECT 226.865 16.760 276.375 16.900 ;
        RECT 226.865 16.715 227.155 16.760 ;
        RECT 276.085 16.715 276.375 16.760 ;
        RECT 323.925 16.900 324.215 16.945 ;
        RECT 358.040 16.900 358.180 17.100 ;
        RECT 375.905 17.055 376.195 17.100 ;
        RECT 323.925 16.760 358.180 16.900 ;
        RECT 323.925 16.715 324.215 16.760 ;
        RECT 375.905 16.220 376.195 16.265 ;
        RECT 414.990 16.220 415.310 16.280 ;
        RECT 375.905 16.080 415.310 16.220 ;
        RECT 375.905 16.035 376.195 16.080 ;
        RECT 414.990 16.020 415.310 16.080 ;
        RECT 186.830 15.200 187.150 15.260 ;
        RECT 226.865 15.200 227.155 15.245 ;
        RECT 186.830 15.060 227.155 15.200 ;
        RECT 186.830 15.000 187.150 15.060 ;
        RECT 226.865 15.015 227.155 15.060 ;
        RECT 276.085 14.180 276.375 14.225 ;
        RECT 323.925 14.180 324.215 14.225 ;
        RECT 276.085 14.040 324.215 14.180 ;
        RECT 276.085 13.995 276.375 14.040 ;
        RECT 323.925 13.995 324.215 14.040 ;
      LAYER via ;
        RECT 415.020 16.020 415.280 16.280 ;
        RECT 186.860 15.000 187.120 15.260 ;
      LAYER met2 ;
        RECT 414.420 1600.450 414.700 1604.000 ;
        RECT 414.420 1600.310 415.220 1600.450 ;
        RECT 414.420 1600.000 414.700 1600.310 ;
        RECT 415.080 16.310 415.220 1600.310 ;
        RECT 415.020 15.990 415.280 16.310 ;
        RECT 186.860 14.970 187.120 15.290 ;
        RECT 186.920 2.400 187.060 14.970 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 206.610 1592.800 206.930 1592.860 ;
        RECT 420.970 1592.800 421.290 1592.860 ;
        RECT 206.610 1592.660 421.290 1592.800 ;
        RECT 206.610 1592.600 206.930 1592.660 ;
        RECT 420.970 1592.600 421.290 1592.660 ;
      LAYER via ;
        RECT 206.640 1592.600 206.900 1592.860 ;
        RECT 421.000 1592.600 421.260 1592.860 ;
      LAYER met2 ;
        RECT 420.860 1600.380 421.140 1604.000 ;
        RECT 420.860 1600.000 421.200 1600.380 ;
        RECT 421.060 1592.890 421.200 1600.000 ;
        RECT 206.640 1592.570 206.900 1592.890 ;
        RECT 421.000 1592.570 421.260 1592.890 ;
        RECT 206.700 17.410 206.840 1592.570 ;
        RECT 204.860 17.270 206.840 17.410 ;
        RECT 204.860 2.400 205.000 17.270 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 311.565 13.685 311.735 15.555 ;
        RECT 323.525 13.685 323.695 16.235 ;
      LAYER mcon ;
        RECT 323.525 16.065 323.695 16.235 ;
        RECT 311.565 15.385 311.735 15.555 ;
      LAYER met1 ;
        RECT 423.270 1545.880 423.590 1545.940 ;
        RECT 425.570 1545.880 425.890 1545.940 ;
        RECT 423.270 1545.740 425.890 1545.880 ;
        RECT 423.270 1545.680 423.590 1545.740 ;
        RECT 425.570 1545.680 425.890 1545.740 ;
        RECT 422.350 1318.080 422.670 1318.140 ;
        RECT 423.270 1318.080 423.590 1318.140 ;
        RECT 422.350 1317.940 423.590 1318.080 ;
        RECT 422.350 1317.880 422.670 1317.940 ;
        RECT 423.270 1317.880 423.590 1317.940 ;
        RECT 422.350 1221.520 422.670 1221.580 ;
        RECT 423.270 1221.520 423.590 1221.580 ;
        RECT 422.350 1221.380 423.590 1221.520 ;
        RECT 422.350 1221.320 422.670 1221.380 ;
        RECT 423.270 1221.320 423.590 1221.380 ;
        RECT 422.350 1124.960 422.670 1125.020 ;
        RECT 423.270 1124.960 423.590 1125.020 ;
        RECT 422.350 1124.820 423.590 1124.960 ;
        RECT 422.350 1124.760 422.670 1124.820 ;
        RECT 423.270 1124.760 423.590 1124.820 ;
        RECT 422.350 1028.400 422.670 1028.460 ;
        RECT 423.270 1028.400 423.590 1028.460 ;
        RECT 422.350 1028.260 423.590 1028.400 ;
        RECT 422.350 1028.200 422.670 1028.260 ;
        RECT 423.270 1028.200 423.590 1028.260 ;
        RECT 422.350 931.840 422.670 931.900 ;
        RECT 423.270 931.840 423.590 931.900 ;
        RECT 422.350 931.700 423.590 931.840 ;
        RECT 422.350 931.640 422.670 931.700 ;
        RECT 423.270 931.640 423.590 931.700 ;
        RECT 422.350 835.280 422.670 835.340 ;
        RECT 423.270 835.280 423.590 835.340 ;
        RECT 422.350 835.140 423.590 835.280 ;
        RECT 422.350 835.080 422.670 835.140 ;
        RECT 423.270 835.080 423.590 835.140 ;
        RECT 422.350 738.380 422.670 738.440 ;
        RECT 423.270 738.380 423.590 738.440 ;
        RECT 422.350 738.240 423.590 738.380 ;
        RECT 422.350 738.180 422.670 738.240 ;
        RECT 423.270 738.180 423.590 738.240 ;
        RECT 422.350 641.820 422.670 641.880 ;
        RECT 423.270 641.820 423.590 641.880 ;
        RECT 422.350 641.680 423.590 641.820 ;
        RECT 422.350 641.620 422.670 641.680 ;
        RECT 423.270 641.620 423.590 641.680 ;
        RECT 422.350 545.260 422.670 545.320 ;
        RECT 423.270 545.260 423.590 545.320 ;
        RECT 422.350 545.120 423.590 545.260 ;
        RECT 422.350 545.060 422.670 545.120 ;
        RECT 423.270 545.060 423.590 545.120 ;
        RECT 422.350 448.700 422.670 448.760 ;
        RECT 423.270 448.700 423.590 448.760 ;
        RECT 422.350 448.560 423.590 448.700 ;
        RECT 422.350 448.500 422.670 448.560 ;
        RECT 423.270 448.500 423.590 448.560 ;
        RECT 422.810 331.400 423.130 331.460 ;
        RECT 423.270 331.400 423.590 331.460 ;
        RECT 422.810 331.260 423.590 331.400 ;
        RECT 422.810 331.200 423.130 331.260 ;
        RECT 423.270 331.200 423.590 331.260 ;
        RECT 422.810 241.640 423.130 241.700 ;
        RECT 423.270 241.640 423.590 241.700 ;
        RECT 422.810 241.500 423.590 241.640 ;
        RECT 422.810 241.440 423.130 241.500 ;
        RECT 423.270 241.440 423.590 241.500 ;
        RECT 423.270 145.420 423.590 145.480 ;
        RECT 422.900 145.280 423.590 145.420 ;
        RECT 422.900 145.140 423.040 145.280 ;
        RECT 423.270 145.220 423.590 145.280 ;
        RECT 422.810 144.880 423.130 145.140 ;
        RECT 422.350 16.560 422.670 16.620 ;
        RECT 358.960 16.420 422.670 16.560 ;
        RECT 323.465 16.220 323.755 16.265 ;
        RECT 358.960 16.220 359.100 16.420 ;
        RECT 422.350 16.360 422.670 16.420 ;
        RECT 323.465 16.080 359.100 16.220 ;
        RECT 323.465 16.035 323.755 16.080 ;
        RECT 222.710 15.880 223.030 15.940 ;
        RECT 222.710 15.740 228.920 15.880 ;
        RECT 222.710 15.680 223.030 15.740 ;
        RECT 228.780 15.540 228.920 15.740 ;
        RECT 311.505 15.540 311.795 15.585 ;
        RECT 228.780 15.400 311.795 15.540 ;
        RECT 311.505 15.355 311.795 15.400 ;
        RECT 311.505 13.840 311.795 13.885 ;
        RECT 323.465 13.840 323.755 13.885 ;
        RECT 311.505 13.700 323.755 13.840 ;
        RECT 311.505 13.655 311.795 13.700 ;
        RECT 323.465 13.655 323.755 13.700 ;
      LAYER via ;
        RECT 423.300 1545.680 423.560 1545.940 ;
        RECT 425.600 1545.680 425.860 1545.940 ;
        RECT 422.380 1317.880 422.640 1318.140 ;
        RECT 423.300 1317.880 423.560 1318.140 ;
        RECT 422.380 1221.320 422.640 1221.580 ;
        RECT 423.300 1221.320 423.560 1221.580 ;
        RECT 422.380 1124.760 422.640 1125.020 ;
        RECT 423.300 1124.760 423.560 1125.020 ;
        RECT 422.380 1028.200 422.640 1028.460 ;
        RECT 423.300 1028.200 423.560 1028.460 ;
        RECT 422.380 931.640 422.640 931.900 ;
        RECT 423.300 931.640 423.560 931.900 ;
        RECT 422.380 835.080 422.640 835.340 ;
        RECT 423.300 835.080 423.560 835.340 ;
        RECT 422.380 738.180 422.640 738.440 ;
        RECT 423.300 738.180 423.560 738.440 ;
        RECT 422.380 641.620 422.640 641.880 ;
        RECT 423.300 641.620 423.560 641.880 ;
        RECT 422.380 545.060 422.640 545.320 ;
        RECT 423.300 545.060 423.560 545.320 ;
        RECT 422.380 448.500 422.640 448.760 ;
        RECT 423.300 448.500 423.560 448.760 ;
        RECT 422.840 331.200 423.100 331.460 ;
        RECT 423.300 331.200 423.560 331.460 ;
        RECT 422.840 241.440 423.100 241.700 ;
        RECT 423.300 241.440 423.560 241.700 ;
        RECT 423.300 145.220 423.560 145.480 ;
        RECT 422.840 144.880 423.100 145.140 ;
        RECT 422.380 16.360 422.640 16.620 ;
        RECT 222.740 15.680 223.000 15.940 ;
      LAYER met2 ;
        RECT 426.840 1600.450 427.120 1604.000 ;
        RECT 425.660 1600.310 427.120 1600.450 ;
        RECT 425.660 1545.970 425.800 1600.310 ;
        RECT 426.840 1600.000 427.120 1600.310 ;
        RECT 423.300 1545.650 423.560 1545.970 ;
        RECT 425.600 1545.650 425.860 1545.970 ;
        RECT 423.360 1521.570 423.500 1545.650 ;
        RECT 422.900 1521.430 423.500 1521.570 ;
        RECT 422.900 1497.090 423.040 1521.430 ;
        RECT 422.900 1496.950 423.500 1497.090 ;
        RECT 423.360 1318.170 423.500 1496.950 ;
        RECT 422.380 1317.850 422.640 1318.170 ;
        RECT 423.300 1317.850 423.560 1318.170 ;
        RECT 422.440 1317.570 422.580 1317.850 ;
        RECT 422.440 1317.430 423.040 1317.570 ;
        RECT 422.900 1269.970 423.040 1317.430 ;
        RECT 422.900 1269.830 423.500 1269.970 ;
        RECT 423.360 1221.610 423.500 1269.830 ;
        RECT 422.380 1221.290 422.640 1221.610 ;
        RECT 423.300 1221.290 423.560 1221.610 ;
        RECT 422.440 1221.010 422.580 1221.290 ;
        RECT 422.440 1220.870 423.040 1221.010 ;
        RECT 422.900 1173.410 423.040 1220.870 ;
        RECT 422.900 1173.270 423.500 1173.410 ;
        RECT 423.360 1125.050 423.500 1173.270 ;
        RECT 422.380 1124.730 422.640 1125.050 ;
        RECT 423.300 1124.730 423.560 1125.050 ;
        RECT 422.440 1124.450 422.580 1124.730 ;
        RECT 422.440 1124.310 423.040 1124.450 ;
        RECT 422.900 1076.850 423.040 1124.310 ;
        RECT 422.900 1076.710 423.500 1076.850 ;
        RECT 423.360 1028.490 423.500 1076.710 ;
        RECT 422.380 1028.170 422.640 1028.490 ;
        RECT 423.300 1028.170 423.560 1028.490 ;
        RECT 422.440 1027.890 422.580 1028.170 ;
        RECT 422.440 1027.750 423.040 1027.890 ;
        RECT 422.900 980.290 423.040 1027.750 ;
        RECT 422.900 980.150 423.500 980.290 ;
        RECT 423.360 931.930 423.500 980.150 ;
        RECT 422.380 931.610 422.640 931.930 ;
        RECT 423.300 931.610 423.560 931.930 ;
        RECT 422.440 931.330 422.580 931.610 ;
        RECT 422.440 931.190 423.040 931.330 ;
        RECT 422.900 895.970 423.040 931.190 ;
        RECT 422.900 895.830 423.500 895.970 ;
        RECT 423.360 835.370 423.500 895.830 ;
        RECT 422.380 835.050 422.640 835.370 ;
        RECT 423.300 835.050 423.560 835.370 ;
        RECT 422.440 834.770 422.580 835.050 ;
        RECT 422.440 834.630 423.040 834.770 ;
        RECT 422.900 796.690 423.040 834.630 ;
        RECT 422.900 796.550 423.500 796.690 ;
        RECT 423.360 738.470 423.500 796.550 ;
        RECT 422.380 738.210 422.640 738.470 ;
        RECT 422.380 738.150 423.040 738.210 ;
        RECT 423.300 738.150 423.560 738.470 ;
        RECT 422.440 738.070 423.040 738.150 ;
        RECT 422.900 700.130 423.040 738.070 ;
        RECT 422.900 699.990 423.960 700.130 ;
        RECT 423.820 689.930 423.960 699.990 ;
        RECT 423.360 689.790 423.960 689.930 ;
        RECT 423.360 641.910 423.500 689.790 ;
        RECT 422.380 641.650 422.640 641.910 ;
        RECT 422.380 641.590 423.040 641.650 ;
        RECT 423.300 641.590 423.560 641.910 ;
        RECT 422.440 641.510 423.040 641.590 ;
        RECT 422.900 603.570 423.040 641.510 ;
        RECT 422.900 603.430 423.960 603.570 ;
        RECT 423.820 593.370 423.960 603.430 ;
        RECT 423.360 593.230 423.960 593.370 ;
        RECT 423.360 545.350 423.500 593.230 ;
        RECT 422.380 545.090 422.640 545.350 ;
        RECT 422.380 545.030 423.040 545.090 ;
        RECT 423.300 545.030 423.560 545.350 ;
        RECT 422.440 544.950 423.040 545.030 ;
        RECT 422.900 507.010 423.040 544.950 ;
        RECT 422.900 506.870 423.500 507.010 ;
        RECT 423.360 448.790 423.500 506.870 ;
        RECT 422.380 448.530 422.640 448.790 ;
        RECT 422.380 448.470 423.040 448.530 ;
        RECT 423.300 448.470 423.560 448.790 ;
        RECT 422.440 448.390 423.040 448.470 ;
        RECT 422.900 400.420 423.040 448.390 ;
        RECT 422.900 400.280 423.500 400.420 ;
        RECT 423.360 331.490 423.500 400.280 ;
        RECT 422.840 331.170 423.100 331.490 ;
        RECT 423.300 331.170 423.560 331.490 ;
        RECT 422.900 303.690 423.040 331.170 ;
        RECT 422.900 303.550 423.500 303.690 ;
        RECT 423.360 241.730 423.500 303.550 ;
        RECT 422.840 241.410 423.100 241.730 ;
        RECT 423.300 241.410 423.560 241.730 ;
        RECT 422.900 207.130 423.040 241.410 ;
        RECT 422.900 206.990 423.500 207.130 ;
        RECT 423.360 145.510 423.500 206.990 ;
        RECT 423.300 145.190 423.560 145.510 ;
        RECT 422.840 144.850 423.100 145.170 ;
        RECT 422.900 110.570 423.040 144.850 ;
        RECT 422.900 110.430 423.500 110.570 ;
        RECT 423.360 62.290 423.500 110.430 ;
        RECT 422.440 62.150 423.500 62.290 ;
        RECT 422.440 16.650 422.580 62.150 ;
        RECT 422.380 16.330 422.640 16.650 ;
        RECT 222.740 15.650 223.000 15.970 ;
        RECT 222.800 2.400 222.940 15.650 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 351.970 1579.880 352.290 1579.940 ;
        RECT 355.190 1579.880 355.510 1579.940 ;
        RECT 351.970 1579.740 355.510 1579.880 ;
        RECT 351.970 1579.680 352.290 1579.740 ;
        RECT 355.190 1579.680 355.510 1579.740 ;
        RECT 20.310 17.240 20.630 17.300 ;
        RECT 351.970 17.240 352.290 17.300 ;
        RECT 20.310 17.100 352.290 17.240 ;
        RECT 20.310 17.040 20.630 17.100 ;
        RECT 351.970 17.040 352.290 17.100 ;
      LAYER via ;
        RECT 352.000 1579.680 352.260 1579.940 ;
        RECT 355.220 1579.680 355.480 1579.940 ;
        RECT 20.340 17.040 20.600 17.300 ;
        RECT 352.000 17.040 352.260 17.300 ;
      LAYER met2 ;
        RECT 356.920 1600.450 357.200 1604.000 ;
        RECT 355.280 1600.310 357.200 1600.450 ;
        RECT 355.280 1579.970 355.420 1600.310 ;
        RECT 356.920 1600.000 357.200 1600.310 ;
        RECT 352.000 1579.650 352.260 1579.970 ;
        RECT 355.220 1579.650 355.480 1579.970 ;
        RECT 352.060 17.330 352.200 1579.650 ;
        RECT 20.340 17.010 20.600 17.330 ;
        RECT 352.000 17.010 352.260 17.330 ;
        RECT 20.400 2.400 20.540 17.010 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 359.330 1579.880 359.650 1579.940 ;
        RECT 363.470 1579.880 363.790 1579.940 ;
        RECT 359.330 1579.740 363.790 1579.880 ;
        RECT 359.330 1579.680 359.650 1579.740 ;
        RECT 363.470 1579.680 363.790 1579.740 ;
        RECT 44.230 17.920 44.550 17.980 ;
        RECT 358.870 17.920 359.190 17.980 ;
        RECT 44.230 17.780 359.190 17.920 ;
        RECT 44.230 17.720 44.550 17.780 ;
        RECT 358.870 17.720 359.190 17.780 ;
      LAYER via ;
        RECT 359.360 1579.680 359.620 1579.940 ;
        RECT 363.500 1579.680 363.760 1579.940 ;
        RECT 44.260 17.720 44.520 17.980 ;
        RECT 358.900 17.720 359.160 17.980 ;
      LAYER met2 ;
        RECT 365.200 1600.450 365.480 1604.000 ;
        RECT 363.560 1600.310 365.480 1600.450 ;
        RECT 363.560 1579.970 363.700 1600.310 ;
        RECT 365.200 1600.000 365.480 1600.310 ;
        RECT 359.360 1579.650 359.620 1579.970 ;
        RECT 363.500 1579.650 363.760 1579.970 ;
        RECT 359.420 20.130 359.560 1579.650 ;
        RECT 358.960 19.990 359.560 20.130 ;
        RECT 358.960 18.010 359.100 19.990 ;
        RECT 44.260 17.690 44.520 18.010 ;
        RECT 358.900 17.690 359.160 18.010 ;
        RECT 44.320 2.400 44.460 17.690 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 248.010 1593.820 248.330 1593.880 ;
        RECT 435.230 1593.820 435.550 1593.880 ;
        RECT 248.010 1593.680 435.550 1593.820 ;
        RECT 248.010 1593.620 248.330 1593.680 ;
        RECT 435.230 1593.620 435.550 1593.680 ;
      LAYER via ;
        RECT 248.040 1593.620 248.300 1593.880 ;
        RECT 435.260 1593.620 435.520 1593.880 ;
      LAYER met2 ;
        RECT 435.120 1600.380 435.400 1604.000 ;
        RECT 435.120 1600.000 435.460 1600.380 ;
        RECT 435.320 1593.910 435.460 1600.000 ;
        RECT 248.040 1593.590 248.300 1593.910 ;
        RECT 435.260 1593.590 435.520 1593.910 ;
        RECT 248.100 17.410 248.240 1593.590 ;
        RECT 246.720 17.270 248.240 17.410 ;
        RECT 246.720 2.400 246.860 17.270 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 348.290 1587.360 348.610 1587.420 ;
        RECT 441.670 1587.360 441.990 1587.420 ;
        RECT 348.290 1587.220 441.990 1587.360 ;
        RECT 348.290 1587.160 348.610 1587.220 ;
        RECT 441.670 1587.160 441.990 1587.220 ;
        RECT 264.110 14.520 264.430 14.580 ;
        RECT 346.910 14.520 347.230 14.580 ;
        RECT 264.110 14.380 347.230 14.520 ;
        RECT 264.110 14.320 264.430 14.380 ;
        RECT 346.910 14.320 347.230 14.380 ;
      LAYER via ;
        RECT 348.320 1587.160 348.580 1587.420 ;
        RECT 441.700 1587.160 441.960 1587.420 ;
        RECT 264.140 14.320 264.400 14.580 ;
        RECT 346.940 14.320 347.200 14.580 ;
      LAYER met2 ;
        RECT 441.560 1600.380 441.840 1604.000 ;
        RECT 441.560 1600.000 441.900 1600.380 ;
        RECT 441.760 1587.450 441.900 1600.000 ;
        RECT 348.320 1587.130 348.580 1587.450 ;
        RECT 441.700 1587.130 441.960 1587.450 ;
        RECT 348.380 15.370 348.520 1587.130 ;
        RECT 347.000 15.230 348.520 15.370 ;
        RECT 347.000 14.610 347.140 15.230 ;
        RECT 264.140 14.290 264.400 14.610 ;
        RECT 346.940 14.290 347.200 14.610 ;
        RECT 264.200 2.400 264.340 14.290 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 1589.400 282.370 1589.460 ;
        RECT 447.650 1589.400 447.970 1589.460 ;
        RECT 282.050 1589.260 447.970 1589.400 ;
        RECT 282.050 1589.200 282.370 1589.260 ;
        RECT 447.650 1589.200 447.970 1589.260 ;
      LAYER via ;
        RECT 282.080 1589.200 282.340 1589.460 ;
        RECT 447.680 1589.200 447.940 1589.460 ;
      LAYER met2 ;
        RECT 447.540 1600.380 447.820 1604.000 ;
        RECT 447.540 1600.000 447.880 1600.380 ;
        RECT 447.740 1589.490 447.880 1600.000 ;
        RECT 282.080 1589.170 282.340 1589.490 ;
        RECT 447.680 1589.170 447.940 1589.490 ;
        RECT 282.140 2.400 282.280 1589.170 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 450.025 1338.665 450.195 1366.715 ;
        RECT 450.025 386.325 450.195 434.435 ;
        RECT 450.025 290.105 450.195 337.875 ;
        RECT 450.025 96.645 450.195 144.755 ;
      LAYER mcon ;
        RECT 450.025 1366.545 450.195 1366.715 ;
        RECT 450.025 434.265 450.195 434.435 ;
        RECT 450.025 337.705 450.195 337.875 ;
        RECT 450.025 144.585 450.195 144.755 ;
      LAYER met1 ;
        RECT 449.950 1491.140 450.270 1491.200 ;
        RECT 450.870 1491.140 451.190 1491.200 ;
        RECT 449.950 1491.000 451.190 1491.140 ;
        RECT 449.950 1490.940 450.270 1491.000 ;
        RECT 450.870 1490.940 451.190 1491.000 ;
        RECT 450.410 1435.380 450.730 1435.440 ;
        RECT 451.330 1435.380 451.650 1435.440 ;
        RECT 450.410 1435.240 451.650 1435.380 ;
        RECT 450.410 1435.180 450.730 1435.240 ;
        RECT 451.330 1435.180 451.650 1435.240 ;
        RECT 449.965 1366.700 450.255 1366.745 ;
        RECT 450.410 1366.700 450.730 1366.760 ;
        RECT 449.965 1366.560 450.730 1366.700 ;
        RECT 449.965 1366.515 450.255 1366.560 ;
        RECT 450.410 1366.500 450.730 1366.560 ;
        RECT 449.950 1338.820 450.270 1338.880 ;
        RECT 449.755 1338.680 450.270 1338.820 ;
        RECT 449.950 1338.620 450.270 1338.680 ;
        RECT 449.950 1304.140 450.270 1304.200 ;
        RECT 450.410 1304.140 450.730 1304.200 ;
        RECT 449.950 1304.000 450.730 1304.140 ;
        RECT 449.950 1303.940 450.270 1304.000 ;
        RECT 450.410 1303.940 450.730 1304.000 ;
        RECT 449.950 1269.600 450.270 1269.860 ;
        RECT 450.040 1269.120 450.180 1269.600 ;
        RECT 450.410 1269.120 450.730 1269.180 ;
        RECT 450.040 1268.980 450.730 1269.120 ;
        RECT 450.410 1268.920 450.730 1268.980 ;
        RECT 449.950 1152.500 450.270 1152.560 ;
        RECT 450.870 1152.500 451.190 1152.560 ;
        RECT 449.950 1152.360 451.190 1152.500 ;
        RECT 449.950 1152.300 450.270 1152.360 ;
        RECT 450.870 1152.300 451.190 1152.360 ;
        RECT 449.950 1028.200 450.270 1028.460 ;
        RECT 450.040 1027.720 450.180 1028.200 ;
        RECT 450.410 1027.720 450.730 1027.780 ;
        RECT 450.040 1027.580 450.730 1027.720 ;
        RECT 450.410 1027.520 450.730 1027.580 ;
        RECT 449.950 869.960 450.270 870.020 ;
        RECT 450.870 869.960 451.190 870.020 ;
        RECT 449.950 869.820 451.190 869.960 ;
        RECT 449.950 869.760 450.270 869.820 ;
        RECT 450.870 869.760 451.190 869.820 ;
        RECT 449.950 787.140 450.270 787.400 ;
        RECT 450.040 786.720 450.180 787.140 ;
        RECT 449.950 786.460 450.270 786.720 ;
        RECT 450.410 627.880 450.730 627.940 ;
        RECT 450.870 627.880 451.190 627.940 ;
        RECT 450.410 627.740 451.190 627.880 ;
        RECT 450.410 627.680 450.730 627.740 ;
        RECT 450.870 627.680 451.190 627.740 ;
        RECT 449.950 579.600 450.270 579.660 ;
        RECT 450.870 579.600 451.190 579.660 ;
        RECT 449.950 579.460 451.190 579.600 ;
        RECT 449.950 579.400 450.270 579.460 ;
        RECT 450.870 579.400 451.190 579.460 ;
        RECT 449.950 434.420 450.270 434.480 ;
        RECT 449.755 434.280 450.270 434.420 ;
        RECT 449.950 434.220 450.270 434.280 ;
        RECT 449.950 386.480 450.270 386.540 ;
        RECT 449.755 386.340 450.270 386.480 ;
        RECT 449.950 386.280 450.270 386.340 ;
        RECT 449.950 337.860 450.270 337.920 ;
        RECT 449.755 337.720 450.270 337.860 ;
        RECT 449.950 337.660 450.270 337.720 ;
        RECT 449.950 290.260 450.270 290.320 ;
        RECT 449.755 290.120 450.270 290.260 ;
        RECT 449.950 290.060 450.270 290.120 ;
        RECT 449.950 206.420 450.270 206.680 ;
        RECT 450.040 206.000 450.180 206.420 ;
        RECT 449.950 205.740 450.270 206.000 ;
        RECT 449.950 144.740 450.270 144.800 ;
        RECT 449.755 144.600 450.270 144.740 ;
        RECT 449.950 144.540 450.270 144.600 ;
        RECT 449.950 96.800 450.270 96.860 ;
        RECT 449.755 96.660 450.270 96.800 ;
        RECT 449.950 96.600 450.270 96.660 ;
        RECT 449.950 15.200 450.270 15.260 ;
        RECT 324.460 15.060 450.270 15.200 ;
        RECT 299.990 14.860 300.310 14.920 ;
        RECT 324.460 14.860 324.600 15.060 ;
        RECT 449.950 15.000 450.270 15.060 ;
        RECT 299.990 14.720 324.600 14.860 ;
        RECT 299.990 14.660 300.310 14.720 ;
      LAYER via ;
        RECT 449.980 1490.940 450.240 1491.200 ;
        RECT 450.900 1490.940 451.160 1491.200 ;
        RECT 450.440 1435.180 450.700 1435.440 ;
        RECT 451.360 1435.180 451.620 1435.440 ;
        RECT 450.440 1366.500 450.700 1366.760 ;
        RECT 449.980 1338.620 450.240 1338.880 ;
        RECT 449.980 1303.940 450.240 1304.200 ;
        RECT 450.440 1303.940 450.700 1304.200 ;
        RECT 449.980 1269.600 450.240 1269.860 ;
        RECT 450.440 1268.920 450.700 1269.180 ;
        RECT 449.980 1152.300 450.240 1152.560 ;
        RECT 450.900 1152.300 451.160 1152.560 ;
        RECT 449.980 1028.200 450.240 1028.460 ;
        RECT 450.440 1027.520 450.700 1027.780 ;
        RECT 449.980 869.760 450.240 870.020 ;
        RECT 450.900 869.760 451.160 870.020 ;
        RECT 449.980 787.140 450.240 787.400 ;
        RECT 449.980 786.460 450.240 786.720 ;
        RECT 450.440 627.680 450.700 627.940 ;
        RECT 450.900 627.680 451.160 627.940 ;
        RECT 449.980 579.400 450.240 579.660 ;
        RECT 450.900 579.400 451.160 579.660 ;
        RECT 449.980 434.220 450.240 434.480 ;
        RECT 449.980 386.280 450.240 386.540 ;
        RECT 449.980 337.660 450.240 337.920 ;
        RECT 449.980 290.060 450.240 290.320 ;
        RECT 449.980 206.420 450.240 206.680 ;
        RECT 449.980 205.740 450.240 206.000 ;
        RECT 449.980 144.540 450.240 144.800 ;
        RECT 449.980 96.600 450.240 96.860 ;
        RECT 300.020 14.660 300.280 14.920 ;
        RECT 449.980 15.000 450.240 15.260 ;
      LAYER met2 ;
        RECT 453.980 1601.130 454.260 1604.000 ;
        RECT 452.340 1600.990 454.260 1601.130 ;
        RECT 452.340 1539.365 452.480 1600.990 ;
        RECT 453.980 1600.000 454.260 1600.990 ;
        RECT 452.270 1538.995 452.550 1539.365 ;
        RECT 450.890 1538.315 451.170 1538.685 ;
        RECT 450.960 1491.230 451.100 1538.315 ;
        RECT 449.980 1490.910 450.240 1491.230 ;
        RECT 450.900 1490.910 451.160 1491.230 ;
        RECT 450.040 1483.605 450.180 1490.910 ;
        RECT 449.970 1483.235 450.250 1483.605 ;
        RECT 451.350 1483.235 451.630 1483.605 ;
        RECT 451.420 1435.470 451.560 1483.235 ;
        RECT 450.440 1435.150 450.700 1435.470 ;
        RECT 451.360 1435.150 451.620 1435.470 ;
        RECT 450.500 1366.790 450.640 1435.150 ;
        RECT 450.440 1366.470 450.700 1366.790 ;
        RECT 449.980 1338.590 450.240 1338.910 ;
        RECT 450.040 1328.450 450.180 1338.590 ;
        RECT 450.040 1328.310 450.640 1328.450 ;
        RECT 450.500 1304.230 450.640 1328.310 ;
        RECT 449.980 1303.910 450.240 1304.230 ;
        RECT 450.440 1303.910 450.700 1304.230 ;
        RECT 450.040 1269.890 450.180 1303.910 ;
        RECT 449.980 1269.570 450.240 1269.890 ;
        RECT 450.440 1268.890 450.700 1269.210 ;
        RECT 450.500 1207.410 450.640 1268.890 ;
        RECT 450.040 1207.270 450.640 1207.410 ;
        RECT 450.040 1200.725 450.180 1207.270 ;
        RECT 449.970 1200.355 450.250 1200.725 ;
        RECT 450.890 1200.355 451.170 1200.725 ;
        RECT 450.960 1152.590 451.100 1200.355 ;
        RECT 449.980 1152.270 450.240 1152.590 ;
        RECT 450.900 1152.270 451.160 1152.590 ;
        RECT 450.040 1135.330 450.180 1152.270 ;
        RECT 450.040 1135.190 451.100 1135.330 ;
        RECT 450.960 1124.450 451.100 1135.190 ;
        RECT 450.500 1124.310 451.100 1124.450 ;
        RECT 450.500 1087.050 450.640 1124.310 ;
        RECT 450.040 1086.910 450.640 1087.050 ;
        RECT 450.040 1028.490 450.180 1086.910 ;
        RECT 449.980 1028.170 450.240 1028.490 ;
        RECT 450.440 1027.490 450.700 1027.810 ;
        RECT 450.500 990.490 450.640 1027.490 ;
        RECT 450.040 990.350 450.640 990.490 ;
        RECT 450.040 966.125 450.180 990.350 ;
        RECT 449.970 965.755 450.250 966.125 ;
        RECT 450.890 965.755 451.170 966.125 ;
        RECT 450.960 870.050 451.100 965.755 ;
        RECT 449.980 869.730 450.240 870.050 ;
        RECT 450.900 869.730 451.160 870.050 ;
        RECT 450.040 787.430 450.180 869.730 ;
        RECT 449.980 787.110 450.240 787.430 ;
        RECT 449.980 786.430 450.240 786.750 ;
        RECT 450.040 677.125 450.180 786.430 ;
        RECT 449.970 676.755 450.250 677.125 ;
        RECT 449.970 676.075 450.250 676.445 ;
        RECT 450.040 628.050 450.180 676.075 ;
        RECT 450.040 627.970 450.640 628.050 ;
        RECT 450.040 627.910 450.700 627.970 ;
        RECT 450.440 627.650 450.700 627.910 ;
        RECT 450.900 627.650 451.160 627.970 ;
        RECT 450.960 579.885 451.100 627.650 ;
        RECT 449.970 579.515 450.250 579.885 ;
        RECT 450.890 579.515 451.170 579.885 ;
        RECT 449.980 579.370 450.240 579.515 ;
        RECT 450.900 579.370 451.160 579.515 ;
        RECT 450.960 483.325 451.100 579.370 ;
        RECT 449.970 482.955 450.250 483.325 ;
        RECT 450.890 482.955 451.170 483.325 ;
        RECT 450.040 434.510 450.180 482.955 ;
        RECT 449.980 434.190 450.240 434.510 ;
        RECT 449.980 386.250 450.240 386.570 ;
        RECT 450.040 337.950 450.180 386.250 ;
        RECT 449.980 337.630 450.240 337.950 ;
        RECT 449.980 290.030 450.240 290.350 ;
        RECT 450.040 206.710 450.180 290.030 ;
        RECT 449.980 206.390 450.240 206.710 ;
        RECT 449.980 205.710 450.240 206.030 ;
        RECT 450.040 144.830 450.180 205.710 ;
        RECT 449.980 144.510 450.240 144.830 ;
        RECT 449.980 96.570 450.240 96.890 ;
        RECT 450.040 15.290 450.180 96.570 ;
        RECT 449.980 14.970 450.240 15.290 ;
        RECT 300.020 14.630 300.280 14.950 ;
        RECT 300.080 2.400 300.220 14.630 ;
        RECT 299.870 -4.800 300.430 2.400 ;
      LAYER via2 ;
        RECT 452.270 1539.040 452.550 1539.320 ;
        RECT 450.890 1538.360 451.170 1538.640 ;
        RECT 449.970 1483.280 450.250 1483.560 ;
        RECT 451.350 1483.280 451.630 1483.560 ;
        RECT 449.970 1200.400 450.250 1200.680 ;
        RECT 450.890 1200.400 451.170 1200.680 ;
        RECT 449.970 965.800 450.250 966.080 ;
        RECT 450.890 965.800 451.170 966.080 ;
        RECT 449.970 676.800 450.250 677.080 ;
        RECT 449.970 676.120 450.250 676.400 ;
        RECT 449.970 579.560 450.250 579.840 ;
        RECT 450.890 579.560 451.170 579.840 ;
        RECT 449.970 483.000 450.250 483.280 ;
        RECT 450.890 483.000 451.170 483.280 ;
      LAYER met3 ;
        RECT 452.245 1539.330 452.575 1539.345 ;
        RECT 451.110 1539.030 452.575 1539.330 ;
        RECT 451.110 1538.665 451.410 1539.030 ;
        RECT 452.245 1539.015 452.575 1539.030 ;
        RECT 450.865 1538.350 451.410 1538.665 ;
        RECT 450.865 1538.335 451.195 1538.350 ;
        RECT 449.945 1483.570 450.275 1483.585 ;
        RECT 451.325 1483.570 451.655 1483.585 ;
        RECT 449.945 1483.270 451.655 1483.570 ;
        RECT 449.945 1483.255 450.275 1483.270 ;
        RECT 451.325 1483.255 451.655 1483.270 ;
        RECT 449.945 1200.690 450.275 1200.705 ;
        RECT 450.865 1200.690 451.195 1200.705 ;
        RECT 449.945 1200.390 451.195 1200.690 ;
        RECT 449.945 1200.375 450.275 1200.390 ;
        RECT 450.865 1200.375 451.195 1200.390 ;
        RECT 449.945 966.090 450.275 966.105 ;
        RECT 450.865 966.090 451.195 966.105 ;
        RECT 449.945 965.790 451.195 966.090 ;
        RECT 449.945 965.775 450.275 965.790 ;
        RECT 450.865 965.775 451.195 965.790 ;
        RECT 449.945 677.090 450.275 677.105 ;
        RECT 449.945 676.775 450.490 677.090 ;
        RECT 450.190 676.425 450.490 676.775 ;
        RECT 449.945 676.110 450.490 676.425 ;
        RECT 449.945 676.095 450.275 676.110 ;
        RECT 449.945 579.850 450.275 579.865 ;
        RECT 450.865 579.850 451.195 579.865 ;
        RECT 449.945 579.550 451.195 579.850 ;
        RECT 449.945 579.535 450.275 579.550 ;
        RECT 450.865 579.535 451.195 579.550 ;
        RECT 449.945 483.290 450.275 483.305 ;
        RECT 450.865 483.290 451.195 483.305 ;
        RECT 449.945 482.990 451.195 483.290 ;
        RECT 449.945 482.975 450.275 482.990 ;
        RECT 450.865 482.975 451.195 482.990 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.450 1587.700 323.770 1587.760 ;
        RECT 460.070 1587.700 460.390 1587.760 ;
        RECT 323.450 1587.560 460.390 1587.700 ;
        RECT 323.450 1587.500 323.770 1587.560 ;
        RECT 460.070 1587.500 460.390 1587.560 ;
        RECT 317.930 15.200 318.250 15.260 ;
        RECT 323.450 15.200 323.770 15.260 ;
        RECT 317.930 15.060 323.770 15.200 ;
        RECT 317.930 15.000 318.250 15.060 ;
        RECT 323.450 15.000 323.770 15.060 ;
      LAYER via ;
        RECT 323.480 1587.500 323.740 1587.760 ;
        RECT 460.100 1587.500 460.360 1587.760 ;
        RECT 317.960 15.000 318.220 15.260 ;
        RECT 323.480 15.000 323.740 15.260 ;
      LAYER met2 ;
        RECT 459.960 1600.380 460.240 1604.000 ;
        RECT 459.960 1600.000 460.300 1600.380 ;
        RECT 460.160 1587.790 460.300 1600.000 ;
        RECT 323.480 1587.470 323.740 1587.790 ;
        RECT 460.100 1587.470 460.360 1587.790 ;
        RECT 323.540 15.290 323.680 1587.470 ;
        RECT 317.960 14.970 318.220 15.290 ;
        RECT 323.480 14.970 323.740 15.290 ;
        RECT 318.020 2.400 318.160 14.970 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 464.285 1538.925 464.455 1587.035 ;
        RECT 463.825 386.325 463.995 434.435 ;
        RECT 463.825 290.105 463.995 337.875 ;
      LAYER mcon ;
        RECT 464.285 1586.865 464.455 1587.035 ;
        RECT 463.825 434.265 463.995 434.435 ;
        RECT 463.825 337.705 463.995 337.875 ;
      LAYER met1 ;
        RECT 464.225 1587.020 464.515 1587.065 ;
        RECT 465.130 1587.020 465.450 1587.080 ;
        RECT 464.225 1586.880 465.450 1587.020 ;
        RECT 464.225 1586.835 464.515 1586.880 ;
        RECT 465.130 1586.820 465.450 1586.880 ;
        RECT 464.210 1539.080 464.530 1539.140 ;
        RECT 464.015 1538.940 464.530 1539.080 ;
        RECT 464.210 1538.880 464.530 1538.940 ;
        RECT 464.210 1497.740 464.530 1498.000 ;
        RECT 464.300 1497.320 464.440 1497.740 ;
        RECT 464.210 1497.060 464.530 1497.320 ;
        RECT 463.750 1345.620 464.070 1345.680 ;
        RECT 464.210 1345.620 464.530 1345.680 ;
        RECT 463.750 1345.480 464.530 1345.620 ;
        RECT 463.750 1345.420 464.070 1345.480 ;
        RECT 464.210 1345.420 464.530 1345.480 ;
        RECT 463.750 1304.280 464.070 1304.540 ;
        RECT 463.840 1303.800 463.980 1304.280 ;
        RECT 464.210 1303.800 464.530 1303.860 ;
        RECT 463.840 1303.660 464.530 1303.800 ;
        RECT 464.210 1303.600 464.530 1303.660 ;
        RECT 463.290 1249.060 463.610 1249.120 ;
        RECT 464.210 1249.060 464.530 1249.120 ;
        RECT 463.290 1248.920 464.530 1249.060 ;
        RECT 463.290 1248.860 463.610 1248.920 ;
        RECT 464.210 1248.860 464.530 1248.920 ;
        RECT 463.750 966.520 464.070 966.580 ;
        RECT 464.670 966.520 464.990 966.580 ;
        RECT 463.750 966.380 464.990 966.520 ;
        RECT 463.750 966.320 464.070 966.380 ;
        RECT 464.670 966.320 464.990 966.380 ;
        RECT 464.210 627.880 464.530 627.940 ;
        RECT 464.670 627.880 464.990 627.940 ;
        RECT 464.210 627.740 464.990 627.880 ;
        RECT 464.210 627.680 464.530 627.740 ;
        RECT 464.670 627.680 464.990 627.740 ;
        RECT 463.750 579.600 464.070 579.660 ;
        RECT 464.670 579.600 464.990 579.660 ;
        RECT 463.750 579.460 464.990 579.600 ;
        RECT 463.750 579.400 464.070 579.460 ;
        RECT 464.670 579.400 464.990 579.460 ;
        RECT 463.750 434.420 464.070 434.480 ;
        RECT 463.555 434.280 464.070 434.420 ;
        RECT 463.750 434.220 464.070 434.280 ;
        RECT 463.750 386.480 464.070 386.540 ;
        RECT 463.555 386.340 464.070 386.480 ;
        RECT 463.750 386.280 464.070 386.340 ;
        RECT 463.750 337.860 464.070 337.920 ;
        RECT 463.555 337.720 464.070 337.860 ;
        RECT 463.750 337.660 464.070 337.720 ;
        RECT 463.750 290.260 464.070 290.320 ;
        RECT 463.555 290.120 464.070 290.260 ;
        RECT 463.750 290.060 464.070 290.120 ;
        RECT 463.750 241.440 464.070 241.700 ;
        RECT 463.840 240.960 463.980 241.440 ;
        RECT 464.210 240.960 464.530 241.020 ;
        RECT 463.840 240.820 464.530 240.960 ;
        RECT 464.210 240.760 464.530 240.820 ;
        RECT 464.210 138.620 464.530 138.680 ;
        RECT 463.840 138.480 464.530 138.620 ;
        RECT 463.840 138.340 463.980 138.480 ;
        RECT 464.210 138.420 464.530 138.480 ;
        RECT 463.750 138.080 464.070 138.340 ;
        RECT 335.870 14.860 336.190 14.920 ;
        RECT 463.750 14.860 464.070 14.920 ;
        RECT 335.870 14.720 464.070 14.860 ;
        RECT 335.870 14.660 336.190 14.720 ;
        RECT 463.750 14.660 464.070 14.720 ;
      LAYER via ;
        RECT 465.160 1586.820 465.420 1587.080 ;
        RECT 464.240 1538.880 464.500 1539.140 ;
        RECT 464.240 1497.740 464.500 1498.000 ;
        RECT 464.240 1497.060 464.500 1497.320 ;
        RECT 463.780 1345.420 464.040 1345.680 ;
        RECT 464.240 1345.420 464.500 1345.680 ;
        RECT 463.780 1304.280 464.040 1304.540 ;
        RECT 464.240 1303.600 464.500 1303.860 ;
        RECT 463.320 1248.860 463.580 1249.120 ;
        RECT 464.240 1248.860 464.500 1249.120 ;
        RECT 463.780 966.320 464.040 966.580 ;
        RECT 464.700 966.320 464.960 966.580 ;
        RECT 464.240 627.680 464.500 627.940 ;
        RECT 464.700 627.680 464.960 627.940 ;
        RECT 463.780 579.400 464.040 579.660 ;
        RECT 464.700 579.400 464.960 579.660 ;
        RECT 463.780 434.220 464.040 434.480 ;
        RECT 463.780 386.280 464.040 386.540 ;
        RECT 463.780 337.660 464.040 337.920 ;
        RECT 463.780 290.060 464.040 290.320 ;
        RECT 463.780 241.440 464.040 241.700 ;
        RECT 464.240 240.760 464.500 241.020 ;
        RECT 464.240 138.420 464.500 138.680 ;
        RECT 463.780 138.080 464.040 138.340 ;
        RECT 335.900 14.660 336.160 14.920 ;
        RECT 463.780 14.660 464.040 14.920 ;
      LAYER met2 ;
        RECT 465.940 1600.450 466.220 1604.000 ;
        RECT 465.220 1600.310 466.220 1600.450 ;
        RECT 465.220 1587.110 465.360 1600.310 ;
        RECT 465.940 1600.000 466.220 1600.310 ;
        RECT 465.160 1586.790 465.420 1587.110 ;
        RECT 464.240 1538.850 464.500 1539.170 ;
        RECT 464.300 1498.030 464.440 1538.850 ;
        RECT 464.240 1497.710 464.500 1498.030 ;
        RECT 464.240 1497.030 464.500 1497.350 ;
        RECT 464.300 1345.710 464.440 1497.030 ;
        RECT 463.780 1345.390 464.040 1345.710 ;
        RECT 464.240 1345.390 464.500 1345.710 ;
        RECT 463.840 1304.570 463.980 1345.390 ;
        RECT 463.780 1304.250 464.040 1304.570 ;
        RECT 464.240 1303.570 464.500 1303.890 ;
        RECT 464.300 1297.170 464.440 1303.570 ;
        RECT 463.380 1297.030 464.440 1297.170 ;
        RECT 463.380 1249.150 463.520 1297.030 ;
        RECT 463.320 1248.830 463.580 1249.150 ;
        RECT 464.240 1248.830 464.500 1249.150 ;
        RECT 464.300 1183.610 464.440 1248.830 ;
        RECT 463.840 1183.470 464.440 1183.610 ;
        RECT 463.840 1135.330 463.980 1183.470 ;
        RECT 463.840 1135.190 464.900 1135.330 ;
        RECT 464.760 1124.450 464.900 1135.190 ;
        RECT 464.300 1124.310 464.900 1124.450 ;
        RECT 464.300 1087.050 464.440 1124.310 ;
        RECT 463.840 1086.910 464.440 1087.050 ;
        RECT 463.840 1062.685 463.980 1086.910 ;
        RECT 463.770 1062.315 464.050 1062.685 ;
        RECT 464.690 1062.315 464.970 1062.685 ;
        RECT 464.760 966.610 464.900 1062.315 ;
        RECT 463.780 966.290 464.040 966.610 ;
        RECT 464.700 966.290 464.960 966.610 ;
        RECT 463.840 787.170 463.980 966.290 ;
        RECT 463.840 787.030 464.440 787.170 ;
        RECT 464.300 786.660 464.440 787.030 ;
        RECT 463.840 786.520 464.440 786.660 ;
        RECT 463.840 677.125 463.980 786.520 ;
        RECT 463.770 676.755 464.050 677.125 ;
        RECT 463.770 676.075 464.050 676.445 ;
        RECT 463.840 628.050 463.980 676.075 ;
        RECT 463.840 627.970 464.440 628.050 ;
        RECT 463.840 627.910 464.500 627.970 ;
        RECT 464.240 627.650 464.500 627.910 ;
        RECT 464.700 627.650 464.960 627.970 ;
        RECT 464.760 579.885 464.900 627.650 ;
        RECT 463.770 579.515 464.050 579.885 ;
        RECT 464.690 579.515 464.970 579.885 ;
        RECT 463.780 579.370 464.040 579.515 ;
        RECT 464.700 579.370 464.960 579.515 ;
        RECT 464.760 483.325 464.900 579.370 ;
        RECT 463.770 482.955 464.050 483.325 ;
        RECT 464.690 482.955 464.970 483.325 ;
        RECT 463.840 434.510 463.980 482.955 ;
        RECT 463.780 434.190 464.040 434.510 ;
        RECT 463.780 386.250 464.040 386.570 ;
        RECT 463.840 337.950 463.980 386.250 ;
        RECT 463.780 337.630 464.040 337.950 ;
        RECT 463.780 290.030 464.040 290.350 ;
        RECT 463.840 241.730 463.980 290.030 ;
        RECT 463.780 241.410 464.040 241.730 ;
        RECT 464.240 240.730 464.500 241.050 ;
        RECT 464.300 138.710 464.440 240.730 ;
        RECT 464.240 138.390 464.500 138.710 ;
        RECT 463.780 138.050 464.040 138.370 ;
        RECT 463.840 14.950 463.980 138.050 ;
        RECT 335.900 14.630 336.160 14.950 ;
        RECT 463.780 14.630 464.040 14.950 ;
        RECT 335.960 2.400 336.100 14.630 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 463.770 1062.360 464.050 1062.640 ;
        RECT 464.690 1062.360 464.970 1062.640 ;
        RECT 463.770 676.800 464.050 677.080 ;
        RECT 463.770 676.120 464.050 676.400 ;
        RECT 463.770 579.560 464.050 579.840 ;
        RECT 464.690 579.560 464.970 579.840 ;
        RECT 463.770 483.000 464.050 483.280 ;
        RECT 464.690 483.000 464.970 483.280 ;
      LAYER met3 ;
        RECT 463.745 1062.650 464.075 1062.665 ;
        RECT 464.665 1062.650 464.995 1062.665 ;
        RECT 463.745 1062.350 464.995 1062.650 ;
        RECT 463.745 1062.335 464.075 1062.350 ;
        RECT 464.665 1062.335 464.995 1062.350 ;
        RECT 463.745 677.090 464.075 677.105 ;
        RECT 463.745 676.775 464.290 677.090 ;
        RECT 463.990 676.425 464.290 676.775 ;
        RECT 463.745 676.110 464.290 676.425 ;
        RECT 463.745 676.095 464.075 676.110 ;
        RECT 463.745 579.850 464.075 579.865 ;
        RECT 464.665 579.850 464.995 579.865 ;
        RECT 463.745 579.550 464.995 579.850 ;
        RECT 463.745 579.535 464.075 579.550 ;
        RECT 464.665 579.535 464.995 579.550 ;
        RECT 463.745 483.290 464.075 483.305 ;
        RECT 464.665 483.290 464.995 483.305 ;
        RECT 463.745 482.990 464.995 483.290 ;
        RECT 463.745 482.975 464.075 482.990 ;
        RECT 464.665 482.975 464.995 482.990 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 368.605 4.845 368.775 18.615 ;
        RECT 399.425 17.255 399.595 18.615 ;
        RECT 399.425 17.085 400.055 17.255 ;
      LAYER mcon ;
        RECT 368.605 18.445 368.775 18.615 ;
        RECT 399.425 18.445 399.595 18.615 ;
        RECT 399.885 17.085 400.055 17.255 ;
      LAYER met1 ;
        RECT 469.270 1579.880 469.590 1579.940 ;
        RECT 471.110 1579.880 471.430 1579.940 ;
        RECT 469.270 1579.740 471.430 1579.880 ;
        RECT 469.270 1579.680 469.590 1579.740 ;
        RECT 471.110 1579.680 471.430 1579.740 ;
        RECT 469.270 385.940 469.590 386.200 ;
        RECT 469.360 385.180 469.500 385.940 ;
        RECT 469.270 384.920 469.590 385.180 ;
        RECT 368.545 18.600 368.835 18.645 ;
        RECT 399.365 18.600 399.655 18.645 ;
        RECT 368.545 18.460 399.655 18.600 ;
        RECT 368.545 18.415 368.835 18.460 ;
        RECT 399.365 18.415 399.655 18.460 ;
        RECT 399.825 17.240 400.115 17.285 ;
        RECT 469.270 17.240 469.590 17.300 ;
        RECT 399.825 17.100 469.590 17.240 ;
        RECT 399.825 17.055 400.115 17.100 ;
        RECT 469.270 17.040 469.590 17.100 ;
        RECT 353.350 5.000 353.670 5.060 ;
        RECT 368.545 5.000 368.835 5.045 ;
        RECT 353.350 4.860 368.835 5.000 ;
        RECT 353.350 4.800 353.670 4.860 ;
        RECT 368.545 4.815 368.835 4.860 ;
      LAYER via ;
        RECT 469.300 1579.680 469.560 1579.940 ;
        RECT 471.140 1579.680 471.400 1579.940 ;
        RECT 469.300 385.940 469.560 386.200 ;
        RECT 469.300 384.920 469.560 385.180 ;
        RECT 469.300 17.040 469.560 17.300 ;
        RECT 353.380 4.800 353.640 5.060 ;
      LAYER met2 ;
        RECT 472.380 1600.450 472.660 1604.000 ;
        RECT 471.200 1600.310 472.660 1600.450 ;
        RECT 471.200 1579.970 471.340 1600.310 ;
        RECT 472.380 1600.000 472.660 1600.310 ;
        RECT 469.300 1579.650 469.560 1579.970 ;
        RECT 471.140 1579.650 471.400 1579.970 ;
        RECT 469.360 386.230 469.500 1579.650 ;
        RECT 469.300 385.910 469.560 386.230 ;
        RECT 469.300 384.890 469.560 385.210 ;
        RECT 469.360 17.330 469.500 384.890 ;
        RECT 469.300 17.010 469.560 17.330 ;
        RECT 353.380 4.770 353.640 5.090 ;
        RECT 353.440 2.400 353.580 4.770 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 371.290 17.920 371.610 17.980 ;
        RECT 477.090 17.920 477.410 17.980 ;
        RECT 371.290 17.780 477.410 17.920 ;
        RECT 371.290 17.720 371.610 17.780 ;
        RECT 477.090 17.720 477.410 17.780 ;
      LAYER via ;
        RECT 371.320 17.720 371.580 17.980 ;
        RECT 477.120 17.720 477.380 17.980 ;
      LAYER met2 ;
        RECT 478.360 1600.450 478.640 1604.000 ;
        RECT 477.180 1600.310 478.640 1600.450 ;
        RECT 477.180 18.010 477.320 1600.310 ;
        RECT 478.360 1600.000 478.640 1600.310 ;
        RECT 371.320 17.690 371.580 18.010 ;
        RECT 477.120 17.690 477.380 18.010 ;
        RECT 371.380 2.400 371.520 17.690 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 458.305 18.785 458.475 20.315 ;
      LAYER mcon ;
        RECT 458.305 20.145 458.475 20.315 ;
      LAYER met1 ;
        RECT 458.245 20.300 458.535 20.345 ;
        RECT 483.530 20.300 483.850 20.360 ;
        RECT 458.245 20.160 483.850 20.300 ;
        RECT 458.245 20.115 458.535 20.160 ;
        RECT 483.530 20.100 483.850 20.160 ;
        RECT 389.230 18.940 389.550 19.000 ;
        RECT 458.245 18.940 458.535 18.985 ;
        RECT 389.230 18.800 458.535 18.940 ;
        RECT 389.230 18.740 389.550 18.800 ;
        RECT 458.245 18.755 458.535 18.800 ;
      LAYER via ;
        RECT 483.560 20.100 483.820 20.360 ;
        RECT 389.260 18.740 389.520 19.000 ;
      LAYER met2 ;
        RECT 484.800 1600.450 485.080 1604.000 ;
        RECT 483.620 1600.310 485.080 1600.450 ;
        RECT 483.620 20.390 483.760 1600.310 ;
        RECT 484.800 1600.000 485.080 1600.310 ;
        RECT 483.560 20.070 483.820 20.390 ;
        RECT 389.260 18.710 389.520 19.030 ;
        RECT 389.320 2.400 389.460 18.710 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 444.890 1592.120 445.210 1592.180 ;
        RECT 490.890 1592.120 491.210 1592.180 ;
        RECT 444.890 1591.980 491.210 1592.120 ;
        RECT 444.890 1591.920 445.210 1591.980 ;
        RECT 490.890 1591.920 491.210 1591.980 ;
        RECT 407.170 19.960 407.490 20.020 ;
        RECT 444.890 19.960 445.210 20.020 ;
        RECT 407.170 19.820 445.210 19.960 ;
        RECT 407.170 19.760 407.490 19.820 ;
        RECT 444.890 19.760 445.210 19.820 ;
      LAYER via ;
        RECT 444.920 1591.920 445.180 1592.180 ;
        RECT 490.920 1591.920 491.180 1592.180 ;
        RECT 407.200 19.760 407.460 20.020 ;
        RECT 444.920 19.760 445.180 20.020 ;
      LAYER met2 ;
        RECT 490.780 1600.380 491.060 1604.000 ;
        RECT 490.780 1600.000 491.120 1600.380 ;
        RECT 490.980 1592.210 491.120 1600.000 ;
        RECT 444.920 1591.890 445.180 1592.210 ;
        RECT 490.920 1591.890 491.180 1592.210 ;
        RECT 444.980 20.050 445.120 1591.890 ;
        RECT 407.200 19.730 407.460 20.050 ;
        RECT 444.920 19.730 445.180 20.050 ;
        RECT 407.260 2.400 407.400 19.730 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 373.480 1600.380 373.760 1604.000 ;
        RECT 373.480 1600.000 373.820 1600.380 ;
        RECT 373.680 1590.365 373.820 1600.000 ;
        RECT 68.630 1589.995 68.910 1590.365 ;
        RECT 373.610 1589.995 373.890 1590.365 ;
        RECT 68.700 17.410 68.840 1589.995 ;
        RECT 68.240 17.270 68.840 17.410 ;
        RECT 68.240 2.400 68.380 17.270 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 68.630 1590.040 68.910 1590.320 ;
        RECT 373.610 1590.040 373.890 1590.320 ;
      LAYER met3 ;
        RECT 68.605 1590.330 68.935 1590.345 ;
        RECT 373.585 1590.330 373.915 1590.345 ;
        RECT 68.605 1590.030 373.915 1590.330 ;
        RECT 68.605 1590.015 68.935 1590.030 ;
        RECT 373.585 1590.015 373.915 1590.030 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 465.590 1592.800 465.910 1592.860 ;
        RECT 497.330 1592.800 497.650 1592.860 ;
        RECT 465.590 1592.660 497.650 1592.800 ;
        RECT 465.590 1592.600 465.910 1592.660 ;
        RECT 497.330 1592.600 497.650 1592.660 ;
        RECT 424.650 16.560 424.970 16.620 ;
        RECT 465.590 16.560 465.910 16.620 ;
        RECT 424.650 16.420 465.910 16.560 ;
        RECT 424.650 16.360 424.970 16.420 ;
        RECT 465.590 16.360 465.910 16.420 ;
      LAYER via ;
        RECT 465.620 1592.600 465.880 1592.860 ;
        RECT 497.360 1592.600 497.620 1592.860 ;
        RECT 424.680 16.360 424.940 16.620 ;
        RECT 465.620 16.360 465.880 16.620 ;
      LAYER met2 ;
        RECT 497.220 1600.380 497.500 1604.000 ;
        RECT 497.220 1600.000 497.560 1600.380 ;
        RECT 497.420 1592.890 497.560 1600.000 ;
        RECT 465.620 1592.570 465.880 1592.890 ;
        RECT 497.360 1592.570 497.620 1592.890 ;
        RECT 465.680 16.650 465.820 1592.570 ;
        RECT 424.680 16.330 424.940 16.650 ;
        RECT 465.620 16.330 465.880 16.650 ;
        RECT 424.740 2.400 424.880 16.330 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 457.385 16.065 457.555 16.915 ;
      LAYER mcon ;
        RECT 457.385 16.745 457.555 16.915 ;
      LAYER met1 ;
        RECT 486.290 1590.760 486.610 1590.820 ;
        RECT 503.310 1590.760 503.630 1590.820 ;
        RECT 486.290 1590.620 503.630 1590.760 ;
        RECT 486.290 1590.560 486.610 1590.620 ;
        RECT 503.310 1590.560 503.630 1590.620 ;
        RECT 442.590 16.900 442.910 16.960 ;
        RECT 457.325 16.900 457.615 16.945 ;
        RECT 442.590 16.760 457.615 16.900 ;
        RECT 442.590 16.700 442.910 16.760 ;
        RECT 457.325 16.715 457.615 16.760 ;
        RECT 457.325 16.220 457.615 16.265 ;
        RECT 486.290 16.220 486.610 16.280 ;
        RECT 457.325 16.080 486.610 16.220 ;
        RECT 457.325 16.035 457.615 16.080 ;
        RECT 486.290 16.020 486.610 16.080 ;
      LAYER via ;
        RECT 486.320 1590.560 486.580 1590.820 ;
        RECT 503.340 1590.560 503.600 1590.820 ;
        RECT 442.620 16.700 442.880 16.960 ;
        RECT 486.320 16.020 486.580 16.280 ;
      LAYER met2 ;
        RECT 503.200 1600.380 503.480 1604.000 ;
        RECT 503.200 1600.000 503.540 1600.380 ;
        RECT 503.400 1590.850 503.540 1600.000 ;
        RECT 486.320 1590.530 486.580 1590.850 ;
        RECT 503.340 1590.530 503.600 1590.850 ;
        RECT 442.620 16.670 442.880 16.990 ;
        RECT 442.680 2.400 442.820 16.670 ;
        RECT 486.380 16.310 486.520 1590.530 ;
        RECT 486.320 15.990 486.580 16.310 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 500.550 1587.360 500.870 1587.420 ;
        RECT 509.750 1587.360 510.070 1587.420 ;
        RECT 500.550 1587.220 510.070 1587.360 ;
        RECT 500.550 1587.160 500.870 1587.220 ;
        RECT 509.750 1587.160 510.070 1587.220 ;
        RECT 460.530 18.600 460.850 18.660 ;
        RECT 500.550 18.600 500.870 18.660 ;
        RECT 460.530 18.460 500.870 18.600 ;
        RECT 460.530 18.400 460.850 18.460 ;
        RECT 500.550 18.400 500.870 18.460 ;
      LAYER via ;
        RECT 500.580 1587.160 500.840 1587.420 ;
        RECT 509.780 1587.160 510.040 1587.420 ;
        RECT 460.560 18.400 460.820 18.660 ;
        RECT 500.580 18.400 500.840 18.660 ;
      LAYER met2 ;
        RECT 509.640 1600.380 509.920 1604.000 ;
        RECT 509.640 1600.000 509.980 1600.380 ;
        RECT 509.840 1587.450 509.980 1600.000 ;
        RECT 500.580 1587.130 500.840 1587.450 ;
        RECT 509.780 1587.130 510.040 1587.450 ;
        RECT 500.640 18.690 500.780 1587.130 ;
        RECT 460.560 18.370 460.820 18.690 ;
        RECT 500.580 18.370 500.840 18.690 ;
        RECT 460.620 2.400 460.760 18.370 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 1589.400 482.930 1589.460 ;
        RECT 515.730 1589.400 516.050 1589.460 ;
        RECT 482.610 1589.260 516.050 1589.400 ;
        RECT 482.610 1589.200 482.930 1589.260 ;
        RECT 515.730 1589.200 516.050 1589.260 ;
        RECT 478.470 17.240 478.790 17.300 ;
        RECT 482.610 17.240 482.930 17.300 ;
        RECT 478.470 17.100 482.930 17.240 ;
        RECT 478.470 17.040 478.790 17.100 ;
        RECT 482.610 17.040 482.930 17.100 ;
      LAYER via ;
        RECT 482.640 1589.200 482.900 1589.460 ;
        RECT 515.760 1589.200 516.020 1589.460 ;
        RECT 478.500 17.040 478.760 17.300 ;
        RECT 482.640 17.040 482.900 17.300 ;
      LAYER met2 ;
        RECT 515.620 1600.380 515.900 1604.000 ;
        RECT 515.620 1600.000 515.960 1600.380 ;
        RECT 515.820 1589.490 515.960 1600.000 ;
        RECT 482.640 1589.170 482.900 1589.490 ;
        RECT 515.760 1589.170 516.020 1589.490 ;
        RECT 482.700 17.330 482.840 1589.170 ;
        RECT 478.500 17.010 478.760 17.330 ;
        RECT 482.640 17.010 482.900 17.330 ;
        RECT 478.560 2.400 478.700 17.010 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 500.090 1588.040 500.410 1588.100 ;
        RECT 521.710 1588.040 522.030 1588.100 ;
        RECT 500.090 1587.900 522.030 1588.040 ;
        RECT 500.090 1587.840 500.410 1587.900 ;
        RECT 521.710 1587.840 522.030 1587.900 ;
        RECT 496.410 17.580 496.730 17.640 ;
        RECT 500.090 17.580 500.410 17.640 ;
        RECT 496.410 17.440 500.410 17.580 ;
        RECT 496.410 17.380 496.730 17.440 ;
        RECT 500.090 17.380 500.410 17.440 ;
      LAYER via ;
        RECT 500.120 1587.840 500.380 1588.100 ;
        RECT 521.740 1587.840 522.000 1588.100 ;
        RECT 496.440 17.380 496.700 17.640 ;
        RECT 500.120 17.380 500.380 17.640 ;
      LAYER met2 ;
        RECT 521.600 1600.380 521.880 1604.000 ;
        RECT 521.600 1600.000 521.940 1600.380 ;
        RECT 521.800 1588.130 521.940 1600.000 ;
        RECT 500.120 1587.810 500.380 1588.130 ;
        RECT 521.740 1587.810 522.000 1588.130 ;
        RECT 500.180 17.670 500.320 1587.810 ;
        RECT 496.440 17.350 496.700 17.670 ;
        RECT 500.120 17.350 500.380 17.670 ;
        RECT 496.500 2.400 496.640 17.350 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.110 1587.700 517.430 1587.760 ;
        RECT 528.150 1587.700 528.470 1587.760 ;
        RECT 517.110 1587.560 528.470 1587.700 ;
        RECT 517.110 1587.500 517.430 1587.560 ;
        RECT 528.150 1587.500 528.470 1587.560 ;
        RECT 513.890 20.640 514.210 20.700 ;
        RECT 517.110 20.640 517.430 20.700 ;
        RECT 513.890 20.500 517.430 20.640 ;
        RECT 513.890 20.440 514.210 20.500 ;
        RECT 517.110 20.440 517.430 20.500 ;
      LAYER via ;
        RECT 517.140 1587.500 517.400 1587.760 ;
        RECT 528.180 1587.500 528.440 1587.760 ;
        RECT 513.920 20.440 514.180 20.700 ;
        RECT 517.140 20.440 517.400 20.700 ;
      LAYER met2 ;
        RECT 528.040 1600.380 528.320 1604.000 ;
        RECT 528.040 1600.000 528.380 1600.380 ;
        RECT 528.240 1587.790 528.380 1600.000 ;
        RECT 517.140 1587.470 517.400 1587.790 ;
        RECT 528.180 1587.470 528.440 1587.790 ;
        RECT 517.200 20.730 517.340 1587.470 ;
        RECT 513.920 20.410 514.180 20.730 ;
        RECT 517.140 20.410 517.400 20.730 ;
        RECT 513.980 2.400 514.120 20.410 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 534.020 1600.450 534.300 1604.000 ;
        RECT 533.300 1600.310 534.300 1600.450 ;
        RECT 533.300 1580.050 533.440 1600.310 ;
        RECT 534.020 1600.000 534.300 1600.310 ;
        RECT 531.920 1579.910 533.440 1580.050 ;
        RECT 531.920 2.400 532.060 1579.910 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 540.570 1587.360 540.890 1587.420 ;
        RECT 544.250 1587.360 544.570 1587.420 ;
        RECT 540.570 1587.220 544.570 1587.360 ;
        RECT 540.570 1587.160 540.890 1587.220 ;
        RECT 544.250 1587.160 544.570 1587.220 ;
        RECT 544.250 16.220 544.570 16.280 ;
        RECT 549.770 16.220 550.090 16.280 ;
        RECT 544.250 16.080 550.090 16.220 ;
        RECT 544.250 16.020 544.570 16.080 ;
        RECT 549.770 16.020 550.090 16.080 ;
      LAYER via ;
        RECT 540.600 1587.160 540.860 1587.420 ;
        RECT 544.280 1587.160 544.540 1587.420 ;
        RECT 544.280 16.020 544.540 16.280 ;
        RECT 549.800 16.020 550.060 16.280 ;
      LAYER met2 ;
        RECT 540.460 1600.380 540.740 1604.000 ;
        RECT 540.460 1600.000 540.800 1600.380 ;
        RECT 540.660 1587.450 540.800 1600.000 ;
        RECT 540.600 1587.130 540.860 1587.450 ;
        RECT 544.280 1587.130 544.540 1587.450 ;
        RECT 544.340 16.310 544.480 1587.130 ;
        RECT 544.280 15.990 544.540 16.310 ;
        RECT 549.800 15.990 550.060 16.310 ;
        RECT 549.860 2.400 550.000 15.990 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 546.550 1589.740 546.870 1589.800 ;
        RECT 551.150 1589.740 551.470 1589.800 ;
        RECT 546.550 1589.600 551.470 1589.740 ;
        RECT 546.550 1589.540 546.870 1589.600 ;
        RECT 551.150 1589.540 551.470 1589.600 ;
        RECT 551.150 17.240 551.470 17.300 ;
        RECT 551.150 17.100 556.440 17.240 ;
        RECT 551.150 17.040 551.470 17.100 ;
        RECT 556.300 16.900 556.440 17.100 ;
        RECT 567.710 16.900 568.030 16.960 ;
        RECT 556.300 16.760 568.030 16.900 ;
        RECT 567.710 16.700 568.030 16.760 ;
      LAYER via ;
        RECT 546.580 1589.540 546.840 1589.800 ;
        RECT 551.180 1589.540 551.440 1589.800 ;
        RECT 551.180 17.040 551.440 17.300 ;
        RECT 567.740 16.700 568.000 16.960 ;
      LAYER met2 ;
        RECT 546.440 1600.380 546.720 1604.000 ;
        RECT 546.440 1600.000 546.780 1600.380 ;
        RECT 546.640 1589.830 546.780 1600.000 ;
        RECT 546.580 1589.510 546.840 1589.830 ;
        RECT 551.180 1589.510 551.440 1589.830 ;
        RECT 551.240 17.330 551.380 1589.510 ;
        RECT 551.180 17.010 551.440 17.330 ;
        RECT 567.740 16.670 568.000 16.990 ;
        RECT 567.800 2.400 567.940 16.670 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 552.990 1587.360 553.310 1587.420 ;
        RECT 569.090 1587.360 569.410 1587.420 ;
        RECT 552.990 1587.220 569.410 1587.360 ;
        RECT 552.990 1587.160 553.310 1587.220 ;
        RECT 569.090 1587.160 569.410 1587.220 ;
        RECT 569.090 17.920 569.410 17.980 ;
        RECT 585.650 17.920 585.970 17.980 ;
        RECT 569.090 17.780 585.970 17.920 ;
        RECT 569.090 17.720 569.410 17.780 ;
        RECT 585.650 17.720 585.970 17.780 ;
      LAYER via ;
        RECT 553.020 1587.160 553.280 1587.420 ;
        RECT 569.120 1587.160 569.380 1587.420 ;
        RECT 569.120 17.720 569.380 17.980 ;
        RECT 585.680 17.720 585.940 17.980 ;
      LAYER met2 ;
        RECT 552.880 1600.380 553.160 1604.000 ;
        RECT 552.880 1600.000 553.220 1600.380 ;
        RECT 553.080 1587.450 553.220 1600.000 ;
        RECT 553.020 1587.130 553.280 1587.450 ;
        RECT 569.120 1587.130 569.380 1587.450 ;
        RECT 569.180 18.010 569.320 1587.130 ;
        RECT 569.120 17.690 569.380 18.010 ;
        RECT 585.680 17.690 585.940 18.010 ;
        RECT 585.740 2.400 585.880 17.690 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.760 1600.450 382.040 1604.000 ;
        RECT 380.580 1600.310 382.040 1600.450 ;
        RECT 380.580 18.205 380.720 1600.310 ;
        RECT 381.760 1600.000 382.040 1600.310 ;
        RECT 91.630 17.835 91.910 18.205 ;
        RECT 380.510 17.835 380.790 18.205 ;
        RECT 91.700 2.400 91.840 17.835 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 91.630 17.880 91.910 18.160 ;
        RECT 380.510 17.880 380.790 18.160 ;
      LAYER met3 ;
        RECT 91.605 18.170 91.935 18.185 ;
        RECT 380.485 18.170 380.815 18.185 ;
        RECT 91.605 17.870 380.815 18.170 ;
        RECT 91.605 17.855 91.935 17.870 ;
        RECT 380.485 17.855 380.815 17.870 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 558.970 1590.420 559.290 1590.480 ;
        RECT 558.970 1590.280 567.020 1590.420 ;
        RECT 558.970 1590.220 559.290 1590.280 ;
        RECT 566.880 1589.740 567.020 1590.280 ;
        RECT 601.290 1589.740 601.610 1589.800 ;
        RECT 566.880 1589.600 601.610 1589.740 ;
        RECT 601.290 1589.540 601.610 1589.600 ;
      LAYER via ;
        RECT 559.000 1590.220 559.260 1590.480 ;
        RECT 601.320 1589.540 601.580 1589.800 ;
      LAYER met2 ;
        RECT 558.860 1600.380 559.140 1604.000 ;
        RECT 558.860 1600.000 559.200 1600.380 ;
        RECT 559.060 1590.510 559.200 1600.000 ;
        RECT 559.000 1590.190 559.260 1590.510 ;
        RECT 601.320 1589.510 601.580 1589.830 ;
        RECT 601.380 3.130 601.520 1589.510 ;
        RECT 601.380 2.990 603.360 3.130 ;
        RECT 603.220 2.400 603.360 2.990 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 1591.100 565.730 1591.160 ;
        RECT 617.390 1591.100 617.710 1591.160 ;
        RECT 565.410 1590.960 617.710 1591.100 ;
        RECT 565.410 1590.900 565.730 1590.960 ;
        RECT 617.390 1590.900 617.710 1590.960 ;
        RECT 617.390 17.580 617.710 17.640 ;
        RECT 621.070 17.580 621.390 17.640 ;
        RECT 617.390 17.440 621.390 17.580 ;
        RECT 617.390 17.380 617.710 17.440 ;
        RECT 621.070 17.380 621.390 17.440 ;
      LAYER via ;
        RECT 565.440 1590.900 565.700 1591.160 ;
        RECT 617.420 1590.900 617.680 1591.160 ;
        RECT 617.420 17.380 617.680 17.640 ;
        RECT 621.100 17.380 621.360 17.640 ;
      LAYER met2 ;
        RECT 565.300 1600.380 565.580 1604.000 ;
        RECT 565.300 1600.000 565.640 1600.380 ;
        RECT 565.500 1591.190 565.640 1600.000 ;
        RECT 565.440 1590.870 565.700 1591.190 ;
        RECT 617.420 1590.870 617.680 1591.190 ;
        RECT 617.480 17.670 617.620 1590.870 ;
        RECT 617.420 17.350 617.680 17.670 ;
        RECT 621.100 17.350 621.360 17.670 ;
        RECT 621.160 2.400 621.300 17.350 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.040 1600.380 390.320 1604.000 ;
        RECT 390.040 1600.000 390.380 1600.380 ;
        RECT 390.240 1593.085 390.380 1600.000 ;
        RECT 116.930 1592.715 117.210 1593.085 ;
        RECT 390.170 1592.715 390.450 1593.085 ;
        RECT 117.000 17.410 117.140 1592.715 ;
        RECT 115.620 17.270 117.140 17.410 ;
        RECT 115.620 2.400 115.760 17.270 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 116.930 1592.760 117.210 1593.040 ;
        RECT 390.170 1592.760 390.450 1593.040 ;
      LAYER met3 ;
        RECT 116.905 1593.050 117.235 1593.065 ;
        RECT 390.145 1593.050 390.475 1593.065 ;
        RECT 116.905 1592.750 390.475 1593.050 ;
        RECT 116.905 1592.735 117.235 1592.750 ;
        RECT 390.145 1592.735 390.475 1592.750 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 394.365 1393.745 394.535 1414.655 ;
        RECT 393.905 1097.265 394.075 1145.375 ;
        RECT 393.905 917.745 394.075 931.855 ;
        RECT 393.905 531.505 394.075 579.615 ;
        RECT 393.445 421.345 393.615 469.115 ;
        RECT 393.445 324.445 393.615 414.035 ;
        RECT 393.905 186.405 394.075 193.375 ;
        RECT 394.365 89.845 394.535 137.955 ;
        RECT 353.425 18.445 353.595 19.635 ;
      LAYER mcon ;
        RECT 394.365 1414.485 394.535 1414.655 ;
        RECT 393.905 1145.205 394.075 1145.375 ;
        RECT 393.905 931.685 394.075 931.855 ;
        RECT 393.905 579.445 394.075 579.615 ;
        RECT 393.445 468.945 393.615 469.115 ;
        RECT 393.445 413.865 393.615 414.035 ;
        RECT 393.905 193.205 394.075 193.375 ;
        RECT 394.365 137.785 394.535 137.955 ;
        RECT 353.425 19.465 353.595 19.635 ;
      LAYER met1 ;
        RECT 394.750 1545.880 395.070 1545.940 ;
        RECT 397.050 1545.880 397.370 1545.940 ;
        RECT 394.750 1545.740 397.370 1545.880 ;
        RECT 394.750 1545.680 395.070 1545.740 ;
        RECT 397.050 1545.680 397.370 1545.740 ;
        RECT 394.750 1449.660 395.070 1449.720 ;
        RECT 394.380 1449.520 395.070 1449.660 ;
        RECT 394.380 1449.380 394.520 1449.520 ;
        RECT 394.750 1449.460 395.070 1449.520 ;
        RECT 394.290 1449.120 394.610 1449.380 ;
        RECT 393.830 1414.640 394.150 1414.700 ;
        RECT 394.305 1414.640 394.595 1414.685 ;
        RECT 393.830 1414.500 394.595 1414.640 ;
        RECT 393.830 1414.440 394.150 1414.500 ;
        RECT 394.305 1414.455 394.595 1414.500 ;
        RECT 394.290 1393.900 394.610 1393.960 ;
        RECT 394.095 1393.760 394.610 1393.900 ;
        RECT 394.290 1393.700 394.610 1393.760 ;
        RECT 393.370 1352.420 393.690 1352.480 ;
        RECT 394.290 1352.420 394.610 1352.480 ;
        RECT 393.370 1352.280 394.610 1352.420 ;
        RECT 393.370 1352.220 393.690 1352.280 ;
        RECT 394.290 1352.220 394.610 1352.280 ;
        RECT 393.830 1242.260 394.150 1242.320 ;
        RECT 394.750 1242.260 395.070 1242.320 ;
        RECT 393.830 1242.120 395.070 1242.260 ;
        RECT 393.830 1242.060 394.150 1242.120 ;
        RECT 394.750 1242.060 395.070 1242.120 ;
        RECT 393.830 1200.580 394.150 1200.840 ;
        RECT 393.920 1200.440 394.060 1200.580 ;
        RECT 394.290 1200.440 394.610 1200.500 ;
        RECT 393.920 1200.300 394.610 1200.440 ;
        RECT 394.290 1200.240 394.610 1200.300 ;
        RECT 393.845 1145.360 394.135 1145.405 ;
        RECT 394.750 1145.360 395.070 1145.420 ;
        RECT 393.845 1145.220 395.070 1145.360 ;
        RECT 393.845 1145.175 394.135 1145.220 ;
        RECT 394.750 1145.160 395.070 1145.220 ;
        RECT 393.830 1097.420 394.150 1097.480 ;
        RECT 393.635 1097.280 394.150 1097.420 ;
        RECT 393.830 1097.220 394.150 1097.280 ;
        RECT 393.370 1055.940 393.690 1056.000 ;
        RECT 393.830 1055.940 394.150 1056.000 ;
        RECT 393.370 1055.800 394.150 1055.940 ;
        RECT 393.370 1055.740 393.690 1055.800 ;
        RECT 393.830 1055.740 394.150 1055.800 ;
        RECT 393.830 931.840 394.150 931.900 ;
        RECT 393.635 931.700 394.150 931.840 ;
        RECT 393.830 931.640 394.150 931.700 ;
        RECT 393.830 917.900 394.150 917.960 ;
        RECT 393.635 917.760 394.150 917.900 ;
        RECT 393.830 917.700 394.150 917.760 ;
        RECT 393.830 869.620 394.150 869.680 ;
        RECT 394.290 869.620 394.610 869.680 ;
        RECT 393.830 869.480 394.610 869.620 ;
        RECT 393.830 869.420 394.150 869.480 ;
        RECT 394.290 869.420 394.610 869.480 ;
        RECT 393.370 838.340 393.690 838.400 ;
        RECT 394.290 838.340 394.610 838.400 ;
        RECT 393.370 838.200 394.610 838.340 ;
        RECT 393.370 838.140 393.690 838.200 ;
        RECT 394.290 838.140 394.610 838.200 ;
        RECT 393.830 765.720 394.150 765.980 ;
        RECT 393.920 765.240 394.060 765.720 ;
        RECT 394.750 765.240 395.070 765.300 ;
        RECT 393.920 765.100 395.070 765.240 ;
        RECT 394.750 765.040 395.070 765.100 ;
        RECT 393.845 579.600 394.135 579.645 ;
        RECT 394.290 579.600 394.610 579.660 ;
        RECT 393.845 579.460 394.610 579.600 ;
        RECT 393.845 579.415 394.135 579.460 ;
        RECT 394.290 579.400 394.610 579.460 ;
        RECT 393.830 531.660 394.150 531.720 ;
        RECT 393.635 531.520 394.150 531.660 ;
        RECT 393.830 531.460 394.150 531.520 ;
        RECT 393.385 469.100 393.675 469.145 ;
        RECT 394.290 469.100 394.610 469.160 ;
        RECT 393.385 468.960 394.610 469.100 ;
        RECT 393.385 468.915 393.675 468.960 ;
        RECT 394.290 468.900 394.610 468.960 ;
        RECT 393.370 421.500 393.690 421.560 ;
        RECT 393.175 421.360 393.690 421.500 ;
        RECT 393.370 421.300 393.690 421.360 ;
        RECT 393.370 420.620 393.690 420.880 ;
        RECT 393.460 420.480 393.600 420.620 ;
        RECT 394.290 420.480 394.610 420.540 ;
        RECT 393.460 420.340 394.610 420.480 ;
        RECT 394.290 420.280 394.610 420.340 ;
        RECT 393.385 414.020 393.675 414.065 ;
        RECT 394.290 414.020 394.610 414.080 ;
        RECT 393.385 413.880 394.610 414.020 ;
        RECT 393.385 413.835 393.675 413.880 ;
        RECT 394.290 413.820 394.610 413.880 ;
        RECT 393.370 324.600 393.690 324.660 ;
        RECT 393.175 324.460 393.690 324.600 ;
        RECT 393.370 324.400 393.690 324.460 ;
        RECT 393.370 307.260 393.690 307.320 ;
        RECT 394.750 307.260 395.070 307.320 ;
        RECT 393.370 307.120 395.070 307.260 ;
        RECT 393.370 307.060 393.690 307.120 ;
        RECT 394.750 307.060 395.070 307.120 ;
        RECT 393.830 241.640 394.150 241.700 ;
        RECT 394.750 241.640 395.070 241.700 ;
        RECT 393.830 241.500 395.070 241.640 ;
        RECT 393.830 241.440 394.150 241.500 ;
        RECT 394.750 241.440 395.070 241.500 ;
        RECT 393.830 193.360 394.150 193.420 ;
        RECT 393.635 193.220 394.150 193.360 ;
        RECT 393.830 193.160 394.150 193.220 ;
        RECT 393.830 186.560 394.150 186.620 ;
        RECT 393.635 186.420 394.150 186.560 ;
        RECT 393.830 186.360 394.150 186.420 ;
        RECT 394.305 137.940 394.595 137.985 ;
        RECT 394.750 137.940 395.070 138.000 ;
        RECT 394.305 137.800 395.070 137.940 ;
        RECT 394.305 137.755 394.595 137.800 ;
        RECT 394.750 137.740 395.070 137.800 ;
        RECT 394.290 90.000 394.610 90.060 ;
        RECT 394.095 89.860 394.610 90.000 ;
        RECT 394.290 89.800 394.610 89.860 ;
        RECT 139.450 19.620 139.770 19.680 ;
        RECT 353.365 19.620 353.655 19.665 ;
        RECT 139.450 19.480 353.655 19.620 ;
        RECT 139.450 19.420 139.770 19.480 ;
        RECT 353.365 19.435 353.655 19.480 ;
        RECT 394.290 19.280 394.610 19.340 ;
        RECT 380.580 19.140 394.610 19.280 ;
        RECT 380.580 18.940 380.720 19.140 ;
        RECT 394.290 19.080 394.610 19.140 ;
        RECT 366.320 18.800 380.720 18.940 ;
        RECT 353.365 18.600 353.655 18.645 ;
        RECT 366.320 18.600 366.460 18.800 ;
        RECT 353.365 18.460 366.460 18.600 ;
        RECT 353.365 18.415 353.655 18.460 ;
      LAYER via ;
        RECT 394.780 1545.680 395.040 1545.940 ;
        RECT 397.080 1545.680 397.340 1545.940 ;
        RECT 394.780 1449.460 395.040 1449.720 ;
        RECT 394.320 1449.120 394.580 1449.380 ;
        RECT 393.860 1414.440 394.120 1414.700 ;
        RECT 394.320 1393.700 394.580 1393.960 ;
        RECT 393.400 1352.220 393.660 1352.480 ;
        RECT 394.320 1352.220 394.580 1352.480 ;
        RECT 393.860 1242.060 394.120 1242.320 ;
        RECT 394.780 1242.060 395.040 1242.320 ;
        RECT 393.860 1200.580 394.120 1200.840 ;
        RECT 394.320 1200.240 394.580 1200.500 ;
        RECT 394.780 1145.160 395.040 1145.420 ;
        RECT 393.860 1097.220 394.120 1097.480 ;
        RECT 393.400 1055.740 393.660 1056.000 ;
        RECT 393.860 1055.740 394.120 1056.000 ;
        RECT 393.860 931.640 394.120 931.900 ;
        RECT 393.860 917.700 394.120 917.960 ;
        RECT 393.860 869.420 394.120 869.680 ;
        RECT 394.320 869.420 394.580 869.680 ;
        RECT 393.400 838.140 393.660 838.400 ;
        RECT 394.320 838.140 394.580 838.400 ;
        RECT 393.860 765.720 394.120 765.980 ;
        RECT 394.780 765.040 395.040 765.300 ;
        RECT 394.320 579.400 394.580 579.660 ;
        RECT 393.860 531.460 394.120 531.720 ;
        RECT 394.320 468.900 394.580 469.160 ;
        RECT 393.400 421.300 393.660 421.560 ;
        RECT 393.400 420.620 393.660 420.880 ;
        RECT 394.320 420.280 394.580 420.540 ;
        RECT 394.320 413.820 394.580 414.080 ;
        RECT 393.400 324.400 393.660 324.660 ;
        RECT 393.400 307.060 393.660 307.320 ;
        RECT 394.780 307.060 395.040 307.320 ;
        RECT 393.860 241.440 394.120 241.700 ;
        RECT 394.780 241.440 395.040 241.700 ;
        RECT 393.860 193.160 394.120 193.420 ;
        RECT 393.860 186.360 394.120 186.620 ;
        RECT 394.780 137.740 395.040 138.000 ;
        RECT 394.320 89.800 394.580 90.060 ;
        RECT 139.480 19.420 139.740 19.680 ;
        RECT 394.320 19.080 394.580 19.340 ;
      LAYER met2 ;
        RECT 398.320 1600.450 398.600 1604.000 ;
        RECT 397.140 1600.310 398.600 1600.450 ;
        RECT 397.140 1545.970 397.280 1600.310 ;
        RECT 398.320 1600.000 398.600 1600.310 ;
        RECT 394.780 1545.650 395.040 1545.970 ;
        RECT 397.080 1545.650 397.340 1545.970 ;
        RECT 394.840 1449.750 394.980 1545.650 ;
        RECT 394.780 1449.430 395.040 1449.750 ;
        RECT 394.320 1449.090 394.580 1449.410 ;
        RECT 394.380 1442.010 394.520 1449.090 ;
        RECT 393.920 1441.870 394.520 1442.010 ;
        RECT 393.920 1414.730 394.060 1441.870 ;
        RECT 393.860 1414.410 394.120 1414.730 ;
        RECT 394.320 1393.670 394.580 1393.990 ;
        RECT 394.380 1352.510 394.520 1393.670 ;
        RECT 393.400 1352.190 393.660 1352.510 ;
        RECT 394.320 1352.190 394.580 1352.510 ;
        RECT 393.460 1338.765 393.600 1352.190 ;
        RECT 393.390 1338.395 393.670 1338.765 ;
        RECT 394.770 1338.395 395.050 1338.765 ;
        RECT 394.840 1242.350 394.980 1338.395 ;
        RECT 393.860 1242.030 394.120 1242.350 ;
        RECT 394.780 1242.030 395.040 1242.350 ;
        RECT 393.920 1200.870 394.060 1242.030 ;
        RECT 393.860 1200.550 394.120 1200.870 ;
        RECT 394.320 1200.210 394.580 1200.530 ;
        RECT 394.380 1145.530 394.520 1200.210 ;
        RECT 394.380 1145.450 394.980 1145.530 ;
        RECT 394.380 1145.390 395.040 1145.450 ;
        RECT 394.780 1145.130 395.040 1145.390 ;
        RECT 394.840 1144.975 394.980 1145.130 ;
        RECT 393.860 1097.190 394.120 1097.510 ;
        RECT 393.920 1056.030 394.060 1097.190 ;
        RECT 393.400 1055.710 393.660 1056.030 ;
        RECT 393.860 1055.710 394.120 1056.030 ;
        RECT 393.460 1017.690 393.600 1055.710 ;
        RECT 393.460 1017.550 394.060 1017.690 ;
        RECT 393.920 1014.405 394.060 1017.550 ;
        RECT 393.850 1014.035 394.130 1014.405 ;
        RECT 394.310 1013.355 394.590 1013.725 ;
        RECT 394.380 966.010 394.520 1013.355 ;
        RECT 393.920 965.870 394.520 966.010 ;
        RECT 393.920 931.930 394.060 965.870 ;
        RECT 393.860 931.610 394.120 931.930 ;
        RECT 393.920 917.990 394.060 918.145 ;
        RECT 393.860 917.730 394.120 917.990 ;
        RECT 393.860 917.670 394.520 917.730 ;
        RECT 393.920 917.590 394.520 917.670 ;
        RECT 394.380 917.050 394.520 917.590 ;
        RECT 393.920 916.910 394.520 917.050 ;
        RECT 393.920 869.710 394.060 916.910 ;
        RECT 393.860 869.390 394.120 869.710 ;
        RECT 394.320 869.390 394.580 869.710 ;
        RECT 394.380 838.430 394.520 869.390 ;
        RECT 393.400 838.110 393.660 838.430 ;
        RECT 394.320 838.110 394.580 838.430 ;
        RECT 393.460 814.370 393.600 838.110 ;
        RECT 393.460 814.230 394.060 814.370 ;
        RECT 393.920 766.010 394.060 814.230 ;
        RECT 393.860 765.690 394.120 766.010 ;
        RECT 394.780 765.010 395.040 765.330 ;
        RECT 394.840 628.165 394.980 765.010 ;
        RECT 393.850 627.795 394.130 628.165 ;
        RECT 394.770 627.795 395.050 628.165 ;
        RECT 393.920 603.570 394.060 627.795 ;
        RECT 393.920 603.430 394.520 603.570 ;
        RECT 394.380 579.690 394.520 603.430 ;
        RECT 394.320 579.370 394.580 579.690 ;
        RECT 393.860 531.430 394.120 531.750 ;
        RECT 393.920 507.010 394.060 531.430 ;
        RECT 393.920 506.870 394.520 507.010 ;
        RECT 394.380 469.190 394.520 506.870 ;
        RECT 394.320 468.870 394.580 469.190 ;
        RECT 393.400 421.270 393.660 421.590 ;
        RECT 393.460 420.910 393.600 421.270 ;
        RECT 393.400 420.590 393.660 420.910 ;
        RECT 394.320 420.250 394.580 420.570 ;
        RECT 394.380 414.110 394.520 420.250 ;
        RECT 394.320 413.790 394.580 414.110 ;
        RECT 393.400 324.370 393.660 324.690 ;
        RECT 393.460 307.350 393.600 324.370 ;
        RECT 393.400 307.030 393.660 307.350 ;
        RECT 394.780 307.030 395.040 307.350 ;
        RECT 394.840 241.730 394.980 307.030 ;
        RECT 393.860 241.410 394.120 241.730 ;
        RECT 394.780 241.410 395.040 241.730 ;
        RECT 393.920 193.450 394.060 241.410 ;
        RECT 393.860 193.130 394.120 193.450 ;
        RECT 393.860 186.330 394.120 186.650 ;
        RECT 393.920 145.250 394.060 186.330 ;
        RECT 393.920 145.110 394.980 145.250 ;
        RECT 394.840 138.030 394.980 145.110 ;
        RECT 394.780 137.710 395.040 138.030 ;
        RECT 394.320 89.770 394.580 90.090 ;
        RECT 139.480 19.390 139.740 19.710 ;
        RECT 139.540 2.400 139.680 19.390 ;
        RECT 394.380 19.370 394.520 89.770 ;
        RECT 394.320 19.050 394.580 19.370 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 393.390 1338.440 393.670 1338.720 ;
        RECT 394.770 1338.440 395.050 1338.720 ;
        RECT 393.850 1014.080 394.130 1014.360 ;
        RECT 394.310 1013.400 394.590 1013.680 ;
        RECT 393.850 627.840 394.130 628.120 ;
        RECT 394.770 627.840 395.050 628.120 ;
      LAYER met3 ;
        RECT 393.365 1338.730 393.695 1338.745 ;
        RECT 394.745 1338.730 395.075 1338.745 ;
        RECT 393.365 1338.430 395.075 1338.730 ;
        RECT 393.365 1338.415 393.695 1338.430 ;
        RECT 394.745 1338.415 395.075 1338.430 ;
        RECT 393.825 1014.370 394.155 1014.385 ;
        RECT 393.150 1014.070 394.155 1014.370 ;
        RECT 393.150 1013.690 393.450 1014.070 ;
        RECT 393.825 1014.055 394.155 1014.070 ;
        RECT 394.285 1013.690 394.615 1013.705 ;
        RECT 393.150 1013.390 394.615 1013.690 ;
        RECT 394.285 1013.375 394.615 1013.390 ;
        RECT 393.825 628.130 394.155 628.145 ;
        RECT 394.745 628.130 395.075 628.145 ;
        RECT 393.825 627.830 395.075 628.130 ;
        RECT 393.825 627.815 394.155 627.830 ;
        RECT 394.745 627.815 395.075 627.830 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 1591.100 158.630 1591.160 ;
        RECT 158.310 1590.960 392.680 1591.100 ;
        RECT 158.310 1590.900 158.630 1590.960 ;
        RECT 392.540 1590.760 392.680 1590.960 ;
        RECT 404.410 1590.760 404.730 1590.820 ;
        RECT 392.540 1590.620 404.730 1590.760 ;
        RECT 404.410 1590.560 404.730 1590.620 ;
      LAYER via ;
        RECT 158.340 1590.900 158.600 1591.160 ;
        RECT 404.440 1590.560 404.700 1590.820 ;
      LAYER met2 ;
        RECT 404.300 1600.380 404.580 1604.000 ;
        RECT 404.300 1600.000 404.640 1600.380 ;
        RECT 158.340 1590.870 158.600 1591.190 ;
        RECT 158.400 17.410 158.540 1590.870 ;
        RECT 404.500 1590.850 404.640 1600.000 ;
        RECT 404.440 1590.530 404.700 1590.850 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 409.545 723.945 409.715 807.075 ;
        RECT 408.625 379.525 408.795 427.635 ;
        RECT 408.625 193.205 408.795 258.995 ;
      LAYER mcon ;
        RECT 409.545 806.905 409.715 807.075 ;
        RECT 408.625 427.465 408.795 427.635 ;
        RECT 408.625 258.825 408.795 258.995 ;
      LAYER met1 ;
        RECT 408.550 1449.320 408.870 1449.380 ;
        RECT 409.010 1449.320 409.330 1449.380 ;
        RECT 408.550 1449.180 409.330 1449.320 ;
        RECT 408.550 1449.120 408.870 1449.180 ;
        RECT 409.010 1449.120 409.330 1449.180 ;
        RECT 408.090 1393.900 408.410 1393.960 ;
        RECT 408.090 1393.760 408.780 1393.900 ;
        RECT 408.090 1393.700 408.410 1393.760 ;
        RECT 408.640 1393.620 408.780 1393.760 ;
        RECT 408.550 1393.360 408.870 1393.620 ;
        RECT 408.550 1379.960 408.870 1380.020 ;
        RECT 409.470 1379.960 409.790 1380.020 ;
        RECT 408.550 1379.820 409.790 1379.960 ;
        RECT 408.550 1379.760 408.870 1379.820 ;
        RECT 409.470 1379.760 409.790 1379.820 ;
        RECT 408.550 1254.980 408.870 1255.240 ;
        RECT 408.640 1254.560 408.780 1254.980 ;
        RECT 408.550 1254.300 408.870 1254.560 ;
        RECT 408.550 1207.380 408.870 1207.640 ;
        RECT 408.640 1207.240 408.780 1207.380 ;
        RECT 409.010 1207.240 409.330 1207.300 ;
        RECT 408.640 1207.100 409.330 1207.240 ;
        RECT 409.010 1207.040 409.330 1207.100 ;
        RECT 409.010 1173.040 409.330 1173.300 ;
        RECT 409.100 1172.620 409.240 1173.040 ;
        RECT 409.010 1172.360 409.330 1172.620 ;
        RECT 408.550 1111.020 408.870 1111.080 ;
        RECT 409.010 1111.020 409.330 1111.080 ;
        RECT 408.550 1110.880 409.330 1111.020 ;
        RECT 408.550 1110.820 408.870 1110.880 ;
        RECT 409.010 1110.820 409.330 1110.880 ;
        RECT 408.550 979.920 408.870 980.180 ;
        RECT 408.640 979.780 408.780 979.920 ;
        RECT 409.010 979.780 409.330 979.840 ;
        RECT 408.640 979.640 409.330 979.780 ;
        RECT 409.010 979.580 409.330 979.640 ;
        RECT 409.010 869.620 409.330 869.680 ;
        RECT 409.470 869.620 409.790 869.680 ;
        RECT 409.010 869.480 409.790 869.620 ;
        RECT 409.010 869.420 409.330 869.480 ;
        RECT 409.470 869.420 409.790 869.480 ;
        RECT 409.010 838.340 409.330 838.400 ;
        RECT 409.930 838.340 410.250 838.400 ;
        RECT 409.010 838.200 410.250 838.340 ;
        RECT 409.010 838.140 409.330 838.200 ;
        RECT 409.930 838.140 410.250 838.200 ;
        RECT 409.470 807.060 409.790 807.120 ;
        RECT 409.275 806.920 409.790 807.060 ;
        RECT 409.470 806.860 409.790 806.920 ;
        RECT 409.470 724.100 409.790 724.160 ;
        RECT 409.275 723.960 409.790 724.100 ;
        RECT 409.470 723.900 409.790 723.960 ;
        RECT 409.470 717.640 409.790 717.700 ;
        RECT 410.390 717.640 410.710 717.700 ;
        RECT 409.470 717.500 410.710 717.640 ;
        RECT 409.470 717.440 409.790 717.500 ;
        RECT 410.390 717.440 410.710 717.500 ;
        RECT 409.010 545.600 409.330 545.660 ;
        RECT 408.640 545.460 409.330 545.600 ;
        RECT 408.640 544.980 408.780 545.460 ;
        RECT 409.010 545.400 409.330 545.460 ;
        RECT 408.550 544.720 408.870 544.980 ;
        RECT 408.550 427.620 408.870 427.680 ;
        RECT 408.355 427.480 408.870 427.620 ;
        RECT 408.550 427.420 408.870 427.480 ;
        RECT 408.565 379.680 408.855 379.725 ;
        RECT 409.010 379.680 409.330 379.740 ;
        RECT 408.565 379.540 409.330 379.680 ;
        RECT 408.565 379.495 408.855 379.540 ;
        RECT 409.010 379.480 409.330 379.540 ;
        RECT 409.010 352.280 409.330 352.540 ;
        RECT 409.100 351.860 409.240 352.280 ;
        RECT 409.010 351.600 409.330 351.860 ;
        RECT 408.565 258.980 408.855 259.025 ;
        RECT 409.010 258.980 409.330 259.040 ;
        RECT 408.565 258.840 409.330 258.980 ;
        RECT 408.565 258.795 408.855 258.840 ;
        RECT 409.010 258.780 409.330 258.840 ;
        RECT 408.565 193.360 408.855 193.405 ;
        RECT 409.010 193.360 409.330 193.420 ;
        RECT 408.565 193.220 409.330 193.360 ;
        RECT 408.565 193.175 408.855 193.220 ;
        RECT 409.010 193.160 409.330 193.220 ;
        RECT 174.870 20.300 175.190 20.360 ;
        RECT 409.010 20.300 409.330 20.360 ;
        RECT 174.870 20.160 409.330 20.300 ;
        RECT 174.870 20.100 175.190 20.160 ;
        RECT 409.010 20.100 409.330 20.160 ;
      LAYER via ;
        RECT 408.580 1449.120 408.840 1449.380 ;
        RECT 409.040 1449.120 409.300 1449.380 ;
        RECT 408.120 1393.700 408.380 1393.960 ;
        RECT 408.580 1393.360 408.840 1393.620 ;
        RECT 408.580 1379.760 408.840 1380.020 ;
        RECT 409.500 1379.760 409.760 1380.020 ;
        RECT 408.580 1254.980 408.840 1255.240 ;
        RECT 408.580 1254.300 408.840 1254.560 ;
        RECT 408.580 1207.380 408.840 1207.640 ;
        RECT 409.040 1207.040 409.300 1207.300 ;
        RECT 409.040 1173.040 409.300 1173.300 ;
        RECT 409.040 1172.360 409.300 1172.620 ;
        RECT 408.580 1110.820 408.840 1111.080 ;
        RECT 409.040 1110.820 409.300 1111.080 ;
        RECT 408.580 979.920 408.840 980.180 ;
        RECT 409.040 979.580 409.300 979.840 ;
        RECT 409.040 869.420 409.300 869.680 ;
        RECT 409.500 869.420 409.760 869.680 ;
        RECT 409.040 838.140 409.300 838.400 ;
        RECT 409.960 838.140 410.220 838.400 ;
        RECT 409.500 806.860 409.760 807.120 ;
        RECT 409.500 723.900 409.760 724.160 ;
        RECT 409.500 717.440 409.760 717.700 ;
        RECT 410.420 717.440 410.680 717.700 ;
        RECT 409.040 545.400 409.300 545.660 ;
        RECT 408.580 544.720 408.840 544.980 ;
        RECT 408.580 427.420 408.840 427.680 ;
        RECT 409.040 379.480 409.300 379.740 ;
        RECT 409.040 352.280 409.300 352.540 ;
        RECT 409.040 351.600 409.300 351.860 ;
        RECT 409.040 258.780 409.300 259.040 ;
        RECT 409.040 193.160 409.300 193.420 ;
        RECT 174.900 20.100 175.160 20.360 ;
        RECT 409.040 20.100 409.300 20.360 ;
      LAYER met2 ;
        RECT 410.280 1601.130 410.560 1604.000 ;
        RECT 409.560 1600.990 410.560 1601.130 ;
        RECT 409.560 1597.050 409.700 1600.990 ;
        RECT 410.280 1600.000 410.560 1600.990 ;
        RECT 409.560 1596.910 410.160 1597.050 ;
        RECT 410.020 1580.050 410.160 1596.910 ;
        RECT 408.180 1579.910 410.160 1580.050 ;
        RECT 408.180 1510.690 408.320 1579.910 ;
        RECT 408.180 1510.550 408.780 1510.690 ;
        RECT 408.640 1449.410 408.780 1510.550 ;
        RECT 408.580 1449.090 408.840 1449.410 ;
        RECT 409.040 1449.090 409.300 1449.410 ;
        RECT 409.100 1435.325 409.240 1449.090 ;
        RECT 408.110 1434.955 408.390 1435.325 ;
        RECT 409.030 1434.955 409.310 1435.325 ;
        RECT 408.180 1393.990 408.320 1434.955 ;
        RECT 408.120 1393.670 408.380 1393.990 ;
        RECT 408.580 1393.330 408.840 1393.650 ;
        RECT 408.640 1380.050 408.780 1393.330 ;
        RECT 408.580 1379.730 408.840 1380.050 ;
        RECT 409.500 1379.730 409.760 1380.050 ;
        RECT 409.560 1290.485 409.700 1379.730 ;
        RECT 408.570 1290.115 408.850 1290.485 ;
        RECT 409.490 1290.115 409.770 1290.485 ;
        RECT 408.640 1255.270 408.780 1290.115 ;
        RECT 408.580 1254.950 408.840 1255.270 ;
        RECT 408.580 1254.270 408.840 1254.590 ;
        RECT 408.640 1207.670 408.780 1254.270 ;
        RECT 408.580 1207.350 408.840 1207.670 ;
        RECT 409.040 1207.010 409.300 1207.330 ;
        RECT 409.100 1173.330 409.240 1207.010 ;
        RECT 409.040 1173.010 409.300 1173.330 ;
        RECT 409.040 1172.330 409.300 1172.650 ;
        RECT 409.100 1111.110 409.240 1172.330 ;
        RECT 408.580 1110.965 408.840 1111.110 ;
        RECT 408.570 1110.595 408.850 1110.965 ;
        RECT 409.040 1110.790 409.300 1111.110 ;
        RECT 409.030 1109.915 409.310 1110.285 ;
        RECT 409.100 1027.890 409.240 1109.915 ;
        RECT 408.640 1027.750 409.240 1027.890 ;
        RECT 408.640 980.210 408.780 1027.750 ;
        RECT 408.580 979.890 408.840 980.210 ;
        RECT 409.040 979.550 409.300 979.870 ;
        RECT 409.100 931.330 409.240 979.550 ;
        RECT 408.640 931.190 409.240 931.330 ;
        RECT 408.640 917.845 408.780 931.190 ;
        RECT 408.570 917.475 408.850 917.845 ;
        RECT 409.490 917.475 409.770 917.845 ;
        RECT 409.560 869.710 409.700 917.475 ;
        RECT 409.040 869.390 409.300 869.710 ;
        RECT 409.500 869.390 409.760 869.710 ;
        RECT 409.100 838.430 409.240 869.390 ;
        RECT 409.040 838.110 409.300 838.430 ;
        RECT 409.960 838.110 410.220 838.430 ;
        RECT 410.020 814.370 410.160 838.110 ;
        RECT 409.560 814.230 410.160 814.370 ;
        RECT 409.560 807.150 409.700 814.230 ;
        RECT 409.500 806.830 409.760 807.150 ;
        RECT 409.500 723.870 409.760 724.190 ;
        RECT 409.560 717.730 409.700 723.870 ;
        RECT 409.500 717.410 409.760 717.730 ;
        RECT 410.420 717.410 410.680 717.730 ;
        RECT 410.480 669.645 410.620 717.410 ;
        RECT 409.490 669.275 409.770 669.645 ;
        RECT 410.410 669.275 410.690 669.645 ;
        RECT 409.560 628.165 409.700 669.275 ;
        RECT 408.570 627.795 408.850 628.165 ;
        RECT 409.490 627.795 409.770 628.165 ;
        RECT 408.640 603.570 408.780 627.795 ;
        RECT 408.640 603.430 409.240 603.570 ;
        RECT 409.100 545.690 409.240 603.430 ;
        RECT 409.040 545.370 409.300 545.690 ;
        RECT 408.580 544.690 408.840 545.010 ;
        RECT 408.640 483.210 408.780 544.690 ;
        RECT 408.640 483.070 409.240 483.210 ;
        RECT 409.100 435.725 409.240 483.070 ;
        RECT 409.030 435.355 409.310 435.725 ;
        RECT 408.570 434.675 408.850 435.045 ;
        RECT 408.640 427.710 408.780 434.675 ;
        RECT 408.580 427.390 408.840 427.710 ;
        RECT 409.040 379.450 409.300 379.770 ;
        RECT 409.100 352.570 409.240 379.450 ;
        RECT 409.040 352.250 409.300 352.570 ;
        RECT 409.040 351.570 409.300 351.890 ;
        RECT 409.100 331.685 409.240 351.570 ;
        RECT 409.030 331.315 409.310 331.685 ;
        RECT 409.030 329.955 409.310 330.325 ;
        RECT 409.100 259.070 409.240 329.955 ;
        RECT 409.040 258.750 409.300 259.070 ;
        RECT 409.040 193.130 409.300 193.450 ;
        RECT 409.100 176.530 409.240 193.130 ;
        RECT 408.640 176.390 409.240 176.530 ;
        RECT 408.640 158.170 408.780 176.390 ;
        RECT 408.640 158.030 409.700 158.170 ;
        RECT 409.560 110.570 409.700 158.030 ;
        RECT 408.640 110.430 409.700 110.570 ;
        RECT 408.640 62.290 408.780 110.430 ;
        RECT 408.640 62.150 409.240 62.290 ;
        RECT 409.100 20.390 409.240 62.150 ;
        RECT 174.900 20.070 175.160 20.390 ;
        RECT 409.040 20.070 409.300 20.390 ;
        RECT 174.960 2.400 175.100 20.070 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 408.110 1435.000 408.390 1435.280 ;
        RECT 409.030 1435.000 409.310 1435.280 ;
        RECT 408.570 1290.160 408.850 1290.440 ;
        RECT 409.490 1290.160 409.770 1290.440 ;
        RECT 408.570 1110.640 408.850 1110.920 ;
        RECT 409.030 1109.960 409.310 1110.240 ;
        RECT 408.570 917.520 408.850 917.800 ;
        RECT 409.490 917.520 409.770 917.800 ;
        RECT 409.490 669.320 409.770 669.600 ;
        RECT 410.410 669.320 410.690 669.600 ;
        RECT 408.570 627.840 408.850 628.120 ;
        RECT 409.490 627.840 409.770 628.120 ;
        RECT 409.030 435.400 409.310 435.680 ;
        RECT 408.570 434.720 408.850 435.000 ;
        RECT 409.030 331.360 409.310 331.640 ;
        RECT 409.030 330.000 409.310 330.280 ;
      LAYER met3 ;
        RECT 408.085 1435.290 408.415 1435.305 ;
        RECT 409.005 1435.290 409.335 1435.305 ;
        RECT 408.085 1434.990 409.335 1435.290 ;
        RECT 408.085 1434.975 408.415 1434.990 ;
        RECT 409.005 1434.975 409.335 1434.990 ;
        RECT 408.545 1290.450 408.875 1290.465 ;
        RECT 409.465 1290.450 409.795 1290.465 ;
        RECT 408.545 1290.150 409.795 1290.450 ;
        RECT 408.545 1290.135 408.875 1290.150 ;
        RECT 409.465 1290.135 409.795 1290.150 ;
        RECT 408.545 1110.930 408.875 1110.945 ;
        RECT 408.545 1110.615 409.090 1110.930 ;
        RECT 408.790 1110.265 409.090 1110.615 ;
        RECT 408.790 1109.950 409.335 1110.265 ;
        RECT 409.005 1109.935 409.335 1109.950 ;
        RECT 408.545 917.810 408.875 917.825 ;
        RECT 409.465 917.810 409.795 917.825 ;
        RECT 408.545 917.510 409.795 917.810 ;
        RECT 408.545 917.495 408.875 917.510 ;
        RECT 409.465 917.495 409.795 917.510 ;
        RECT 409.465 669.610 409.795 669.625 ;
        RECT 410.385 669.610 410.715 669.625 ;
        RECT 409.465 669.310 410.715 669.610 ;
        RECT 409.465 669.295 409.795 669.310 ;
        RECT 410.385 669.295 410.715 669.310 ;
        RECT 408.545 628.130 408.875 628.145 ;
        RECT 409.465 628.130 409.795 628.145 ;
        RECT 408.545 627.830 409.795 628.130 ;
        RECT 408.545 627.815 408.875 627.830 ;
        RECT 409.465 627.815 409.795 627.830 ;
        RECT 409.005 435.690 409.335 435.705 ;
        RECT 408.790 435.375 409.335 435.690 ;
        RECT 408.790 435.025 409.090 435.375 ;
        RECT 408.545 434.710 409.090 435.025 ;
        RECT 408.545 434.695 408.875 434.710 ;
        RECT 409.005 331.650 409.335 331.665 ;
        RECT 407.870 331.350 409.335 331.650 ;
        RECT 407.870 330.290 408.170 331.350 ;
        RECT 409.005 331.335 409.335 331.350 ;
        RECT 409.005 330.290 409.335 330.305 ;
        RECT 407.870 329.990 409.335 330.290 ;
        RECT 409.005 329.975 409.335 329.990 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 375.505 1590.265 375.675 1592.475 ;
      LAYER mcon ;
        RECT 375.505 1592.305 375.675 1592.475 ;
      LAYER met1 ;
        RECT 192.810 1592.460 193.130 1592.520 ;
        RECT 375.445 1592.460 375.735 1592.505 ;
        RECT 192.810 1592.320 375.735 1592.460 ;
        RECT 192.810 1592.260 193.130 1592.320 ;
        RECT 375.445 1592.275 375.735 1592.320 ;
        RECT 375.445 1590.420 375.735 1590.465 ;
        RECT 416.830 1590.420 417.150 1590.480 ;
        RECT 375.445 1590.280 417.150 1590.420 ;
        RECT 375.445 1590.235 375.735 1590.280 ;
        RECT 416.830 1590.220 417.150 1590.280 ;
      LAYER via ;
        RECT 192.840 1592.260 193.100 1592.520 ;
        RECT 416.860 1590.220 417.120 1590.480 ;
      LAYER met2 ;
        RECT 416.720 1600.380 417.000 1604.000 ;
        RECT 416.720 1600.000 417.060 1600.380 ;
        RECT 192.840 1592.230 193.100 1592.550 ;
        RECT 192.900 2.400 193.040 1592.230 ;
        RECT 416.920 1590.510 417.060 1600.000 ;
        RECT 416.860 1590.190 417.120 1590.510 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 422.700 1600.450 422.980 1604.000 ;
        RECT 421.520 1600.310 422.980 1600.450 ;
        RECT 421.520 20.245 421.660 1600.310 ;
        RECT 422.700 1600.000 422.980 1600.310 ;
        RECT 210.770 19.875 211.050 20.245 ;
        RECT 421.450 19.875 421.730 20.245 ;
        RECT 210.840 2.400 210.980 19.875 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 210.770 19.920 211.050 20.200 ;
        RECT 421.450 19.920 421.730 20.200 ;
      LAYER met3 ;
        RECT 210.745 20.210 211.075 20.225 ;
        RECT 421.425 20.210 421.755 20.225 ;
        RECT 210.745 19.910 421.755 20.210 ;
        RECT 210.745 19.895 211.075 19.910 ;
        RECT 421.425 19.895 421.755 19.910 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 234.210 1593.480 234.530 1593.540 ;
        RECT 429.250 1593.480 429.570 1593.540 ;
        RECT 234.210 1593.340 429.570 1593.480 ;
        RECT 234.210 1593.280 234.530 1593.340 ;
        RECT 429.250 1593.280 429.570 1593.340 ;
        RECT 228.690 16.220 229.010 16.280 ;
        RECT 234.210 16.220 234.530 16.280 ;
        RECT 228.690 16.080 234.530 16.220 ;
        RECT 228.690 16.020 229.010 16.080 ;
        RECT 234.210 16.020 234.530 16.080 ;
      LAYER via ;
        RECT 234.240 1593.280 234.500 1593.540 ;
        RECT 429.280 1593.280 429.540 1593.540 ;
        RECT 228.720 16.020 228.980 16.280 ;
        RECT 234.240 16.020 234.500 16.280 ;
      LAYER met2 ;
        RECT 429.140 1600.380 429.420 1604.000 ;
        RECT 429.140 1600.000 429.480 1600.380 ;
        RECT 429.340 1593.570 429.480 1600.000 ;
        RECT 234.240 1593.250 234.500 1593.570 ;
        RECT 429.280 1593.250 429.540 1593.570 ;
        RECT 234.300 16.310 234.440 1593.250 ;
        RECT 228.720 15.990 228.980 16.310 ;
        RECT 234.240 15.990 234.500 16.310 ;
        RECT 228.780 2.400 228.920 15.990 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 367.225 1207.425 367.395 1263.015 ;
        RECT 367.225 724.285 367.395 765.935 ;
        RECT 367.685 657.645 367.855 717.315 ;
        RECT 367.685 476.085 367.855 531.335 ;
        RECT 367.225 379.525 367.395 427.635 ;
        RECT 367.225 186.405 367.395 234.515 ;
        RECT 367.225 144.925 367.395 181.475 ;
        RECT 366.765 41.565 366.935 89.675 ;
      LAYER mcon ;
        RECT 367.225 1262.845 367.395 1263.015 ;
        RECT 367.225 765.765 367.395 765.935 ;
        RECT 367.685 717.145 367.855 717.315 ;
        RECT 367.685 531.165 367.855 531.335 ;
        RECT 367.225 427.465 367.395 427.635 ;
        RECT 367.225 234.345 367.395 234.515 ;
        RECT 367.225 181.305 367.395 181.475 ;
        RECT 366.765 89.505 366.935 89.675 ;
      LAYER met1 ;
        RECT 367.610 1539.080 367.930 1539.140 ;
        RECT 368.070 1539.080 368.390 1539.140 ;
        RECT 367.610 1538.940 368.390 1539.080 ;
        RECT 367.610 1538.880 367.930 1538.940 ;
        RECT 368.070 1538.880 368.390 1538.940 ;
        RECT 367.150 1497.260 367.470 1497.320 ;
        RECT 367.610 1497.260 367.930 1497.320 ;
        RECT 367.150 1497.120 367.930 1497.260 ;
        RECT 367.150 1497.060 367.470 1497.120 ;
        RECT 367.610 1497.060 367.930 1497.120 ;
        RECT 367.150 1490.460 367.470 1490.520 ;
        RECT 367.610 1490.460 367.930 1490.520 ;
        RECT 367.150 1490.320 367.930 1490.460 ;
        RECT 367.150 1490.260 367.470 1490.320 ;
        RECT 367.610 1490.260 367.930 1490.320 ;
        RECT 367.150 1394.240 367.470 1394.300 ;
        RECT 367.610 1394.240 367.930 1394.300 ;
        RECT 367.150 1394.100 367.930 1394.240 ;
        RECT 367.150 1394.040 367.470 1394.100 ;
        RECT 367.610 1394.040 367.930 1394.100 ;
        RECT 367.150 1338.820 367.470 1338.880 ;
        RECT 368.070 1338.820 368.390 1338.880 ;
        RECT 367.150 1338.680 368.390 1338.820 ;
        RECT 367.150 1338.620 367.470 1338.680 ;
        RECT 368.070 1338.620 368.390 1338.680 ;
        RECT 367.150 1317.880 367.470 1318.140 ;
        RECT 367.240 1317.400 367.380 1317.880 ;
        RECT 367.610 1317.400 367.930 1317.460 ;
        RECT 367.240 1317.260 367.930 1317.400 ;
        RECT 367.610 1317.200 367.930 1317.260 ;
        RECT 367.165 1263.000 367.455 1263.045 ;
        RECT 367.610 1263.000 367.930 1263.060 ;
        RECT 367.165 1262.860 367.930 1263.000 ;
        RECT 367.165 1262.815 367.455 1262.860 ;
        RECT 367.610 1262.800 367.930 1262.860 ;
        RECT 367.165 1207.580 367.455 1207.625 ;
        RECT 368.530 1207.580 368.850 1207.640 ;
        RECT 367.165 1207.440 368.850 1207.580 ;
        RECT 367.165 1207.395 367.455 1207.440 ;
        RECT 368.530 1207.380 368.850 1207.440 ;
        RECT 367.150 1159.300 367.470 1159.360 ;
        RECT 368.530 1159.300 368.850 1159.360 ;
        RECT 367.150 1159.160 368.850 1159.300 ;
        RECT 367.150 1159.100 367.470 1159.160 ;
        RECT 368.530 1159.100 368.850 1159.160 ;
        RECT 367.150 1062.740 367.470 1062.800 ;
        RECT 368.530 1062.740 368.850 1062.800 ;
        RECT 367.150 1062.600 368.850 1062.740 ;
        RECT 367.150 1062.540 367.470 1062.600 ;
        RECT 368.530 1062.540 368.850 1062.600 ;
        RECT 367.150 966.180 367.470 966.240 ;
        RECT 368.530 966.180 368.850 966.240 ;
        RECT 367.150 966.040 368.850 966.180 ;
        RECT 367.150 965.980 367.470 966.040 ;
        RECT 368.530 965.980 368.850 966.040 ;
        RECT 366.690 959.040 367.010 959.100 ;
        RECT 367.150 959.040 367.470 959.100 ;
        RECT 366.690 958.900 367.470 959.040 ;
        RECT 366.690 958.840 367.010 958.900 ;
        RECT 367.150 958.840 367.470 958.900 ;
        RECT 367.150 869.620 367.470 869.680 ;
        RECT 368.070 869.620 368.390 869.680 ;
        RECT 367.150 869.480 368.390 869.620 ;
        RECT 367.150 869.420 367.470 869.480 ;
        RECT 368.070 869.420 368.390 869.480 ;
        RECT 366.690 862.480 367.010 862.540 ;
        RECT 367.150 862.480 367.470 862.540 ;
        RECT 366.690 862.340 367.470 862.480 ;
        RECT 366.690 862.280 367.010 862.340 ;
        RECT 367.150 862.280 367.470 862.340 ;
        RECT 367.610 773.060 367.930 773.120 ;
        RECT 368.070 773.060 368.390 773.120 ;
        RECT 367.610 772.920 368.390 773.060 ;
        RECT 367.610 772.860 367.930 772.920 ;
        RECT 368.070 772.860 368.390 772.920 ;
        RECT 367.150 765.920 367.470 765.980 ;
        RECT 366.955 765.780 367.470 765.920 ;
        RECT 367.150 765.720 367.470 765.780 ;
        RECT 367.150 724.440 367.470 724.500 ;
        RECT 366.955 724.300 367.470 724.440 ;
        RECT 367.150 724.240 367.470 724.300 ;
        RECT 367.610 717.300 367.930 717.360 ;
        RECT 367.415 717.160 367.930 717.300 ;
        RECT 367.610 717.100 367.930 717.160 ;
        RECT 367.625 657.800 367.915 657.845 ;
        RECT 368.070 657.800 368.390 657.860 ;
        RECT 367.625 657.660 368.390 657.800 ;
        RECT 367.625 657.615 367.915 657.660 ;
        RECT 368.070 657.600 368.390 657.660 ;
        RECT 367.150 572.800 367.470 572.860 ;
        RECT 367.610 572.800 367.930 572.860 ;
        RECT 367.150 572.660 367.930 572.800 ;
        RECT 367.150 572.600 367.470 572.660 ;
        RECT 367.610 572.600 367.930 572.660 ;
        RECT 367.610 531.320 367.930 531.380 ;
        RECT 367.415 531.180 367.930 531.320 ;
        RECT 367.610 531.120 367.930 531.180 ;
        RECT 367.625 476.240 367.915 476.285 ;
        RECT 368.070 476.240 368.390 476.300 ;
        RECT 367.625 476.100 368.390 476.240 ;
        RECT 367.625 476.055 367.915 476.100 ;
        RECT 368.070 476.040 368.390 476.100 ;
        RECT 367.150 427.620 367.470 427.680 ;
        RECT 366.955 427.480 367.470 427.620 ;
        RECT 367.150 427.420 367.470 427.480 ;
        RECT 367.165 379.680 367.455 379.725 ;
        RECT 367.610 379.680 367.930 379.740 ;
        RECT 367.165 379.540 367.930 379.680 ;
        RECT 367.165 379.495 367.455 379.540 ;
        RECT 367.610 379.480 367.930 379.540 ;
        RECT 367.150 241.780 367.470 242.040 ;
        RECT 367.240 241.640 367.380 241.780 ;
        RECT 367.610 241.640 367.930 241.700 ;
        RECT 367.240 241.500 367.930 241.640 ;
        RECT 367.610 241.440 367.930 241.500 ;
        RECT 367.165 234.500 367.455 234.545 ;
        RECT 367.610 234.500 367.930 234.560 ;
        RECT 367.165 234.360 367.930 234.500 ;
        RECT 367.165 234.315 367.455 234.360 ;
        RECT 367.610 234.300 367.930 234.360 ;
        RECT 367.150 186.560 367.470 186.620 ;
        RECT 366.955 186.420 367.470 186.560 ;
        RECT 367.150 186.360 367.470 186.420 ;
        RECT 367.150 181.460 367.470 181.520 ;
        RECT 366.955 181.320 367.470 181.460 ;
        RECT 367.150 181.260 367.470 181.320 ;
        RECT 367.165 145.080 367.455 145.125 ;
        RECT 367.610 145.080 367.930 145.140 ;
        RECT 367.165 144.940 367.930 145.080 ;
        RECT 367.165 144.895 367.455 144.940 ;
        RECT 367.610 144.880 367.930 144.940 ;
        RECT 366.705 89.660 366.995 89.705 ;
        RECT 367.150 89.660 367.470 89.720 ;
        RECT 366.705 89.520 367.470 89.660 ;
        RECT 366.705 89.475 366.995 89.520 ;
        RECT 367.150 89.460 367.470 89.520 ;
        RECT 366.690 41.720 367.010 41.780 ;
        RECT 366.495 41.580 367.010 41.720 ;
        RECT 366.690 41.520 367.010 41.580 ;
      LAYER via ;
        RECT 367.640 1538.880 367.900 1539.140 ;
        RECT 368.100 1538.880 368.360 1539.140 ;
        RECT 367.180 1497.060 367.440 1497.320 ;
        RECT 367.640 1497.060 367.900 1497.320 ;
        RECT 367.180 1490.260 367.440 1490.520 ;
        RECT 367.640 1490.260 367.900 1490.520 ;
        RECT 367.180 1394.040 367.440 1394.300 ;
        RECT 367.640 1394.040 367.900 1394.300 ;
        RECT 367.180 1338.620 367.440 1338.880 ;
        RECT 368.100 1338.620 368.360 1338.880 ;
        RECT 367.180 1317.880 367.440 1318.140 ;
        RECT 367.640 1317.200 367.900 1317.460 ;
        RECT 367.640 1262.800 367.900 1263.060 ;
        RECT 368.560 1207.380 368.820 1207.640 ;
        RECT 367.180 1159.100 367.440 1159.360 ;
        RECT 368.560 1159.100 368.820 1159.360 ;
        RECT 367.180 1062.540 367.440 1062.800 ;
        RECT 368.560 1062.540 368.820 1062.800 ;
        RECT 367.180 965.980 367.440 966.240 ;
        RECT 368.560 965.980 368.820 966.240 ;
        RECT 366.720 958.840 366.980 959.100 ;
        RECT 367.180 958.840 367.440 959.100 ;
        RECT 367.180 869.420 367.440 869.680 ;
        RECT 368.100 869.420 368.360 869.680 ;
        RECT 366.720 862.280 366.980 862.540 ;
        RECT 367.180 862.280 367.440 862.540 ;
        RECT 367.640 772.860 367.900 773.120 ;
        RECT 368.100 772.860 368.360 773.120 ;
        RECT 367.180 765.720 367.440 765.980 ;
        RECT 367.180 724.240 367.440 724.500 ;
        RECT 367.640 717.100 367.900 717.360 ;
        RECT 368.100 657.600 368.360 657.860 ;
        RECT 367.180 572.600 367.440 572.860 ;
        RECT 367.640 572.600 367.900 572.860 ;
        RECT 367.640 531.120 367.900 531.380 ;
        RECT 368.100 476.040 368.360 476.300 ;
        RECT 367.180 427.420 367.440 427.680 ;
        RECT 367.640 379.480 367.900 379.740 ;
        RECT 367.180 241.780 367.440 242.040 ;
        RECT 367.640 241.440 367.900 241.700 ;
        RECT 367.640 234.300 367.900 234.560 ;
        RECT 367.180 186.360 367.440 186.620 ;
        RECT 367.180 181.260 367.440 181.520 ;
        RECT 367.640 144.880 367.900 145.140 ;
        RECT 367.180 89.460 367.440 89.720 ;
        RECT 366.720 41.520 366.980 41.780 ;
      LAYER met2 ;
        RECT 367.040 1600.450 367.320 1604.000 ;
        RECT 367.040 1600.310 367.840 1600.450 ;
        RECT 367.040 1600.000 367.320 1600.310 ;
        RECT 367.700 1552.850 367.840 1600.310 ;
        RECT 367.700 1552.710 368.300 1552.850 ;
        RECT 368.160 1539.170 368.300 1552.710 ;
        RECT 367.640 1538.850 367.900 1539.170 ;
        RECT 368.100 1538.850 368.360 1539.170 ;
        RECT 367.700 1497.350 367.840 1538.850 ;
        RECT 367.180 1497.030 367.440 1497.350 ;
        RECT 367.640 1497.030 367.900 1497.350 ;
        RECT 367.240 1490.550 367.380 1497.030 ;
        RECT 367.180 1490.230 367.440 1490.550 ;
        RECT 367.640 1490.230 367.900 1490.550 ;
        RECT 367.700 1394.330 367.840 1490.230 ;
        RECT 367.180 1394.010 367.440 1394.330 ;
        RECT 367.640 1394.010 367.900 1394.330 ;
        RECT 367.240 1387.045 367.380 1394.010 ;
        RECT 367.170 1386.675 367.450 1387.045 ;
        RECT 368.090 1386.675 368.370 1387.045 ;
        RECT 368.160 1338.910 368.300 1386.675 ;
        RECT 367.180 1338.590 367.440 1338.910 ;
        RECT 368.100 1338.590 368.360 1338.910 ;
        RECT 367.240 1318.170 367.380 1338.590 ;
        RECT 367.180 1317.850 367.440 1318.170 ;
        RECT 367.640 1317.170 367.900 1317.490 ;
        RECT 367.700 1263.090 367.840 1317.170 ;
        RECT 367.640 1262.770 367.900 1263.090 ;
        RECT 368.560 1207.350 368.820 1207.670 ;
        RECT 368.620 1159.390 368.760 1207.350 ;
        RECT 367.180 1159.245 367.440 1159.390 ;
        RECT 368.560 1159.245 368.820 1159.390 ;
        RECT 367.170 1158.875 367.450 1159.245 ;
        RECT 368.550 1158.875 368.830 1159.245 ;
        RECT 368.620 1062.830 368.760 1158.875 ;
        RECT 367.180 1062.685 367.440 1062.830 ;
        RECT 368.560 1062.685 368.820 1062.830 ;
        RECT 367.170 1062.315 367.450 1062.685 ;
        RECT 368.550 1062.315 368.830 1062.685 ;
        RECT 368.620 966.270 368.760 1062.315 ;
        RECT 367.180 965.950 367.440 966.270 ;
        RECT 368.560 965.950 368.820 966.270 ;
        RECT 367.240 959.130 367.380 965.950 ;
        RECT 366.720 958.810 366.980 959.130 ;
        RECT 367.180 958.810 367.440 959.130 ;
        RECT 366.780 911.045 366.920 958.810 ;
        RECT 366.710 910.675 366.990 911.045 ;
        RECT 368.090 910.675 368.370 911.045 ;
        RECT 368.160 869.710 368.300 910.675 ;
        RECT 367.180 869.390 367.440 869.710 ;
        RECT 368.100 869.390 368.360 869.710 ;
        RECT 367.240 862.570 367.380 869.390 ;
        RECT 366.720 862.250 366.980 862.570 ;
        RECT 367.180 862.250 367.440 862.570 ;
        RECT 366.780 814.485 366.920 862.250 ;
        RECT 366.710 814.115 366.990 814.485 ;
        RECT 368.090 814.115 368.370 814.485 ;
        RECT 368.160 773.150 368.300 814.115 ;
        RECT 367.640 772.890 367.900 773.150 ;
        RECT 367.240 772.830 367.900 772.890 ;
        RECT 368.100 772.830 368.360 773.150 ;
        RECT 367.240 772.750 367.840 772.830 ;
        RECT 367.240 766.010 367.380 772.750 ;
        RECT 367.180 765.690 367.440 766.010 ;
        RECT 367.180 724.210 367.440 724.530 ;
        RECT 367.240 717.810 367.380 724.210 ;
        RECT 367.240 717.670 367.840 717.810 ;
        RECT 367.700 717.390 367.840 717.670 ;
        RECT 367.640 717.070 367.900 717.390 ;
        RECT 368.100 657.570 368.360 657.890 ;
        RECT 368.160 580.450 368.300 657.570 ;
        RECT 367.700 580.310 368.300 580.450 ;
        RECT 367.700 572.890 367.840 580.310 ;
        RECT 367.180 572.570 367.440 572.890 ;
        RECT 367.640 572.570 367.900 572.890 ;
        RECT 367.240 544.410 367.380 572.570 ;
        RECT 367.240 544.270 367.840 544.410 ;
        RECT 367.700 531.410 367.840 544.270 ;
        RECT 367.640 531.090 367.900 531.410 ;
        RECT 368.100 476.010 368.360 476.330 ;
        RECT 368.160 435.045 368.300 476.010 ;
        RECT 367.170 434.675 367.450 435.045 ;
        RECT 368.090 434.675 368.370 435.045 ;
        RECT 367.240 427.710 367.380 434.675 ;
        RECT 367.180 427.390 367.440 427.710 ;
        RECT 367.640 379.450 367.900 379.770 ;
        RECT 367.700 313.890 367.840 379.450 ;
        RECT 367.240 313.750 367.840 313.890 ;
        RECT 367.240 242.070 367.380 313.750 ;
        RECT 367.180 241.750 367.440 242.070 ;
        RECT 367.640 241.410 367.900 241.730 ;
        RECT 367.700 234.590 367.840 241.410 ;
        RECT 367.640 234.270 367.900 234.590 ;
        RECT 367.180 186.330 367.440 186.650 ;
        RECT 367.240 181.550 367.380 186.330 ;
        RECT 367.180 181.230 367.440 181.550 ;
        RECT 367.640 144.850 367.900 145.170 ;
        RECT 367.700 113.290 367.840 144.850 ;
        RECT 367.240 113.150 367.840 113.290 ;
        RECT 367.240 89.750 367.380 113.150 ;
        RECT 367.180 89.430 367.440 89.750 ;
        RECT 366.720 41.490 366.980 41.810 ;
        RECT 366.780 17.525 366.920 41.490 ;
        RECT 50.230 17.155 50.510 17.525 ;
        RECT 366.710 17.155 366.990 17.525 ;
        RECT 50.300 2.400 50.440 17.155 ;
        RECT 50.090 -4.800 50.650 2.400 ;
      LAYER via2 ;
        RECT 367.170 1386.720 367.450 1387.000 ;
        RECT 368.090 1386.720 368.370 1387.000 ;
        RECT 367.170 1158.920 367.450 1159.200 ;
        RECT 368.550 1158.920 368.830 1159.200 ;
        RECT 367.170 1062.360 367.450 1062.640 ;
        RECT 368.550 1062.360 368.830 1062.640 ;
        RECT 366.710 910.720 366.990 911.000 ;
        RECT 368.090 910.720 368.370 911.000 ;
        RECT 366.710 814.160 366.990 814.440 ;
        RECT 368.090 814.160 368.370 814.440 ;
        RECT 367.170 434.720 367.450 435.000 ;
        RECT 368.090 434.720 368.370 435.000 ;
        RECT 50.230 17.200 50.510 17.480 ;
        RECT 366.710 17.200 366.990 17.480 ;
      LAYER met3 ;
        RECT 367.145 1387.010 367.475 1387.025 ;
        RECT 368.065 1387.010 368.395 1387.025 ;
        RECT 367.145 1386.710 368.395 1387.010 ;
        RECT 367.145 1386.695 367.475 1386.710 ;
        RECT 368.065 1386.695 368.395 1386.710 ;
        RECT 367.145 1159.210 367.475 1159.225 ;
        RECT 368.525 1159.210 368.855 1159.225 ;
        RECT 367.145 1158.910 368.855 1159.210 ;
        RECT 367.145 1158.895 367.475 1158.910 ;
        RECT 368.525 1158.895 368.855 1158.910 ;
        RECT 367.145 1062.650 367.475 1062.665 ;
        RECT 368.525 1062.650 368.855 1062.665 ;
        RECT 367.145 1062.350 368.855 1062.650 ;
        RECT 367.145 1062.335 367.475 1062.350 ;
        RECT 368.525 1062.335 368.855 1062.350 ;
        RECT 366.685 911.010 367.015 911.025 ;
        RECT 368.065 911.010 368.395 911.025 ;
        RECT 366.685 910.710 368.395 911.010 ;
        RECT 366.685 910.695 367.015 910.710 ;
        RECT 368.065 910.695 368.395 910.710 ;
        RECT 366.685 814.450 367.015 814.465 ;
        RECT 368.065 814.450 368.395 814.465 ;
        RECT 366.685 814.150 368.395 814.450 ;
        RECT 366.685 814.135 367.015 814.150 ;
        RECT 368.065 814.135 368.395 814.150 ;
        RECT 367.145 435.010 367.475 435.025 ;
        RECT 368.065 435.010 368.395 435.025 ;
        RECT 367.145 434.710 368.395 435.010 ;
        RECT 367.145 434.695 367.475 434.710 ;
        RECT 368.065 434.695 368.395 434.710 ;
        RECT 50.205 17.490 50.535 17.505 ;
        RECT 366.685 17.490 367.015 17.505 ;
        RECT 50.205 17.190 367.015 17.490 ;
        RECT 50.205 17.175 50.535 17.190 ;
        RECT 366.685 17.175 367.015 17.190 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 1589.740 255.230 1589.800 ;
        RECT 437.530 1589.740 437.850 1589.800 ;
        RECT 254.910 1589.600 437.850 1589.740 ;
        RECT 254.910 1589.540 255.230 1589.600 ;
        RECT 437.530 1589.540 437.850 1589.600 ;
        RECT 252.610 16.220 252.930 16.280 ;
        RECT 254.910 16.220 255.230 16.280 ;
        RECT 252.610 16.080 255.230 16.220 ;
        RECT 252.610 16.020 252.930 16.080 ;
        RECT 254.910 16.020 255.230 16.080 ;
      LAYER via ;
        RECT 254.940 1589.540 255.200 1589.800 ;
        RECT 437.560 1589.540 437.820 1589.800 ;
        RECT 252.640 16.020 252.900 16.280 ;
        RECT 254.940 16.020 255.200 16.280 ;
      LAYER met2 ;
        RECT 437.420 1600.380 437.700 1604.000 ;
        RECT 437.420 1600.000 437.760 1600.380 ;
        RECT 437.620 1589.830 437.760 1600.000 ;
        RECT 254.940 1589.510 255.200 1589.830 ;
        RECT 437.560 1589.510 437.820 1589.830 ;
        RECT 255.000 16.310 255.140 1589.510 ;
        RECT 252.640 15.990 252.900 16.310 ;
        RECT 254.940 15.990 255.200 16.310 ;
        RECT 252.700 2.400 252.840 15.990 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 412.690 16.900 413.010 16.960 ;
        RECT 442.130 16.900 442.450 16.960 ;
        RECT 412.690 16.760 442.450 16.900 ;
        RECT 412.690 16.700 413.010 16.760 ;
        RECT 442.130 16.700 442.450 16.760 ;
        RECT 270.090 15.880 270.410 15.940 ;
        RECT 400.730 15.880 401.050 15.940 ;
        RECT 270.090 15.740 401.050 15.880 ;
        RECT 270.090 15.680 270.410 15.740 ;
        RECT 400.730 15.680 401.050 15.740 ;
      LAYER via ;
        RECT 412.720 16.700 412.980 16.960 ;
        RECT 442.160 16.700 442.420 16.960 ;
        RECT 270.120 15.680 270.380 15.940 ;
        RECT 400.760 15.680 401.020 15.940 ;
      LAYER met2 ;
        RECT 443.400 1600.450 443.680 1604.000 ;
        RECT 442.680 1600.310 443.680 1600.450 ;
        RECT 442.680 17.410 442.820 1600.310 ;
        RECT 443.400 1600.000 443.680 1600.310 ;
        RECT 442.220 17.270 442.820 17.410 ;
        RECT 442.220 16.990 442.360 17.270 ;
        RECT 412.720 16.845 412.980 16.990 ;
        RECT 400.750 16.475 401.030 16.845 ;
        RECT 412.710 16.475 412.990 16.845 ;
        RECT 442.160 16.670 442.420 16.990 ;
        RECT 400.820 15.970 400.960 16.475 ;
        RECT 270.120 15.650 270.380 15.970 ;
        RECT 400.760 15.650 401.020 15.970 ;
        RECT 270.180 2.400 270.320 15.650 ;
        RECT 269.970 -4.800 270.530 2.400 ;
      LAYER via2 ;
        RECT 400.750 16.520 401.030 16.800 ;
        RECT 412.710 16.520 412.990 16.800 ;
      LAYER met3 ;
        RECT 400.725 16.810 401.055 16.825 ;
        RECT 412.685 16.810 413.015 16.825 ;
        RECT 400.725 16.510 413.015 16.810 ;
        RECT 400.725 16.495 401.055 16.510 ;
        RECT 412.685 16.495 413.015 16.510 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 1589.060 289.730 1589.120 ;
        RECT 289.410 1588.920 424.420 1589.060 ;
        RECT 289.410 1588.860 289.730 1588.920 ;
        RECT 424.280 1588.720 424.420 1588.920 ;
        RECT 449.950 1588.720 450.270 1588.780 ;
        RECT 424.280 1588.580 450.270 1588.720 ;
        RECT 449.950 1588.520 450.270 1588.580 ;
      LAYER via ;
        RECT 289.440 1588.860 289.700 1589.120 ;
        RECT 449.980 1588.520 450.240 1588.780 ;
      LAYER met2 ;
        RECT 449.840 1600.380 450.120 1604.000 ;
        RECT 449.840 1600.000 450.180 1600.380 ;
        RECT 289.440 1588.830 289.700 1589.150 ;
        RECT 289.500 17.410 289.640 1588.830 ;
        RECT 450.040 1588.810 450.180 1600.000 ;
        RECT 449.980 1588.490 450.240 1588.810 ;
        RECT 288.120 17.270 289.640 17.410 ;
        RECT 288.120 2.400 288.260 17.270 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 456.390 15.540 456.710 15.600 ;
        RECT 317.560 15.400 456.710 15.540 ;
        RECT 305.970 15.200 306.290 15.260 ;
        RECT 317.560 15.200 317.700 15.400 ;
        RECT 456.390 15.340 456.710 15.400 ;
        RECT 305.970 15.060 317.700 15.200 ;
        RECT 305.970 15.000 306.290 15.060 ;
      LAYER via ;
        RECT 306.000 15.000 306.260 15.260 ;
        RECT 456.420 15.340 456.680 15.600 ;
      LAYER met2 ;
        RECT 455.820 1600.450 456.100 1604.000 ;
        RECT 455.820 1600.310 456.620 1600.450 ;
        RECT 455.820 1600.000 456.100 1600.310 ;
        RECT 456.480 15.630 456.620 1600.310 ;
        RECT 456.420 15.310 456.680 15.630 ;
        RECT 306.000 14.970 306.260 15.290 ;
        RECT 306.060 2.400 306.200 14.970 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 423.805 1587.885 423.975 1588.735 ;
      LAYER mcon ;
        RECT 423.805 1588.565 423.975 1588.735 ;
      LAYER met1 ;
        RECT 323.910 1588.720 324.230 1588.780 ;
        RECT 423.745 1588.720 424.035 1588.765 ;
        RECT 323.910 1588.580 424.035 1588.720 ;
        RECT 323.910 1588.520 324.230 1588.580 ;
        RECT 423.745 1588.535 424.035 1588.580 ;
        RECT 423.745 1588.040 424.035 1588.085 ;
        RECT 462.370 1588.040 462.690 1588.100 ;
        RECT 423.745 1587.900 462.690 1588.040 ;
        RECT 423.745 1587.855 424.035 1587.900 ;
        RECT 462.370 1587.840 462.690 1587.900 ;
      LAYER via ;
        RECT 323.940 1588.520 324.200 1588.780 ;
        RECT 462.400 1587.840 462.660 1588.100 ;
      LAYER met2 ;
        RECT 462.260 1600.380 462.540 1604.000 ;
        RECT 462.260 1600.000 462.600 1600.380 ;
        RECT 323.940 1588.490 324.200 1588.810 ;
        RECT 324.000 2.400 324.140 1588.490 ;
        RECT 462.460 1588.130 462.600 1600.000 ;
        RECT 462.400 1587.810 462.660 1588.130 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 462.830 1579.880 463.150 1579.940 ;
        RECT 466.510 1579.880 466.830 1579.940 ;
        RECT 462.830 1579.740 466.830 1579.880 ;
        RECT 462.830 1579.680 463.150 1579.740 ;
        RECT 466.510 1579.680 466.830 1579.740 ;
        RECT 341.390 14.180 341.710 14.240 ;
        RECT 462.830 14.180 463.150 14.240 ;
        RECT 341.390 14.040 463.150 14.180 ;
        RECT 341.390 13.980 341.710 14.040 ;
        RECT 462.830 13.980 463.150 14.040 ;
      LAYER via ;
        RECT 462.860 1579.680 463.120 1579.940 ;
        RECT 466.540 1579.680 466.800 1579.940 ;
        RECT 341.420 13.980 341.680 14.240 ;
        RECT 462.860 13.980 463.120 14.240 ;
      LAYER met2 ;
        RECT 468.240 1600.450 468.520 1604.000 ;
        RECT 466.600 1600.310 468.520 1600.450 ;
        RECT 466.600 1579.970 466.740 1600.310 ;
        RECT 468.240 1600.000 468.520 1600.310 ;
        RECT 462.860 1579.650 463.120 1579.970 ;
        RECT 466.540 1579.650 466.800 1579.970 ;
        RECT 462.920 14.270 463.060 1579.650 ;
        RECT 341.420 13.950 341.680 14.270 ;
        RECT 462.860 13.950 463.120 14.270 ;
        RECT 341.480 2.400 341.620 13.950 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 399.885 18.445 400.055 19.635 ;
      LAYER mcon ;
        RECT 399.885 19.465 400.055 19.635 ;
      LAYER met1 ;
        RECT 469.730 1580.220 470.050 1580.280 ;
        RECT 472.950 1580.220 473.270 1580.280 ;
        RECT 469.730 1580.080 473.270 1580.220 ;
        RECT 469.730 1580.020 470.050 1580.080 ;
        RECT 472.950 1580.020 473.270 1580.080 ;
        RECT 469.730 385.940 470.050 386.200 ;
        RECT 469.820 385.520 469.960 385.940 ;
        RECT 469.730 385.260 470.050 385.520 ;
        RECT 359.330 19.620 359.650 19.680 ;
        RECT 399.825 19.620 400.115 19.665 ;
        RECT 359.330 19.480 400.115 19.620 ;
        RECT 359.330 19.420 359.650 19.480 ;
        RECT 399.825 19.435 400.115 19.480 ;
        RECT 469.730 18.940 470.050 19.000 ;
        RECT 459.240 18.800 470.050 18.940 ;
        RECT 399.825 18.600 400.115 18.645 ;
        RECT 459.240 18.600 459.380 18.800 ;
        RECT 469.730 18.740 470.050 18.800 ;
        RECT 399.825 18.460 459.380 18.600 ;
        RECT 399.825 18.415 400.115 18.460 ;
      LAYER via ;
        RECT 469.760 1580.020 470.020 1580.280 ;
        RECT 472.980 1580.020 473.240 1580.280 ;
        RECT 469.760 385.940 470.020 386.200 ;
        RECT 469.760 385.260 470.020 385.520 ;
        RECT 359.360 19.420 359.620 19.680 ;
        RECT 469.760 18.740 470.020 19.000 ;
      LAYER met2 ;
        RECT 474.220 1600.450 474.500 1604.000 ;
        RECT 473.040 1600.310 474.500 1600.450 ;
        RECT 473.040 1580.310 473.180 1600.310 ;
        RECT 474.220 1600.000 474.500 1600.310 ;
        RECT 469.760 1579.990 470.020 1580.310 ;
        RECT 472.980 1579.990 473.240 1580.310 ;
        RECT 469.820 386.230 469.960 1579.990 ;
        RECT 469.760 385.910 470.020 386.230 ;
        RECT 469.760 385.230 470.020 385.550 ;
        RECT 359.360 19.390 359.620 19.710 ;
        RECT 359.420 2.400 359.560 19.390 ;
        RECT 469.820 19.030 469.960 385.230 ;
        RECT 469.760 18.710 470.020 19.030 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 476.170 1580.560 476.490 1580.620 ;
        RECT 479.390 1580.560 479.710 1580.620 ;
        RECT 476.170 1580.420 479.710 1580.560 ;
        RECT 476.170 1580.360 476.490 1580.420 ;
        RECT 479.390 1580.360 479.710 1580.420 ;
        RECT 377.270 18.260 377.590 18.320 ;
        RECT 476.170 18.260 476.490 18.320 ;
        RECT 377.270 18.120 476.490 18.260 ;
        RECT 377.270 18.060 377.590 18.120 ;
        RECT 476.170 18.060 476.490 18.120 ;
      LAYER via ;
        RECT 476.200 1580.360 476.460 1580.620 ;
        RECT 479.420 1580.360 479.680 1580.620 ;
        RECT 377.300 18.060 377.560 18.320 ;
        RECT 476.200 18.060 476.460 18.320 ;
      LAYER met2 ;
        RECT 480.660 1600.450 480.940 1604.000 ;
        RECT 479.480 1600.310 480.940 1600.450 ;
        RECT 479.480 1580.650 479.620 1600.310 ;
        RECT 480.660 1600.000 480.940 1600.310 ;
        RECT 476.200 1580.330 476.460 1580.650 ;
        RECT 479.420 1580.330 479.680 1580.650 ;
        RECT 476.260 18.350 476.400 1580.330 ;
        RECT 377.300 18.030 377.560 18.350 ;
        RECT 476.200 18.030 476.460 18.350 ;
        RECT 377.360 2.400 377.500 18.030 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 484.985 235.025 485.155 282.795 ;
        RECT 484.985 186.405 485.155 234.515 ;
        RECT 484.985 109.565 485.155 144.755 ;
      LAYER mcon ;
        RECT 484.985 282.625 485.155 282.795 ;
        RECT 484.985 234.345 485.155 234.515 ;
        RECT 484.985 144.585 485.155 144.755 ;
      LAYER met1 ;
        RECT 484.910 282.780 485.230 282.840 ;
        RECT 484.715 282.640 485.230 282.780 ;
        RECT 484.910 282.580 485.230 282.640 ;
        RECT 484.910 235.180 485.230 235.240 ;
        RECT 484.715 235.040 485.230 235.180 ;
        RECT 484.910 234.980 485.230 235.040 ;
        RECT 484.910 234.500 485.230 234.560 ;
        RECT 484.715 234.360 485.230 234.500 ;
        RECT 484.910 234.300 485.230 234.360 ;
        RECT 484.910 186.560 485.230 186.620 ;
        RECT 484.715 186.420 485.230 186.560 ;
        RECT 484.910 186.360 485.230 186.420 ;
        RECT 484.910 144.740 485.230 144.800 ;
        RECT 484.715 144.600 485.230 144.740 ;
        RECT 484.910 144.540 485.230 144.600 ;
        RECT 484.910 109.720 485.230 109.780 ;
        RECT 484.715 109.580 485.230 109.720 ;
        RECT 484.910 109.520 485.230 109.580 ;
        RECT 484.910 19.620 485.230 19.680 ;
        RECT 409.100 19.480 485.230 19.620 ;
        RECT 395.210 19.280 395.530 19.340 ;
        RECT 409.100 19.280 409.240 19.480 ;
        RECT 484.910 19.420 485.230 19.480 ;
        RECT 395.210 19.140 409.240 19.280 ;
        RECT 395.210 19.080 395.530 19.140 ;
      LAYER via ;
        RECT 484.940 282.580 485.200 282.840 ;
        RECT 484.940 234.980 485.200 235.240 ;
        RECT 484.940 234.300 485.200 234.560 ;
        RECT 484.940 186.360 485.200 186.620 ;
        RECT 484.940 144.540 485.200 144.800 ;
        RECT 484.940 109.520 485.200 109.780 ;
        RECT 395.240 19.080 395.500 19.340 ;
        RECT 484.940 19.420 485.200 19.680 ;
      LAYER met2 ;
        RECT 486.640 1600.450 486.920 1604.000 ;
        RECT 485.920 1600.310 486.920 1600.450 ;
        RECT 485.920 1580.050 486.060 1600.310 ;
        RECT 486.640 1600.000 486.920 1600.310 ;
        RECT 485.000 1579.910 486.060 1580.050 ;
        RECT 485.000 1512.050 485.140 1579.910 ;
        RECT 484.540 1511.910 485.140 1512.050 ;
        RECT 484.540 1511.370 484.680 1511.910 ;
        RECT 484.080 1511.230 484.680 1511.370 ;
        RECT 484.080 1510.690 484.220 1511.230 ;
        RECT 484.080 1510.550 485.140 1510.690 ;
        RECT 485.000 1366.530 485.140 1510.550 ;
        RECT 484.080 1366.390 485.140 1366.530 ;
        RECT 484.080 1365.850 484.220 1366.390 ;
        RECT 484.080 1365.710 485.140 1365.850 ;
        RECT 485.000 1269.970 485.140 1365.710 ;
        RECT 484.080 1269.830 485.140 1269.970 ;
        RECT 484.080 1269.290 484.220 1269.830 ;
        RECT 484.080 1269.150 485.140 1269.290 ;
        RECT 485.000 1173.410 485.140 1269.150 ;
        RECT 484.080 1173.270 485.140 1173.410 ;
        RECT 484.080 1172.730 484.220 1173.270 ;
        RECT 484.080 1172.590 485.140 1172.730 ;
        RECT 485.000 1076.850 485.140 1172.590 ;
        RECT 484.080 1076.710 485.140 1076.850 ;
        RECT 484.080 1076.170 484.220 1076.710 ;
        RECT 484.080 1076.030 485.140 1076.170 ;
        RECT 485.000 980.290 485.140 1076.030 ;
        RECT 484.080 980.150 485.140 980.290 ;
        RECT 484.080 979.610 484.220 980.150 ;
        RECT 484.080 979.470 485.140 979.610 ;
        RECT 485.000 883.730 485.140 979.470 ;
        RECT 484.080 883.590 485.140 883.730 ;
        RECT 484.080 883.050 484.220 883.590 ;
        RECT 484.080 882.910 485.140 883.050 ;
        RECT 485.000 787.170 485.140 882.910 ;
        RECT 484.080 787.030 485.140 787.170 ;
        RECT 484.080 786.490 484.220 787.030 ;
        RECT 484.080 786.350 484.680 786.490 ;
        RECT 484.540 785.810 484.680 786.350 ;
        RECT 484.540 785.670 485.140 785.810 ;
        RECT 485.000 303.805 485.140 785.670 ;
        RECT 484.930 303.435 485.210 303.805 ;
        RECT 484.930 283.035 485.210 283.405 ;
        RECT 485.000 282.870 485.140 283.035 ;
        RECT 484.940 282.550 485.200 282.870 ;
        RECT 484.940 234.950 485.200 235.270 ;
        RECT 485.000 234.590 485.140 234.950 ;
        RECT 484.940 234.270 485.200 234.590 ;
        RECT 484.940 186.330 485.200 186.650 ;
        RECT 485.000 144.830 485.140 186.330 ;
        RECT 484.940 144.510 485.200 144.830 ;
        RECT 484.940 109.490 485.200 109.810 ;
        RECT 485.000 19.710 485.140 109.490 ;
        RECT 484.940 19.390 485.200 19.710 ;
        RECT 395.240 19.050 395.500 19.370 ;
        RECT 395.300 2.400 395.440 19.050 ;
        RECT 395.090 -4.800 395.650 2.400 ;
      LAYER via2 ;
        RECT 484.930 303.480 485.210 303.760 ;
        RECT 484.930 283.080 485.210 283.360 ;
      LAYER met3 ;
        RECT 484.905 303.780 485.235 303.785 ;
        RECT 484.905 303.770 485.490 303.780 ;
        RECT 484.905 303.470 485.690 303.770 ;
        RECT 484.905 303.460 485.490 303.470 ;
        RECT 484.905 303.455 485.235 303.460 ;
        RECT 484.905 283.380 485.235 283.385 ;
        RECT 484.905 283.370 485.490 283.380 ;
        RECT 484.905 283.070 485.690 283.370 ;
        RECT 484.905 283.060 485.490 283.070 ;
        RECT 484.905 283.055 485.235 283.060 ;
      LAYER via3 ;
        RECT 485.140 303.460 485.460 303.780 ;
        RECT 485.140 283.060 485.460 283.380 ;
      LAYER met4 ;
        RECT 485.135 303.455 485.465 303.785 ;
        RECT 485.150 283.385 485.450 303.455 ;
        RECT 485.135 283.055 485.465 283.385 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 424.650 1589.060 424.970 1589.120 ;
        RECT 424.650 1588.920 460.760 1589.060 ;
        RECT 424.650 1588.860 424.970 1588.920 ;
        RECT 460.620 1588.720 460.760 1588.920 ;
        RECT 493.190 1588.720 493.510 1588.780 ;
        RECT 460.620 1588.580 493.510 1588.720 ;
        RECT 493.190 1588.520 493.510 1588.580 ;
        RECT 413.150 20.640 413.470 20.700 ;
        RECT 424.190 20.640 424.510 20.700 ;
        RECT 413.150 20.500 424.510 20.640 ;
        RECT 413.150 20.440 413.470 20.500 ;
        RECT 424.190 20.440 424.510 20.500 ;
      LAYER via ;
        RECT 424.680 1588.860 424.940 1589.120 ;
        RECT 493.220 1588.520 493.480 1588.780 ;
        RECT 413.180 20.440 413.440 20.700 ;
        RECT 424.220 20.440 424.480 20.700 ;
      LAYER met2 ;
        RECT 493.080 1600.380 493.360 1604.000 ;
        RECT 493.080 1600.000 493.420 1600.380 ;
        RECT 424.680 1589.060 424.940 1589.150 ;
        RECT 424.280 1588.920 424.940 1589.060 ;
        RECT 424.280 20.730 424.420 1588.920 ;
        RECT 424.680 1588.830 424.940 1588.920 ;
        RECT 493.280 1588.810 493.420 1600.000 ;
        RECT 493.220 1588.490 493.480 1588.810 ;
        RECT 413.180 20.410 413.440 20.730 ;
        RECT 424.220 20.410 424.480 20.730 ;
        RECT 413.240 2.400 413.380 20.410 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 375.320 1600.380 375.600 1604.000 ;
        RECT 375.320 1600.000 375.660 1600.380 ;
        RECT 375.520 1591.045 375.660 1600.000 ;
        RECT 75.530 1590.675 75.810 1591.045 ;
        RECT 375.450 1590.675 375.730 1591.045 ;
        RECT 75.600 17.410 75.740 1590.675 ;
        RECT 74.220 17.270 75.740 17.410 ;
        RECT 74.220 2.400 74.360 17.270 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 75.530 1590.720 75.810 1591.000 ;
        RECT 375.450 1590.720 375.730 1591.000 ;
      LAYER met3 ;
        RECT 75.505 1591.010 75.835 1591.025 ;
        RECT 375.425 1591.010 375.755 1591.025 ;
        RECT 75.505 1590.710 375.755 1591.010 ;
        RECT 75.505 1590.695 75.835 1590.710 ;
        RECT 375.425 1590.695 375.755 1590.710 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.350 1591.440 445.670 1591.500 ;
        RECT 499.170 1591.440 499.490 1591.500 ;
        RECT 445.350 1591.300 499.490 1591.440 ;
        RECT 445.350 1591.240 445.670 1591.300 ;
        RECT 499.170 1591.240 499.490 1591.300 ;
        RECT 430.630 20.300 430.950 20.360 ;
        RECT 445.350 20.300 445.670 20.360 ;
        RECT 430.630 20.160 445.670 20.300 ;
        RECT 430.630 20.100 430.950 20.160 ;
        RECT 445.350 20.100 445.670 20.160 ;
      LAYER via ;
        RECT 445.380 1591.240 445.640 1591.500 ;
        RECT 499.200 1591.240 499.460 1591.500 ;
        RECT 430.660 20.100 430.920 20.360 ;
        RECT 445.380 20.100 445.640 20.360 ;
      LAYER met2 ;
        RECT 499.060 1600.380 499.340 1604.000 ;
        RECT 499.060 1600.000 499.400 1600.380 ;
        RECT 499.260 1591.530 499.400 1600.000 ;
        RECT 445.380 1591.210 445.640 1591.530 ;
        RECT 499.200 1591.210 499.460 1591.530 ;
        RECT 445.440 20.390 445.580 1591.210 ;
        RECT 430.660 20.070 430.920 20.390 ;
        RECT 445.380 20.070 445.640 20.390 ;
        RECT 430.720 2.400 430.860 20.070 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 458.690 1591.780 459.010 1591.840 ;
        RECT 505.610 1591.780 505.930 1591.840 ;
        RECT 458.690 1591.640 505.930 1591.780 ;
        RECT 458.690 1591.580 459.010 1591.640 ;
        RECT 505.610 1591.580 505.930 1591.640 ;
        RECT 448.570 20.640 448.890 20.700 ;
        RECT 458.690 20.640 459.010 20.700 ;
        RECT 448.570 20.500 459.010 20.640 ;
        RECT 448.570 20.440 448.890 20.500 ;
        RECT 458.690 20.440 459.010 20.500 ;
      LAYER via ;
        RECT 458.720 1591.580 458.980 1591.840 ;
        RECT 505.640 1591.580 505.900 1591.840 ;
        RECT 448.600 20.440 448.860 20.700 ;
        RECT 458.720 20.440 458.980 20.700 ;
      LAYER met2 ;
        RECT 505.500 1600.380 505.780 1604.000 ;
        RECT 505.500 1600.000 505.840 1600.380 ;
        RECT 505.700 1591.870 505.840 1600.000 ;
        RECT 458.720 1591.550 458.980 1591.870 ;
        RECT 505.640 1591.550 505.900 1591.870 ;
        RECT 458.780 20.730 458.920 1591.550 ;
        RECT 448.600 20.410 448.860 20.730 ;
        RECT 458.720 20.410 458.980 20.730 ;
        RECT 448.660 2.400 448.800 20.410 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.810 1592.460 469.130 1592.520 ;
        RECT 511.590 1592.460 511.910 1592.520 ;
        RECT 468.810 1592.320 511.910 1592.460 ;
        RECT 468.810 1592.260 469.130 1592.320 ;
        RECT 511.590 1592.260 511.910 1592.320 ;
        RECT 466.510 20.640 466.830 20.700 ;
        RECT 468.810 20.640 469.130 20.700 ;
        RECT 466.510 20.500 469.130 20.640 ;
        RECT 466.510 20.440 466.830 20.500 ;
        RECT 468.810 20.440 469.130 20.500 ;
      LAYER via ;
        RECT 468.840 1592.260 469.100 1592.520 ;
        RECT 511.620 1592.260 511.880 1592.520 ;
        RECT 466.540 20.440 466.800 20.700 ;
        RECT 468.840 20.440 469.100 20.700 ;
      LAYER met2 ;
        RECT 511.480 1600.380 511.760 1604.000 ;
        RECT 511.480 1600.000 511.820 1600.380 ;
        RECT 511.680 1592.550 511.820 1600.000 ;
        RECT 468.840 1592.230 469.100 1592.550 ;
        RECT 511.620 1592.230 511.880 1592.550 ;
        RECT 468.900 20.730 469.040 1592.230 ;
        RECT 466.540 20.410 466.800 20.730 ;
        RECT 468.840 20.410 469.100 20.730 ;
        RECT 466.600 2.400 466.740 20.410 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 489.510 1588.380 489.830 1588.440 ;
        RECT 518.030 1588.380 518.350 1588.440 ;
        RECT 489.510 1588.240 518.350 1588.380 ;
        RECT 489.510 1588.180 489.830 1588.240 ;
        RECT 518.030 1588.180 518.350 1588.240 ;
        RECT 484.450 20.640 484.770 20.700 ;
        RECT 489.510 20.640 489.830 20.700 ;
        RECT 484.450 20.500 489.830 20.640 ;
        RECT 484.450 20.440 484.770 20.500 ;
        RECT 489.510 20.440 489.830 20.500 ;
      LAYER via ;
        RECT 489.540 1588.180 489.800 1588.440 ;
        RECT 518.060 1588.180 518.320 1588.440 ;
        RECT 484.480 20.440 484.740 20.700 ;
        RECT 489.540 20.440 489.800 20.700 ;
      LAYER met2 ;
        RECT 517.920 1600.380 518.200 1604.000 ;
        RECT 517.920 1600.000 518.260 1600.380 ;
        RECT 518.120 1588.470 518.260 1600.000 ;
        RECT 489.540 1588.150 489.800 1588.470 ;
        RECT 518.060 1588.150 518.320 1588.470 ;
        RECT 489.600 20.730 489.740 1588.150 ;
        RECT 484.480 20.410 484.740 20.730 ;
        RECT 489.540 20.410 489.800 20.730 ;
        RECT 484.540 2.400 484.680 20.410 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 502.390 19.620 502.710 19.680 ;
        RECT 518.490 19.620 518.810 19.680 ;
        RECT 502.390 19.480 518.810 19.620 ;
        RECT 502.390 19.420 502.710 19.480 ;
        RECT 518.490 19.420 518.810 19.480 ;
      LAYER via ;
        RECT 502.420 19.420 502.680 19.680 ;
        RECT 518.520 19.420 518.780 19.680 ;
      LAYER met2 ;
        RECT 523.900 1601.130 524.180 1604.000 ;
        RECT 522.260 1600.990 524.180 1601.130 ;
        RECT 522.260 1580.050 522.400 1600.990 ;
        RECT 523.900 1600.000 524.180 1600.990 ;
        RECT 518.580 1579.910 522.400 1580.050 ;
        RECT 518.580 19.710 518.720 1579.910 ;
        RECT 502.420 19.390 502.680 19.710 ;
        RECT 518.520 19.390 518.780 19.710 ;
        RECT 502.480 2.400 502.620 19.390 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 524.010 1587.360 524.330 1587.420 ;
        RECT 529.990 1587.360 530.310 1587.420 ;
        RECT 524.010 1587.220 530.310 1587.360 ;
        RECT 524.010 1587.160 524.330 1587.220 ;
        RECT 529.990 1587.160 530.310 1587.220 ;
        RECT 519.870 17.580 520.190 17.640 ;
        RECT 524.010 17.580 524.330 17.640 ;
        RECT 519.870 17.440 524.330 17.580 ;
        RECT 519.870 17.380 520.190 17.440 ;
        RECT 524.010 17.380 524.330 17.440 ;
      LAYER via ;
        RECT 524.040 1587.160 524.300 1587.420 ;
        RECT 530.020 1587.160 530.280 1587.420 ;
        RECT 519.900 17.380 520.160 17.640 ;
        RECT 524.040 17.380 524.300 17.640 ;
      LAYER met2 ;
        RECT 529.880 1600.380 530.160 1604.000 ;
        RECT 529.880 1600.000 530.220 1600.380 ;
        RECT 530.080 1587.450 530.220 1600.000 ;
        RECT 524.040 1587.130 524.300 1587.450 ;
        RECT 530.020 1587.130 530.280 1587.450 ;
        RECT 524.100 17.670 524.240 1587.130 ;
        RECT 519.900 17.350 520.160 17.670 ;
        RECT 524.040 17.350 524.300 17.670 ;
        RECT 519.960 2.400 520.100 17.350 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 533.285 1366.205 533.455 1400.715 ;
        RECT 534.205 1304.325 534.375 1352.435 ;
        RECT 532.365 1104.405 532.535 1152.175 ;
        RECT 533.285 786.505 533.455 821.015 ;
        RECT 533.285 689.605 533.455 724.455 ;
        RECT 532.365 572.985 532.535 620.415 ;
        RECT 533.285 469.285 533.455 517.395 ;
        RECT 533.285 427.805 533.455 449.055 ;
        RECT 532.365 331.585 532.535 379.355 ;
        RECT 534.205 157.845 534.375 193.035 ;
      LAYER mcon ;
        RECT 533.285 1400.545 533.455 1400.715 ;
        RECT 534.205 1352.265 534.375 1352.435 ;
        RECT 532.365 1152.005 532.535 1152.175 ;
        RECT 533.285 820.845 533.455 821.015 ;
        RECT 533.285 724.285 533.455 724.455 ;
        RECT 532.365 620.245 532.535 620.415 ;
        RECT 533.285 517.225 533.455 517.395 ;
        RECT 533.285 448.885 533.455 449.055 ;
        RECT 532.365 379.185 532.535 379.355 ;
        RECT 534.205 192.865 534.375 193.035 ;
      LAYER met1 ;
        RECT 532.750 1511.200 533.070 1511.260 ;
        RECT 533.670 1511.200 533.990 1511.260 ;
        RECT 532.750 1511.060 533.990 1511.200 ;
        RECT 532.750 1511.000 533.070 1511.060 ;
        RECT 533.670 1511.000 533.990 1511.060 ;
        RECT 532.750 1414.640 533.070 1414.700 ;
        RECT 533.670 1414.640 533.990 1414.700 ;
        RECT 532.750 1414.500 533.990 1414.640 ;
        RECT 532.750 1414.440 533.070 1414.500 ;
        RECT 533.670 1414.440 533.990 1414.500 ;
        RECT 533.210 1400.700 533.530 1400.760 ;
        RECT 533.015 1400.560 533.530 1400.700 ;
        RECT 533.210 1400.500 533.530 1400.560 ;
        RECT 533.225 1366.360 533.515 1366.405 ;
        RECT 534.130 1366.360 534.450 1366.420 ;
        RECT 533.225 1366.220 534.450 1366.360 ;
        RECT 533.225 1366.175 533.515 1366.220 ;
        RECT 534.130 1366.160 534.450 1366.220 ;
        RECT 534.130 1352.420 534.450 1352.480 ;
        RECT 533.935 1352.280 534.450 1352.420 ;
        RECT 534.130 1352.220 534.450 1352.280 ;
        RECT 534.145 1304.480 534.435 1304.525 ;
        RECT 534.590 1304.480 534.910 1304.540 ;
        RECT 534.145 1304.340 534.910 1304.480 ;
        RECT 534.145 1304.295 534.435 1304.340 ;
        RECT 534.590 1304.280 534.910 1304.340 ;
        RECT 534.590 1270.140 534.910 1270.200 ;
        RECT 534.220 1270.000 534.910 1270.140 ;
        RECT 534.220 1269.520 534.360 1270.000 ;
        RECT 534.590 1269.940 534.910 1270.000 ;
        RECT 534.130 1269.260 534.450 1269.520 ;
        RECT 532.305 1152.160 532.595 1152.205 ;
        RECT 532.750 1152.160 533.070 1152.220 ;
        RECT 532.305 1152.020 533.070 1152.160 ;
        RECT 532.305 1151.975 532.595 1152.020 ;
        RECT 532.750 1151.960 533.070 1152.020 ;
        RECT 532.290 1104.560 532.610 1104.620 ;
        RECT 532.095 1104.420 532.610 1104.560 ;
        RECT 532.290 1104.360 532.610 1104.420 ;
        RECT 532.290 1103.880 532.610 1103.940 ;
        RECT 533.210 1103.880 533.530 1103.940 ;
        RECT 532.290 1103.740 533.530 1103.880 ;
        RECT 532.290 1103.680 532.610 1103.740 ;
        RECT 533.210 1103.680 533.530 1103.740 ;
        RECT 532.750 1014.460 533.070 1014.520 ;
        RECT 533.670 1014.460 533.990 1014.520 ;
        RECT 532.750 1014.320 533.990 1014.460 ;
        RECT 532.750 1014.260 533.070 1014.320 ;
        RECT 533.670 1014.260 533.990 1014.320 ;
        RECT 533.670 979.920 533.990 980.180 ;
        RECT 533.760 979.780 533.900 979.920 ;
        RECT 534.130 979.780 534.450 979.840 ;
        RECT 533.760 979.640 534.450 979.780 ;
        RECT 534.130 979.580 534.450 979.640 ;
        RECT 533.210 917.900 533.530 917.960 ;
        RECT 534.590 917.900 534.910 917.960 ;
        RECT 533.210 917.760 534.910 917.900 ;
        RECT 533.210 917.700 533.530 917.760 ;
        RECT 534.590 917.700 534.910 917.760 ;
        RECT 533.670 869.620 533.990 869.680 ;
        RECT 534.590 869.620 534.910 869.680 ;
        RECT 533.670 869.480 534.910 869.620 ;
        RECT 533.670 869.420 533.990 869.480 ;
        RECT 534.590 869.420 534.910 869.480 ;
        RECT 533.210 821.000 533.530 821.060 ;
        RECT 533.015 820.860 533.530 821.000 ;
        RECT 533.210 820.800 533.530 820.860 ;
        RECT 533.210 786.660 533.530 786.720 ;
        RECT 533.015 786.520 533.530 786.660 ;
        RECT 533.210 786.460 533.530 786.520 ;
        RECT 532.750 738.380 533.070 738.440 ;
        RECT 533.670 738.380 533.990 738.440 ;
        RECT 532.750 738.240 533.990 738.380 ;
        RECT 532.750 738.180 533.070 738.240 ;
        RECT 533.670 738.180 533.990 738.240 ;
        RECT 533.210 724.440 533.530 724.500 ;
        RECT 533.015 724.300 533.530 724.440 ;
        RECT 533.210 724.240 533.530 724.300 ;
        RECT 533.210 689.760 533.530 689.820 ;
        RECT 533.015 689.620 533.530 689.760 ;
        RECT 533.210 689.560 533.530 689.620 ;
        RECT 532.290 621.080 532.610 621.140 ;
        RECT 533.670 621.080 533.990 621.140 ;
        RECT 532.290 620.940 533.990 621.080 ;
        RECT 532.290 620.880 532.610 620.940 ;
        RECT 533.670 620.880 533.990 620.940 ;
        RECT 532.290 620.400 532.610 620.460 ;
        RECT 532.095 620.260 532.610 620.400 ;
        RECT 532.290 620.200 532.610 620.260 ;
        RECT 532.305 573.140 532.595 573.185 ;
        RECT 532.750 573.140 533.070 573.200 ;
        RECT 532.305 573.000 533.070 573.140 ;
        RECT 532.305 572.955 532.595 573.000 ;
        RECT 532.750 572.940 533.070 573.000 ;
        RECT 532.750 545.400 533.070 545.660 ;
        RECT 532.840 544.980 532.980 545.400 ;
        RECT 532.750 544.720 533.070 544.980 ;
        RECT 533.210 517.380 533.530 517.440 ;
        RECT 533.210 517.240 533.725 517.380 ;
        RECT 533.210 517.180 533.530 517.240 ;
        RECT 532.750 469.440 533.070 469.500 ;
        RECT 533.225 469.440 533.515 469.485 ;
        RECT 532.750 469.300 533.515 469.440 ;
        RECT 532.750 469.240 533.070 469.300 ;
        RECT 533.225 469.255 533.515 469.300 ;
        RECT 532.750 449.040 533.070 449.100 ;
        RECT 533.225 449.040 533.515 449.085 ;
        RECT 532.750 448.900 533.515 449.040 ;
        RECT 532.750 448.840 533.070 448.900 ;
        RECT 533.225 448.855 533.515 448.900 ;
        RECT 533.210 427.960 533.530 428.020 ;
        RECT 533.015 427.820 533.530 427.960 ;
        RECT 533.210 427.760 533.530 427.820 ;
        RECT 532.305 379.340 532.595 379.385 ;
        RECT 532.750 379.340 533.070 379.400 ;
        RECT 532.305 379.200 533.070 379.340 ;
        RECT 532.305 379.155 532.595 379.200 ;
        RECT 532.750 379.140 533.070 379.200 ;
        RECT 532.290 331.740 532.610 331.800 ;
        RECT 532.095 331.600 532.610 331.740 ;
        RECT 532.290 331.540 532.610 331.600 ;
        RECT 532.290 331.060 532.610 331.120 ;
        RECT 532.750 331.060 533.070 331.120 ;
        RECT 532.290 330.920 533.070 331.060 ;
        RECT 532.290 330.860 532.610 330.920 ;
        RECT 532.750 330.860 533.070 330.920 ;
        RECT 532.750 255.240 533.070 255.300 ;
        RECT 533.670 255.240 533.990 255.300 ;
        RECT 532.750 255.100 533.990 255.240 ;
        RECT 532.750 255.040 533.070 255.100 ;
        RECT 533.670 255.040 533.990 255.100 ;
        RECT 534.130 193.020 534.450 193.080 ;
        RECT 533.935 192.880 534.450 193.020 ;
        RECT 534.130 192.820 534.450 192.880 ;
        RECT 534.130 158.000 534.450 158.060 ;
        RECT 533.935 157.860 534.450 158.000 ;
        RECT 534.130 157.800 534.450 157.860 ;
        RECT 534.130 20.640 534.450 20.700 ;
        RECT 537.810 20.640 538.130 20.700 ;
        RECT 534.130 20.500 538.130 20.640 ;
        RECT 534.130 20.440 534.450 20.500 ;
        RECT 537.810 20.440 538.130 20.500 ;
      LAYER via ;
        RECT 532.780 1511.000 533.040 1511.260 ;
        RECT 533.700 1511.000 533.960 1511.260 ;
        RECT 532.780 1414.440 533.040 1414.700 ;
        RECT 533.700 1414.440 533.960 1414.700 ;
        RECT 533.240 1400.500 533.500 1400.760 ;
        RECT 534.160 1366.160 534.420 1366.420 ;
        RECT 534.160 1352.220 534.420 1352.480 ;
        RECT 534.620 1304.280 534.880 1304.540 ;
        RECT 534.620 1269.940 534.880 1270.200 ;
        RECT 534.160 1269.260 534.420 1269.520 ;
        RECT 532.780 1151.960 533.040 1152.220 ;
        RECT 532.320 1104.360 532.580 1104.620 ;
        RECT 532.320 1103.680 532.580 1103.940 ;
        RECT 533.240 1103.680 533.500 1103.940 ;
        RECT 532.780 1014.260 533.040 1014.520 ;
        RECT 533.700 1014.260 533.960 1014.520 ;
        RECT 533.700 979.920 533.960 980.180 ;
        RECT 534.160 979.580 534.420 979.840 ;
        RECT 533.240 917.700 533.500 917.960 ;
        RECT 534.620 917.700 534.880 917.960 ;
        RECT 533.700 869.420 533.960 869.680 ;
        RECT 534.620 869.420 534.880 869.680 ;
        RECT 533.240 820.800 533.500 821.060 ;
        RECT 533.240 786.460 533.500 786.720 ;
        RECT 532.780 738.180 533.040 738.440 ;
        RECT 533.700 738.180 533.960 738.440 ;
        RECT 533.240 724.240 533.500 724.500 ;
        RECT 533.240 689.560 533.500 689.820 ;
        RECT 532.320 620.880 532.580 621.140 ;
        RECT 533.700 620.880 533.960 621.140 ;
        RECT 532.320 620.200 532.580 620.460 ;
        RECT 532.780 572.940 533.040 573.200 ;
        RECT 532.780 545.400 533.040 545.660 ;
        RECT 532.780 544.720 533.040 544.980 ;
        RECT 533.240 517.180 533.500 517.440 ;
        RECT 532.780 469.240 533.040 469.500 ;
        RECT 532.780 448.840 533.040 449.100 ;
        RECT 533.240 427.760 533.500 428.020 ;
        RECT 532.780 379.140 533.040 379.400 ;
        RECT 532.320 331.540 532.580 331.800 ;
        RECT 532.320 330.860 532.580 331.120 ;
        RECT 532.780 330.860 533.040 331.120 ;
        RECT 532.780 255.040 533.040 255.300 ;
        RECT 533.700 255.040 533.960 255.300 ;
        RECT 534.160 192.820 534.420 193.080 ;
        RECT 534.160 157.800 534.420 158.060 ;
        RECT 534.160 20.440 534.420 20.700 ;
        RECT 537.840 20.440 538.100 20.700 ;
      LAYER met2 ;
        RECT 536.320 1600.450 536.600 1604.000 ;
        RECT 535.140 1600.310 536.600 1600.450 ;
        RECT 535.140 1580.050 535.280 1600.310 ;
        RECT 536.320 1600.000 536.600 1600.310 ;
        RECT 533.760 1579.910 535.280 1580.050 ;
        RECT 533.760 1511.290 533.900 1579.910 ;
        RECT 532.780 1510.970 533.040 1511.290 ;
        RECT 533.700 1510.970 533.960 1511.290 ;
        RECT 532.840 1510.690 532.980 1510.970 ;
        RECT 532.840 1510.550 533.440 1510.690 ;
        RECT 533.300 1463.090 533.440 1510.550 ;
        RECT 533.300 1462.950 533.900 1463.090 ;
        RECT 533.760 1414.730 533.900 1462.950 ;
        RECT 532.780 1414.410 533.040 1414.730 ;
        RECT 533.700 1414.410 533.960 1414.730 ;
        RECT 532.840 1414.130 532.980 1414.410 ;
        RECT 532.840 1413.990 533.440 1414.130 ;
        RECT 533.300 1400.790 533.440 1413.990 ;
        RECT 533.240 1400.470 533.500 1400.790 ;
        RECT 534.160 1366.130 534.420 1366.450 ;
        RECT 534.220 1352.510 534.360 1366.130 ;
        RECT 534.160 1352.190 534.420 1352.510 ;
        RECT 534.620 1304.250 534.880 1304.570 ;
        RECT 534.680 1270.230 534.820 1304.250 ;
        RECT 534.620 1269.910 534.880 1270.230 ;
        RECT 534.160 1269.230 534.420 1269.550 ;
        RECT 534.220 1221.010 534.360 1269.230 ;
        RECT 533.300 1220.870 534.360 1221.010 ;
        RECT 533.300 1207.525 533.440 1220.870 ;
        RECT 533.230 1207.155 533.510 1207.525 ;
        RECT 532.770 1176.555 533.050 1176.925 ;
        RECT 532.840 1152.250 532.980 1176.555 ;
        RECT 532.780 1151.930 533.040 1152.250 ;
        RECT 532.320 1104.330 532.580 1104.650 ;
        RECT 532.380 1103.970 532.520 1104.330 ;
        RECT 532.320 1103.650 532.580 1103.970 ;
        RECT 533.240 1103.650 533.500 1103.970 ;
        RECT 533.300 1076.170 533.440 1103.650 ;
        RECT 532.840 1076.030 533.440 1076.170 ;
        RECT 532.840 1014.550 532.980 1076.030 ;
        RECT 532.780 1014.230 533.040 1014.550 ;
        RECT 533.700 1014.230 533.960 1014.550 ;
        RECT 533.760 980.210 533.900 1014.230 ;
        RECT 533.700 979.890 533.960 980.210 ;
        RECT 534.160 979.550 534.420 979.870 ;
        RECT 534.220 966.125 534.360 979.550 ;
        RECT 533.230 965.755 533.510 966.125 ;
        RECT 534.150 965.755 534.430 966.125 ;
        RECT 533.300 917.990 533.440 965.755 ;
        RECT 533.240 917.670 533.500 917.990 ;
        RECT 534.620 917.670 534.880 917.990 ;
        RECT 534.680 869.710 534.820 917.670 ;
        RECT 533.700 869.565 533.960 869.710 ;
        RECT 532.310 869.195 532.590 869.565 ;
        RECT 533.690 869.195 533.970 869.565 ;
        RECT 534.620 869.390 534.880 869.710 ;
        RECT 532.380 821.285 532.520 869.195 ;
        RECT 532.310 820.915 532.590 821.285 ;
        RECT 533.230 820.915 533.510 821.285 ;
        RECT 533.240 820.770 533.500 820.915 ;
        RECT 533.240 786.430 533.500 786.750 ;
        RECT 533.300 772.890 533.440 786.430 ;
        RECT 533.300 772.750 533.900 772.890 ;
        RECT 533.760 738.470 533.900 772.750 ;
        RECT 532.780 738.210 533.040 738.470 ;
        RECT 532.780 738.150 533.440 738.210 ;
        RECT 533.700 738.150 533.960 738.470 ;
        RECT 532.840 738.070 533.440 738.150 ;
        RECT 533.300 724.530 533.440 738.070 ;
        RECT 533.240 724.210 533.500 724.530 ;
        RECT 533.240 689.530 533.500 689.850 ;
        RECT 533.300 676.330 533.440 689.530 ;
        RECT 533.300 676.190 533.900 676.330 ;
        RECT 533.760 621.170 533.900 676.190 ;
        RECT 532.320 620.850 532.580 621.170 ;
        RECT 533.700 620.850 533.960 621.170 ;
        RECT 532.380 620.490 532.520 620.850 ;
        RECT 532.320 620.170 532.580 620.490 ;
        RECT 532.780 572.910 533.040 573.230 ;
        RECT 532.840 545.690 532.980 572.910 ;
        RECT 532.780 545.370 533.040 545.690 ;
        RECT 532.780 544.690 533.040 545.010 ;
        RECT 532.840 524.690 532.980 544.690 ;
        RECT 532.840 524.550 533.440 524.690 ;
        RECT 533.300 517.470 533.440 524.550 ;
        RECT 533.240 517.150 533.500 517.470 ;
        RECT 532.780 469.210 533.040 469.530 ;
        RECT 532.840 449.130 532.980 469.210 ;
        RECT 532.780 448.810 533.040 449.130 ;
        RECT 533.240 427.730 533.500 428.050 ;
        RECT 533.300 379.850 533.440 427.730 ;
        RECT 532.840 379.710 533.440 379.850 ;
        RECT 532.840 379.430 532.980 379.710 ;
        RECT 532.780 379.110 533.040 379.430 ;
        RECT 532.320 331.510 532.580 331.830 ;
        RECT 532.380 331.150 532.520 331.510 ;
        RECT 532.320 330.830 532.580 331.150 ;
        RECT 532.780 330.830 533.040 331.150 ;
        RECT 532.840 255.330 532.980 330.830 ;
        RECT 532.780 255.010 533.040 255.330 ;
        RECT 533.700 255.010 533.960 255.330 ;
        RECT 533.760 217.330 533.900 255.010 ;
        RECT 533.760 217.190 534.360 217.330 ;
        RECT 534.220 193.110 534.360 217.190 ;
        RECT 534.160 192.790 534.420 193.110 ;
        RECT 534.160 157.770 534.420 158.090 ;
        RECT 534.220 20.730 534.360 157.770 ;
        RECT 534.160 20.410 534.420 20.730 ;
        RECT 537.840 20.410 538.100 20.730 ;
        RECT 537.900 2.400 538.040 20.410 ;
        RECT 537.690 -4.800 538.250 2.400 ;
      LAYER via2 ;
        RECT 533.230 1207.200 533.510 1207.480 ;
        RECT 532.770 1176.600 533.050 1176.880 ;
        RECT 533.230 965.800 533.510 966.080 ;
        RECT 534.150 965.800 534.430 966.080 ;
        RECT 532.310 869.240 532.590 869.520 ;
        RECT 533.690 869.240 533.970 869.520 ;
        RECT 532.310 820.960 532.590 821.240 ;
        RECT 533.230 820.960 533.510 821.240 ;
      LAYER met3 ;
        RECT 533.205 1207.500 533.535 1207.505 ;
        RECT 532.950 1207.490 533.535 1207.500 ;
        RECT 532.750 1207.190 533.535 1207.490 ;
        RECT 532.950 1207.180 533.535 1207.190 ;
        RECT 533.205 1207.175 533.535 1207.180 ;
        RECT 532.745 1176.900 533.075 1176.905 ;
        RECT 532.745 1176.890 533.330 1176.900 ;
        RECT 532.520 1176.590 533.330 1176.890 ;
        RECT 532.745 1176.580 533.330 1176.590 ;
        RECT 532.745 1176.575 533.075 1176.580 ;
        RECT 533.205 966.090 533.535 966.105 ;
        RECT 534.125 966.090 534.455 966.105 ;
        RECT 533.205 965.790 534.455 966.090 ;
        RECT 533.205 965.775 533.535 965.790 ;
        RECT 534.125 965.775 534.455 965.790 ;
        RECT 532.285 869.530 532.615 869.545 ;
        RECT 533.665 869.530 533.995 869.545 ;
        RECT 532.285 869.230 533.995 869.530 ;
        RECT 532.285 869.215 532.615 869.230 ;
        RECT 533.665 869.215 533.995 869.230 ;
        RECT 532.285 821.250 532.615 821.265 ;
        RECT 533.205 821.250 533.535 821.265 ;
        RECT 532.285 820.950 533.535 821.250 ;
        RECT 532.285 820.935 532.615 820.950 ;
        RECT 533.205 820.935 533.535 820.950 ;
      LAYER via3 ;
        RECT 532.980 1207.180 533.300 1207.500 ;
        RECT 532.980 1176.580 533.300 1176.900 ;
      LAYER met4 ;
        RECT 532.975 1207.175 533.305 1207.505 ;
        RECT 532.990 1176.905 533.290 1207.175 ;
        RECT 532.975 1176.575 533.305 1176.905 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 544.710 16.900 545.030 16.960 ;
        RECT 555.750 16.900 556.070 16.960 ;
        RECT 544.710 16.760 556.070 16.900 ;
        RECT 544.710 16.700 545.030 16.760 ;
        RECT 555.750 16.700 556.070 16.760 ;
      LAYER via ;
        RECT 544.740 16.700 545.000 16.960 ;
        RECT 555.780 16.700 556.040 16.960 ;
      LAYER met2 ;
        RECT 542.300 1600.450 542.580 1604.000 ;
        RECT 542.300 1600.310 544.020 1600.450 ;
        RECT 542.300 1600.000 542.580 1600.310 ;
        RECT 543.880 1588.210 544.020 1600.310 ;
        RECT 543.880 1588.070 544.940 1588.210 ;
        RECT 544.800 16.990 544.940 1588.070 ;
        RECT 544.740 16.670 545.000 16.990 ;
        RECT 555.780 16.670 556.040 16.990 ;
        RECT 555.840 2.400 555.980 16.670 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 551.610 19.960 551.930 20.020 ;
        RECT 573.690 19.960 574.010 20.020 ;
        RECT 551.610 19.820 574.010 19.960 ;
        RECT 551.610 19.760 551.930 19.820 ;
        RECT 573.690 19.760 574.010 19.820 ;
      LAYER via ;
        RECT 551.640 19.760 551.900 20.020 ;
        RECT 573.720 19.760 573.980 20.020 ;
      LAYER met2 ;
        RECT 548.740 1600.450 549.020 1604.000 ;
        RECT 548.740 1600.310 550.000 1600.450 ;
        RECT 548.740 1600.000 549.020 1600.310 ;
        RECT 549.860 1590.250 550.000 1600.310 ;
        RECT 549.860 1590.110 551.840 1590.250 ;
        RECT 551.700 20.050 551.840 1590.110 ;
        RECT 551.640 19.730 551.900 20.050 ;
        RECT 573.720 19.730 573.980 20.050 ;
        RECT 573.780 2.400 573.920 19.730 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 554.830 1590.080 555.150 1590.140 ;
        RECT 558.510 1590.080 558.830 1590.140 ;
        RECT 554.830 1589.940 558.830 1590.080 ;
        RECT 554.830 1589.880 555.150 1589.940 ;
        RECT 558.510 1589.880 558.830 1589.940 ;
        RECT 558.510 17.240 558.830 17.300 ;
        RECT 591.170 17.240 591.490 17.300 ;
        RECT 558.510 17.100 591.490 17.240 ;
        RECT 558.510 17.040 558.830 17.100 ;
        RECT 591.170 17.040 591.490 17.100 ;
      LAYER via ;
        RECT 554.860 1589.880 555.120 1590.140 ;
        RECT 558.540 1589.880 558.800 1590.140 ;
        RECT 558.540 17.040 558.800 17.300 ;
        RECT 591.200 17.040 591.460 17.300 ;
      LAYER met2 ;
        RECT 554.720 1600.380 555.000 1604.000 ;
        RECT 554.720 1600.000 555.060 1600.380 ;
        RECT 554.920 1590.170 555.060 1600.000 ;
        RECT 554.860 1589.850 555.120 1590.170 ;
        RECT 558.540 1589.850 558.800 1590.170 ;
        RECT 558.600 17.330 558.740 1589.850 ;
        RECT 558.540 17.010 558.800 17.330 ;
        RECT 591.200 17.010 591.460 17.330 ;
        RECT 591.260 2.400 591.400 17.010 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 379.570 1580.220 379.890 1580.280 ;
        RECT 382.330 1580.220 382.650 1580.280 ;
        RECT 379.570 1580.080 382.650 1580.220 ;
        RECT 379.570 1580.020 379.890 1580.080 ;
        RECT 382.330 1580.020 382.650 1580.080 ;
      LAYER via ;
        RECT 379.600 1580.020 379.860 1580.280 ;
        RECT 382.360 1580.020 382.620 1580.280 ;
      LAYER met2 ;
        RECT 383.600 1600.450 383.880 1604.000 ;
        RECT 382.420 1600.310 383.880 1600.450 ;
        RECT 382.420 1580.310 382.560 1600.310 ;
        RECT 383.600 1600.000 383.880 1600.310 ;
        RECT 379.600 1579.990 379.860 1580.310 ;
        RECT 382.360 1579.990 382.620 1580.310 ;
        RECT 379.660 18.885 379.800 1579.990 ;
        RECT 97.610 18.515 97.890 18.885 ;
        RECT 379.590 18.515 379.870 18.885 ;
        RECT 97.680 2.400 97.820 18.515 ;
        RECT 97.470 -4.800 98.030 2.400 ;
      LAYER via2 ;
        RECT 97.610 18.560 97.890 18.840 ;
        RECT 379.590 18.560 379.870 18.840 ;
      LAYER met3 ;
        RECT 97.585 18.850 97.915 18.865 ;
        RECT 379.565 18.850 379.895 18.865 ;
        RECT 97.585 18.550 379.895 18.850 ;
        RECT 97.585 18.535 97.915 18.550 ;
        RECT 379.565 18.535 379.895 18.550 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 561.270 1590.760 561.590 1590.820 ;
        RECT 582.890 1590.760 583.210 1590.820 ;
        RECT 561.270 1590.620 583.210 1590.760 ;
        RECT 561.270 1590.560 561.590 1590.620 ;
        RECT 582.890 1590.560 583.210 1590.620 ;
        RECT 582.890 16.560 583.210 16.620 ;
        RECT 609.110 16.560 609.430 16.620 ;
        RECT 582.890 16.420 609.430 16.560 ;
        RECT 582.890 16.360 583.210 16.420 ;
        RECT 609.110 16.360 609.430 16.420 ;
      LAYER via ;
        RECT 561.300 1590.560 561.560 1590.820 ;
        RECT 582.920 1590.560 583.180 1590.820 ;
        RECT 582.920 16.360 583.180 16.620 ;
        RECT 609.140 16.360 609.400 16.620 ;
      LAYER met2 ;
        RECT 561.160 1600.380 561.440 1604.000 ;
        RECT 561.160 1600.000 561.500 1600.380 ;
        RECT 561.360 1590.850 561.500 1600.000 ;
        RECT 561.300 1590.530 561.560 1590.850 ;
        RECT 582.920 1590.530 583.180 1590.850 ;
        RECT 582.980 16.650 583.120 1590.530 ;
        RECT 582.920 16.330 583.180 16.650 ;
        RECT 609.140 16.330 609.400 16.650 ;
        RECT 609.200 2.400 609.340 16.330 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 610.105 15.725 610.275 16.915 ;
      LAYER mcon ;
        RECT 610.105 16.745 610.275 16.915 ;
      LAYER met1 ;
        RECT 567.250 1590.080 567.570 1590.140 ;
        RECT 572.310 1590.080 572.630 1590.140 ;
        RECT 567.250 1589.940 572.630 1590.080 ;
        RECT 567.250 1589.880 567.570 1589.940 ;
        RECT 572.310 1589.880 572.630 1589.940 ;
        RECT 610.045 16.900 610.335 16.945 ;
        RECT 627.050 16.900 627.370 16.960 ;
        RECT 610.045 16.760 627.370 16.900 ;
        RECT 610.045 16.715 610.335 16.760 ;
        RECT 627.050 16.700 627.370 16.760 ;
        RECT 572.310 15.880 572.630 15.940 ;
        RECT 610.045 15.880 610.335 15.925 ;
        RECT 572.310 15.740 610.335 15.880 ;
        RECT 572.310 15.680 572.630 15.740 ;
        RECT 610.045 15.695 610.335 15.740 ;
      LAYER via ;
        RECT 567.280 1589.880 567.540 1590.140 ;
        RECT 572.340 1589.880 572.600 1590.140 ;
        RECT 627.080 16.700 627.340 16.960 ;
        RECT 572.340 15.680 572.600 15.940 ;
      LAYER met2 ;
        RECT 567.140 1600.380 567.420 1604.000 ;
        RECT 567.140 1600.000 567.480 1600.380 ;
        RECT 567.340 1590.170 567.480 1600.000 ;
        RECT 567.280 1589.850 567.540 1590.170 ;
        RECT 572.340 1589.850 572.600 1590.170 ;
        RECT 572.400 15.970 572.540 1589.850 ;
        RECT 627.080 16.670 627.340 16.990 ;
        RECT 572.340 15.650 572.600 15.970 ;
        RECT 627.140 2.400 627.280 16.670 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 371.825 1590.605 372.915 1590.775 ;
        RECT 371.825 1590.265 371.995 1590.605 ;
      LAYER mcon ;
        RECT 372.745 1590.605 372.915 1590.775 ;
      LAYER met1 ;
        RECT 372.685 1590.760 372.975 1590.805 ;
        RECT 391.990 1590.760 392.310 1590.820 ;
        RECT 372.685 1590.620 392.310 1590.760 ;
        RECT 372.685 1590.575 372.975 1590.620 ;
        RECT 391.990 1590.560 392.310 1590.620 ;
        RECT 123.810 1590.420 124.130 1590.480 ;
        RECT 371.765 1590.420 372.055 1590.465 ;
        RECT 123.810 1590.280 372.055 1590.420 ;
        RECT 123.810 1590.220 124.130 1590.280 ;
        RECT 371.765 1590.235 372.055 1590.280 ;
        RECT 121.510 16.900 121.830 16.960 ;
        RECT 123.810 16.900 124.130 16.960 ;
        RECT 121.510 16.760 124.130 16.900 ;
        RECT 121.510 16.700 121.830 16.760 ;
        RECT 123.810 16.700 124.130 16.760 ;
      LAYER via ;
        RECT 392.020 1590.560 392.280 1590.820 ;
        RECT 123.840 1590.220 124.100 1590.480 ;
        RECT 121.540 16.700 121.800 16.960 ;
        RECT 123.840 16.700 124.100 16.960 ;
      LAYER met2 ;
        RECT 391.880 1600.380 392.160 1604.000 ;
        RECT 391.880 1600.000 392.220 1600.380 ;
        RECT 392.080 1590.850 392.220 1600.000 ;
        RECT 392.020 1590.530 392.280 1590.850 ;
        RECT 123.840 1590.190 124.100 1590.510 ;
        RECT 123.900 16.990 124.040 1590.190 ;
        RECT 121.540 16.670 121.800 16.990 ;
        RECT 123.840 16.670 124.100 16.990 ;
        RECT 121.600 2.400 121.740 16.670 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 400.160 1600.450 400.440 1604.000 ;
        RECT 400.160 1600.310 400.960 1600.450 ;
        RECT 400.160 1600.000 400.440 1600.310 ;
        RECT 400.820 19.565 400.960 1600.310 ;
        RECT 145.450 19.195 145.730 19.565 ;
        RECT 400.750 19.195 401.030 19.565 ;
        RECT 145.520 2.400 145.660 19.195 ;
        RECT 145.310 -4.800 145.870 2.400 ;
      LAYER via2 ;
        RECT 145.450 19.240 145.730 19.520 ;
        RECT 400.750 19.240 401.030 19.520 ;
      LAYER met3 ;
        RECT 145.425 19.530 145.755 19.545 ;
        RECT 400.725 19.530 401.055 19.545 ;
        RECT 145.425 19.230 401.055 19.530 ;
        RECT 145.425 19.215 145.755 19.230 ;
        RECT 400.725 19.215 401.055 19.230 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 406.710 1592.120 407.030 1592.180 ;
        RECT 394.840 1591.980 407.030 1592.120 ;
        RECT 165.210 1591.780 165.530 1591.840 ;
        RECT 394.840 1591.780 394.980 1591.980 ;
        RECT 406.710 1591.920 407.030 1591.980 ;
        RECT 165.210 1591.640 394.980 1591.780 ;
        RECT 165.210 1591.580 165.530 1591.640 ;
      LAYER via ;
        RECT 165.240 1591.580 165.500 1591.840 ;
        RECT 406.740 1591.920 407.000 1592.180 ;
      LAYER met2 ;
        RECT 406.600 1600.380 406.880 1604.000 ;
        RECT 406.600 1600.000 406.940 1600.380 ;
        RECT 406.800 1592.210 406.940 1600.000 ;
        RECT 406.740 1591.890 407.000 1592.210 ;
        RECT 165.240 1591.550 165.500 1591.870 ;
        RECT 165.300 17.410 165.440 1591.550 ;
        RECT 163.460 17.270 165.440 17.410 ;
        RECT 163.460 2.400 163.600 17.270 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 407.630 1579.880 407.950 1579.940 ;
        RECT 411.310 1579.880 411.630 1579.940 ;
        RECT 407.630 1579.740 411.630 1579.880 ;
        RECT 407.630 1579.680 407.950 1579.740 ;
        RECT 411.310 1579.680 411.630 1579.740 ;
        RECT 180.850 20.640 181.170 20.700 ;
        RECT 407.630 20.640 407.950 20.700 ;
        RECT 180.850 20.500 407.950 20.640 ;
        RECT 180.850 20.440 181.170 20.500 ;
        RECT 407.630 20.440 407.950 20.500 ;
      LAYER via ;
        RECT 407.660 1579.680 407.920 1579.940 ;
        RECT 411.340 1579.680 411.600 1579.940 ;
        RECT 180.880 20.440 181.140 20.700 ;
        RECT 407.660 20.440 407.920 20.700 ;
      LAYER met2 ;
        RECT 412.580 1600.450 412.860 1604.000 ;
        RECT 411.400 1600.310 412.860 1600.450 ;
        RECT 411.400 1579.970 411.540 1600.310 ;
        RECT 412.580 1600.000 412.860 1600.310 ;
        RECT 407.660 1579.650 407.920 1579.970 ;
        RECT 411.340 1579.650 411.600 1579.970 ;
        RECT 407.720 20.730 407.860 1579.650 ;
        RECT 180.880 20.410 181.140 20.730 ;
        RECT 407.660 20.410 407.920 20.730 ;
        RECT 180.940 2.400 181.080 20.410 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 199.710 1593.140 200.030 1593.200 ;
        RECT 418.670 1593.140 418.990 1593.200 ;
        RECT 199.710 1593.000 418.990 1593.140 ;
        RECT 199.710 1592.940 200.030 1593.000 ;
        RECT 418.670 1592.940 418.990 1593.000 ;
      LAYER via ;
        RECT 199.740 1592.940 200.000 1593.200 ;
        RECT 418.700 1592.940 418.960 1593.200 ;
      LAYER met2 ;
        RECT 418.560 1600.380 418.840 1604.000 ;
        RECT 418.560 1600.000 418.900 1600.380 ;
        RECT 418.760 1593.230 418.900 1600.000 ;
        RECT 199.740 1592.910 200.000 1593.230 ;
        RECT 418.700 1592.910 418.960 1593.230 ;
        RECT 199.800 17.410 199.940 1592.910 ;
        RECT 198.880 17.270 199.940 17.410 ;
        RECT 198.880 2.400 199.020 17.270 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 408.165 19.465 408.335 20.655 ;
        RECT 227.385 15.385 227.555 16.575 ;
        RECT 276.605 15.045 276.775 16.575 ;
        RECT 305.585 13.345 305.755 15.215 ;
        RECT 323.065 13.345 323.235 16.575 ;
      LAYER mcon ;
        RECT 408.165 20.485 408.335 20.655 ;
        RECT 227.385 16.405 227.555 16.575 ;
        RECT 276.605 16.405 276.775 16.575 ;
        RECT 323.065 16.405 323.235 16.575 ;
        RECT 305.585 15.045 305.755 15.215 ;
      LAYER met1 ;
        RECT 408.105 20.640 408.395 20.685 ;
        RECT 408.105 20.500 409.700 20.640 ;
        RECT 408.105 20.455 408.395 20.500 ;
        RECT 409.560 20.300 409.700 20.500 ;
        RECT 421.890 20.300 422.210 20.360 ;
        RECT 409.560 20.160 422.210 20.300 ;
        RECT 421.890 20.100 422.210 20.160 ;
        RECT 400.270 19.620 400.590 19.680 ;
        RECT 408.105 19.620 408.395 19.665 ;
        RECT 400.270 19.480 408.395 19.620 ;
        RECT 400.270 19.420 400.590 19.480 ;
        RECT 408.105 19.435 408.395 19.480 ;
        RECT 398.890 16.900 399.210 16.960 ;
        RECT 358.500 16.760 399.210 16.900 ;
        RECT 227.325 16.560 227.615 16.605 ;
        RECT 276.545 16.560 276.835 16.605 ;
        RECT 227.325 16.420 276.835 16.560 ;
        RECT 227.325 16.375 227.615 16.420 ;
        RECT 276.545 16.375 276.835 16.420 ;
        RECT 323.005 16.560 323.295 16.605 ;
        RECT 358.500 16.560 358.640 16.760 ;
        RECT 398.890 16.700 399.210 16.760 ;
        RECT 323.005 16.420 358.640 16.560 ;
        RECT 323.005 16.375 323.295 16.420 ;
        RECT 216.730 15.540 217.050 15.600 ;
        RECT 227.325 15.540 227.615 15.585 ;
        RECT 216.730 15.400 227.615 15.540 ;
        RECT 216.730 15.340 217.050 15.400 ;
        RECT 227.325 15.355 227.615 15.400 ;
        RECT 276.545 15.200 276.835 15.245 ;
        RECT 305.525 15.200 305.815 15.245 ;
        RECT 276.545 15.060 305.815 15.200 ;
        RECT 276.545 15.015 276.835 15.060 ;
        RECT 305.525 15.015 305.815 15.060 ;
        RECT 305.525 13.500 305.815 13.545 ;
        RECT 323.005 13.500 323.295 13.545 ;
        RECT 305.525 13.360 323.295 13.500 ;
        RECT 305.525 13.315 305.815 13.360 ;
        RECT 323.005 13.315 323.295 13.360 ;
      LAYER via ;
        RECT 421.920 20.100 422.180 20.360 ;
        RECT 400.300 19.420 400.560 19.680 ;
        RECT 398.920 16.700 399.180 16.960 ;
        RECT 216.760 15.340 217.020 15.600 ;
      LAYER met2 ;
        RECT 425.000 1600.450 425.280 1604.000 ;
        RECT 423.360 1600.310 425.280 1600.450 ;
        RECT 423.360 1580.050 423.500 1600.310 ;
        RECT 425.000 1600.000 425.280 1600.310 ;
        RECT 421.980 1579.910 423.500 1580.050 ;
        RECT 421.980 20.390 422.120 1579.910 ;
        RECT 421.920 20.070 422.180 20.390 ;
        RECT 400.300 19.390 400.560 19.710 ;
        RECT 398.920 16.670 399.180 16.990 ;
        RECT 398.980 16.165 399.120 16.670 ;
        RECT 400.360 16.165 400.500 19.390 ;
        RECT 398.910 15.795 399.190 16.165 ;
        RECT 400.290 15.795 400.570 16.165 ;
        RECT 216.760 15.310 217.020 15.630 ;
        RECT 216.820 2.400 216.960 15.310 ;
        RECT 216.610 -4.800 217.170 2.400 ;
      LAYER via2 ;
        RECT 398.910 15.840 399.190 16.120 ;
        RECT 400.290 15.840 400.570 16.120 ;
      LAYER met3 ;
        RECT 398.885 16.130 399.215 16.145 ;
        RECT 400.265 16.130 400.595 16.145 ;
        RECT 398.885 15.830 400.595 16.130 ;
        RECT 398.885 15.815 399.215 15.830 ;
        RECT 400.265 15.815 400.595 15.830 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 431.090 1590.420 431.410 1590.480 ;
        RECT 417.380 1590.280 431.410 1590.420 ;
        RECT 240.650 1590.080 240.970 1590.140 ;
        RECT 417.380 1590.080 417.520 1590.280 ;
        RECT 431.090 1590.220 431.410 1590.280 ;
        RECT 240.650 1589.940 417.520 1590.080 ;
        RECT 240.650 1589.880 240.970 1589.940 ;
        RECT 234.670 16.220 234.990 16.280 ;
        RECT 240.650 16.220 240.970 16.280 ;
        RECT 234.670 16.080 240.970 16.220 ;
        RECT 234.670 16.020 234.990 16.080 ;
        RECT 240.650 16.020 240.970 16.080 ;
      LAYER via ;
        RECT 240.680 1589.880 240.940 1590.140 ;
        RECT 431.120 1590.220 431.380 1590.480 ;
        RECT 234.700 16.020 234.960 16.280 ;
        RECT 240.680 16.020 240.940 16.280 ;
      LAYER met2 ;
        RECT 430.980 1600.380 431.260 1604.000 ;
        RECT 430.980 1600.000 431.320 1600.380 ;
        RECT 431.180 1590.510 431.320 1600.000 ;
        RECT 431.120 1590.190 431.380 1590.510 ;
        RECT 240.680 1589.850 240.940 1590.170 ;
        RECT 240.740 16.310 240.880 1589.850 ;
        RECT 234.700 15.990 234.960 16.310 ;
        RECT 240.680 15.990 240.940 16.310 ;
        RECT 234.760 2.400 234.900 15.990 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 351.585 18.445 352.215 18.615 ;
        RECT 351.585 18.105 351.755 18.445 ;
        RECT 352.045 18.105 352.215 18.445 ;
      LAYER met1 ;
        RECT 366.230 1576.480 366.550 1576.540 ;
        RECT 368.070 1576.480 368.390 1576.540 ;
        RECT 366.230 1576.340 368.390 1576.480 ;
        RECT 366.230 1576.280 366.550 1576.340 ;
        RECT 368.070 1576.280 368.390 1576.340 ;
        RECT 56.190 18.260 56.510 18.320 ;
        RECT 351.525 18.260 351.815 18.305 ;
        RECT 56.190 18.120 351.815 18.260 ;
        RECT 56.190 18.060 56.510 18.120 ;
        RECT 351.525 18.075 351.815 18.120 ;
        RECT 351.985 18.260 352.275 18.305 ;
        RECT 366.230 18.260 366.550 18.320 ;
        RECT 351.985 18.120 366.550 18.260 ;
        RECT 351.985 18.075 352.275 18.120 ;
        RECT 366.230 18.060 366.550 18.120 ;
      LAYER via ;
        RECT 366.260 1576.280 366.520 1576.540 ;
        RECT 368.100 1576.280 368.360 1576.540 ;
        RECT 56.220 18.060 56.480 18.320 ;
        RECT 366.260 18.060 366.520 18.320 ;
      LAYER met2 ;
        RECT 369.340 1600.450 369.620 1604.000 ;
        RECT 368.160 1600.310 369.620 1600.450 ;
        RECT 368.160 1576.570 368.300 1600.310 ;
        RECT 369.340 1600.000 369.620 1600.310 ;
        RECT 366.260 1576.250 366.520 1576.570 ;
        RECT 368.100 1576.250 368.360 1576.570 ;
        RECT 366.320 18.350 366.460 1576.250 ;
        RECT 56.220 18.030 56.480 18.350 ;
        RECT 366.260 18.030 366.520 18.350 ;
        RECT 56.280 2.400 56.420 18.030 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 80.110 16.900 80.430 16.960 ;
        RECT 82.410 16.900 82.730 16.960 ;
        RECT 80.110 16.760 82.730 16.900 ;
        RECT 80.110 16.700 80.430 16.760 ;
        RECT 82.410 16.700 82.730 16.760 ;
      LAYER via ;
        RECT 80.140 16.700 80.400 16.960 ;
        RECT 82.440 16.700 82.700 16.960 ;
      LAYER met2 ;
        RECT 377.620 1600.380 377.900 1604.000 ;
        RECT 377.620 1600.000 377.960 1600.380 ;
        RECT 377.820 1591.725 377.960 1600.000 ;
        RECT 82.430 1591.355 82.710 1591.725 ;
        RECT 377.750 1591.355 378.030 1591.725 ;
        RECT 82.500 16.990 82.640 1591.355 ;
        RECT 80.140 16.670 80.400 16.990 ;
        RECT 82.440 16.670 82.700 16.990 ;
        RECT 80.200 2.400 80.340 16.670 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 82.430 1591.400 82.710 1591.680 ;
        RECT 377.750 1591.400 378.030 1591.680 ;
      LAYER met3 ;
        RECT 82.405 1591.690 82.735 1591.705 ;
        RECT 377.725 1591.690 378.055 1591.705 ;
        RECT 82.405 1591.390 378.055 1591.690 ;
        RECT 82.405 1591.375 82.735 1591.390 ;
        RECT 377.725 1591.375 378.055 1591.390 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 380.030 1579.880 380.350 1579.940 ;
        RECT 384.630 1579.880 384.950 1579.940 ;
        RECT 380.030 1579.740 384.950 1579.880 ;
        RECT 380.030 1579.680 380.350 1579.740 ;
        RECT 384.630 1579.680 384.950 1579.740 ;
        RECT 103.570 19.280 103.890 19.340 ;
        RECT 380.030 19.280 380.350 19.340 ;
        RECT 103.570 19.140 380.350 19.280 ;
        RECT 103.570 19.080 103.890 19.140 ;
        RECT 380.030 19.080 380.350 19.140 ;
      LAYER via ;
        RECT 380.060 1579.680 380.320 1579.940 ;
        RECT 384.660 1579.680 384.920 1579.940 ;
        RECT 103.600 19.080 103.860 19.340 ;
        RECT 380.060 19.080 380.320 19.340 ;
      LAYER met2 ;
        RECT 385.900 1600.450 386.180 1604.000 ;
        RECT 384.720 1600.310 386.180 1600.450 ;
        RECT 384.720 1579.970 384.860 1600.310 ;
        RECT 385.900 1600.000 386.180 1600.310 ;
        RECT 380.060 1579.650 380.320 1579.970 ;
        RECT 384.660 1579.650 384.920 1579.970 ;
        RECT 380.120 19.370 380.260 1579.650 ;
        RECT 103.600 19.050 103.860 19.370 ;
        RECT 380.060 19.050 380.320 19.370 ;
        RECT 103.660 2.400 103.800 19.050 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 375.045 1590.095 375.215 1590.435 ;
        RECT 376.425 1590.095 376.595 1592.135 ;
        RECT 375.045 1589.925 376.595 1590.095 ;
      LAYER mcon ;
        RECT 376.425 1591.965 376.595 1592.135 ;
        RECT 375.045 1590.265 375.215 1590.435 ;
      LAYER met1 ;
        RECT 376.365 1592.120 376.655 1592.165 ;
        RECT 394.290 1592.120 394.610 1592.180 ;
        RECT 376.365 1591.980 394.610 1592.120 ;
        RECT 376.365 1591.935 376.655 1591.980 ;
        RECT 394.290 1591.920 394.610 1591.980 ;
        RECT 130.710 1590.760 131.030 1590.820 ;
        RECT 130.710 1590.620 372.440 1590.760 ;
        RECT 130.710 1590.560 131.030 1590.620 ;
        RECT 372.300 1590.420 372.440 1590.620 ;
        RECT 374.985 1590.420 375.275 1590.465 ;
        RECT 372.300 1590.280 375.275 1590.420 ;
        RECT 374.985 1590.235 375.275 1590.280 ;
        RECT 127.490 16.900 127.810 16.960 ;
        RECT 130.710 16.900 131.030 16.960 ;
        RECT 127.490 16.760 131.030 16.900 ;
        RECT 127.490 16.700 127.810 16.760 ;
        RECT 130.710 16.700 131.030 16.760 ;
      LAYER via ;
        RECT 394.320 1591.920 394.580 1592.180 ;
        RECT 130.740 1590.560 131.000 1590.820 ;
        RECT 127.520 16.700 127.780 16.960 ;
        RECT 130.740 16.700 131.000 16.960 ;
      LAYER met2 ;
        RECT 394.180 1600.380 394.460 1604.000 ;
        RECT 394.180 1600.000 394.520 1600.380 ;
        RECT 394.380 1592.210 394.520 1600.000 ;
        RECT 394.320 1591.890 394.580 1592.210 ;
        RECT 130.740 1590.530 131.000 1590.850 ;
        RECT 130.800 16.990 130.940 1590.530 ;
        RECT 127.520 16.670 127.780 16.990 ;
        RECT 130.740 16.670 131.000 16.990 ;
        RECT 127.580 2.400 127.720 16.670 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 358.760 1600.380 359.040 1604.000 ;
        RECT 358.760 1600.000 359.100 1600.380 ;
        RECT 358.960 20.810 359.100 1600.000 ;
        RECT 358.500 20.670 359.100 20.810 ;
        RECT 358.500 16.845 358.640 20.670 ;
        RECT 26.310 16.475 26.590 16.845 ;
        RECT 358.430 16.475 358.710 16.845 ;
        RECT 26.380 2.400 26.520 16.475 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 26.310 16.520 26.590 16.800 ;
        RECT 358.430 16.520 358.710 16.800 ;
      LAYER met3 ;
        RECT 26.285 16.810 26.615 16.825 ;
        RECT 358.405 16.810 358.735 16.825 ;
        RECT 26.285 16.510 358.735 16.810 ;
        RECT 26.285 16.495 26.615 16.510 ;
        RECT 358.405 16.495 358.735 16.510 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 17.580 32.590 17.640 ;
        RECT 359.790 17.580 360.110 17.640 ;
        RECT 32.270 17.440 360.110 17.580 ;
        RECT 32.270 17.380 32.590 17.440 ;
        RECT 359.790 17.380 360.110 17.440 ;
      LAYER via ;
        RECT 32.300 17.380 32.560 17.640 ;
        RECT 359.820 17.380 360.080 17.640 ;
      LAYER met2 ;
        RECT 361.060 1600.450 361.340 1604.000 ;
        RECT 359.880 1600.310 361.340 1600.450 ;
        RECT 359.880 17.670 360.020 1600.310 ;
        RECT 361.060 1600.000 361.340 1600.310 ;
        RECT 32.300 17.350 32.560 17.670 ;
        RECT 359.820 17.350 360.080 17.670 ;
        RECT 32.360 2.400 32.500 17.350 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 584.345 2836.365 584.515 2841.295 ;
      LAYER mcon ;
        RECT 584.345 2841.125 584.515 2841.295 ;
      LAYER met1 ;
        RECT 551.610 2842.300 551.930 2842.360 ;
        RECT 679.490 2842.300 679.810 2842.360 ;
        RECT 551.610 2842.160 679.810 2842.300 ;
        RECT 551.610 2842.100 551.930 2842.160 ;
        RECT 679.490 2842.100 679.810 2842.160 ;
        RECT 503.310 2841.280 503.630 2841.340 ;
        RECT 545.170 2841.280 545.490 2841.340 ;
        RECT 584.285 2841.280 584.575 2841.325 ;
        RECT 503.310 2841.140 584.575 2841.280 ;
        RECT 503.310 2841.080 503.630 2841.140 ;
        RECT 545.170 2841.080 545.490 2841.140 ;
        RECT 584.285 2841.095 584.575 2841.140 ;
        RECT 638.090 2837.200 638.410 2837.260 ;
        RECT 624.840 2837.060 638.410 2837.200 ;
        RECT 624.840 2836.860 624.980 2837.060 ;
        RECT 638.090 2837.000 638.410 2837.060 ;
        RECT 603.680 2836.720 624.980 2836.860 ;
        RECT 584.285 2836.520 584.575 2836.565 ;
        RECT 591.630 2836.520 591.950 2836.580 ;
        RECT 603.680 2836.520 603.820 2836.720 ;
        RECT 584.285 2836.380 603.820 2836.520 ;
        RECT 584.285 2836.335 584.575 2836.380 ;
        RECT 591.630 2836.320 591.950 2836.380 ;
        RECT 1089.810 2619.260 1090.130 2619.320 ;
        RECT 1173.990 2619.260 1174.310 2619.320 ;
        RECT 1089.810 2619.120 1174.310 2619.260 ;
        RECT 1089.810 2619.060 1090.130 2619.120 ;
        RECT 1173.990 2619.060 1174.310 2619.120 ;
        RECT 638.090 2617.560 638.410 2617.620 ;
        RECT 735.610 2617.560 735.930 2617.620 ;
        RECT 638.090 2617.420 735.930 2617.560 ;
        RECT 638.090 2617.360 638.410 2617.420 ;
        RECT 735.610 2617.360 735.930 2617.420 ;
        RECT 679.490 2615.860 679.810 2615.920 ;
        RECT 888.330 2615.860 888.650 2615.920 ;
        RECT 679.490 2615.720 888.650 2615.860 ;
        RECT 679.490 2615.660 679.810 2615.720 ;
        RECT 888.330 2615.660 888.650 2615.720 ;
      LAYER via ;
        RECT 551.640 2842.100 551.900 2842.360 ;
        RECT 679.520 2842.100 679.780 2842.360 ;
        RECT 503.340 2841.080 503.600 2841.340 ;
        RECT 545.200 2841.080 545.460 2841.340 ;
        RECT 638.120 2837.000 638.380 2837.260 ;
        RECT 591.660 2836.320 591.920 2836.580 ;
        RECT 1089.840 2619.060 1090.100 2619.320 ;
        RECT 1174.020 2619.060 1174.280 2619.320 ;
        RECT 638.120 2617.360 638.380 2617.620 ;
        RECT 735.640 2617.360 735.900 2617.620 ;
        RECT 679.520 2615.660 679.780 2615.920 ;
        RECT 888.360 2615.660 888.620 2615.920 ;
      LAYER met2 ;
        RECT 545.190 2850.715 545.470 2851.085 ;
        RECT 503.330 2841.195 503.610 2841.565 ;
        RECT 545.260 2841.370 545.400 2850.715 ;
        RECT 591.650 2848.675 591.930 2849.045 ;
        RECT 551.630 2842.555 551.910 2842.925 ;
        RECT 551.700 2842.390 551.840 2842.555 ;
        RECT 551.640 2842.070 551.900 2842.390 ;
        RECT 503.340 2841.050 503.600 2841.195 ;
        RECT 545.200 2841.050 545.460 2841.370 ;
        RECT 591.720 2836.610 591.860 2848.675 ;
        RECT 679.520 2842.070 679.780 2842.390 ;
        RECT 638.120 2836.970 638.380 2837.290 ;
        RECT 591.660 2836.290 591.920 2836.610 ;
        RECT 638.180 2836.125 638.320 2836.970 ;
        RECT 638.110 2835.755 638.390 2836.125 ;
        RECT 638.180 2617.650 638.320 2835.755 ;
        RECT 638.120 2617.330 638.380 2617.650 ;
        RECT 679.580 2615.950 679.720 2842.070 ;
        RECT 1089.830 2836.435 1090.110 2836.805 ;
        RECT 1089.900 2619.350 1090.040 2836.435 ;
        RECT 1089.840 2619.030 1090.100 2619.350 ;
        RECT 1174.020 2619.030 1174.280 2619.350 ;
        RECT 735.640 2617.330 735.900 2617.650 ;
        RECT 679.520 2615.630 679.780 2615.950 ;
        RECT 735.700 2610.000 735.840 2617.330 ;
        RECT 888.360 2615.630 888.620 2615.950 ;
        RECT 888.420 2610.000 888.560 2615.630 ;
        RECT 1174.080 2610.000 1174.220 2619.030 ;
        RECT 735.500 2609.500 735.840 2610.000 ;
        RECT 888.220 2609.500 888.560 2610.000 ;
        RECT 1173.880 2609.500 1174.220 2610.000 ;
        RECT 735.500 2606.000 735.780 2609.500 ;
        RECT 888.220 2606.000 888.500 2609.500 ;
        RECT 1173.880 2606.000 1174.160 2609.500 ;
      LAYER via2 ;
        RECT 545.190 2850.760 545.470 2851.040 ;
        RECT 503.330 2841.240 503.610 2841.520 ;
        RECT 591.650 2848.720 591.930 2849.000 ;
        RECT 551.630 2842.600 551.910 2842.880 ;
        RECT 638.110 2835.800 638.390 2836.080 ;
        RECT 1089.830 2836.480 1090.110 2836.760 ;
      LAYER met3 ;
        RECT 543.990 2851.050 544.370 2851.060 ;
        RECT 545.165 2851.050 545.495 2851.065 ;
        RECT 543.990 2850.750 545.495 2851.050 ;
        RECT 543.990 2850.740 544.370 2850.750 ;
        RECT 545.165 2850.735 545.495 2850.750 ;
        RECT 591.625 2849.020 591.955 2849.025 ;
        RECT 591.625 2849.010 592.030 2849.020 ;
        RECT 591.625 2848.710 592.410 2849.010 ;
        RECT 591.625 2848.700 592.030 2848.710 ;
        RECT 591.625 2848.695 591.955 2848.700 ;
        RECT 548.590 2842.890 548.970 2842.900 ;
        RECT 551.605 2842.890 551.935 2842.905 ;
        RECT 548.590 2842.590 551.935 2842.890 ;
        RECT 548.590 2842.580 548.970 2842.590 ;
        RECT 551.605 2842.575 551.935 2842.590 ;
        RECT 497.990 2841.530 498.370 2841.540 ;
        RECT 503.305 2841.530 503.635 2841.545 ;
        RECT 497.990 2841.230 503.635 2841.530 ;
        RECT 497.990 2841.220 498.370 2841.230 ;
        RECT 503.305 2841.215 503.635 2841.230 ;
        RECT 1087.710 2836.770 1088.090 2836.780 ;
        RECT 1089.805 2836.770 1090.135 2836.785 ;
        RECT 1087.710 2836.470 1090.135 2836.770 ;
        RECT 1087.710 2836.460 1088.090 2836.470 ;
        RECT 1089.805 2836.455 1090.135 2836.470 ;
        RECT 638.085 2836.090 638.415 2836.105 ;
        RECT 638.750 2836.090 639.130 2836.100 ;
        RECT 638.085 2835.790 639.130 2836.090 ;
        RECT 638.085 2835.775 638.415 2835.790 ;
        RECT 638.750 2835.780 639.130 2835.790 ;
      LAYER via3 ;
        RECT 544.020 2850.740 544.340 2851.060 ;
        RECT 591.680 2848.700 592.000 2849.020 ;
        RECT 548.620 2842.580 548.940 2842.900 ;
        RECT 498.020 2841.220 498.340 2841.540 ;
        RECT 1087.740 2836.460 1088.060 2836.780 ;
        RECT 638.780 2835.780 639.100 2836.100 ;
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 364.020 -9.320 367.020 3529.000 ;
        RECT 544.020 3306.235 547.020 3529.000 ;
        RECT 724.020 3306.235 727.020 3529.000 ;
        RECT 543.945 3301.635 544.245 3306.235 ;
        RECT 498.250 2851.050 498.550 2854.600 ;
        RECT 498.030 2850.000 498.550 2851.050 ;
        RECT 544.015 2851.050 544.345 2851.065 ;
        RECT 544.970 2851.050 545.270 2854.600 ;
        RECT 544.015 2850.750 545.270 2851.050 ;
        RECT 544.015 2850.735 544.345 2850.750 ;
        RECT 544.970 2850.000 545.270 2850.750 ;
        RECT 545.590 2851.050 545.890 2854.600 ;
        RECT 545.590 2850.750 548.930 2851.050 ;
        RECT 545.590 2850.000 545.890 2850.750 ;
        RECT 498.030 2841.545 498.330 2850.000 ;
        RECT 498.015 2841.215 498.345 2841.545 ;
        RECT 544.020 -9.320 547.020 2850.000 ;
        RECT 548.630 2842.905 548.930 2850.750 ;
        RECT 591.690 2849.025 591.990 2854.600 ;
        RECT 591.675 2848.695 592.005 2849.025 ;
        RECT 638.410 2847.650 638.710 2854.600 ;
        RECT 638.410 2847.350 639.090 2847.650 ;
        RECT 548.615 2842.575 548.945 2842.905 ;
        RECT 638.790 2836.105 639.090 2847.350 ;
        RECT 638.775 2835.775 639.105 2836.105 ;
        RECT 724.020 -9.320 727.020 2850.000 ;
        RECT 904.020 -9.320 907.020 3529.000 ;
        RECT 1084.020 3306.235 1087.020 3529.000 ;
        RECT 1264.020 3306.235 1267.020 3529.000 ;
        RECT 1083.910 2851.050 1084.210 2854.600 ;
        RECT 1083.910 2850.750 1088.050 2851.050 ;
        RECT 1083.910 2850.000 1084.210 2850.750 ;
        RECT 1084.020 -9.320 1087.020 2850.000 ;
        RECT 1087.750 2836.785 1088.050 2850.750 ;
        RECT 1087.735 2836.455 1088.065 2836.785 ;
        RECT 1264.020 -9.320 1267.020 2850.000 ;
        RECT 1444.020 -9.320 1447.020 3529.000 ;
        RECT 1624.020 2586.480 1627.020 3529.000 ;
        RECT 1804.020 2586.480 1807.020 3529.000 ;
        RECT 1984.020 2586.480 1987.020 3529.000 ;
        RECT 1624.020 1986.480 1627.020 2200.000 ;
        RECT 1804.020 1986.480 1807.020 2200.000 ;
        RECT 1984.020 1986.480 1987.020 2200.000 ;
        RECT 1624.020 -9.320 1627.020 1600.000 ;
        RECT 1804.020 -9.320 1807.020 1600.000 ;
        RECT 1984.020 -9.320 1987.020 1600.000 ;
        RECT 2164.020 -9.320 2167.020 3529.000 ;
        RECT 2344.020 -9.320 2347.020 3529.000 ;
        RECT 2524.020 -9.320 2527.020 3529.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1085.670 2841.620 1085.990 2841.680 ;
        RECT 1129.370 2841.620 1129.690 2841.680 ;
        RECT 1173.070 2841.620 1173.390 2841.680 ;
        RECT 1085.670 2841.480 1173.390 2841.620 ;
        RECT 1085.670 2841.420 1085.990 2841.480 ;
        RECT 1129.370 2841.420 1129.690 2841.480 ;
        RECT 1173.070 2841.420 1173.390 2841.480 ;
        RECT 1041.510 2839.240 1041.830 2839.300 ;
        RECT 1085.670 2839.240 1085.990 2839.300 ;
        RECT 1041.510 2839.100 1085.990 2839.240 ;
        RECT 1041.510 2839.040 1041.830 2839.100 ;
        RECT 1085.670 2839.040 1085.990 2839.100 ;
        RECT 641.310 2837.200 641.630 2837.260 ;
        RECT 1035.070 2837.200 1035.390 2837.260 ;
        RECT 1041.510 2837.200 1041.830 2837.260 ;
        RECT 641.310 2837.060 1041.830 2837.200 ;
        RECT 641.310 2837.000 641.630 2837.060 ;
        RECT 1035.070 2837.000 1035.390 2837.060 ;
        RECT 1041.510 2837.000 1041.830 2837.060 ;
      LAYER via ;
        RECT 1085.700 2841.420 1085.960 2841.680 ;
        RECT 1129.400 2841.420 1129.660 2841.680 ;
        RECT 1173.100 2841.420 1173.360 2841.680 ;
        RECT 1041.540 2839.040 1041.800 2839.300 ;
        RECT 1085.700 2839.040 1085.960 2839.300 ;
        RECT 641.340 2837.000 641.600 2837.260 ;
        RECT 1035.100 2837.000 1035.360 2837.260 ;
        RECT 1041.540 2837.000 1041.800 2837.260 ;
      LAYER met2 ;
        RECT 1035.090 2842.555 1035.370 2842.925 ;
        RECT 1085.690 2842.555 1085.970 2842.925 ;
        RECT 1129.390 2842.555 1129.670 2842.925 ;
        RECT 365.330 2839.155 365.610 2839.525 ;
        RECT 363.820 2609.570 364.100 2610.000 ;
        RECT 365.400 2609.570 365.540 2839.155 ;
        RECT 1035.160 2837.290 1035.300 2842.555 ;
        RECT 1085.760 2841.710 1085.900 2842.555 ;
        RECT 1129.460 2841.710 1129.600 2842.555 ;
        RECT 1173.090 2841.875 1173.370 2842.245 ;
        RECT 1173.160 2841.710 1173.300 2841.875 ;
        RECT 1085.700 2841.390 1085.960 2841.710 ;
        RECT 1129.400 2841.390 1129.660 2841.710 ;
        RECT 1173.100 2841.390 1173.360 2841.710 ;
        RECT 1085.760 2839.330 1085.900 2841.390 ;
        RECT 1041.540 2839.010 1041.800 2839.330 ;
        RECT 1085.700 2839.010 1085.960 2839.330 ;
        RECT 1041.600 2837.290 1041.740 2839.010 ;
        RECT 641.340 2836.970 641.600 2837.290 ;
        RECT 1035.100 2836.970 1035.360 2837.290 ;
        RECT 1041.540 2836.970 1041.800 2837.290 ;
        RECT 363.820 2609.430 365.540 2609.570 ;
        RECT 640.280 2609.570 640.560 2610.000 ;
        RECT 641.400 2609.570 641.540 2836.970 ;
        RECT 640.280 2609.430 641.540 2609.570 ;
        RECT 363.820 2606.000 364.100 2609.430 ;
        RECT 640.280 2606.000 640.560 2609.430 ;
      LAYER via2 ;
        RECT 1035.090 2842.600 1035.370 2842.880 ;
        RECT 1085.690 2842.600 1085.970 2842.880 ;
        RECT 1129.390 2842.600 1129.670 2842.880 ;
        RECT 365.330 2839.200 365.610 2839.480 ;
        RECT 1173.090 2841.920 1173.370 2842.200 ;
      LAYER met3 ;
        RECT 1035.065 2842.900 1035.395 2842.905 ;
        RECT 1035.065 2842.890 1035.650 2842.900 ;
        RECT 1083.110 2842.890 1083.490 2842.900 ;
        RECT 1085.665 2842.890 1085.995 2842.905 ;
        RECT 1129.365 2842.900 1129.695 2842.905 ;
        RECT 1129.110 2842.890 1129.695 2842.900 ;
        RECT 1035.065 2842.590 1035.850 2842.890 ;
        RECT 1083.110 2842.590 1085.995 2842.890 ;
        RECT 1128.910 2842.590 1129.695 2842.890 ;
        RECT 1035.065 2842.580 1035.650 2842.590 ;
        RECT 1083.110 2842.580 1083.490 2842.590 ;
        RECT 1035.065 2842.575 1035.395 2842.580 ;
        RECT 1085.665 2842.575 1085.995 2842.590 ;
        RECT 1129.110 2842.580 1129.695 2842.590 ;
        RECT 1129.365 2842.575 1129.695 2842.580 ;
        RECT 1173.065 2842.220 1173.395 2842.225 ;
        RECT 1173.065 2842.210 1173.650 2842.220 ;
        RECT 1172.840 2841.910 1173.650 2842.210 ;
        RECT 1173.065 2841.900 1173.650 2841.910 ;
        RECT 1173.065 2841.895 1173.395 2841.900 ;
        RECT 365.305 2839.490 365.635 2839.505 ;
        RECT 997.550 2839.490 997.930 2839.500 ;
        RECT 365.305 2839.190 997.930 2839.490 ;
        RECT 365.305 2839.175 365.635 2839.190 ;
        RECT 997.550 2839.180 997.930 2839.190 ;
      LAYER via3 ;
        RECT 1035.300 2842.580 1035.620 2842.900 ;
        RECT 1083.140 2842.580 1083.460 2842.900 ;
        RECT 1129.140 2842.580 1129.460 2842.900 ;
        RECT 1173.300 2841.900 1173.620 2842.220 ;
        RECT 997.580 2839.180 997.900 2839.500 ;
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 454.020 3306.235 457.020 3529.000 ;
        RECT 634.020 3306.235 637.020 3529.000 ;
        RECT 454.020 -9.320 457.020 2850.000 ;
        RECT 634.020 -9.320 637.020 2850.000 ;
        RECT 814.020 -9.320 817.020 3529.000 ;
        RECT 994.020 3306.235 997.020 3529.000 ;
        RECT 1174.020 3306.235 1177.020 3529.000 ;
        RECT 1175.065 3301.635 1175.365 3306.235 ;
        RECT 995.690 2851.050 995.990 2854.600 ;
        RECT 1036.570 2852.750 1036.870 2854.600 ;
        RECT 1035.310 2852.450 1036.870 2852.750 ;
        RECT 995.690 2850.750 997.890 2851.050 ;
        RECT 995.690 2850.000 995.990 2850.750 ;
        RECT 994.020 -9.320 997.020 2850.000 ;
        RECT 997.590 2839.505 997.890 2850.750 ;
        RECT 1035.310 2842.905 1035.610 2852.450 ;
        RECT 1036.570 2850.000 1036.870 2852.450 ;
        RECT 1083.290 2851.050 1083.590 2854.600 ;
        RECT 1130.010 2851.050 1130.310 2854.600 ;
        RECT 1176.730 2851.050 1177.030 2854.600 ;
        RECT 1083.150 2850.000 1083.590 2851.050 ;
        RECT 1129.150 2850.750 1130.310 2851.050 ;
        RECT 1083.150 2842.905 1083.450 2850.000 ;
        RECT 1129.150 2842.905 1129.450 2850.750 ;
        RECT 1130.010 2850.000 1130.310 2850.750 ;
        RECT 1173.310 2850.750 1177.030 2851.050 ;
        RECT 1035.295 2842.575 1035.625 2842.905 ;
        RECT 1083.135 2842.575 1083.465 2842.905 ;
        RECT 1129.135 2842.575 1129.465 2842.905 ;
        RECT 1173.310 2842.225 1173.610 2850.750 ;
        RECT 1176.730 2850.000 1177.030 2850.750 ;
        RECT 1173.295 2841.895 1173.625 2842.225 ;
        RECT 997.575 2839.175 997.905 2839.505 ;
        RECT 1174.020 -9.320 1177.020 2850.000 ;
        RECT 1354.020 -9.320 1357.020 3529.000 ;
        RECT 1534.020 -9.320 1537.020 3529.000 ;
        RECT 1714.020 2586.480 1717.020 3529.000 ;
        RECT 1894.020 2586.480 1897.020 3529.000 ;
        RECT 1714.020 1986.480 1717.020 2200.000 ;
        RECT 1894.020 1986.480 1897.020 2200.000 ;
        RECT 1714.020 -9.320 1717.020 1600.000 ;
        RECT 1894.020 -9.320 1897.020 1600.000 ;
        RECT 2074.020 -9.320 2077.020 3529.000 ;
        RECT 2254.020 -9.320 2257.020 3529.000 ;
        RECT 2434.020 -9.320 2437.020 3529.000 ;
        RECT 2614.020 -9.320 2617.020 3529.000 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 576.985 2836.705 577.155 2840.275 ;
      LAYER mcon ;
        RECT 576.985 2840.105 577.155 2840.275 ;
      LAYER met1 ;
        RECT 475.710 2842.640 476.030 2842.700 ;
        RECT 515.730 2842.640 516.050 2842.700 ;
        RECT 475.710 2842.500 516.050 2842.640 ;
        RECT 475.710 2842.440 476.030 2842.500 ;
        RECT 515.730 2842.440 516.050 2842.500 ;
        RECT 589.790 2841.960 590.110 2842.020 ;
        RECT 686.390 2841.960 686.710 2842.020 ;
        RECT 589.790 2841.820 686.710 2841.960 ;
        RECT 589.790 2841.760 590.110 2841.820 ;
        RECT 686.390 2841.760 686.710 2841.820 ;
        RECT 515.730 2840.260 516.050 2840.320 ;
        RECT 561.270 2840.260 561.590 2840.320 ;
        RECT 576.925 2840.260 577.215 2840.305 ;
        RECT 515.730 2840.120 577.215 2840.260 ;
        RECT 515.730 2840.060 516.050 2840.120 ;
        RECT 561.270 2840.060 561.590 2840.120 ;
        RECT 576.925 2840.075 577.215 2840.120 ;
        RECT 576.925 2836.860 577.215 2836.905 ;
        RECT 603.130 2836.860 603.450 2836.920 ;
        RECT 576.925 2836.720 603.450 2836.860 ;
        RECT 576.925 2836.675 577.215 2836.720 ;
        RECT 603.130 2836.660 603.450 2836.720 ;
        RECT 686.390 2616.540 686.710 2616.600 ;
        RECT 916.850 2616.540 917.170 2616.600 ;
        RECT 686.390 2616.400 917.170 2616.540 ;
        RECT 686.390 2616.340 686.710 2616.400 ;
        RECT 916.850 2616.340 917.170 2616.400 ;
        RECT 610.490 2616.200 610.810 2616.260 ;
        RECT 688.230 2616.200 688.550 2616.260 ;
        RECT 610.490 2616.060 688.550 2616.200 ;
        RECT 610.490 2616.000 610.810 2616.060 ;
        RECT 688.230 2616.000 688.550 2616.060 ;
      LAYER via ;
        RECT 475.740 2842.440 476.000 2842.700 ;
        RECT 515.760 2842.440 516.020 2842.700 ;
        RECT 589.820 2841.760 590.080 2842.020 ;
        RECT 686.420 2841.760 686.680 2842.020 ;
        RECT 515.760 2840.060 516.020 2840.320 ;
        RECT 561.300 2840.060 561.560 2840.320 ;
        RECT 603.160 2836.660 603.420 2836.920 ;
        RECT 686.420 2616.340 686.680 2616.600 ;
        RECT 916.880 2616.340 917.140 2616.600 ;
        RECT 610.520 2616.000 610.780 2616.260 ;
        RECT 688.260 2616.000 688.520 2616.260 ;
      LAYER met2 ;
        RECT 561.290 2850.715 561.570 2851.085 ;
        RECT 589.810 2850.715 590.090 2851.085 ;
        RECT 475.730 2842.555 476.010 2842.925 ;
        RECT 515.750 2842.555 516.030 2842.925 ;
        RECT 475.740 2842.410 476.000 2842.555 ;
        RECT 515.760 2842.410 516.020 2842.555 ;
        RECT 515.820 2840.350 515.960 2842.410 ;
        RECT 561.360 2840.350 561.500 2850.715 ;
        RECT 589.880 2842.050 590.020 2850.715 ;
        RECT 589.820 2841.730 590.080 2842.050 ;
        RECT 686.420 2841.730 686.680 2842.050 ;
        RECT 515.760 2840.030 516.020 2840.350 ;
        RECT 561.300 2840.030 561.560 2840.350 ;
        RECT 603.160 2836.805 603.420 2836.950 ;
        RECT 603.150 2836.435 603.430 2836.805 ;
        RECT 610.510 2830.315 610.790 2830.685 ;
        RECT 610.580 2616.290 610.720 2830.315 ;
        RECT 686.480 2616.630 686.620 2841.730 ;
        RECT 686.420 2616.310 686.680 2616.630 ;
        RECT 916.880 2616.310 917.140 2616.630 ;
        RECT 610.520 2615.970 610.780 2616.290 ;
        RECT 688.260 2615.970 688.520 2616.290 ;
        RECT 688.320 2610.000 688.460 2615.970 ;
        RECT 916.940 2610.000 917.080 2616.310 ;
        RECT 688.120 2609.500 688.460 2610.000 ;
        RECT 916.740 2609.500 917.080 2610.000 ;
        RECT 688.120 2606.000 688.400 2609.500 ;
        RECT 916.740 2606.000 917.020 2609.500 ;
      LAYER via2 ;
        RECT 561.290 2850.760 561.570 2851.040 ;
        RECT 589.810 2850.760 590.090 2851.040 ;
        RECT 475.730 2842.600 476.010 2842.880 ;
        RECT 515.750 2842.600 516.030 2842.880 ;
        RECT 603.150 2836.480 603.430 2836.760 ;
        RECT 610.510 2830.360 610.790 2830.640 ;
      LAYER met3 ;
        RECT 561.265 2851.060 561.595 2851.065 ;
        RECT 561.265 2851.050 561.850 2851.060 ;
        RECT 566.070 2851.050 566.450 2851.060 ;
        RECT 589.785 2851.050 590.115 2851.065 ;
        RECT 561.265 2850.750 562.050 2851.050 ;
        RECT 566.070 2850.750 590.115 2851.050 ;
        RECT 561.265 2850.740 561.850 2850.750 ;
        RECT 566.070 2850.740 566.450 2850.750 ;
        RECT 561.265 2850.735 561.595 2850.740 ;
        RECT 589.785 2850.735 590.115 2850.750 ;
        RECT 469.470 2842.890 469.850 2842.900 ;
        RECT 475.705 2842.890 476.035 2842.905 ;
        RECT 515.725 2842.900 516.055 2842.905 ;
        RECT 469.470 2842.590 476.035 2842.890 ;
        RECT 469.470 2842.580 469.850 2842.590 ;
        RECT 475.705 2842.575 476.035 2842.590 ;
        RECT 515.470 2842.890 516.055 2842.900 ;
        RECT 515.470 2842.590 516.280 2842.890 ;
        RECT 515.470 2842.580 516.055 2842.590 ;
        RECT 515.725 2842.575 516.055 2842.580 ;
        RECT 603.125 2836.770 603.455 2836.785 ;
        RECT 607.470 2836.770 607.850 2836.780 ;
        RECT 603.125 2836.470 607.850 2836.770 ;
        RECT 603.125 2836.455 603.455 2836.470 ;
        RECT 607.470 2836.460 607.850 2836.470 ;
        RECT 607.470 2830.650 607.850 2830.660 ;
        RECT 610.485 2830.650 610.815 2830.665 ;
        RECT 607.470 2830.350 610.815 2830.650 ;
        RECT 607.470 2830.340 607.850 2830.350 ;
        RECT 610.485 2830.335 610.815 2830.350 ;
      LAYER via3 ;
        RECT 561.500 2850.740 561.820 2851.060 ;
        RECT 566.100 2850.740 566.420 2851.060 ;
        RECT 469.500 2842.580 469.820 2842.900 ;
        RECT 515.500 2842.580 515.820 2842.900 ;
        RECT 607.500 2836.460 607.820 2836.780 ;
        RECT 607.500 2830.340 607.820 2830.660 ;
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 382.020 -18.720 385.020 3538.400 ;
        RECT 562.020 3306.235 565.020 3538.400 ;
        RECT 742.020 3306.235 745.020 3538.400 ;
        RECT 562.665 3301.635 562.965 3306.235 ;
        RECT 742.890 3301.635 743.190 3306.235 ;
        RECT 469.050 2847.650 469.350 2854.600 ;
        RECT 515.770 2851.050 516.070 2854.600 ;
        RECT 515.510 2850.000 516.070 2851.050 ;
        RECT 561.495 2851.050 561.825 2851.065 ;
        RECT 562.490 2851.050 562.790 2854.600 ;
        RECT 561.495 2850.750 562.790 2851.050 ;
        RECT 561.495 2850.735 561.825 2850.750 ;
        RECT 562.490 2850.000 562.790 2850.750 ;
        RECT 563.110 2851.050 563.410 2854.600 ;
        RECT 566.095 2851.050 566.425 2851.065 ;
        RECT 609.210 2851.050 609.510 2854.600 ;
        RECT 563.110 2850.750 566.425 2851.050 ;
        RECT 563.110 2850.000 563.410 2850.750 ;
        RECT 566.095 2850.735 566.425 2850.750 ;
        RECT 607.510 2850.750 609.510 2851.050 ;
        RECT 469.050 2847.350 469.810 2847.650 ;
        RECT 469.510 2842.905 469.810 2847.350 ;
        RECT 515.510 2842.905 515.810 2850.000 ;
        RECT 469.495 2842.575 469.825 2842.905 ;
        RECT 515.495 2842.575 515.825 2842.905 ;
        RECT 562.020 -18.720 565.020 2850.000 ;
        RECT 607.510 2836.785 607.810 2850.750 ;
        RECT 609.210 2850.000 609.510 2850.750 ;
        RECT 607.495 2836.455 607.825 2836.785 ;
        RECT 607.510 2830.665 607.810 2836.455 ;
        RECT 607.495 2830.335 607.825 2830.665 ;
        RECT 742.020 -18.720 745.020 2850.000 ;
        RECT 922.020 -18.720 925.020 3538.400 ;
        RECT 1102.020 3306.235 1105.020 3538.400 ;
        RECT 1282.020 3306.235 1285.020 3538.400 ;
        RECT 1102.020 -18.720 1105.020 2850.000 ;
        RECT 1282.020 -18.720 1285.020 2850.000 ;
        RECT 1462.020 -18.720 1465.020 3538.400 ;
        RECT 1642.020 2586.480 1645.020 3538.400 ;
        RECT 1822.020 2586.480 1825.020 3538.400 ;
        RECT 2002.020 2586.480 2005.020 3538.400 ;
        RECT 1642.020 1986.480 1645.020 2200.000 ;
        RECT 1822.020 1986.480 1825.020 2200.000 ;
        RECT 2002.020 1986.480 2005.020 2200.000 ;
        RECT 1642.020 -18.720 1645.020 1600.000 ;
        RECT 1822.020 -18.720 1825.020 1600.000 ;
        RECT 2002.020 -18.720 2005.020 1600.000 ;
        RECT 2182.020 -18.720 2185.020 3538.400 ;
        RECT 2362.020 -18.720 2365.020 3538.400 ;
        RECT 2542.020 -18.720 2545.020 3538.400 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1217.305 2618.255 1217.475 2619.275 ;
        RECT 1218.685 2618.255 1218.855 2618.595 ;
        RECT 1217.305 2618.085 1218.855 2618.255 ;
      LAYER mcon ;
        RECT 1217.305 2619.105 1217.475 2619.275 ;
        RECT 1218.685 2618.425 1218.855 2618.595 ;
      LAYER met1 ;
        RECT 617.390 2840.600 617.710 2840.660 ;
        RECT 589.880 2840.460 617.710 2840.600 ;
        RECT 474.330 2839.240 474.650 2839.300 ;
        RECT 520.330 2839.240 520.650 2839.300 ;
        RECT 568.170 2839.240 568.490 2839.300 ;
        RECT 589.880 2839.240 590.020 2840.460 ;
        RECT 617.390 2840.400 617.710 2840.460 ;
        RECT 1011.150 2840.260 1011.470 2840.320 ;
        RECT 1059.450 2840.260 1059.770 2840.320 ;
        RECT 1107.290 2840.260 1107.610 2840.320 ;
        RECT 1152.370 2840.260 1152.690 2840.320 ;
        RECT 1011.150 2840.120 1152.690 2840.260 ;
        RECT 1011.150 2840.060 1011.470 2840.120 ;
        RECT 1059.450 2840.060 1059.770 2840.120 ;
        RECT 1107.290 2840.060 1107.610 2840.120 ;
        RECT 1152.370 2840.060 1152.690 2840.120 ;
        RECT 474.330 2839.100 590.020 2839.240 ;
        RECT 1100.390 2839.240 1100.710 2839.300 ;
        RECT 1146.850 2839.240 1147.170 2839.300 ;
        RECT 1193.770 2839.240 1194.090 2839.300 ;
        RECT 1100.390 2839.100 1194.090 2839.240 ;
        RECT 474.330 2839.040 474.650 2839.100 ;
        RECT 520.330 2839.040 520.650 2839.100 ;
        RECT 568.170 2839.040 568.490 2839.100 ;
        RECT 1100.390 2839.040 1100.710 2839.100 ;
        RECT 1146.850 2839.040 1147.170 2839.100 ;
        RECT 1193.770 2839.040 1194.090 2839.100 ;
        RECT 606.350 2836.520 606.670 2836.580 ;
        RECT 1011.150 2836.520 1011.470 2836.580 ;
        RECT 606.350 2836.380 1011.470 2836.520 ;
        RECT 606.350 2836.320 606.670 2836.380 ;
        RECT 1011.150 2836.320 1011.470 2836.380 ;
        RECT 1052.090 2836.520 1052.410 2836.580 ;
        RECT 1100.390 2836.520 1100.710 2836.580 ;
        RECT 1052.090 2836.380 1100.710 2836.520 ;
        RECT 1052.090 2836.320 1052.410 2836.380 ;
        RECT 1100.390 2836.320 1100.710 2836.380 ;
        RECT 602.210 2620.280 602.530 2620.340 ;
        RECT 606.350 2620.280 606.670 2620.340 ;
        RECT 602.210 2620.140 606.670 2620.280 ;
        RECT 602.210 2620.080 602.530 2620.140 ;
        RECT 606.350 2620.080 606.670 2620.140 ;
        RECT 1013.910 2619.600 1014.230 2619.660 ;
        RECT 1059.910 2619.600 1060.230 2619.660 ;
        RECT 1013.910 2619.460 1060.230 2619.600 ;
        RECT 1013.910 2619.400 1014.230 2619.460 ;
        RECT 1059.910 2619.400 1060.230 2619.460 ;
        RECT 668.910 2619.260 669.230 2619.320 ;
        RECT 1052.090 2619.260 1052.410 2619.320 ;
        RECT 668.910 2619.120 1052.410 2619.260 ;
        RECT 668.910 2619.060 669.230 2619.120 ;
        RECT 1052.090 2619.060 1052.410 2619.120 ;
        RECT 1200.210 2619.260 1200.530 2619.320 ;
        RECT 1217.245 2619.260 1217.535 2619.305 ;
        RECT 1200.210 2619.120 1217.535 2619.260 ;
        RECT 1200.210 2619.060 1200.530 2619.120 ;
        RECT 1217.245 2619.075 1217.535 2619.120 ;
        RECT 1218.625 2618.580 1218.915 2618.625 ;
        RECT 1355.230 2618.580 1355.550 2618.640 ;
        RECT 1218.625 2618.440 1355.550 2618.580 ;
        RECT 1218.625 2618.395 1218.915 2618.440 ;
        RECT 1355.230 2618.380 1355.550 2618.440 ;
        RECT 617.390 2618.240 617.710 2618.300 ;
        RECT 697.430 2618.240 697.750 2618.300 ;
        RECT 617.390 2618.100 697.750 2618.240 ;
        RECT 617.390 2618.040 617.710 2618.100 ;
        RECT 697.430 2618.040 697.750 2618.100 ;
      LAYER via ;
        RECT 474.360 2839.040 474.620 2839.300 ;
        RECT 520.360 2839.040 520.620 2839.300 ;
        RECT 568.200 2839.040 568.460 2839.300 ;
        RECT 617.420 2840.400 617.680 2840.660 ;
        RECT 1011.180 2840.060 1011.440 2840.320 ;
        RECT 1059.480 2840.060 1059.740 2840.320 ;
        RECT 1107.320 2840.060 1107.580 2840.320 ;
        RECT 1152.400 2840.060 1152.660 2840.320 ;
        RECT 1100.420 2839.040 1100.680 2839.300 ;
        RECT 1146.880 2839.040 1147.140 2839.300 ;
        RECT 1193.800 2839.040 1194.060 2839.300 ;
        RECT 606.380 2836.320 606.640 2836.580 ;
        RECT 1011.180 2836.320 1011.440 2836.580 ;
        RECT 1052.120 2836.320 1052.380 2836.580 ;
        RECT 1100.420 2836.320 1100.680 2836.580 ;
        RECT 602.240 2620.080 602.500 2620.340 ;
        RECT 606.380 2620.080 606.640 2620.340 ;
        RECT 1013.940 2619.400 1014.200 2619.660 ;
        RECT 1059.940 2619.400 1060.200 2619.660 ;
        RECT 668.940 2619.060 669.200 2619.320 ;
        RECT 1052.120 2619.060 1052.380 2619.320 ;
        RECT 1200.240 2619.060 1200.500 2619.320 ;
        RECT 1355.260 2618.380 1355.520 2618.640 ;
        RECT 617.420 2618.040 617.680 2618.300 ;
        RECT 697.460 2618.040 697.720 2618.300 ;
      LAYER met2 ;
        RECT 474.350 2850.715 474.630 2851.085 ;
        RECT 1013.930 2850.715 1014.210 2851.085 ;
        RECT 1193.790 2850.715 1194.070 2851.085 ;
        RECT 474.420 2839.330 474.560 2850.715 ;
        RECT 568.190 2848.675 568.470 2849.045 ;
        RECT 520.350 2842.555 520.630 2842.925 ;
        RECT 520.420 2839.330 520.560 2842.555 ;
        RECT 568.260 2839.330 568.400 2848.675 ;
        RECT 1011.170 2842.555 1011.450 2842.925 ;
        RECT 617.420 2840.370 617.680 2840.690 ;
        RECT 474.360 2839.010 474.620 2839.330 ;
        RECT 520.360 2839.010 520.620 2839.330 ;
        RECT 568.200 2839.010 568.460 2839.330 ;
        RECT 606.380 2836.290 606.640 2836.610 ;
        RECT 606.440 2620.370 606.580 2836.290 ;
        RECT 617.480 2836.125 617.620 2840.370 ;
        RECT 1011.240 2840.350 1011.380 2842.555 ;
        RECT 1011.180 2840.030 1011.440 2840.350 ;
        RECT 1011.240 2836.610 1011.380 2840.030 ;
        RECT 1011.180 2836.290 1011.440 2836.610 ;
        RECT 617.410 2835.755 617.690 2836.125 ;
        RECT 602.240 2620.050 602.500 2620.370 ;
        RECT 606.380 2620.050 606.640 2620.370 ;
        RECT 602.300 2610.000 602.440 2620.050 ;
        RECT 617.480 2618.330 617.620 2835.755 ;
        RECT 1014.000 2619.690 1014.140 2850.715 ;
        RECT 1059.470 2842.555 1059.750 2842.925 ;
        RECT 1107.310 2842.555 1107.590 2842.925 ;
        RECT 1146.870 2842.555 1147.150 2842.925 ;
        RECT 1059.540 2840.350 1059.680 2842.555 ;
        RECT 1100.410 2841.875 1100.690 2842.245 ;
        RECT 1059.480 2840.030 1059.740 2840.350 ;
        RECT 1100.480 2839.330 1100.620 2841.875 ;
        RECT 1107.380 2840.350 1107.520 2842.555 ;
        RECT 1107.320 2840.030 1107.580 2840.350 ;
        RECT 1146.940 2839.330 1147.080 2842.555 ;
        RECT 1152.390 2840.515 1152.670 2840.885 ;
        RECT 1152.460 2840.350 1152.600 2840.515 ;
        RECT 1152.400 2840.030 1152.660 2840.350 ;
        RECT 1193.860 2839.330 1194.000 2850.715 ;
        RECT 1200.230 2842.555 1200.510 2842.925 ;
        RECT 1100.420 2839.010 1100.680 2839.330 ;
        RECT 1146.880 2839.010 1147.140 2839.330 ;
        RECT 1193.800 2839.010 1194.060 2839.330 ;
        RECT 1100.480 2836.610 1100.620 2839.010 ;
        RECT 1052.120 2836.290 1052.380 2836.610 ;
        RECT 1100.420 2836.290 1100.680 2836.610 ;
        RECT 1052.180 2836.125 1052.320 2836.290 ;
        RECT 1052.110 2835.755 1052.390 2836.125 ;
        RECT 1013.940 2619.370 1014.200 2619.690 ;
        RECT 1052.180 2619.350 1052.320 2835.755 ;
        RECT 1059.940 2619.370 1060.200 2619.690 ;
        RECT 668.940 2619.030 669.200 2619.350 ;
        RECT 1052.120 2619.030 1052.380 2619.350 ;
        RECT 617.420 2618.010 617.680 2618.330 ;
        RECT 669.000 2610.000 669.140 2619.030 ;
        RECT 697.460 2618.010 697.720 2618.330 ;
        RECT 697.520 2610.000 697.660 2618.010 ;
        RECT 1060.000 2610.000 1060.140 2619.370 ;
        RECT 1200.300 2619.350 1200.440 2842.555 ;
        RECT 1200.240 2619.030 1200.500 2619.350 ;
        RECT 1355.260 2618.350 1355.520 2618.670 ;
        RECT 1355.320 2610.000 1355.460 2618.350 ;
        RECT 602.100 2609.500 602.440 2610.000 ;
        RECT 668.800 2609.500 669.140 2610.000 ;
        RECT 697.320 2609.500 697.660 2610.000 ;
        RECT 1059.800 2609.500 1060.140 2610.000 ;
        RECT 1355.120 2609.500 1355.460 2610.000 ;
        RECT 602.100 2606.000 602.380 2609.500 ;
        RECT 668.800 2606.000 669.080 2609.500 ;
        RECT 697.320 2606.000 697.600 2609.500 ;
        RECT 1059.800 2606.000 1060.080 2609.500 ;
        RECT 1355.120 2606.000 1355.400 2609.500 ;
      LAYER via2 ;
        RECT 474.350 2850.760 474.630 2851.040 ;
        RECT 1013.930 2850.760 1014.210 2851.040 ;
        RECT 1193.790 2850.760 1194.070 2851.040 ;
        RECT 568.190 2848.720 568.470 2849.000 ;
        RECT 520.350 2842.600 520.630 2842.880 ;
        RECT 1011.170 2842.600 1011.450 2842.880 ;
        RECT 617.410 2835.800 617.690 2836.080 ;
        RECT 1059.470 2842.600 1059.750 2842.880 ;
        RECT 1107.310 2842.600 1107.590 2842.880 ;
        RECT 1146.870 2842.600 1147.150 2842.880 ;
        RECT 1100.410 2841.920 1100.690 2842.200 ;
        RECT 1152.390 2840.560 1152.670 2840.840 ;
        RECT 1200.230 2842.600 1200.510 2842.880 ;
        RECT 1052.110 2835.800 1052.390 2836.080 ;
      LAYER met3 ;
        RECT 474.325 2851.060 474.655 2851.065 ;
        RECT 474.070 2851.050 474.655 2851.060 ;
        RECT 1013.905 2851.050 1014.235 2851.065 ;
        RECT 1193.765 2851.060 1194.095 2851.065 ;
        RECT 1015.030 2851.050 1015.410 2851.060 ;
        RECT 474.070 2850.750 474.880 2851.050 ;
        RECT 1013.905 2850.750 1015.410 2851.050 ;
        RECT 474.070 2850.740 474.655 2850.750 ;
        RECT 474.325 2850.735 474.655 2850.740 ;
        RECT 1013.905 2850.735 1014.235 2850.750 ;
        RECT 1015.030 2850.740 1015.410 2850.750 ;
        RECT 1193.510 2851.050 1194.095 2851.060 ;
        RECT 1193.510 2850.750 1194.320 2851.050 ;
        RECT 1193.510 2850.740 1194.095 2850.750 ;
        RECT 1193.765 2850.735 1194.095 2850.740 ;
        RECT 568.165 2849.020 568.495 2849.025 ;
        RECT 568.165 2849.010 568.670 2849.020 ;
        RECT 568.165 2848.710 568.950 2849.010 ;
        RECT 568.165 2848.700 568.670 2848.710 ;
        RECT 568.165 2848.695 568.495 2848.700 ;
        RECT 520.325 2842.900 520.655 2842.905 ;
        RECT 520.070 2842.890 520.655 2842.900 ;
        RECT 519.870 2842.590 520.655 2842.890 ;
        RECT 520.070 2842.580 520.655 2842.590 ;
        RECT 520.325 2842.575 520.655 2842.580 ;
        RECT 1011.145 2842.900 1011.475 2842.905 ;
        RECT 1059.445 2842.900 1059.775 2842.905 ;
        RECT 1107.285 2842.900 1107.615 2842.905 ;
        RECT 1146.845 2842.900 1147.175 2842.905 ;
        RECT 1011.145 2842.890 1011.730 2842.900 ;
        RECT 1059.190 2842.890 1059.775 2842.900 ;
        RECT 1107.030 2842.890 1107.615 2842.900 ;
        RECT 1146.590 2842.890 1147.175 2842.900 ;
        RECT 1011.145 2842.590 1011.930 2842.890 ;
        RECT 1058.990 2842.590 1059.775 2842.890 ;
        RECT 1106.830 2842.590 1107.615 2842.890 ;
        RECT 1146.390 2842.590 1147.175 2842.890 ;
        RECT 1011.145 2842.580 1011.730 2842.590 ;
        RECT 1059.190 2842.580 1059.775 2842.590 ;
        RECT 1107.030 2842.580 1107.615 2842.590 ;
        RECT 1146.590 2842.580 1147.175 2842.590 ;
        RECT 1198.110 2842.890 1198.490 2842.900 ;
        RECT 1200.205 2842.890 1200.535 2842.905 ;
        RECT 1198.110 2842.590 1200.535 2842.890 ;
        RECT 1198.110 2842.580 1198.490 2842.590 ;
        RECT 1011.145 2842.575 1011.475 2842.580 ;
        RECT 1059.445 2842.575 1059.775 2842.580 ;
        RECT 1107.285 2842.575 1107.615 2842.580 ;
        RECT 1146.845 2842.575 1147.175 2842.580 ;
        RECT 1200.205 2842.575 1200.535 2842.590 ;
        RECT 1100.385 2842.220 1100.715 2842.225 ;
        RECT 1100.385 2842.210 1100.970 2842.220 ;
        RECT 1100.385 2841.910 1101.170 2842.210 ;
        RECT 1100.385 2841.900 1100.970 2841.910 ;
        RECT 1100.385 2841.895 1100.715 2841.900 ;
        RECT 1152.365 2840.850 1152.695 2840.865 ;
        RECT 1153.030 2840.850 1153.410 2840.860 ;
        RECT 1152.365 2840.550 1153.410 2840.850 ;
        RECT 1152.365 2840.535 1152.695 2840.550 ;
        RECT 1153.030 2840.540 1153.410 2840.550 ;
        RECT 614.830 2836.090 615.210 2836.100 ;
        RECT 617.385 2836.090 617.715 2836.105 ;
        RECT 614.830 2835.790 617.715 2836.090 ;
        RECT 614.830 2835.780 615.210 2835.790 ;
        RECT 617.385 2835.775 617.715 2835.790 ;
        RECT 1052.085 2836.090 1052.415 2836.105 ;
        RECT 1052.750 2836.090 1053.130 2836.100 ;
        RECT 1052.085 2835.790 1053.130 2836.090 ;
        RECT 1052.085 2835.775 1052.415 2835.790 ;
        RECT 1052.750 2835.780 1053.130 2835.790 ;
      LAYER via3 ;
        RECT 474.100 2850.740 474.420 2851.060 ;
        RECT 1015.060 2850.740 1015.380 2851.060 ;
        RECT 1193.540 2850.740 1193.860 2851.060 ;
        RECT 568.320 2848.700 568.640 2849.020 ;
        RECT 520.100 2842.580 520.420 2842.900 ;
        RECT 1011.380 2842.580 1011.700 2842.900 ;
        RECT 1059.220 2842.580 1059.540 2842.900 ;
        RECT 1107.060 2842.580 1107.380 2842.900 ;
        RECT 1146.620 2842.580 1146.940 2842.900 ;
        RECT 1198.140 2842.580 1198.460 2842.900 ;
        RECT 1100.620 2841.900 1100.940 2842.220 ;
        RECT 1153.060 2840.540 1153.380 2840.860 ;
        RECT 614.860 2835.780 615.180 2836.100 ;
        RECT 1052.780 2835.780 1053.100 2836.100 ;
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 292.020 -18.720 295.020 3538.400 ;
        RECT 472.020 3306.235 475.020 3538.400 ;
        RECT 652.020 3306.235 655.020 3538.400 ;
        RECT 474.095 2851.050 474.425 2851.065 ;
        RECT 474.890 2851.050 475.190 2854.600 ;
        RECT 521.610 2852.750 521.910 2854.600 ;
        RECT 474.095 2850.750 475.190 2851.050 ;
        RECT 474.095 2850.735 474.425 2850.750 ;
        RECT 474.890 2850.000 475.190 2850.750 ;
        RECT 520.110 2852.450 521.910 2852.750 ;
        RECT 472.020 -18.720 475.020 2850.000 ;
        RECT 520.110 2842.905 520.410 2852.450 ;
        RECT 521.610 2850.000 521.910 2852.450 ;
        RECT 568.330 2849.025 568.630 2854.600 ;
        RECT 615.050 2851.050 615.350 2854.600 ;
        RECT 614.870 2850.000 615.350 2851.050 ;
        RECT 568.315 2848.695 568.645 2849.025 ;
        RECT 520.095 2842.575 520.425 2842.905 ;
        RECT 614.870 2836.105 615.170 2850.000 ;
        RECT 614.855 2835.775 615.185 2836.105 ;
        RECT 652.020 -18.720 655.020 2850.000 ;
        RECT 832.020 -18.720 835.020 3538.400 ;
        RECT 1012.020 3306.235 1015.020 3538.400 ;
        RECT 1192.020 3306.235 1195.020 3538.400 ;
        RECT 1193.785 3301.635 1194.085 3306.235 ;
        RECT 1013.210 2851.050 1013.510 2854.600 ;
        RECT 1011.390 2850.750 1013.510 2851.050 ;
        RECT 1011.390 2842.905 1011.690 2850.750 ;
        RECT 1013.210 2850.000 1013.510 2850.750 ;
        RECT 1013.830 2851.050 1014.130 2854.600 ;
        RECT 1015.055 2851.050 1015.385 2851.065 ;
        RECT 1054.090 2851.050 1054.390 2854.600 ;
        RECT 1059.930 2851.050 1060.230 2854.600 ;
        RECT 1100.810 2851.050 1101.110 2854.600 ;
        RECT 1013.830 2850.750 1015.385 2851.050 ;
        RECT 1013.830 2850.000 1014.130 2850.750 ;
        RECT 1015.055 2850.735 1015.385 2850.750 ;
        RECT 1052.790 2850.750 1054.390 2851.050 ;
        RECT 1011.375 2842.575 1011.705 2842.905 ;
        RECT 1012.020 -18.720 1015.020 2850.000 ;
        RECT 1052.790 2836.105 1053.090 2850.750 ;
        RECT 1054.090 2850.000 1054.390 2850.750 ;
        RECT 1059.230 2850.750 1060.230 2851.050 ;
        RECT 1059.230 2842.905 1059.530 2850.750 ;
        RECT 1059.930 2850.000 1060.230 2850.750 ;
        RECT 1100.630 2850.000 1101.110 2851.050 ;
        RECT 1059.215 2842.575 1059.545 2842.905 ;
        RECT 1100.630 2842.225 1100.930 2850.000 ;
        RECT 1106.650 2847.650 1106.950 2854.600 ;
        RECT 1147.530 2851.050 1147.830 2854.600 ;
        RECT 1153.370 2851.050 1153.670 2854.600 ;
        RECT 1146.630 2850.750 1147.830 2851.050 ;
        RECT 1106.650 2847.350 1107.370 2847.650 ;
        RECT 1107.070 2842.905 1107.370 2847.350 ;
        RECT 1146.630 2842.905 1146.930 2850.750 ;
        RECT 1147.530 2850.000 1147.830 2850.750 ;
        RECT 1153.070 2850.000 1153.670 2851.050 ;
        RECT 1193.535 2851.050 1193.865 2851.065 ;
        RECT 1194.250 2851.050 1194.550 2854.600 ;
        RECT 1193.535 2850.750 1194.550 2851.050 ;
        RECT 1193.535 2850.735 1193.865 2850.750 ;
        RECT 1194.250 2850.000 1194.550 2850.750 ;
        RECT 1194.870 2851.050 1195.170 2854.600 ;
        RECT 1194.870 2850.750 1198.450 2851.050 ;
        RECT 1194.870 2850.000 1195.170 2850.750 ;
        RECT 1107.055 2842.575 1107.385 2842.905 ;
        RECT 1146.615 2842.575 1146.945 2842.905 ;
        RECT 1100.615 2841.895 1100.945 2842.225 ;
        RECT 1153.070 2840.865 1153.370 2850.000 ;
        RECT 1153.055 2840.535 1153.385 2840.865 ;
        RECT 1052.775 2835.775 1053.105 2836.105 ;
        RECT 1192.020 -18.720 1195.020 2850.000 ;
        RECT 1198.150 2842.905 1198.450 2850.750 ;
        RECT 1198.135 2842.575 1198.465 2842.905 ;
        RECT 1372.020 -18.720 1375.020 3538.400 ;
        RECT 1552.020 -18.720 1555.020 3538.400 ;
        RECT 1732.020 2586.480 1735.020 3538.400 ;
        RECT 1912.020 2586.480 1915.020 3538.400 ;
        RECT 1732.020 1986.480 1735.020 2200.000 ;
        RECT 1912.020 1986.480 1915.020 2200.000 ;
        RECT 1732.020 -18.720 1735.020 1600.000 ;
        RECT 1912.020 -18.720 1915.020 1600.000 ;
        RECT 2092.020 -18.720 2095.020 3538.400 ;
        RECT 2272.020 -18.720 2275.020 3538.400 ;
        RECT 2452.020 -18.720 2455.020 3538.400 ;
        RECT 2632.020 -18.720 2635.020 3538.400 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 584.805 2837.045 584.975 2840.955 ;
        RECT 737.525 2616.045 737.695 2616.895 ;
      LAYER mcon ;
        RECT 584.805 2840.785 584.975 2840.955 ;
        RECT 737.525 2616.725 737.695 2616.895 ;
      LAYER met1 ;
        RECT 489.510 2840.940 489.830 2841.000 ;
        RECT 533.210 2840.940 533.530 2841.000 ;
        RECT 579.210 2840.940 579.530 2841.000 ;
        RECT 584.745 2840.940 585.035 2840.985 ;
        RECT 489.510 2840.800 585.035 2840.940 ;
        RECT 489.510 2840.740 489.830 2840.800 ;
        RECT 533.210 2840.740 533.530 2840.800 ;
        RECT 579.210 2840.740 579.530 2840.800 ;
        RECT 584.745 2840.755 585.035 2840.800 ;
        RECT 596.230 2839.920 596.550 2839.980 ;
        RECT 714.450 2839.920 714.770 2839.980 ;
        RECT 596.230 2839.780 714.770 2839.920 ;
        RECT 596.230 2839.720 596.550 2839.780 ;
        RECT 714.450 2839.720 714.770 2839.780 ;
        RECT 584.745 2837.200 585.035 2837.245 ;
        RECT 624.290 2837.200 624.610 2837.260 ;
        RECT 584.745 2837.060 624.610 2837.200 ;
        RECT 584.745 2837.015 585.035 2837.060 ;
        RECT 624.290 2837.000 624.610 2837.060 ;
        RECT 624.290 2617.220 624.610 2617.280 ;
        RECT 716.750 2617.220 717.070 2617.280 ;
        RECT 624.290 2617.080 717.070 2617.220 ;
        RECT 624.290 2617.020 624.610 2617.080 ;
        RECT 716.750 2617.020 717.070 2617.080 ;
        RECT 737.465 2616.880 737.755 2616.925 ;
        RECT 945.370 2616.880 945.690 2616.940 ;
        RECT 737.465 2616.740 945.690 2616.880 ;
        RECT 737.465 2616.695 737.755 2616.740 ;
        RECT 945.370 2616.680 945.690 2616.740 ;
        RECT 714.450 2616.200 714.770 2616.260 ;
        RECT 737.465 2616.200 737.755 2616.245 ;
        RECT 714.450 2616.060 737.755 2616.200 ;
        RECT 714.450 2616.000 714.770 2616.060 ;
        RECT 737.465 2616.015 737.755 2616.060 ;
      LAYER via ;
        RECT 489.540 2840.740 489.800 2841.000 ;
        RECT 533.240 2840.740 533.500 2841.000 ;
        RECT 579.240 2840.740 579.500 2841.000 ;
        RECT 596.260 2839.720 596.520 2839.980 ;
        RECT 714.480 2839.720 714.740 2839.980 ;
        RECT 624.320 2837.000 624.580 2837.260 ;
        RECT 624.320 2617.020 624.580 2617.280 ;
        RECT 716.780 2617.020 717.040 2617.280 ;
        RECT 945.400 2616.680 945.660 2616.940 ;
        RECT 714.480 2616.000 714.740 2616.260 ;
      LAYER met2 ;
        RECT 596.250 2844.595 596.530 2844.965 ;
        RECT 533.230 2842.555 533.510 2842.925 ;
        RECT 579.230 2842.555 579.510 2842.925 ;
        RECT 489.530 2841.195 489.810 2841.565 ;
        RECT 489.600 2841.030 489.740 2841.195 ;
        RECT 533.300 2841.030 533.440 2842.555 ;
        RECT 579.300 2841.030 579.440 2842.555 ;
        RECT 489.540 2840.710 489.800 2841.030 ;
        RECT 533.240 2840.710 533.500 2841.030 ;
        RECT 579.240 2840.710 579.500 2841.030 ;
        RECT 596.320 2840.010 596.460 2844.595 ;
        RECT 596.260 2839.690 596.520 2840.010 ;
        RECT 714.480 2839.690 714.740 2840.010 ;
        RECT 624.310 2838.475 624.590 2838.845 ;
        RECT 624.380 2837.290 624.520 2838.475 ;
        RECT 624.320 2836.970 624.580 2837.290 ;
        RECT 624.380 2617.310 624.520 2836.970 ;
        RECT 624.320 2616.990 624.580 2617.310 ;
        RECT 714.540 2616.290 714.680 2839.690 ;
        RECT 716.780 2616.990 717.040 2617.310 ;
        RECT 714.480 2615.970 714.740 2616.290 ;
        RECT 716.840 2610.000 716.980 2616.990 ;
        RECT 945.400 2616.650 945.660 2616.970 ;
        RECT 945.460 2610.000 945.600 2616.650 ;
        RECT 716.640 2609.500 716.980 2610.000 ;
        RECT 945.260 2609.500 945.600 2610.000 ;
        RECT 716.640 2606.000 716.920 2609.500 ;
        RECT 945.260 2606.000 945.540 2609.500 ;
      LAYER via2 ;
        RECT 596.250 2844.640 596.530 2844.920 ;
        RECT 533.230 2842.600 533.510 2842.880 ;
        RECT 579.230 2842.600 579.510 2842.880 ;
        RECT 489.530 2841.240 489.810 2841.520 ;
        RECT 624.310 2838.520 624.590 2838.800 ;
      LAYER met3 ;
        RECT 583.550 2844.930 583.930 2844.940 ;
        RECT 596.225 2844.930 596.555 2844.945 ;
        RECT 583.550 2844.630 596.555 2844.930 ;
        RECT 583.550 2844.620 583.930 2844.630 ;
        RECT 596.225 2844.615 596.555 2844.630 ;
        RECT 533.205 2842.900 533.535 2842.905 ;
        RECT 579.205 2842.900 579.535 2842.905 ;
        RECT 532.950 2842.890 533.535 2842.900 ;
        RECT 578.950 2842.890 579.535 2842.900 ;
        RECT 532.750 2842.590 533.535 2842.890 ;
        RECT 578.750 2842.590 579.535 2842.890 ;
        RECT 532.950 2842.580 533.535 2842.590 ;
        RECT 578.950 2842.580 579.535 2842.590 ;
        RECT 533.205 2842.575 533.535 2842.580 ;
        RECT 579.205 2842.575 579.535 2842.580 ;
        RECT 486.950 2841.530 487.330 2841.540 ;
        RECT 489.505 2841.530 489.835 2841.545 ;
        RECT 486.950 2841.230 489.835 2841.530 ;
        RECT 486.950 2841.220 487.330 2841.230 ;
        RECT 489.505 2841.215 489.835 2841.230 ;
        RECT 624.285 2838.810 624.615 2838.825 ;
        RECT 624.950 2838.810 625.330 2838.820 ;
        RECT 624.285 2838.510 625.330 2838.810 ;
        RECT 624.285 2838.495 624.615 2838.510 ;
        RECT 624.950 2838.500 625.330 2838.510 ;
      LAYER via3 ;
        RECT 583.580 2844.620 583.900 2844.940 ;
        RECT 532.980 2842.580 533.300 2842.900 ;
        RECT 578.980 2842.580 579.300 2842.900 ;
        RECT 486.980 2841.220 487.300 2841.540 ;
        RECT 624.980 2838.500 625.300 2838.820 ;
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 400.020 3306.235 403.020 3547.800 ;
        RECT 580.020 3306.235 583.020 3547.800 ;
        RECT 760.020 3306.235 763.020 3547.800 ;
        RECT 581.385 3301.635 581.685 3306.235 ;
        RECT 400.020 -28.120 403.020 2850.000 ;
        RECT 486.570 2847.650 486.870 2854.600 ;
        RECT 533.290 2851.050 533.590 2854.600 ;
        RECT 580.010 2851.050 580.310 2854.600 ;
        RECT 532.990 2850.000 533.590 2851.050 ;
        RECT 578.990 2850.750 580.310 2851.050 ;
        RECT 486.570 2847.350 487.290 2847.650 ;
        RECT 486.990 2841.545 487.290 2847.350 ;
        RECT 532.990 2842.905 533.290 2850.000 ;
        RECT 578.990 2842.905 579.290 2850.750 ;
        RECT 580.010 2850.000 580.310 2850.750 ;
        RECT 580.630 2851.050 580.930 2854.600 ;
        RECT 626.730 2851.050 627.030 2854.600 ;
        RECT 580.630 2850.750 583.890 2851.050 ;
        RECT 580.630 2850.000 580.930 2850.750 ;
        RECT 532.975 2842.575 533.305 2842.905 ;
        RECT 578.975 2842.575 579.305 2842.905 ;
        RECT 486.975 2841.215 487.305 2841.545 ;
        RECT 580.020 -28.120 583.020 2850.000 ;
        RECT 583.590 2844.945 583.890 2850.750 ;
        RECT 624.990 2850.750 627.030 2851.050 ;
        RECT 583.575 2844.615 583.905 2844.945 ;
        RECT 624.990 2838.825 625.290 2850.750 ;
        RECT 626.730 2850.000 627.030 2850.750 ;
        RECT 624.975 2838.495 625.305 2838.825 ;
        RECT 760.020 -28.120 763.020 2850.000 ;
        RECT 940.020 -28.120 943.020 3547.800 ;
        RECT 1120.020 3306.235 1123.020 3547.800 ;
        RECT 1300.020 3306.235 1303.020 3547.800 ;
        RECT 1120.020 -28.120 1123.020 2850.000 ;
        RECT 1300.020 -28.120 1303.020 2850.000 ;
        RECT 1480.020 -28.120 1483.020 3547.800 ;
        RECT 1660.020 2586.480 1663.020 3547.800 ;
        RECT 1840.020 2586.480 1843.020 3547.800 ;
        RECT 2020.020 2586.480 2023.020 3547.800 ;
        RECT 1660.020 1986.480 1663.020 2200.000 ;
        RECT 1840.020 1986.480 1843.020 2200.000 ;
        RECT 2020.020 1986.480 2023.020 2200.000 ;
        RECT 1660.020 -28.120 1663.020 1600.000 ;
        RECT 1840.020 -28.120 1843.020 1600.000 ;
        RECT 2020.020 -28.120 2023.020 1600.000 ;
        RECT 2200.020 -28.120 2203.020 3547.800 ;
        RECT 2380.020 -28.120 2383.020 3547.800 ;
        RECT 2560.020 -28.120 2563.020 3547.800 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 491.810 2841.620 492.130 2841.680 ;
        RECT 538.730 2841.620 539.050 2841.680 ;
        RECT 585.650 2841.620 585.970 2841.680 ;
        RECT 491.810 2841.480 585.970 2841.620 ;
        RECT 491.810 2841.420 492.130 2841.480 ;
        RECT 538.730 2841.420 539.050 2841.480 ;
        RECT 585.650 2841.420 585.970 2841.480 ;
        RECT 633.030 2841.280 633.350 2841.340 ;
        RECT 724.570 2841.280 724.890 2841.340 ;
        RECT 622.540 2841.140 724.890 2841.280 ;
        RECT 585.650 2840.940 585.970 2841.000 ;
        RECT 622.540 2840.940 622.680 2841.140 ;
        RECT 633.030 2841.080 633.350 2841.140 ;
        RECT 724.570 2841.080 724.890 2841.140 ;
        RECT 1077.850 2841.280 1078.170 2841.340 ;
        RECT 1123.850 2841.280 1124.170 2841.340 ;
        RECT 1166.170 2841.280 1166.490 2841.340 ;
        RECT 1077.850 2841.140 1166.490 2841.280 ;
        RECT 1077.850 2841.080 1078.170 2841.140 ;
        RECT 1123.850 2841.080 1124.170 2841.140 ;
        RECT 1166.170 2841.080 1166.490 2841.140 ;
        RECT 585.650 2840.800 622.680 2840.940 ;
        RECT 585.650 2840.740 585.970 2840.800 ;
        RECT 1031.390 2836.180 1031.710 2836.240 ;
        RECT 1077.850 2836.180 1078.170 2836.240 ;
        RECT 1031.390 2836.040 1078.170 2836.180 ;
        RECT 1031.390 2835.980 1031.710 2836.040 ;
        RECT 1077.850 2835.980 1078.170 2836.040 ;
        RECT 630.730 2618.580 631.050 2618.640 ;
        RECT 1031.390 2618.580 1031.710 2618.640 ;
        RECT 630.730 2618.440 1031.710 2618.580 ;
        RECT 630.730 2618.380 631.050 2618.440 ;
        RECT 1031.390 2618.380 1031.710 2618.440 ;
        RECT 1034.610 2618.580 1034.930 2618.640 ;
        RECT 1088.430 2618.580 1088.750 2618.640 ;
        RECT 1034.610 2618.440 1088.750 2618.580 ;
        RECT 1034.610 2618.380 1034.930 2618.440 ;
        RECT 1088.430 2618.380 1088.750 2618.440 ;
      LAYER via ;
        RECT 491.840 2841.420 492.100 2841.680 ;
        RECT 538.760 2841.420 539.020 2841.680 ;
        RECT 585.680 2841.420 585.940 2841.680 ;
        RECT 585.680 2840.740 585.940 2841.000 ;
        RECT 633.060 2841.080 633.320 2841.340 ;
        RECT 724.600 2841.080 724.860 2841.340 ;
        RECT 1077.880 2841.080 1078.140 2841.340 ;
        RECT 1123.880 2841.080 1124.140 2841.340 ;
        RECT 1166.200 2841.080 1166.460 2841.340 ;
        RECT 1031.420 2835.980 1031.680 2836.240 ;
        RECT 1077.880 2835.980 1078.140 2836.240 ;
        RECT 630.760 2618.380 631.020 2618.640 ;
        RECT 1031.420 2618.380 1031.680 2618.640 ;
        RECT 1034.640 2618.380 1034.900 2618.640 ;
        RECT 1088.460 2618.380 1088.720 2618.640 ;
      LAYER met2 ;
        RECT 491.830 2850.715 492.110 2851.085 ;
        RECT 491.900 2841.710 492.040 2850.715 ;
        RECT 585.670 2847.995 585.950 2848.365 ;
        RECT 538.750 2842.555 539.030 2842.925 ;
        RECT 538.820 2841.710 538.960 2842.555 ;
        RECT 585.740 2841.710 585.880 2847.995 ;
        RECT 633.050 2842.555 633.330 2842.925 ;
        RECT 1077.870 2842.555 1078.150 2842.925 ;
        RECT 491.840 2841.390 492.100 2841.710 ;
        RECT 538.760 2841.390 539.020 2841.710 ;
        RECT 585.680 2841.390 585.940 2841.710 ;
        RECT 585.740 2841.030 585.880 2841.390 ;
        RECT 633.120 2841.370 633.260 2842.555 ;
        RECT 1077.940 2841.370 1078.080 2842.555 ;
        RECT 633.060 2841.050 633.320 2841.370 ;
        RECT 724.600 2841.050 724.860 2841.370 ;
        RECT 1077.880 2841.050 1078.140 2841.370 ;
        RECT 1123.870 2841.195 1124.150 2841.565 ;
        RECT 1166.190 2841.195 1166.470 2841.565 ;
        RECT 1123.880 2841.050 1124.140 2841.195 ;
        RECT 1166.200 2841.050 1166.460 2841.195 ;
        RECT 585.680 2840.710 585.940 2841.030 ;
        RECT 630.760 2618.350 631.020 2618.670 ;
        RECT 630.820 2610.000 630.960 2618.350 ;
        RECT 630.620 2609.500 630.960 2610.000 ;
        RECT 724.660 2609.570 724.800 2841.050 ;
        RECT 1031.480 2836.270 1031.620 2836.425 ;
        RECT 1077.940 2836.270 1078.080 2841.050 ;
        RECT 1031.420 2836.125 1031.680 2836.270 ;
        RECT 1031.410 2835.755 1031.690 2836.125 ;
        RECT 1034.630 2835.755 1034.910 2836.125 ;
        RECT 1077.880 2835.950 1078.140 2836.270 ;
        RECT 1031.480 2618.670 1031.620 2835.755 ;
        RECT 1034.700 2618.670 1034.840 2835.755 ;
        RECT 1031.420 2618.350 1031.680 2618.670 ;
        RECT 1034.640 2618.350 1034.900 2618.670 ;
        RECT 1088.460 2618.350 1088.720 2618.670 ;
        RECT 1088.520 2610.000 1088.660 2618.350 ;
        RECT 725.840 2609.570 726.120 2610.000 ;
        RECT 630.620 2606.000 630.900 2609.500 ;
        RECT 724.660 2609.430 726.120 2609.570 ;
        RECT 725.840 2606.000 726.120 2609.430 ;
        RECT 1088.320 2609.500 1088.660 2610.000 ;
        RECT 1088.320 2606.000 1088.600 2609.500 ;
      LAYER via2 ;
        RECT 491.830 2850.760 492.110 2851.040 ;
        RECT 585.670 2848.040 585.950 2848.320 ;
        RECT 538.750 2842.600 539.030 2842.880 ;
        RECT 633.050 2842.600 633.330 2842.880 ;
        RECT 1077.870 2842.600 1078.150 2842.880 ;
        RECT 1123.870 2841.240 1124.150 2841.520 ;
        RECT 1166.190 2841.240 1166.470 2841.520 ;
        RECT 1031.410 2835.800 1031.690 2836.080 ;
        RECT 1034.630 2835.800 1034.910 2836.080 ;
      LAYER met3 ;
        RECT 491.805 2851.060 492.135 2851.065 ;
        RECT 491.550 2851.050 492.135 2851.060 ;
        RECT 491.550 2850.750 492.360 2851.050 ;
        RECT 491.550 2850.740 492.135 2850.750 ;
        RECT 491.805 2850.735 492.135 2850.740 ;
        RECT 585.645 2848.340 585.975 2848.345 ;
        RECT 585.645 2848.330 586.190 2848.340 ;
        RECT 585.380 2848.030 586.190 2848.330 ;
        RECT 585.645 2848.020 586.190 2848.030 ;
        RECT 585.645 2848.015 585.975 2848.020 ;
        RECT 538.725 2842.900 539.055 2842.905 ;
        RECT 538.470 2842.890 539.055 2842.900 ;
        RECT 632.310 2842.890 632.690 2842.900 ;
        RECT 633.025 2842.890 633.355 2842.905 ;
        RECT 1077.845 2842.900 1078.175 2842.905 ;
        RECT 1077.590 2842.890 1078.175 2842.900 ;
        RECT 538.470 2842.590 539.280 2842.890 ;
        RECT 632.310 2842.590 633.355 2842.890 ;
        RECT 1077.390 2842.590 1078.175 2842.890 ;
        RECT 538.470 2842.580 539.055 2842.590 ;
        RECT 632.310 2842.580 632.690 2842.590 ;
        RECT 538.725 2842.575 539.055 2842.580 ;
        RECT 633.025 2842.575 633.355 2842.590 ;
        RECT 1077.590 2842.580 1078.175 2842.590 ;
        RECT 1077.845 2842.575 1078.175 2842.580 ;
        RECT 1123.845 2841.540 1124.175 2841.545 ;
        RECT 1123.590 2841.530 1124.175 2841.540 ;
        RECT 1166.165 2841.530 1166.495 2841.545 ;
        RECT 1167.750 2841.530 1168.130 2841.540 ;
        RECT 1123.590 2841.230 1124.400 2841.530 ;
        RECT 1166.165 2841.230 1168.130 2841.530 ;
        RECT 1123.590 2841.220 1124.175 2841.230 ;
        RECT 1123.845 2841.215 1124.175 2841.220 ;
        RECT 1166.165 2841.215 1166.495 2841.230 ;
        RECT 1167.750 2841.220 1168.130 2841.230 ;
        RECT 1028.830 2836.090 1029.210 2836.100 ;
        RECT 1031.385 2836.090 1031.715 2836.105 ;
        RECT 1034.605 2836.100 1034.935 2836.105 ;
        RECT 1028.830 2835.790 1031.715 2836.090 ;
        RECT 1028.830 2835.780 1029.210 2835.790 ;
        RECT 1031.385 2835.775 1031.715 2835.790 ;
        RECT 1034.350 2836.090 1034.935 2836.100 ;
        RECT 1034.350 2835.790 1035.160 2836.090 ;
        RECT 1034.350 2835.780 1034.935 2835.790 ;
        RECT 1034.605 2835.775 1034.935 2835.780 ;
      LAYER via3 ;
        RECT 491.580 2850.740 491.900 2851.060 ;
        RECT 585.840 2848.020 586.160 2848.340 ;
        RECT 538.500 2842.580 538.820 2842.900 ;
        RECT 632.340 2842.580 632.660 2842.900 ;
        RECT 1077.620 2842.580 1077.940 2842.900 ;
        RECT 1123.620 2841.220 1123.940 2841.540 ;
        RECT 1167.780 2841.220 1168.100 2841.540 ;
        RECT 1028.860 2835.780 1029.180 2836.100 ;
        RECT 1034.380 2835.780 1034.700 2836.100 ;
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 310.020 -28.120 313.020 3547.800 ;
        RECT 490.020 3306.235 493.020 3547.800 ;
        RECT 670.020 3306.235 673.020 3547.800 ;
        RECT 491.575 2851.050 491.905 2851.065 ;
        RECT 492.410 2851.050 492.710 2854.600 ;
        RECT 539.130 2851.050 539.430 2854.600 ;
        RECT 491.575 2850.750 492.710 2851.050 ;
        RECT 491.575 2850.735 491.905 2850.750 ;
        RECT 492.410 2850.000 492.710 2850.750 ;
        RECT 538.510 2850.750 539.430 2851.050 ;
        RECT 490.020 -28.120 493.020 2850.000 ;
        RECT 538.510 2842.905 538.810 2850.750 ;
        RECT 539.130 2850.000 539.430 2850.750 ;
        RECT 585.850 2848.345 586.150 2854.600 ;
        RECT 632.570 2851.050 632.870 2854.600 ;
        RECT 632.350 2850.000 632.870 2851.050 ;
        RECT 585.835 2848.015 586.165 2848.345 ;
        RECT 632.350 2842.905 632.650 2850.000 ;
        RECT 538.495 2842.575 538.825 2842.905 ;
        RECT 632.335 2842.575 632.665 2842.905 ;
        RECT 670.020 -28.120 673.020 2850.000 ;
        RECT 850.020 -28.120 853.020 3547.800 ;
        RECT 1030.020 3306.235 1033.020 3547.800 ;
        RECT 1210.020 3306.235 1213.020 3547.800 ;
        RECT 1212.505 3301.635 1212.805 3306.235 ;
        RECT 1030.730 2851.050 1031.030 2854.600 ;
        RECT 1028.870 2850.750 1031.030 2851.050 ;
        RECT 1028.870 2836.105 1029.170 2850.750 ;
        RECT 1030.730 2850.000 1031.030 2850.750 ;
        RECT 1031.350 2851.050 1031.650 2854.600 ;
        RECT 1031.350 2850.750 1034.690 2851.050 ;
        RECT 1031.350 2850.000 1031.650 2850.750 ;
        RECT 1028.855 2835.775 1029.185 2836.105 ;
        RECT 1030.020 -28.120 1033.020 2850.000 ;
        RECT 1034.390 2836.105 1034.690 2850.750 ;
        RECT 1077.450 2847.650 1077.750 2854.600 ;
        RECT 1124.170 2847.650 1124.470 2854.600 ;
        RECT 1170.890 2851.050 1171.190 2854.600 ;
        RECT 1077.450 2847.350 1077.930 2847.650 ;
        RECT 1077.630 2842.905 1077.930 2847.350 ;
        RECT 1123.630 2847.350 1124.470 2847.650 ;
        RECT 1167.790 2850.750 1171.190 2851.050 ;
        RECT 1077.615 2842.575 1077.945 2842.905 ;
        RECT 1123.630 2841.545 1123.930 2847.350 ;
        RECT 1167.790 2841.545 1168.090 2850.750 ;
        RECT 1170.890 2850.000 1171.190 2850.750 ;
        RECT 1123.615 2841.215 1123.945 2841.545 ;
        RECT 1167.775 2841.215 1168.105 2841.545 ;
        RECT 1034.375 2835.775 1034.705 2836.105 ;
        RECT 1210.020 -28.120 1213.020 2850.000 ;
        RECT 1390.020 -28.120 1393.020 3547.800 ;
        RECT 1570.020 -28.120 1573.020 3547.800 ;
        RECT 1750.020 2586.480 1753.020 3547.800 ;
        RECT 1930.020 2586.480 1933.020 3547.800 ;
        RECT 1750.020 1986.480 1753.020 2200.000 ;
        RECT 1930.020 1986.480 1933.020 2200.000 ;
        RECT 1750.020 -28.120 1753.020 1600.000 ;
        RECT 1930.020 -28.120 1933.020 1600.000 ;
        RECT 2110.020 -28.120 2113.020 3547.800 ;
        RECT 2290.020 -28.120 2293.020 3547.800 ;
        RECT 2470.020 -28.120 2473.020 3547.800 ;
        RECT 2650.020 -28.120 2653.020 3547.800 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 795.945 2621.485 797.035 2621.655 ;
      LAYER mcon ;
        RECT 796.865 2621.485 797.035 2621.655 ;
      LAYER met1 ;
        RECT 662.010 2842.640 662.330 2842.700 ;
        RECT 1047.950 2842.640 1048.270 2842.700 ;
        RECT 662.010 2842.500 1048.270 2842.640 ;
        RECT 662.010 2842.440 662.330 2842.500 ;
        RECT 1047.950 2842.440 1048.270 2842.500 ;
        RECT 1047.950 2840.940 1048.270 2841.000 ;
        RECT 1094.870 2840.940 1095.190 2841.000 ;
        RECT 1141.790 2840.940 1142.110 2841.000 ;
        RECT 1186.870 2840.940 1187.190 2841.000 ;
        RECT 1047.950 2840.800 1187.190 2840.940 ;
        RECT 1047.950 2840.740 1048.270 2840.800 ;
        RECT 1094.870 2840.740 1095.190 2840.800 ;
        RECT 1141.790 2840.740 1142.110 2840.800 ;
        RECT 1186.870 2840.740 1187.190 2840.800 ;
        RECT 468.810 2840.600 469.130 2840.660 ;
        RECT 508.830 2840.600 509.150 2840.660 ;
        RECT 553.450 2840.600 553.770 2840.660 ;
        RECT 468.810 2840.460 553.770 2840.600 ;
        RECT 468.810 2840.400 469.130 2840.460 ;
        RECT 508.830 2840.400 509.150 2840.460 ;
        RECT 553.450 2840.400 553.770 2840.460 ;
        RECT 514.810 2838.900 515.130 2838.960 ;
        RECT 783.450 2838.900 783.770 2838.960 ;
        RECT 514.810 2838.760 783.770 2838.900 ;
        RECT 514.810 2838.700 515.130 2838.760 ;
        RECT 783.450 2838.700 783.770 2838.760 ;
        RECT 553.450 2836.180 553.770 2836.240 ;
        RECT 603.590 2836.180 603.910 2836.240 ;
        RECT 553.450 2836.040 603.910 2836.180 ;
        RECT 553.450 2835.980 553.770 2836.040 ;
        RECT 603.590 2835.980 603.910 2836.040 ;
        RECT 783.450 2621.640 783.770 2621.700 ;
        RECT 795.885 2621.640 796.175 2621.685 ;
        RECT 783.450 2621.500 796.175 2621.640 ;
        RECT 783.450 2621.440 783.770 2621.500 ;
        RECT 795.885 2621.455 796.175 2621.500 ;
        RECT 796.805 2621.640 797.095 2621.685 ;
        RECT 830.830 2621.640 831.150 2621.700 ;
        RECT 796.805 2621.500 831.150 2621.640 ;
        RECT 796.805 2621.455 797.095 2621.500 ;
        RECT 830.830 2621.440 831.150 2621.500 ;
        RECT 1055.310 2621.640 1055.630 2621.700 ;
        RECT 1116.950 2621.640 1117.270 2621.700 ;
        RECT 1055.310 2621.500 1117.270 2621.640 ;
        RECT 1055.310 2621.440 1055.630 2621.500 ;
        RECT 1116.950 2621.440 1117.270 2621.500 ;
        RECT 603.590 2616.540 603.910 2616.600 ;
        RECT 678.570 2616.540 678.890 2616.600 ;
        RECT 603.590 2616.400 678.890 2616.540 ;
        RECT 603.590 2616.340 603.910 2616.400 ;
        RECT 678.570 2616.340 678.890 2616.400 ;
      LAYER via ;
        RECT 662.040 2842.440 662.300 2842.700 ;
        RECT 1047.980 2842.440 1048.240 2842.700 ;
        RECT 1047.980 2840.740 1048.240 2841.000 ;
        RECT 1094.900 2840.740 1095.160 2841.000 ;
        RECT 1141.820 2840.740 1142.080 2841.000 ;
        RECT 1186.900 2840.740 1187.160 2841.000 ;
        RECT 468.840 2840.400 469.100 2840.660 ;
        RECT 508.860 2840.400 509.120 2840.660 ;
        RECT 553.480 2840.400 553.740 2840.660 ;
        RECT 514.840 2838.700 515.100 2838.960 ;
        RECT 783.480 2838.700 783.740 2838.960 ;
        RECT 553.480 2835.980 553.740 2836.240 ;
        RECT 603.620 2835.980 603.880 2836.240 ;
        RECT 783.480 2621.440 783.740 2621.700 ;
        RECT 830.860 2621.440 831.120 2621.700 ;
        RECT 1055.340 2621.440 1055.600 2621.700 ;
        RECT 1116.980 2621.440 1117.240 2621.700 ;
        RECT 603.620 2616.340 603.880 2616.600 ;
        RECT 678.600 2616.340 678.860 2616.600 ;
      LAYER met2 ;
        RECT 508.850 2850.715 509.130 2851.085 ;
        RECT 468.830 2841.195 469.110 2841.565 ;
        RECT 468.900 2840.690 469.040 2841.195 ;
        RECT 508.920 2840.690 509.060 2850.715 ;
        RECT 603.610 2848.675 603.890 2849.045 ;
        RECT 514.830 2842.555 515.110 2842.925 ;
        RECT 553.470 2842.555 553.750 2842.925 ;
        RECT 468.840 2840.370 469.100 2840.690 ;
        RECT 508.860 2840.370 509.120 2840.690 ;
        RECT 514.900 2838.990 515.040 2842.555 ;
        RECT 553.540 2840.690 553.680 2842.555 ;
        RECT 553.480 2840.370 553.740 2840.690 ;
        RECT 514.840 2838.670 515.100 2838.990 ;
        RECT 553.540 2836.270 553.680 2840.370 ;
        RECT 603.680 2836.270 603.820 2848.675 ;
        RECT 662.040 2842.410 662.300 2842.730 ;
        RECT 1047.970 2842.555 1048.250 2842.925 ;
        RECT 1094.890 2842.555 1095.170 2842.925 ;
        RECT 1141.810 2842.555 1142.090 2842.925 ;
        RECT 1047.980 2842.410 1048.240 2842.555 ;
        RECT 553.480 2835.950 553.740 2836.270 ;
        RECT 603.620 2835.950 603.880 2836.270 ;
        RECT 603.680 2616.630 603.820 2835.950 ;
        RECT 603.620 2616.310 603.880 2616.630 ;
        RECT 659.140 2609.570 659.420 2610.000 ;
        RECT 662.100 2609.570 662.240 2842.410 ;
        RECT 1048.040 2841.030 1048.180 2842.410 ;
        RECT 1094.960 2841.030 1095.100 2842.555 ;
        RECT 1141.880 2841.030 1142.020 2842.555 ;
        RECT 1186.890 2841.195 1187.170 2841.565 ;
        RECT 1186.960 2841.030 1187.100 2841.195 ;
        RECT 1047.980 2840.710 1048.240 2841.030 ;
        RECT 1094.900 2840.710 1095.160 2841.030 ;
        RECT 1141.820 2840.710 1142.080 2841.030 ;
        RECT 1186.900 2840.710 1187.160 2841.030 ;
        RECT 783.480 2838.670 783.740 2838.990 ;
        RECT 783.540 2621.730 783.680 2838.670 ;
        RECT 1055.330 2836.435 1055.610 2836.805 ;
        RECT 1055.400 2621.730 1055.540 2836.435 ;
        RECT 783.480 2621.410 783.740 2621.730 ;
        RECT 830.860 2621.410 831.120 2621.730 ;
        RECT 1055.340 2621.410 1055.600 2621.730 ;
        RECT 1116.980 2621.410 1117.240 2621.730 ;
        RECT 678.600 2616.310 678.860 2616.630 ;
        RECT 678.660 2610.000 678.800 2616.310 ;
        RECT 830.920 2610.000 831.060 2621.410 ;
        RECT 1117.040 2610.000 1117.180 2621.410 ;
        RECT 659.140 2609.430 662.240 2609.570 ;
        RECT 678.460 2609.500 678.800 2610.000 ;
        RECT 830.720 2609.500 831.060 2610.000 ;
        RECT 1116.840 2609.500 1117.180 2610.000 ;
        RECT 659.140 2606.000 659.420 2609.430 ;
        RECT 678.460 2606.000 678.740 2609.500 ;
        RECT 830.720 2606.000 831.000 2609.500 ;
        RECT 1116.840 2606.000 1117.120 2609.500 ;
      LAYER via2 ;
        RECT 508.850 2850.760 509.130 2851.040 ;
        RECT 468.830 2841.240 469.110 2841.520 ;
        RECT 603.610 2848.720 603.890 2849.000 ;
        RECT 514.830 2842.600 515.110 2842.880 ;
        RECT 553.470 2842.600 553.750 2842.880 ;
        RECT 1047.970 2842.600 1048.250 2842.880 ;
        RECT 1094.890 2842.600 1095.170 2842.880 ;
        RECT 1141.810 2842.600 1142.090 2842.880 ;
        RECT 1186.890 2841.240 1187.170 2841.520 ;
        RECT 1055.330 2836.480 1055.610 2836.760 ;
      LAYER met3 ;
        RECT 508.825 2851.060 509.155 2851.065 ;
        RECT 508.825 2851.050 509.410 2851.060 ;
        RECT 508.825 2850.750 509.610 2851.050 ;
        RECT 508.825 2850.740 509.410 2850.750 ;
        RECT 508.825 2850.735 509.155 2850.740 ;
        RECT 603.585 2849.020 603.915 2849.025 ;
        RECT 603.330 2849.010 603.915 2849.020 ;
        RECT 603.330 2848.710 604.140 2849.010 ;
        RECT 603.330 2848.700 603.915 2848.710 ;
        RECT 603.585 2848.695 603.915 2848.700 ;
        RECT 513.630 2842.890 514.010 2842.900 ;
        RECT 514.805 2842.890 515.135 2842.905 ;
        RECT 513.630 2842.590 515.135 2842.890 ;
        RECT 513.630 2842.580 514.010 2842.590 ;
        RECT 514.805 2842.575 515.135 2842.590 ;
        RECT 553.445 2842.890 553.775 2842.905 ;
        RECT 554.110 2842.890 554.490 2842.900 ;
        RECT 553.445 2842.590 554.490 2842.890 ;
        RECT 553.445 2842.575 553.775 2842.590 ;
        RECT 554.110 2842.580 554.490 2842.590 ;
        RECT 1047.230 2842.890 1047.610 2842.900 ;
        RECT 1047.945 2842.890 1048.275 2842.905 ;
        RECT 1047.230 2842.590 1048.275 2842.890 ;
        RECT 1047.230 2842.580 1047.610 2842.590 ;
        RECT 1047.945 2842.575 1048.275 2842.590 ;
        RECT 1094.150 2842.890 1094.530 2842.900 ;
        RECT 1094.865 2842.890 1095.195 2842.905 ;
        RECT 1094.150 2842.590 1095.195 2842.890 ;
        RECT 1094.150 2842.580 1094.530 2842.590 ;
        RECT 1094.865 2842.575 1095.195 2842.590 ;
        RECT 1141.785 2842.900 1142.115 2842.905 ;
        RECT 1141.785 2842.890 1142.370 2842.900 ;
        RECT 1141.785 2842.590 1142.570 2842.890 ;
        RECT 1141.785 2842.580 1142.370 2842.590 ;
        RECT 1141.785 2842.575 1142.115 2842.580 ;
        RECT 463.030 2841.530 463.410 2841.540 ;
        RECT 468.805 2841.530 469.135 2841.545 ;
        RECT 1186.865 2841.540 1187.195 2841.545 ;
        RECT 1186.865 2841.530 1187.450 2841.540 ;
        RECT 463.030 2841.230 469.135 2841.530 ;
        RECT 1186.640 2841.230 1187.450 2841.530 ;
        RECT 463.030 2841.220 463.410 2841.230 ;
        RECT 468.805 2841.215 469.135 2841.230 ;
        RECT 1186.865 2841.220 1187.450 2841.230 ;
        RECT 1186.865 2841.215 1187.195 2841.220 ;
        RECT 1051.830 2836.770 1052.210 2836.780 ;
        RECT 1055.305 2836.770 1055.635 2836.785 ;
        RECT 1051.830 2836.470 1055.635 2836.770 ;
        RECT 1051.830 2836.460 1052.210 2836.470 ;
        RECT 1055.305 2836.455 1055.635 2836.470 ;
      LAYER via3 ;
        RECT 509.060 2850.740 509.380 2851.060 ;
        RECT 603.360 2848.700 603.680 2849.020 ;
        RECT 513.660 2842.580 513.980 2842.900 ;
        RECT 554.140 2842.580 554.460 2842.900 ;
        RECT 1047.260 2842.580 1047.580 2842.900 ;
        RECT 1094.180 2842.580 1094.500 2842.900 ;
        RECT 1142.020 2842.580 1142.340 2842.900 ;
        RECT 463.060 2841.220 463.380 2841.540 ;
        RECT 1187.100 2841.220 1187.420 2841.540 ;
        RECT 1051.860 2836.460 1052.180 2836.780 ;
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 328.020 -37.520 331.020 3557.200 ;
        RECT 508.020 3306.235 511.020 3557.200 ;
        RECT 688.020 3306.235 691.020 3557.200 ;
        RECT 463.210 2851.050 463.510 2854.600 ;
        RECT 463.070 2850.000 463.510 2851.050 ;
        RECT 509.055 2851.050 509.385 2851.065 ;
        RECT 509.930 2851.050 510.230 2854.600 ;
        RECT 509.055 2850.750 510.230 2851.050 ;
        RECT 509.055 2850.735 509.385 2850.750 ;
        RECT 509.930 2850.000 510.230 2850.750 ;
        RECT 510.550 2851.050 510.850 2854.600 ;
        RECT 556.650 2851.050 556.950 2854.600 ;
        RECT 510.550 2850.750 513.970 2851.050 ;
        RECT 510.550 2850.000 510.850 2850.750 ;
        RECT 463.070 2841.545 463.370 2850.000 ;
        RECT 463.055 2841.215 463.385 2841.545 ;
        RECT 508.020 -37.520 511.020 2850.000 ;
        RECT 513.670 2842.905 513.970 2850.750 ;
        RECT 554.150 2850.750 556.950 2851.050 ;
        RECT 554.150 2842.905 554.450 2850.750 ;
        RECT 556.650 2850.000 556.950 2850.750 ;
        RECT 603.370 2849.025 603.670 2854.600 ;
        RECT 603.355 2848.695 603.685 2849.025 ;
        RECT 513.655 2842.575 513.985 2842.905 ;
        RECT 554.135 2842.575 554.465 2842.905 ;
        RECT 688.020 -37.520 691.020 2850.000 ;
        RECT 868.020 -37.520 871.020 3557.200 ;
        RECT 1048.020 3306.235 1051.020 3557.200 ;
        RECT 1228.020 3306.235 1231.020 3557.200 ;
        RECT 1050.265 3301.635 1050.565 3306.235 ;
        RECT 1048.250 2851.050 1048.550 2854.600 ;
        RECT 1047.270 2850.750 1048.550 2851.050 ;
        RECT 1047.270 2842.905 1047.570 2850.750 ;
        RECT 1048.250 2850.000 1048.550 2850.750 ;
        RECT 1048.870 2851.050 1049.170 2854.600 ;
        RECT 1094.970 2851.050 1095.270 2854.600 ;
        RECT 1048.870 2850.750 1052.170 2851.050 ;
        RECT 1048.870 2850.000 1049.170 2850.750 ;
        RECT 1047.255 2842.575 1047.585 2842.905 ;
        RECT 1048.020 -37.520 1051.020 2850.000 ;
        RECT 1051.870 2836.785 1052.170 2850.750 ;
        RECT 1094.190 2850.750 1095.270 2851.050 ;
        RECT 1094.190 2842.905 1094.490 2850.750 ;
        RECT 1094.970 2850.000 1095.270 2850.750 ;
        RECT 1141.690 2847.650 1141.990 2854.600 ;
        RECT 1188.410 2851.050 1188.710 2854.600 ;
        RECT 1187.110 2850.750 1188.710 2851.050 ;
        RECT 1141.690 2847.350 1142.330 2847.650 ;
        RECT 1142.030 2842.905 1142.330 2847.350 ;
        RECT 1094.175 2842.575 1094.505 2842.905 ;
        RECT 1142.015 2842.575 1142.345 2842.905 ;
        RECT 1187.110 2841.545 1187.410 2850.750 ;
        RECT 1188.410 2850.000 1188.710 2850.750 ;
        RECT 1187.095 2841.215 1187.425 2841.545 ;
        RECT 1051.855 2836.455 1052.185 2836.785 ;
        RECT 1228.020 -37.520 1231.020 2850.000 ;
        RECT 1408.020 -37.520 1411.020 3557.200 ;
        RECT 1588.020 -37.520 1591.020 3557.200 ;
        RECT 1768.020 2586.480 1771.020 3557.200 ;
        RECT 1948.020 2586.480 1951.020 3557.200 ;
        RECT 1768.020 1986.480 1771.020 2200.000 ;
        RECT 1948.020 1986.480 1951.020 2200.000 ;
        RECT 1768.020 -37.520 1771.020 1600.000 ;
        RECT 1948.020 -37.520 1951.020 1600.000 ;
        RECT 2128.020 -37.520 2131.020 3557.200 ;
        RECT 2308.020 -37.520 2311.020 3557.200 ;
        RECT 2488.020 -37.520 2491.020 3557.200 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 405.000 2855.000 781.480 3301.235 ;
        RECT 955.000 2855.000 1331.480 3301.235 ;
      LAYER li1 ;
        RECT 583.425 2839.425 583.595 2842.655 ;
        RECT 515.805 2621.485 517.355 2621.655 ;
        RECT 515.805 2621.145 515.975 2621.485 ;
        RECT 541.565 2620.125 541.735 2621.315 ;
        RECT 528.685 2617.405 528.855 2619.615 ;
        RECT 565.945 2618.085 566.115 2621.655 ;
        RECT 589.865 2619.105 590.035 2620.295 ;
        RECT 606.885 2619.445 607.055 2620.295 ;
        RECT 613.325 2619.105 613.495 2621.315 ;
        RECT 613.785 2618.085 613.955 2621.655 ;
        RECT 662.545 2615.025 662.715 2621.655 ;
        RECT 663.005 2615.365 663.175 2621.315 ;
        RECT 688.765 2615.365 688.935 2616.215 ;
        RECT 709.925 2616.045 710.095 2621.315 ;
        RECT 710.385 2615.025 710.555 2621.655 ;
        RECT 780.765 2617.745 780.935 2621.315 ;
        RECT 1070.105 2619.105 1070.275 2620.635 ;
        RECT 1217.765 2619.105 1217.935 2619.955 ;
        RECT 1218.225 2618.425 1218.395 2619.955 ;
        RECT 737.985 2615.025 738.155 2616.215 ;
      LAYER li1 ;
        RECT 355.450 1610.795 1354.110 2598.325 ;
      LAYER li1 ;
        RECT 1400.845 2512.345 1401.015 2513.195 ;
        RECT 1448.225 2511.665 1448.395 2513.195 ;
        RECT 1449.145 2511.665 1449.315 2513.535 ;
        RECT 1497.445 2513.365 1497.615 2514.215 ;
        RECT 1545.285 2513.025 1545.455 2514.215 ;
        RECT 1559.085 2513.025 1559.715 2513.195 ;
        RECT 1603.245 2449.445 1603.415 2477.495 ;
        RECT 1604.165 2436.185 1604.335 2449.275 ;
        RECT 1602.325 2401.505 1602.495 2414.255 ;
        RECT 1604.165 2394.705 1604.335 2397.255 ;
        RECT 1601.865 2337.925 1602.035 2339.115 ;
        RECT 1603.705 2337.585 1603.875 2380.255 ;
        RECT 1604.165 2336.905 1604.335 2378.895 ;
        RECT 1600.945 2233.885 1601.115 2261.595 ;
        RECT 1601.405 2234.225 1601.575 2287.435 ;
        RECT 1601.865 2283.185 1602.035 2284.715 ;
        RECT 1603.245 2263.125 1603.415 2286.755 ;
        RECT 1601.865 2234.905 1602.035 2236.775 ;
        RECT 1603.245 2234.565 1603.415 2249.355 ;
        RECT 1603.705 2235.585 1603.875 2287.435 ;
        RECT 1604.165 2282.505 1604.335 2284.715 ;
        RECT 1604.165 2235.245 1604.335 2263.295 ;
      LAYER li1 ;
        RECT 1605.000 2205.000 2051.235 2581.480 ;
      LAYER li1 ;
        RECT 1603.245 1891.505 1603.415 1898.815 ;
        RECT 1603.705 1897.625 1603.875 1906.975 ;
        RECT 1448.685 1883.345 1449.315 1883.515 ;
        RECT 1490.545 1883.005 1490.715 1883.855 ;
        RECT 1514.465 1882.665 1514.635 1883.855 ;
        RECT 1600.485 1864.645 1600.655 1873.315 ;
        RECT 1604.165 1873.145 1604.335 1901.535 ;
        RECT 1601.405 1839.145 1601.575 1855.295 ;
        RECT 1462.945 1834.555 1463.115 1834.895 ;
        RECT 1462.485 1834.385 1463.115 1834.555 ;
        RECT 1490.545 1834.385 1490.715 1835.235 ;
        RECT 1538.845 1834.045 1539.015 1834.895 ;
        RECT 1587.145 1831.325 1587.315 1834.895 ;
        RECT 1601.405 1779.305 1601.575 1800.895 ;
        RECT 1601.865 1799.365 1602.035 1843.055 ;
        RECT 1602.325 1818.745 1602.495 1864.815 ;
        RECT 1604.165 1852.405 1604.335 1858.015 ;
      LAYER li1 ;
        RECT 1605.000 1605.000 2051.235 1981.480 ;
      LAYER mcon ;
        RECT 583.425 2842.485 583.595 2842.655 ;
        RECT 517.185 2621.485 517.355 2621.655 ;
        RECT 565.945 2621.485 566.115 2621.655 ;
        RECT 541.565 2621.145 541.735 2621.315 ;
        RECT 528.685 2619.445 528.855 2619.615 ;
        RECT 613.785 2621.485 613.955 2621.655 ;
        RECT 613.325 2621.145 613.495 2621.315 ;
        RECT 589.865 2620.125 590.035 2620.295 ;
        RECT 606.885 2620.125 607.055 2620.295 ;
        RECT 662.545 2621.485 662.715 2621.655 ;
        RECT 710.385 2621.485 710.555 2621.655 ;
        RECT 663.005 2621.145 663.175 2621.315 ;
        RECT 709.925 2621.145 710.095 2621.315 ;
        RECT 688.765 2616.045 688.935 2616.215 ;
        RECT 780.765 2621.145 780.935 2621.315 ;
        RECT 1070.105 2620.465 1070.275 2620.635 ;
        RECT 1217.765 2619.785 1217.935 2619.955 ;
        RECT 1218.225 2619.785 1218.395 2619.955 ;
        RECT 737.985 2616.045 738.155 2616.215 ;
        RECT 1497.445 2514.045 1497.615 2514.215 ;
        RECT 1449.145 2513.365 1449.315 2513.535 ;
        RECT 1545.285 2514.045 1545.455 2514.215 ;
        RECT 1400.845 2513.025 1401.015 2513.195 ;
        RECT 1448.225 2513.025 1448.395 2513.195 ;
        RECT 1559.545 2513.025 1559.715 2513.195 ;
        RECT 1603.245 2477.325 1603.415 2477.495 ;
        RECT 1603.245 2454.545 1603.415 2454.715 ;
        RECT 1604.165 2449.105 1604.335 2449.275 ;
        RECT 1602.325 2414.085 1602.495 2414.255 ;
        RECT 1604.165 2397.085 1604.335 2397.255 ;
        RECT 1603.705 2380.085 1603.875 2380.255 ;
        RECT 1603.705 2352.205 1603.875 2352.375 ;
        RECT 1601.865 2338.945 1602.035 2339.115 ;
        RECT 1604.165 2378.725 1604.335 2378.895 ;
        RECT 1601.405 2287.265 1601.575 2287.435 ;
        RECT 1600.945 2261.425 1601.115 2261.595 ;
        RECT 1603.705 2287.265 1603.875 2287.435 ;
        RECT 1603.245 2286.585 1603.415 2286.755 ;
        RECT 1601.865 2284.545 1602.035 2284.715 ;
        RECT 1603.245 2249.185 1603.415 2249.355 ;
        RECT 1601.865 2236.605 1602.035 2236.775 ;
        RECT 1604.165 2284.545 1604.335 2284.715 ;
        RECT 1604.165 2263.125 1604.335 2263.295 ;
        RECT 1603.705 1906.805 1603.875 1906.975 ;
        RECT 1603.245 1898.645 1603.415 1898.815 ;
        RECT 1604.165 1901.365 1604.335 1901.535 ;
        RECT 1490.545 1883.685 1490.715 1883.855 ;
        RECT 1449.145 1883.345 1449.315 1883.515 ;
        RECT 1514.465 1883.685 1514.635 1883.855 ;
        RECT 1600.485 1873.145 1600.655 1873.315 ;
        RECT 1602.325 1864.645 1602.495 1864.815 ;
        RECT 1601.405 1855.125 1601.575 1855.295 ;
        RECT 1601.865 1842.885 1602.035 1843.055 ;
        RECT 1490.545 1835.065 1490.715 1835.235 ;
        RECT 1462.945 1834.725 1463.115 1834.895 ;
        RECT 1538.845 1834.725 1539.015 1834.895 ;
        RECT 1587.145 1834.725 1587.315 1834.895 ;
        RECT 1604.165 1857.845 1604.335 1858.015 ;
        RECT 1601.865 1813.305 1602.035 1813.475 ;
        RECT 1601.405 1800.725 1601.575 1800.895 ;
      LAYER met1 ;
        RECT 405.000 2855.000 781.480 3301.235 ;
      LAYER met1 ;
        RECT 782.990 3277.840 783.310 3277.900 ;
        RECT 938.470 3277.840 938.790 3277.900 ;
        RECT 782.990 3277.700 938.790 3277.840 ;
        RECT 782.990 3277.640 783.310 3277.700 ;
        RECT 938.470 3277.640 938.790 3277.700 ;
      LAYER met1 ;
        RECT 955.000 2855.000 1331.480 3301.235 ;
      LAYER met1 ;
        RECT 583.365 2842.640 583.655 2842.685 ;
        RECT 597.150 2842.640 597.470 2842.700 ;
        RECT 642.230 2842.640 642.550 2842.700 ;
        RECT 583.365 2842.500 642.550 2842.640 ;
        RECT 583.365 2842.455 583.655 2842.500 ;
        RECT 597.150 2842.440 597.470 2842.500 ;
        RECT 642.230 2842.440 642.550 2842.500 ;
        RECT 604.970 2841.620 605.290 2841.680 ;
        RECT 700.190 2841.620 700.510 2841.680 ;
        RECT 604.970 2841.480 700.510 2841.620 ;
        RECT 604.970 2841.420 605.290 2841.480 ;
        RECT 700.190 2841.420 700.510 2841.480 ;
        RECT 621.530 2841.280 621.850 2841.340 ;
        RECT 585.280 2841.140 621.850 2841.280 ;
        RECT 482.610 2839.920 482.930 2839.980 ;
        RECT 526.310 2839.920 526.630 2839.980 ;
        RECT 573.690 2839.920 574.010 2839.980 ;
        RECT 585.280 2839.920 585.420 2841.140 ;
        RECT 621.530 2841.080 621.850 2841.140 ;
        RECT 642.230 2840.940 642.550 2841.000 ;
        RECT 745.270 2840.940 745.590 2841.000 ;
        RECT 642.230 2840.800 745.590 2840.940 ;
        RECT 642.230 2840.740 642.550 2840.800 ;
        RECT 745.270 2840.740 745.590 2840.800 ;
        RECT 620.610 2840.600 620.930 2840.660 ;
        RECT 734.690 2840.600 735.010 2840.660 ;
        RECT 620.610 2840.460 735.010 2840.600 ;
        RECT 620.610 2840.400 620.930 2840.460 ;
        RECT 734.690 2840.400 735.010 2840.460 ;
        RECT 1089.350 2840.600 1089.670 2840.660 ;
        RECT 1135.810 2840.600 1136.130 2840.660 ;
        RECT 1179.970 2840.600 1180.290 2840.660 ;
        RECT 1089.350 2840.460 1180.290 2840.600 ;
        RECT 1089.350 2840.400 1089.670 2840.460 ;
        RECT 1135.810 2840.400 1136.130 2840.460 ;
        RECT 1179.970 2840.400 1180.290 2840.460 ;
        RECT 600.370 2840.260 600.690 2840.320 ;
        RECT 720.890 2840.260 721.210 2840.320 ;
        RECT 600.370 2840.120 721.210 2840.260 ;
        RECT 600.370 2840.060 600.690 2840.120 ;
        RECT 720.890 2840.060 721.210 2840.120 ;
        RECT 482.610 2839.780 585.420 2839.920 ;
        RECT 1018.510 2839.920 1018.830 2839.980 ;
        RECT 1065.430 2839.920 1065.750 2839.980 ;
        RECT 1111.890 2839.920 1112.210 2839.980 ;
        RECT 1159.270 2839.920 1159.590 2839.980 ;
        RECT 1018.510 2839.780 1159.590 2839.920 ;
        RECT 482.610 2839.720 482.930 2839.780 ;
        RECT 526.310 2839.720 526.630 2839.780 ;
        RECT 573.690 2839.720 574.010 2839.780 ;
        RECT 1018.510 2839.720 1018.830 2839.780 ;
        RECT 1065.430 2839.720 1065.750 2839.780 ;
        RECT 1111.890 2839.720 1112.210 2839.780 ;
        RECT 1159.270 2839.720 1159.590 2839.780 ;
        RECT 510.210 2839.580 510.530 2839.640 ;
        RECT 549.310 2839.580 549.630 2839.640 ;
        RECT 583.365 2839.580 583.655 2839.625 ;
        RECT 510.210 2839.440 583.655 2839.580 ;
        RECT 510.210 2839.380 510.530 2839.440 ;
        RECT 549.310 2839.380 549.630 2839.440 ;
        RECT 583.365 2839.395 583.655 2839.440 ;
        RECT 627.510 2839.580 627.830 2839.640 ;
        RECT 762.290 2839.580 762.610 2839.640 ;
        RECT 627.510 2839.440 762.610 2839.580 ;
        RECT 627.510 2839.380 627.830 2839.440 ;
        RECT 762.290 2839.380 762.610 2839.440 ;
        RECT 1024.030 2839.580 1024.350 2839.640 ;
        RECT 1070.490 2839.580 1070.810 2839.640 ;
        RECT 1118.330 2839.580 1118.650 2839.640 ;
        RECT 1159.730 2839.580 1160.050 2839.640 ;
        RECT 1024.030 2839.440 1160.050 2839.580 ;
        RECT 1024.030 2839.380 1024.350 2839.440 ;
        RECT 1070.490 2839.380 1070.810 2839.440 ;
        RECT 1118.330 2839.380 1118.650 2839.440 ;
        RECT 1159.730 2839.380 1160.050 2839.440 ;
        RECT 590.250 2839.240 590.570 2839.300 ;
        RECT 713.990 2839.240 714.310 2839.300 ;
        RECT 590.250 2839.100 714.310 2839.240 ;
        RECT 590.250 2839.040 590.570 2839.100 ;
        RECT 713.990 2839.040 714.310 2839.100 ;
        RECT 427.410 2838.560 427.730 2838.620 ;
        RECT 455.470 2838.560 455.790 2838.620 ;
        RECT 427.410 2838.420 455.790 2838.560 ;
        RECT 427.410 2838.360 427.730 2838.420 ;
        RECT 455.470 2838.360 455.790 2838.420 ;
        RECT 503.310 2838.560 503.630 2838.620 ;
        RECT 783.910 2838.560 784.230 2838.620 ;
        RECT 503.310 2838.420 784.230 2838.560 ;
        RECT 503.310 2838.360 503.630 2838.420 ;
        RECT 783.910 2838.360 784.230 2838.420 ;
        RECT 489.510 2838.220 489.830 2838.280 ;
        RECT 776.090 2838.220 776.410 2838.280 ;
        RECT 489.510 2838.080 776.410 2838.220 ;
        RECT 489.510 2838.020 489.830 2838.080 ;
        RECT 776.090 2838.020 776.410 2838.080 ;
        RECT 475.710 2837.880 476.030 2837.940 ;
        RECT 769.190 2837.880 769.510 2837.940 ;
        RECT 475.710 2837.740 769.510 2837.880 ;
        RECT 475.710 2837.680 476.030 2837.740 ;
        RECT 769.190 2837.680 769.510 2837.740 ;
        RECT 551.610 2837.540 551.930 2837.600 ;
        RECT 693.290 2837.540 693.610 2837.600 ;
        RECT 551.610 2837.400 693.610 2837.540 ;
        RECT 551.610 2837.340 551.930 2837.400 ;
        RECT 693.290 2837.340 693.610 2837.400 ;
        RECT 406.710 2836.860 407.030 2836.920 ;
        RECT 441.670 2836.860 441.990 2836.920 ;
        RECT 406.710 2836.720 441.990 2836.860 ;
        RECT 406.710 2836.660 407.030 2836.720 ;
        RECT 441.670 2836.660 441.990 2836.720 ;
        RECT 627.050 2836.860 627.370 2836.920 ;
        RECT 1024.030 2836.860 1024.350 2836.920 ;
        RECT 627.050 2836.720 1024.350 2836.860 ;
        RECT 627.050 2836.660 627.370 2836.720 ;
        RECT 1024.030 2836.660 1024.350 2836.720 ;
        RECT 1045.190 2836.860 1045.510 2836.920 ;
        RECT 1089.350 2836.860 1089.670 2836.920 ;
        RECT 1045.190 2836.720 1089.670 2836.860 ;
        RECT 1045.190 2836.660 1045.510 2836.720 ;
        RECT 1089.350 2836.660 1089.670 2836.720 ;
        RECT 413.610 2836.520 413.930 2836.580 ;
        RECT 449.950 2836.520 450.270 2836.580 ;
        RECT 413.610 2836.380 450.270 2836.520 ;
        RECT 413.610 2836.320 413.930 2836.380 ;
        RECT 449.950 2836.320 450.270 2836.380 ;
        RECT 390.610 2836.180 390.930 2836.240 ;
        RECT 434.770 2836.180 435.090 2836.240 ;
        RECT 390.610 2836.040 435.090 2836.180 ;
        RECT 390.610 2835.980 390.930 2836.040 ;
        RECT 434.770 2835.980 435.090 2836.040 ;
        RECT 613.250 2836.180 613.570 2836.240 ;
        RECT 1018.510 2836.180 1018.830 2836.240 ;
        RECT 613.250 2836.040 1018.830 2836.180 ;
        RECT 613.250 2835.980 613.570 2836.040 ;
        RECT 1018.510 2835.980 1018.830 2836.040 ;
        RECT 558.510 2628.780 558.830 2628.840 ;
        RECT 907.190 2628.780 907.510 2628.840 ;
        RECT 558.510 2628.640 907.510 2628.780 ;
        RECT 558.510 2628.580 558.830 2628.640 ;
        RECT 907.190 2628.580 907.510 2628.640 ;
        RECT 640.850 2628.100 641.170 2628.160 ;
        RECT 1040.590 2628.100 1040.910 2628.160 ;
        RECT 640.850 2627.960 1040.910 2628.100 ;
        RECT 640.850 2627.900 641.170 2627.960 ;
        RECT 1040.590 2627.900 1040.910 2627.960 ;
        RECT 506.990 2627.760 507.310 2627.820 ;
        RECT 941.690 2627.760 942.010 2627.820 ;
        RECT 506.990 2627.620 942.010 2627.760 ;
        RECT 506.990 2627.560 507.310 2627.620 ;
        RECT 941.690 2627.560 942.010 2627.620 ;
        RECT 497.330 2627.420 497.650 2627.480 ;
        RECT 942.150 2627.420 942.470 2627.480 ;
        RECT 497.330 2627.280 942.470 2627.420 ;
        RECT 497.330 2627.220 497.650 2627.280 ;
        RECT 942.150 2627.220 942.470 2627.280 ;
        RECT 488.130 2627.080 488.450 2627.140 ;
        RECT 942.610 2627.080 942.930 2627.140 ;
        RECT 488.130 2626.940 942.930 2627.080 ;
        RECT 488.130 2626.880 488.450 2626.940 ;
        RECT 942.610 2626.880 942.930 2626.940 ;
        RECT 478.470 2626.740 478.790 2626.800 ;
        RECT 943.070 2626.740 943.390 2626.800 ;
        RECT 478.470 2626.600 943.390 2626.740 ;
        RECT 478.470 2626.540 478.790 2626.600 ;
        RECT 943.070 2626.540 943.390 2626.600 ;
        RECT 468.810 2626.400 469.130 2626.460 ;
        RECT 943.530 2626.400 943.850 2626.460 ;
        RECT 468.810 2626.260 943.850 2626.400 ;
        RECT 468.810 2626.200 469.130 2626.260 ;
        RECT 943.530 2626.200 943.850 2626.260 ;
        RECT 459.150 2626.060 459.470 2626.120 ;
        RECT 943.990 2626.060 944.310 2626.120 ;
        RECT 459.150 2625.920 944.310 2626.060 ;
        RECT 459.150 2625.860 459.470 2625.920 ;
        RECT 943.990 2625.860 944.310 2625.920 ;
        RECT 430.630 2625.720 430.950 2625.780 ;
        RECT 944.450 2625.720 944.770 2625.780 ;
        RECT 430.630 2625.580 944.770 2625.720 ;
        RECT 430.630 2625.520 430.950 2625.580 ;
        RECT 944.450 2625.520 944.770 2625.580 ;
        RECT 449.950 2625.380 450.270 2625.440 ;
        RECT 979.870 2625.380 980.190 2625.440 ;
        RECT 449.950 2625.240 980.190 2625.380 ;
        RECT 449.950 2625.180 450.270 2625.240 ;
        RECT 979.870 2625.180 980.190 2625.240 ;
        RECT 544.710 2625.040 545.030 2625.100 ;
        RECT 878.670 2625.040 878.990 2625.100 ;
        RECT 544.710 2624.900 878.990 2625.040 ;
        RECT 544.710 2624.840 545.030 2624.900 ;
        RECT 878.670 2624.840 878.990 2624.900 ;
        RECT 537.810 2624.700 538.130 2624.760 ;
        RECT 869.010 2624.700 869.330 2624.760 ;
        RECT 537.810 2624.560 869.330 2624.700 ;
        RECT 537.810 2624.500 538.130 2624.560 ;
        RECT 869.010 2624.500 869.330 2624.560 ;
        RECT 524.010 2624.360 524.330 2624.420 ;
        RECT 850.150 2624.360 850.470 2624.420 ;
        RECT 524.010 2624.220 850.470 2624.360 ;
        RECT 524.010 2624.160 524.330 2624.220 ;
        RECT 850.150 2624.160 850.470 2624.220 ;
        RECT 530.910 2624.020 531.230 2624.080 ;
        RECT 859.810 2624.020 860.130 2624.080 ;
        RECT 530.910 2623.880 860.130 2624.020 ;
        RECT 530.910 2623.820 531.230 2623.880 ;
        RECT 859.810 2623.820 860.130 2623.880 ;
        RECT 468.350 2623.680 468.670 2623.740 ;
        RECT 754.930 2623.680 755.250 2623.740 ;
        RECT 468.350 2623.540 755.250 2623.680 ;
        RECT 468.350 2623.480 468.670 2623.540 ;
        RECT 754.930 2623.480 755.250 2623.540 ;
        RECT 373.590 2621.980 373.910 2622.040 ;
        RECT 379.110 2621.980 379.430 2622.040 ;
        RECT 373.590 2621.840 379.430 2621.980 ;
        RECT 373.590 2621.780 373.910 2621.840 ;
        RECT 379.110 2621.780 379.430 2621.840 ;
        RECT 402.110 2621.980 402.430 2622.040 ;
        RECT 406.710 2621.980 407.030 2622.040 ;
        RECT 402.110 2621.840 407.030 2621.980 ;
        RECT 402.110 2621.780 402.430 2621.840 ;
        RECT 406.710 2621.780 407.030 2621.840 ;
        RECT 421.430 2621.980 421.750 2622.040 ;
        RECT 427.410 2621.980 427.730 2622.040 ;
        RECT 421.430 2621.840 427.730 2621.980 ;
        RECT 421.430 2621.780 421.750 2621.840 ;
        RECT 427.410 2621.780 427.730 2621.840 ;
        RECT 475.250 2621.980 475.570 2622.040 ;
        RECT 764.130 2621.980 764.450 2622.040 ;
        RECT 475.250 2621.840 764.450 2621.980 ;
        RECT 475.250 2621.780 475.570 2621.840 ;
        RECT 764.130 2621.780 764.450 2621.840 ;
        RECT 769.190 2621.980 769.510 2622.040 ;
        RECT 773.790 2621.980 774.110 2622.040 ;
        RECT 769.190 2621.840 774.110 2621.980 ;
        RECT 769.190 2621.780 769.510 2621.840 ;
        RECT 773.790 2621.780 774.110 2621.840 ;
        RECT 776.090 2621.980 776.410 2622.040 ;
        RECT 792.650 2621.980 792.970 2622.040 ;
        RECT 811.970 2621.980 812.290 2622.040 ;
        RECT 776.090 2621.840 792.970 2621.980 ;
        RECT 776.090 2621.780 776.410 2621.840 ;
        RECT 792.650 2621.780 792.970 2621.840 ;
        RECT 796.420 2621.840 812.290 2621.980 ;
        RECT 495.950 2621.640 496.270 2621.700 ;
        RECT 517.125 2621.640 517.415 2621.685 ;
        RECT 565.885 2621.640 566.175 2621.685 ;
        RECT 495.950 2621.500 516.420 2621.640 ;
        RECT 495.950 2621.440 496.270 2621.500 ;
        RECT 482.150 2621.300 482.470 2621.360 ;
        RECT 515.745 2621.300 516.035 2621.345 ;
        RECT 482.150 2621.160 516.035 2621.300 ;
        RECT 516.280 2621.300 516.420 2621.500 ;
        RECT 517.125 2621.500 566.175 2621.640 ;
        RECT 517.125 2621.455 517.415 2621.500 ;
        RECT 565.885 2621.455 566.175 2621.500 ;
        RECT 613.725 2621.640 614.015 2621.685 ;
        RECT 662.485 2621.640 662.775 2621.685 ;
        RECT 613.725 2621.500 662.775 2621.640 ;
        RECT 613.725 2621.455 614.015 2621.500 ;
        RECT 662.485 2621.455 662.775 2621.500 ;
        RECT 710.325 2621.640 710.615 2621.685 ;
        RECT 782.070 2621.640 782.390 2621.700 ;
        RECT 710.325 2621.500 782.390 2621.640 ;
        RECT 710.325 2621.455 710.615 2621.500 ;
        RECT 782.070 2621.440 782.390 2621.500 ;
        RECT 541.505 2621.300 541.795 2621.345 ;
        RECT 516.280 2621.160 541.795 2621.300 ;
        RECT 482.150 2621.100 482.470 2621.160 ;
        RECT 515.745 2621.115 516.035 2621.160 ;
        RECT 541.505 2621.115 541.795 2621.160 ;
        RECT 613.265 2621.300 613.555 2621.345 ;
        RECT 662.945 2621.300 663.235 2621.345 ;
        RECT 613.265 2621.160 663.235 2621.300 ;
        RECT 613.265 2621.115 613.555 2621.160 ;
        RECT 662.945 2621.115 663.235 2621.160 ;
        RECT 709.865 2621.300 710.155 2621.345 ;
        RECT 780.705 2621.300 780.995 2621.345 ;
        RECT 709.865 2621.160 780.995 2621.300 ;
        RECT 709.865 2621.115 710.155 2621.160 ;
        RECT 780.705 2621.115 780.995 2621.160 ;
        RECT 783.910 2621.300 784.230 2621.360 ;
        RECT 796.420 2621.300 796.560 2621.840 ;
        RECT 811.970 2621.780 812.290 2621.840 ;
        RECT 1041.510 2621.980 1041.830 2622.040 ;
        RECT 1097.630 2621.980 1097.950 2622.040 ;
        RECT 1041.510 2621.840 1097.950 2621.980 ;
        RECT 1041.510 2621.780 1041.830 2621.840 ;
        RECT 1097.630 2621.780 1097.950 2621.840 ;
        RECT 1145.010 2621.980 1145.330 2622.040 ;
        RECT 1269.210 2621.980 1269.530 2622.040 ;
        RECT 1145.010 2621.840 1269.530 2621.980 ;
        RECT 1145.010 2621.780 1145.330 2621.840 ;
        RECT 1269.210 2621.780 1269.530 2621.840 ;
        RECT 1138.110 2621.640 1138.430 2621.700 ;
        RECT 1260.010 2621.640 1260.330 2621.700 ;
        RECT 1138.110 2621.500 1260.330 2621.640 ;
        RECT 1138.110 2621.440 1138.430 2621.500 ;
        RECT 1260.010 2621.440 1260.330 2621.500 ;
        RECT 783.910 2621.160 796.560 2621.300 ;
        RECT 1048.410 2621.300 1048.730 2621.360 ;
        RECT 1107.290 2621.300 1107.610 2621.360 ;
        RECT 1048.410 2621.160 1107.610 2621.300 ;
        RECT 783.910 2621.100 784.230 2621.160 ;
        RECT 1048.410 2621.100 1048.730 2621.160 ;
        RECT 1107.290 2621.100 1107.610 2621.160 ;
        RECT 1158.810 2621.300 1159.130 2621.360 ;
        RECT 1288.530 2621.300 1288.850 2621.360 ;
        RECT 1158.810 2621.160 1288.850 2621.300 ;
        RECT 1158.810 2621.100 1159.130 2621.160 ;
        RECT 1288.530 2621.100 1288.850 2621.160 ;
        RECT 509.750 2620.960 510.070 2621.020 ;
        RECT 821.630 2620.960 821.950 2621.020 ;
        RECT 509.750 2620.820 821.950 2620.960 ;
        RECT 509.750 2620.760 510.070 2620.820 ;
        RECT 821.630 2620.760 821.950 2620.820 ;
        RECT 1062.210 2620.960 1062.530 2621.020 ;
        RECT 1135.810 2620.960 1136.130 2621.020 ;
        RECT 1062.210 2620.820 1136.130 2620.960 ;
        RECT 1062.210 2620.760 1062.530 2620.820 ;
        RECT 1135.810 2620.760 1136.130 2620.820 ;
        RECT 1151.910 2620.960 1152.230 2621.020 ;
        RECT 1278.870 2620.960 1279.190 2621.020 ;
        RECT 1151.910 2620.820 1279.190 2620.960 ;
        RECT 1151.910 2620.760 1152.230 2620.820 ;
        RECT 1278.870 2620.760 1279.190 2620.820 ;
        RECT 394.290 2620.620 394.610 2620.680 ;
        RECT 440.290 2620.620 440.610 2620.680 ;
        RECT 394.290 2620.480 440.610 2620.620 ;
        RECT 394.290 2620.420 394.610 2620.480 ;
        RECT 440.290 2620.420 440.610 2620.480 ;
        RECT 516.650 2620.620 516.970 2620.680 ;
        RECT 840.490 2620.620 840.810 2620.680 ;
        RECT 516.650 2620.480 840.810 2620.620 ;
        RECT 516.650 2620.420 516.970 2620.480 ;
        RECT 840.490 2620.420 840.810 2620.480 ;
        RECT 1070.045 2620.620 1070.335 2620.665 ;
        RECT 1126.610 2620.620 1126.930 2620.680 ;
        RECT 1070.045 2620.480 1126.930 2620.620 ;
        RECT 1070.045 2620.435 1070.335 2620.480 ;
        RECT 1126.610 2620.420 1126.930 2620.480 ;
        RECT 1165.710 2620.620 1166.030 2620.680 ;
        RECT 1297.730 2620.620 1298.050 2620.680 ;
        RECT 1165.710 2620.480 1298.050 2620.620 ;
        RECT 1165.710 2620.420 1166.030 2620.480 ;
        RECT 1297.730 2620.420 1298.050 2620.480 ;
        RECT 393.830 2620.280 394.150 2620.340 ;
        RECT 541.505 2620.280 541.795 2620.325 ;
        RECT 589.805 2620.280 590.095 2620.325 ;
        RECT 393.830 2620.140 531.600 2620.280 ;
        RECT 393.830 2620.080 394.150 2620.140 ;
        RECT 393.370 2619.940 393.690 2620.000 ;
        RECT 531.460 2619.940 531.600 2620.140 ;
        RECT 541.505 2620.140 590.095 2620.280 ;
        RECT 541.505 2620.095 541.795 2620.140 ;
        RECT 589.805 2620.095 590.095 2620.140 ;
        RECT 606.825 2620.280 607.115 2620.325 ;
        RECT 926.510 2620.280 926.830 2620.340 ;
        RECT 606.825 2620.140 926.830 2620.280 ;
        RECT 606.825 2620.095 607.115 2620.140 ;
        RECT 926.510 2620.080 926.830 2620.140 ;
        RECT 1020.810 2620.280 1021.130 2620.340 ;
        RECT 1069.110 2620.280 1069.430 2620.340 ;
        RECT 1020.810 2620.140 1069.430 2620.280 ;
        RECT 1020.810 2620.080 1021.130 2620.140 ;
        RECT 1069.110 2620.080 1069.430 2620.140 ;
        RECT 1069.570 2620.280 1069.890 2620.340 ;
        RECT 1145.470 2620.280 1145.790 2620.340 ;
        RECT 1069.570 2620.140 1145.790 2620.280 ;
        RECT 1069.570 2620.080 1069.890 2620.140 ;
        RECT 1145.470 2620.080 1145.790 2620.140 ;
        RECT 1172.610 2620.280 1172.930 2620.340 ;
        RECT 1317.050 2620.280 1317.370 2620.340 ;
        RECT 1172.610 2620.140 1317.370 2620.280 ;
        RECT 1172.610 2620.080 1172.930 2620.140 ;
        RECT 1317.050 2620.080 1317.370 2620.140 ;
        RECT 545.170 2619.940 545.490 2620.000 ;
        RECT 393.370 2619.800 529.300 2619.940 ;
        RECT 531.460 2619.800 545.490 2619.940 ;
        RECT 393.370 2619.740 393.690 2619.800 ;
        RECT 391.530 2619.600 391.850 2619.660 ;
        RECT 528.625 2619.600 528.915 2619.645 ;
        RECT 391.530 2619.460 528.915 2619.600 ;
        RECT 529.160 2619.600 529.300 2619.800 ;
        RECT 545.170 2619.740 545.490 2619.800 ;
        RECT 592.550 2619.940 592.870 2620.000 ;
        RECT 955.030 2619.940 955.350 2620.000 ;
        RECT 592.550 2619.800 955.350 2619.940 ;
        RECT 592.550 2619.740 592.870 2619.800 ;
        RECT 955.030 2619.740 955.350 2619.800 ;
        RECT 1027.710 2619.940 1028.030 2620.000 ;
        RECT 1078.770 2619.940 1079.090 2620.000 ;
        RECT 1027.710 2619.800 1079.090 2619.940 ;
        RECT 1027.710 2619.740 1028.030 2619.800 ;
        RECT 1078.770 2619.740 1079.090 2619.800 ;
        RECT 1082.910 2619.940 1083.230 2620.000 ;
        RECT 1164.330 2619.940 1164.650 2620.000 ;
        RECT 1082.910 2619.800 1164.650 2619.940 ;
        RECT 1082.910 2619.740 1083.230 2619.800 ;
        RECT 1164.330 2619.740 1164.650 2619.800 ;
        RECT 1179.510 2619.940 1179.830 2620.000 ;
        RECT 1217.705 2619.940 1217.995 2619.985 ;
        RECT 1179.510 2619.800 1217.995 2619.940 ;
        RECT 1179.510 2619.740 1179.830 2619.800 ;
        RECT 1217.705 2619.755 1217.995 2619.800 ;
        RECT 1218.165 2619.940 1218.455 2619.985 ;
        RECT 1307.390 2619.940 1307.710 2620.000 ;
        RECT 1218.165 2619.800 1307.710 2619.940 ;
        RECT 1218.165 2619.755 1218.455 2619.800 ;
        RECT 1307.390 2619.740 1307.710 2619.800 ;
        RECT 554.830 2619.600 555.150 2619.660 ;
        RECT 529.160 2619.460 555.150 2619.600 ;
        RECT 391.530 2619.400 391.850 2619.460 ;
        RECT 528.625 2619.415 528.915 2619.460 ;
        RECT 554.830 2619.400 555.150 2619.460 ;
        RECT 572.310 2619.600 572.630 2619.660 ;
        RECT 606.825 2619.600 607.115 2619.645 ;
        RECT 572.310 2619.460 607.115 2619.600 ;
        RECT 572.310 2619.400 572.630 2619.460 ;
        RECT 606.825 2619.415 607.115 2619.460 ;
        RECT 613.710 2619.600 614.030 2619.660 ;
        RECT 993.210 2619.600 993.530 2619.660 ;
        RECT 613.710 2619.460 993.530 2619.600 ;
        RECT 613.710 2619.400 614.030 2619.460 ;
        RECT 993.210 2619.400 993.530 2619.460 ;
        RECT 1076.010 2619.600 1076.330 2619.660 ;
        RECT 1155.130 2619.600 1155.450 2619.660 ;
        RECT 1076.010 2619.460 1155.450 2619.600 ;
        RECT 1076.010 2619.400 1076.330 2619.460 ;
        RECT 1155.130 2619.400 1155.450 2619.460 ;
        RECT 1165.250 2619.600 1165.570 2619.660 ;
        RECT 1186.410 2619.600 1186.730 2619.660 ;
        RECT 1335.910 2619.600 1336.230 2619.660 ;
        RECT 1165.250 2619.460 1175.140 2619.600 ;
        RECT 1165.250 2619.400 1165.570 2619.460 ;
        RECT 391.990 2619.260 392.310 2619.320 ;
        RECT 573.690 2619.260 574.010 2619.320 ;
        RECT 391.990 2619.120 574.010 2619.260 ;
        RECT 391.990 2619.060 392.310 2619.120 ;
        RECT 573.690 2619.060 574.010 2619.120 ;
        RECT 589.805 2619.260 590.095 2619.305 ;
        RECT 613.265 2619.260 613.555 2619.305 ;
        RECT 589.805 2619.120 613.555 2619.260 ;
        RECT 589.805 2619.075 590.095 2619.120 ;
        RECT 613.265 2619.075 613.555 2619.120 ;
        RECT 621.530 2619.260 621.850 2619.320 ;
        RECT 627.050 2619.260 627.370 2619.320 ;
        RECT 621.530 2619.120 627.370 2619.260 ;
        RECT 621.530 2619.060 621.850 2619.120 ;
        RECT 627.050 2619.060 627.370 2619.120 ;
        RECT 1054.850 2619.260 1055.170 2619.320 ;
        RECT 1070.045 2619.260 1070.335 2619.305 ;
        RECT 1054.850 2619.120 1070.335 2619.260 ;
        RECT 1175.000 2619.260 1175.140 2619.460 ;
        RECT 1186.410 2619.460 1336.230 2619.600 ;
        RECT 1186.410 2619.400 1186.730 2619.460 ;
        RECT 1335.910 2619.400 1336.230 2619.460 ;
        RECT 1193.310 2619.260 1193.630 2619.320 ;
        RECT 1217.705 2619.260 1217.995 2619.305 ;
        RECT 1326.710 2619.260 1327.030 2619.320 ;
        RECT 1175.000 2619.120 1192.160 2619.260 ;
        RECT 1054.850 2619.060 1055.170 2619.120 ;
        RECT 1070.045 2619.075 1070.335 2619.120 ;
        RECT 392.450 2618.920 392.770 2618.980 ;
        RECT 583.350 2618.920 583.670 2618.980 ;
        RECT 392.450 2618.780 583.670 2618.920 ;
        RECT 392.450 2618.720 392.770 2618.780 ;
        RECT 583.350 2618.720 583.670 2618.780 ;
        RECT 650.050 2618.920 650.370 2618.980 ;
        RECT 1045.190 2618.920 1045.510 2618.980 ;
        RECT 650.050 2618.780 1045.510 2618.920 ;
        RECT 650.050 2618.720 650.370 2618.780 ;
        RECT 1045.190 2618.720 1045.510 2618.780 ;
        RECT 1096.710 2618.920 1097.030 2618.980 ;
        RECT 1191.470 2618.920 1191.790 2618.980 ;
        RECT 1096.710 2618.780 1191.790 2618.920 ;
        RECT 1096.710 2618.720 1097.030 2618.780 ;
        RECT 1191.470 2618.720 1191.790 2618.780 ;
        RECT 392.910 2618.580 393.230 2618.640 ;
        RECT 592.550 2618.580 592.870 2618.640 ;
        RECT 392.910 2618.440 592.870 2618.580 ;
        RECT 392.910 2618.380 393.230 2618.440 ;
        RECT 592.550 2618.380 592.870 2618.440 ;
        RECT 1089.350 2618.580 1089.670 2618.640 ;
        RECT 1183.650 2618.580 1183.970 2618.640 ;
        RECT 1089.350 2618.440 1183.970 2618.580 ;
        RECT 1192.020 2618.580 1192.160 2619.120 ;
        RECT 1193.310 2619.120 1199.980 2619.260 ;
        RECT 1193.310 2619.060 1193.630 2619.120 ;
        RECT 1199.840 2618.920 1199.980 2619.120 ;
        RECT 1217.705 2619.120 1327.030 2619.260 ;
        RECT 1217.705 2619.075 1217.995 2619.120 ;
        RECT 1326.710 2619.060 1327.030 2619.120 ;
        RECT 1345.570 2618.920 1345.890 2618.980 ;
        RECT 1199.840 2618.780 1345.890 2618.920 ;
        RECT 1345.570 2618.720 1345.890 2618.780 ;
        RECT 1218.165 2618.580 1218.455 2618.625 ;
        RECT 1192.020 2618.440 1218.455 2618.580 ;
        RECT 1089.350 2618.380 1089.670 2618.440 ;
        RECT 1183.650 2618.380 1183.970 2618.440 ;
        RECT 1218.165 2618.395 1218.455 2618.440 ;
        RECT 391.070 2618.240 391.390 2618.300 ;
        RECT 535.510 2618.240 535.830 2618.300 ;
        RECT 391.070 2618.100 535.830 2618.240 ;
        RECT 391.070 2618.040 391.390 2618.100 ;
        RECT 535.510 2618.040 535.830 2618.100 ;
        RECT 565.885 2618.240 566.175 2618.285 ;
        RECT 613.725 2618.240 614.015 2618.285 ;
        RECT 565.885 2618.100 614.015 2618.240 ;
        RECT 565.885 2618.055 566.175 2618.100 ;
        RECT 613.725 2618.055 614.015 2618.100 ;
        RECT 700.190 2618.240 700.510 2618.300 ;
        RECT 983.550 2618.240 983.870 2618.300 ;
        RECT 700.190 2618.100 983.870 2618.240 ;
        RECT 700.190 2618.040 700.510 2618.100 ;
        RECT 983.550 2618.040 983.870 2618.100 ;
        RECT 1131.210 2618.240 1131.530 2618.300 ;
        RECT 1250.350 2618.240 1250.670 2618.300 ;
        RECT 1131.210 2618.100 1250.670 2618.240 ;
        RECT 1131.210 2618.040 1131.530 2618.100 ;
        RECT 1250.350 2618.040 1250.670 2618.100 ;
        RECT 516.650 2617.900 516.970 2617.960 ;
        RECT 779.770 2617.900 780.090 2617.960 ;
        RECT 516.650 2617.760 780.090 2617.900 ;
        RECT 516.650 2617.700 516.970 2617.760 ;
        RECT 779.770 2617.700 780.090 2617.760 ;
        RECT 780.705 2617.900 780.995 2617.945 ;
        RECT 802.310 2617.900 802.630 2617.960 ;
        RECT 780.705 2617.760 802.630 2617.900 ;
        RECT 780.705 2617.715 780.995 2617.760 ;
        RECT 802.310 2617.700 802.630 2617.760 ;
        RECT 1130.750 2617.900 1131.070 2617.960 ;
        RECT 1240.690 2617.900 1241.010 2617.960 ;
        RECT 1130.750 2617.760 1241.010 2617.900 ;
        RECT 1130.750 2617.700 1131.070 2617.760 ;
        RECT 1240.690 2617.700 1241.010 2617.760 ;
        RECT 433.850 2617.560 434.170 2617.620 ;
        RECT 525.850 2617.560 526.170 2617.620 ;
        RECT 433.850 2617.420 526.170 2617.560 ;
        RECT 433.850 2617.360 434.170 2617.420 ;
        RECT 525.850 2617.360 526.170 2617.420 ;
        RECT 528.625 2617.560 528.915 2617.605 ;
        RECT 564.030 2617.560 564.350 2617.620 ;
        RECT 1002.410 2617.560 1002.730 2617.620 ;
        RECT 528.625 2617.420 564.350 2617.560 ;
        RECT 528.625 2617.375 528.915 2617.420 ;
        RECT 564.030 2617.360 564.350 2617.420 ;
        RECT 736.620 2617.420 1002.730 2617.560 ;
        RECT 734.690 2617.220 735.010 2617.280 ;
        RECT 736.620 2617.220 736.760 2617.420 ;
        RECT 1002.410 2617.360 1002.730 2617.420 ;
        RECT 1117.410 2617.560 1117.730 2617.620 ;
        RECT 1221.830 2617.560 1222.150 2617.620 ;
        RECT 1117.410 2617.420 1222.150 2617.560 ;
        RECT 1117.410 2617.360 1117.730 2617.420 ;
        RECT 1221.830 2617.360 1222.150 2617.420 ;
        RECT 964.230 2617.220 964.550 2617.280 ;
        RECT 734.690 2617.080 736.760 2617.220 ;
        RECT 737.080 2617.080 964.550 2617.220 ;
        RECT 734.690 2617.020 735.010 2617.080 ;
        RECT 625.210 2616.880 625.530 2616.940 ;
        RECT 707.090 2616.880 707.410 2616.940 ;
        RECT 625.210 2616.740 707.410 2616.880 ;
        RECT 625.210 2616.680 625.530 2616.740 ;
        RECT 707.090 2616.680 707.410 2616.740 ;
        RECT 720.890 2616.880 721.210 2616.940 ;
        RECT 737.080 2616.880 737.220 2617.080 ;
        RECT 964.230 2617.020 964.550 2617.080 ;
        RECT 1124.310 2617.220 1124.630 2617.280 ;
        RECT 1231.030 2617.220 1231.350 2617.280 ;
        RECT 1124.310 2617.080 1231.350 2617.220 ;
        RECT 1124.310 2617.020 1124.630 2617.080 ;
        RECT 1231.030 2617.020 1231.350 2617.080 ;
        RECT 720.890 2616.740 737.220 2616.880 ;
        RECT 1110.510 2616.880 1110.830 2616.940 ;
        RECT 1212.170 2616.880 1212.490 2616.940 ;
        RECT 1110.510 2616.740 1212.490 2616.880 ;
        RECT 720.890 2616.680 721.210 2616.740 ;
        RECT 1110.510 2616.680 1110.830 2616.740 ;
        RECT 1212.170 2616.680 1212.490 2616.740 ;
        RECT 1103.610 2616.540 1103.930 2616.600 ;
        RECT 1202.510 2616.540 1202.830 2616.600 ;
        RECT 1103.610 2616.400 1202.830 2616.540 ;
        RECT 1103.610 2616.340 1103.930 2616.400 ;
        RECT 1202.510 2616.340 1202.830 2616.400 ;
        RECT 688.705 2616.200 688.995 2616.245 ;
        RECT 709.865 2616.200 710.155 2616.245 ;
        RECT 688.705 2616.060 710.155 2616.200 ;
        RECT 688.705 2616.015 688.995 2616.060 ;
        RECT 709.865 2616.015 710.155 2616.060 ;
        RECT 737.925 2616.200 738.215 2616.245 ;
        RECT 935.710 2616.200 936.030 2616.260 ;
        RECT 737.925 2616.060 936.030 2616.200 ;
        RECT 737.925 2616.015 738.215 2616.060 ;
        RECT 935.710 2616.000 936.030 2616.060 ;
        RECT 662.945 2615.520 663.235 2615.565 ;
        RECT 688.705 2615.520 688.995 2615.565 ;
        RECT 662.945 2615.380 688.995 2615.520 ;
        RECT 662.945 2615.335 663.235 2615.380 ;
        RECT 688.705 2615.335 688.995 2615.380 ;
        RECT 693.290 2615.520 693.610 2615.580 ;
        RECT 897.530 2615.520 897.850 2615.580 ;
        RECT 693.290 2615.380 897.850 2615.520 ;
        RECT 693.290 2615.320 693.610 2615.380 ;
        RECT 897.530 2615.320 897.850 2615.380 ;
        RECT 662.485 2615.180 662.775 2615.225 ;
        RECT 710.325 2615.180 710.615 2615.225 ;
        RECT 662.485 2615.040 710.615 2615.180 ;
        RECT 662.485 2614.995 662.775 2615.040 ;
        RECT 710.325 2614.995 710.615 2615.040 ;
        RECT 713.990 2615.180 714.310 2615.240 ;
        RECT 737.925 2615.180 738.215 2615.225 ;
        RECT 713.990 2615.040 738.215 2615.180 ;
        RECT 713.990 2614.980 714.310 2615.040 ;
        RECT 737.925 2614.995 738.215 2615.040 ;
      LAYER met1 ;
        RECT 350.000 1606.500 1357.260 2605.680 ;
      LAYER met1 ;
        RECT 1371.330 2594.780 1371.650 2594.840 ;
        RECT 1507.490 2594.780 1507.810 2594.840 ;
        RECT 1371.330 2594.640 1507.810 2594.780 ;
        RECT 1371.330 2594.580 1371.650 2594.640 ;
        RECT 1507.490 2594.580 1507.810 2594.640 ;
        RECT 1369.490 2583.900 1369.810 2583.960 ;
        RECT 1688.730 2583.900 1689.050 2583.960 ;
        RECT 1369.490 2583.760 1689.050 2583.900 ;
        RECT 1369.490 2583.700 1369.810 2583.760 ;
        RECT 1688.730 2583.700 1689.050 2583.760 ;
        RECT 1691.950 2583.900 1692.270 2583.960 ;
        RECT 1704.370 2583.900 1704.690 2583.960 ;
        RECT 1691.950 2583.760 1704.690 2583.900 ;
        RECT 1691.950 2583.700 1692.270 2583.760 ;
        RECT 1704.370 2583.700 1704.690 2583.760 ;
        RECT 1376.850 2583.560 1377.170 2583.620 ;
        RECT 1994.170 2583.560 1994.490 2583.620 ;
        RECT 1376.850 2583.420 1994.490 2583.560 ;
        RECT 1376.850 2583.360 1377.170 2583.420 ;
        RECT 1994.170 2583.360 1994.490 2583.420 ;
        RECT 1377.310 2583.220 1377.630 2583.280 ;
        RECT 2001.070 2583.220 2001.390 2583.280 ;
        RECT 1377.310 2583.080 2001.390 2583.220 ;
        RECT 1377.310 2583.020 1377.630 2583.080 ;
        RECT 2001.070 2583.020 2001.390 2583.080 ;
        RECT 1371.790 2582.880 1372.110 2582.940 ;
        RECT 2007.970 2582.880 2008.290 2582.940 ;
        RECT 1371.790 2582.740 2008.290 2582.880 ;
        RECT 1371.790 2582.680 1372.110 2582.740 ;
        RECT 2007.970 2582.680 2008.290 2582.740 ;
        RECT 1372.250 2582.540 1372.570 2582.600 ;
        RECT 2016.710 2582.540 2017.030 2582.600 ;
        RECT 1372.250 2582.400 2017.030 2582.540 ;
        RECT 1372.250 2582.340 1372.570 2582.400 ;
        RECT 2016.710 2582.340 2017.030 2582.400 ;
        RECT 1372.710 2582.200 1373.030 2582.260 ;
        RECT 2021.770 2582.200 2022.090 2582.260 ;
        RECT 1372.710 2582.060 2022.090 2582.200 ;
        RECT 1372.710 2582.000 1373.030 2582.060 ;
        RECT 2021.770 2582.000 2022.090 2582.060 ;
        RECT 2030.050 2582.000 2030.370 2582.260 ;
        RECT 1369.030 2581.860 1369.350 2581.920 ;
        RECT 2030.140 2581.860 2030.280 2582.000 ;
        RECT 1369.030 2581.720 2030.280 2581.860 ;
        RECT 1369.030 2581.660 1369.350 2581.720 ;
        RECT 1368.110 2574.040 1368.430 2574.100 ;
        RECT 1493.690 2574.040 1494.010 2574.100 ;
        RECT 1368.110 2573.900 1494.010 2574.040 ;
        RECT 1368.110 2573.840 1368.430 2573.900 ;
        RECT 1493.690 2573.840 1494.010 2573.900 ;
        RECT 1376.390 2560.100 1376.710 2560.160 ;
        RECT 1600.870 2560.100 1601.190 2560.160 ;
        RECT 1376.390 2559.960 1601.190 2560.100 ;
        RECT 1376.390 2559.900 1376.710 2559.960 ;
        RECT 1600.870 2559.900 1601.190 2559.960 ;
        RECT 1367.650 2553.300 1367.970 2553.360 ;
        RECT 1486.790 2553.300 1487.110 2553.360 ;
        RECT 1367.650 2553.160 1487.110 2553.300 ;
        RECT 1367.650 2553.100 1367.970 2553.160 ;
        RECT 1486.790 2553.100 1487.110 2553.160 ;
        RECT 1397.090 2546.500 1397.410 2546.560 ;
        RECT 1601.790 2546.500 1602.110 2546.560 ;
        RECT 1397.090 2546.360 1602.110 2546.500 ;
        RECT 1397.090 2546.300 1397.410 2546.360 ;
        RECT 1601.790 2546.300 1602.110 2546.360 ;
        RECT 1514.390 2539.360 1514.710 2539.420 ;
        RECT 1600.870 2539.360 1601.190 2539.420 ;
        RECT 1514.390 2539.220 1601.190 2539.360 ;
        RECT 1514.390 2539.160 1514.710 2539.220 ;
        RECT 1600.870 2539.160 1601.190 2539.220 ;
        RECT 1368.570 2532.900 1368.890 2532.960 ;
        RECT 1472.990 2532.900 1473.310 2532.960 ;
        RECT 1368.570 2532.760 1473.310 2532.900 ;
        RECT 1368.570 2532.700 1368.890 2532.760 ;
        RECT 1472.990 2532.700 1473.310 2532.760 ;
        RECT 1377.770 2532.560 1378.090 2532.620 ;
        RECT 1599.030 2532.560 1599.350 2532.620 ;
        RECT 1377.770 2532.420 1599.350 2532.560 ;
        RECT 1377.770 2532.360 1378.090 2532.420 ;
        RECT 1599.030 2532.360 1599.350 2532.420 ;
        RECT 1367.650 2526.100 1367.970 2526.160 ;
        RECT 1459.190 2526.100 1459.510 2526.160 ;
        RECT 1367.650 2525.960 1459.510 2526.100 ;
        RECT 1367.650 2525.900 1367.970 2525.960 ;
        RECT 1459.190 2525.900 1459.510 2525.960 ;
        RECT 1378.230 2525.760 1378.550 2525.820 ;
        RECT 1600.870 2525.760 1601.190 2525.820 ;
        RECT 1378.230 2525.620 1601.190 2525.760 ;
        RECT 1378.230 2525.560 1378.550 2525.620 ;
        RECT 1600.870 2525.560 1601.190 2525.620 ;
        RECT 1383.290 2518.620 1383.610 2518.680 ;
        RECT 1599.950 2518.620 1600.270 2518.680 ;
        RECT 1383.290 2518.480 1600.270 2518.620 ;
        RECT 1383.290 2518.420 1383.610 2518.480 ;
        RECT 1599.950 2518.420 1600.270 2518.480 ;
        RECT 1497.385 2514.200 1497.675 2514.245 ;
        RECT 1545.225 2514.200 1545.515 2514.245 ;
        RECT 1497.385 2514.060 1545.515 2514.200 ;
        RECT 1497.385 2514.015 1497.675 2514.060 ;
        RECT 1545.225 2514.015 1545.515 2514.060 ;
        RECT 1449.085 2513.520 1449.375 2513.565 ;
        RECT 1497.385 2513.520 1497.675 2513.565 ;
        RECT 1449.085 2513.380 1497.675 2513.520 ;
        RECT 1449.085 2513.335 1449.375 2513.380 ;
        RECT 1497.385 2513.335 1497.675 2513.380 ;
        RECT 1400.785 2513.180 1401.075 2513.225 ;
        RECT 1448.165 2513.180 1448.455 2513.225 ;
        RECT 1400.785 2513.040 1448.455 2513.180 ;
        RECT 1400.785 2512.995 1401.075 2513.040 ;
        RECT 1448.165 2512.995 1448.455 2513.040 ;
        RECT 1545.225 2513.180 1545.515 2513.225 ;
        RECT 1559.025 2513.180 1559.315 2513.225 ;
        RECT 1545.225 2513.040 1559.315 2513.180 ;
        RECT 1545.225 2512.995 1545.515 2513.040 ;
        RECT 1559.025 2512.995 1559.315 2513.040 ;
        RECT 1559.485 2513.180 1559.775 2513.225 ;
        RECT 1559.485 2513.040 1560.620 2513.180 ;
        RECT 1559.485 2512.995 1559.775 2513.040 ;
        RECT 1560.480 2512.840 1560.620 2513.040 ;
        RECT 1601.330 2512.840 1601.650 2512.900 ;
        RECT 1560.480 2512.700 1601.650 2512.840 ;
        RECT 1601.330 2512.640 1601.650 2512.700 ;
        RECT 1383.750 2512.500 1384.070 2512.560 ;
        RECT 1400.785 2512.500 1401.075 2512.545 ;
        RECT 1383.750 2512.360 1401.075 2512.500 ;
        RECT 1383.750 2512.300 1384.070 2512.360 ;
        RECT 1400.785 2512.315 1401.075 2512.360 ;
        RECT 1448.165 2511.820 1448.455 2511.865 ;
        RECT 1449.085 2511.820 1449.375 2511.865 ;
        RECT 1448.165 2511.680 1449.375 2511.820 ;
        RECT 1448.165 2511.635 1448.455 2511.680 ;
        RECT 1449.085 2511.635 1449.375 2511.680 ;
        RECT 1368.110 2505.360 1368.430 2505.420 ;
        RECT 1452.290 2505.360 1452.610 2505.420 ;
        RECT 1368.110 2505.220 1452.610 2505.360 ;
        RECT 1368.110 2505.160 1368.430 2505.220 ;
        RECT 1452.290 2505.160 1452.610 2505.220 ;
        RECT 1384.210 2505.020 1384.530 2505.080 ;
        RECT 1599.030 2505.020 1599.350 2505.080 ;
        RECT 1384.210 2504.880 1599.350 2505.020 ;
        RECT 1384.210 2504.820 1384.530 2504.880 ;
        RECT 1599.030 2504.820 1599.350 2504.880 ;
        RECT 1368.570 2498.220 1368.890 2498.280 ;
        RECT 1438.490 2498.220 1438.810 2498.280 ;
        RECT 1368.570 2498.080 1438.810 2498.220 ;
        RECT 1368.570 2498.020 1368.890 2498.080 ;
        RECT 1438.490 2498.020 1438.810 2498.080 ;
        RECT 1384.670 2497.880 1384.990 2497.940 ;
        RECT 1600.870 2497.880 1601.190 2497.940 ;
        RECT 1384.670 2497.740 1601.190 2497.880 ;
        RECT 1384.670 2497.680 1384.990 2497.740 ;
        RECT 1600.870 2497.680 1601.190 2497.740 ;
        RECT 1385.130 2491.080 1385.450 2491.140 ;
        RECT 1599.030 2491.080 1599.350 2491.140 ;
        RECT 1385.130 2490.940 1599.350 2491.080 ;
        RECT 1385.130 2490.880 1385.450 2490.940 ;
        RECT 1599.030 2490.880 1599.350 2490.940 ;
        RECT 1368.570 2484.620 1368.890 2484.680 ;
        RECT 1431.590 2484.620 1431.910 2484.680 ;
        RECT 1368.570 2484.480 1431.910 2484.620 ;
        RECT 1368.570 2484.420 1368.890 2484.480 ;
        RECT 1431.590 2484.420 1431.910 2484.480 ;
        RECT 1392.950 2484.280 1393.270 2484.340 ;
        RECT 1600.870 2484.280 1601.190 2484.340 ;
        RECT 1392.950 2484.140 1601.190 2484.280 ;
        RECT 1392.950 2484.080 1393.270 2484.140 ;
        RECT 1600.870 2484.080 1601.190 2484.140 ;
        RECT 1368.570 2478.160 1368.890 2478.220 ;
        RECT 1424.690 2478.160 1425.010 2478.220 ;
        RECT 1368.570 2478.020 1425.010 2478.160 ;
        RECT 1368.570 2477.960 1368.890 2478.020 ;
        RECT 1424.690 2477.960 1425.010 2478.020 ;
        RECT 1397.550 2477.820 1397.870 2477.880 ;
        RECT 1599.030 2477.820 1599.350 2477.880 ;
        RECT 1397.550 2477.680 1599.350 2477.820 ;
        RECT 1397.550 2477.620 1397.870 2477.680 ;
        RECT 1599.030 2477.620 1599.350 2477.680 ;
        RECT 1378.690 2477.480 1379.010 2477.540 ;
        RECT 1599.950 2477.480 1600.270 2477.540 ;
        RECT 1603.170 2477.480 1603.490 2477.540 ;
        RECT 1378.690 2477.340 1600.270 2477.480 ;
        RECT 1602.975 2477.340 1603.490 2477.480 ;
        RECT 1378.690 2477.280 1379.010 2477.340 ;
        RECT 1599.950 2477.280 1600.270 2477.340 ;
        RECT 1603.170 2477.280 1603.490 2477.340 ;
        RECT 1368.110 2470.680 1368.430 2470.740 ;
        RECT 1390.190 2470.680 1390.510 2470.740 ;
        RECT 1368.110 2470.540 1390.510 2470.680 ;
        RECT 1368.110 2470.480 1368.430 2470.540 ;
        RECT 1390.190 2470.480 1390.510 2470.540 ;
        RECT 1379.150 2470.340 1379.470 2470.400 ;
        RECT 1599.030 2470.340 1599.350 2470.400 ;
        RECT 1379.150 2470.200 1599.350 2470.340 ;
        RECT 1379.150 2470.140 1379.470 2470.200 ;
        RECT 1599.030 2470.140 1599.350 2470.200 ;
        RECT 1379.610 2463.540 1379.930 2463.600 ;
        RECT 1600.870 2463.540 1601.190 2463.600 ;
        RECT 1379.610 2463.400 1601.190 2463.540 ;
        RECT 1379.610 2463.340 1379.930 2463.400 ;
        RECT 1600.870 2463.340 1601.190 2463.400 ;
        RECT 1603.630 2461.640 1603.950 2461.900 ;
        RECT 1604.090 2461.640 1604.410 2461.900 ;
        RECT 1603.720 2460.880 1603.860 2461.640 ;
        RECT 1604.180 2460.880 1604.320 2461.640 ;
        RECT 1603.630 2460.620 1603.950 2460.880 ;
        RECT 1604.090 2460.620 1604.410 2460.880 ;
        RECT 1368.110 2457.080 1368.430 2457.140 ;
        RECT 1417.790 2457.080 1418.110 2457.140 ;
        RECT 1368.110 2456.940 1418.110 2457.080 ;
        RECT 1368.110 2456.880 1368.430 2456.940 ;
        RECT 1417.790 2456.880 1418.110 2456.940 ;
        RECT 1375.930 2456.740 1376.250 2456.800 ;
        RECT 1599.030 2456.740 1599.350 2456.800 ;
        RECT 1375.930 2456.600 1599.350 2456.740 ;
        RECT 1375.930 2456.540 1376.250 2456.600 ;
        RECT 1599.030 2456.540 1599.350 2456.600 ;
        RECT 1603.170 2454.700 1603.490 2454.760 ;
        RECT 1602.975 2454.560 1603.490 2454.700 ;
        RECT 1603.170 2454.500 1603.490 2454.560 ;
        RECT 1367.190 2449.940 1367.510 2450.000 ;
        RECT 1403.990 2449.940 1404.310 2450.000 ;
        RECT 1367.190 2449.800 1404.310 2449.940 ;
        RECT 1367.190 2449.740 1367.510 2449.800 ;
        RECT 1403.990 2449.740 1404.310 2449.800 ;
        RECT 1375.470 2449.600 1375.790 2449.660 ;
        RECT 1600.870 2449.600 1601.190 2449.660 ;
        RECT 1603.170 2449.600 1603.490 2449.660 ;
        RECT 1375.470 2449.460 1601.190 2449.600 ;
        RECT 1602.975 2449.460 1603.490 2449.600 ;
        RECT 1375.470 2449.400 1375.790 2449.460 ;
        RECT 1600.870 2449.400 1601.190 2449.460 ;
        RECT 1603.170 2449.400 1603.490 2449.460 ;
        RECT 1600.410 2449.260 1600.730 2449.320 ;
        RECT 1603.630 2449.260 1603.950 2449.320 ;
        RECT 1600.410 2449.120 1603.950 2449.260 ;
        RECT 1600.410 2449.060 1600.730 2449.120 ;
        RECT 1603.630 2449.060 1603.950 2449.120 ;
        RECT 1604.090 2449.260 1604.410 2449.320 ;
        RECT 1604.090 2449.120 1604.605 2449.260 ;
        RECT 1604.090 2449.060 1604.410 2449.120 ;
        RECT 1603.720 2448.580 1603.860 2449.060 ;
        RECT 1603.720 2448.440 1604.320 2448.580 ;
        RECT 1604.180 2447.280 1604.320 2448.440 ;
        RECT 1604.090 2447.020 1604.410 2447.280 ;
        RECT 1368.110 2443.480 1368.430 2443.540 ;
        RECT 1390.650 2443.480 1390.970 2443.540 ;
        RECT 1368.110 2443.340 1390.970 2443.480 ;
        RECT 1368.110 2443.280 1368.430 2443.340 ;
        RECT 1390.650 2443.280 1390.970 2443.340 ;
        RECT 1375.010 2443.140 1375.330 2443.200 ;
        RECT 1599.030 2443.140 1599.350 2443.200 ;
        RECT 1375.010 2443.000 1599.350 2443.140 ;
        RECT 1375.010 2442.940 1375.330 2443.000 ;
        RECT 1599.030 2442.940 1599.350 2443.000 ;
        RECT 1374.550 2442.800 1374.870 2442.860 ;
        RECT 1598.570 2442.800 1598.890 2442.860 ;
        RECT 1374.550 2442.660 1598.890 2442.800 ;
        RECT 1374.550 2442.600 1374.870 2442.660 ;
        RECT 1598.570 2442.600 1598.890 2442.660 ;
        RECT 1602.250 2436.340 1602.570 2436.400 ;
        RECT 1604.105 2436.340 1604.395 2436.385 ;
        RECT 1602.250 2436.200 1604.395 2436.340 ;
        RECT 1602.250 2436.140 1602.570 2436.200 ;
        RECT 1604.105 2436.155 1604.395 2436.200 ;
        RECT 1374.090 2436.000 1374.410 2436.060 ;
        RECT 1600.870 2436.000 1601.190 2436.060 ;
        RECT 1374.090 2435.860 1601.190 2436.000 ;
        RECT 1374.090 2435.800 1374.410 2435.860 ;
        RECT 1600.870 2435.800 1601.190 2435.860 ;
        RECT 1602.710 2431.040 1603.030 2431.300 ;
        RECT 1603.170 2431.040 1603.490 2431.300 ;
        RECT 1602.800 2430.280 1602.940 2431.040 ;
        RECT 1603.260 2430.280 1603.400 2431.040 ;
        RECT 1602.710 2430.020 1603.030 2430.280 ;
        RECT 1603.170 2430.020 1603.490 2430.280 ;
        RECT 1367.650 2429.540 1367.970 2429.600 ;
        RECT 1391.110 2429.540 1391.430 2429.600 ;
        RECT 1367.650 2429.400 1391.430 2429.540 ;
        RECT 1367.650 2429.340 1367.970 2429.400 ;
        RECT 1391.110 2429.340 1391.430 2429.400 ;
        RECT 1373.630 2429.200 1373.950 2429.260 ;
        RECT 1599.030 2429.200 1599.350 2429.260 ;
        RECT 1373.630 2429.060 1599.350 2429.200 ;
        RECT 1373.630 2429.000 1373.950 2429.060 ;
        RECT 1599.030 2429.000 1599.350 2429.060 ;
        RECT 1368.110 2422.400 1368.430 2422.460 ;
        RECT 1391.570 2422.400 1391.890 2422.460 ;
        RECT 1368.110 2422.260 1391.890 2422.400 ;
        RECT 1368.110 2422.200 1368.430 2422.260 ;
        RECT 1391.570 2422.200 1391.890 2422.260 ;
        RECT 1373.170 2422.060 1373.490 2422.120 ;
        RECT 1600.870 2422.060 1601.190 2422.120 ;
        RECT 1373.170 2421.920 1601.190 2422.060 ;
        RECT 1373.170 2421.860 1373.490 2421.920 ;
        RECT 1600.870 2421.860 1601.190 2421.920 ;
        RECT 1386.050 2415.260 1386.370 2415.320 ;
        RECT 1599.030 2415.260 1599.350 2415.320 ;
        RECT 1386.050 2415.120 1599.350 2415.260 ;
        RECT 1386.050 2415.060 1386.370 2415.120 ;
        RECT 1599.030 2415.060 1599.350 2415.120 ;
        RECT 1602.250 2414.240 1602.570 2414.300 ;
        RECT 1602.055 2414.100 1602.570 2414.240 ;
        RECT 1602.250 2414.040 1602.570 2414.100 ;
        RECT 1602.250 2413.560 1602.570 2413.620 ;
        RECT 1603.170 2413.560 1603.490 2413.620 ;
        RECT 1602.250 2413.420 1603.490 2413.560 ;
        RECT 1602.250 2413.360 1602.570 2413.420 ;
        RECT 1603.170 2413.360 1603.490 2413.420 ;
        RECT 1604.090 2413.360 1604.410 2413.620 ;
        RECT 1602.710 2411.860 1603.030 2411.920 ;
        RECT 1604.180 2411.860 1604.320 2413.360 ;
        RECT 1602.710 2411.720 1604.320 2411.860 ;
        RECT 1602.710 2411.660 1603.030 2411.720 ;
        RECT 1368.110 2408.800 1368.430 2408.860 ;
        RECT 1392.030 2408.800 1392.350 2408.860 ;
        RECT 1368.110 2408.660 1392.350 2408.800 ;
        RECT 1368.110 2408.600 1368.430 2408.660 ;
        RECT 1392.030 2408.600 1392.350 2408.660 ;
        RECT 1386.510 2408.460 1386.830 2408.520 ;
        RECT 1600.870 2408.460 1601.190 2408.520 ;
        RECT 1386.510 2408.320 1601.190 2408.460 ;
        RECT 1386.510 2408.260 1386.830 2408.320 ;
        RECT 1600.870 2408.260 1601.190 2408.320 ;
        RECT 1601.330 2402.340 1601.650 2402.400 ;
        RECT 1604.090 2402.340 1604.410 2402.400 ;
        RECT 1601.330 2402.200 1604.410 2402.340 ;
        RECT 1601.330 2402.140 1601.650 2402.200 ;
        RECT 1604.090 2402.140 1604.410 2402.200 ;
        RECT 1368.110 2401.660 1368.430 2401.720 ;
        RECT 1392.490 2401.660 1392.810 2401.720 ;
        RECT 1368.110 2401.520 1392.810 2401.660 ;
        RECT 1368.110 2401.460 1368.430 2401.520 ;
        RECT 1392.490 2401.460 1392.810 2401.520 ;
        RECT 1601.330 2401.660 1601.650 2401.720 ;
        RECT 1602.265 2401.660 1602.555 2401.705 ;
        RECT 1601.330 2401.520 1602.555 2401.660 ;
        RECT 1601.330 2401.460 1601.650 2401.520 ;
        RECT 1602.265 2401.475 1602.555 2401.520 ;
        RECT 1382.830 2401.320 1383.150 2401.380 ;
        RECT 1599.030 2401.320 1599.350 2401.380 ;
        RECT 1382.830 2401.180 1599.350 2401.320 ;
        RECT 1382.830 2401.120 1383.150 2401.180 ;
        RECT 1599.030 2401.120 1599.350 2401.180 ;
        RECT 1604.090 2397.240 1604.410 2397.300 ;
        RECT 1603.895 2397.100 1604.410 2397.240 ;
        RECT 1604.090 2397.040 1604.410 2397.100 ;
        RECT 1600.870 2396.560 1601.190 2396.620 ;
        RECT 1604.090 2396.560 1604.410 2396.620 ;
        RECT 1600.870 2396.420 1604.410 2396.560 ;
        RECT 1600.870 2396.360 1601.190 2396.420 ;
        RECT 1604.090 2396.360 1604.410 2396.420 ;
        RECT 1603.170 2394.860 1603.490 2394.920 ;
        RECT 1604.105 2394.860 1604.395 2394.905 ;
        RECT 1603.170 2394.720 1604.395 2394.860 ;
        RECT 1603.170 2394.660 1603.490 2394.720 ;
        RECT 1604.105 2394.675 1604.395 2394.720 ;
        RECT 1368.110 2394.520 1368.430 2394.580 ;
        RECT 1576.490 2394.520 1576.810 2394.580 ;
        RECT 1368.110 2394.380 1576.810 2394.520 ;
        RECT 1368.110 2394.320 1368.430 2394.380 ;
        RECT 1576.490 2394.320 1576.810 2394.380 ;
        RECT 1602.250 2385.000 1602.570 2385.060 ;
        RECT 1603.170 2385.000 1603.490 2385.060 ;
        RECT 1602.250 2384.860 1603.490 2385.000 ;
        RECT 1602.250 2384.800 1602.570 2384.860 ;
        RECT 1603.170 2384.800 1603.490 2384.860 ;
        RECT 1600.870 2384.120 1601.190 2384.380 ;
        RECT 1600.960 2383.300 1601.100 2384.120 ;
        RECT 1601.330 2383.300 1601.650 2383.360 ;
        RECT 1600.960 2383.160 1601.650 2383.300 ;
        RECT 1601.330 2383.100 1601.650 2383.160 ;
        RECT 1368.110 2380.580 1368.430 2380.640 ;
        RECT 1562.690 2380.580 1563.010 2380.640 ;
        RECT 1368.110 2380.440 1563.010 2380.580 ;
        RECT 1368.110 2380.380 1368.430 2380.440 ;
        RECT 1562.690 2380.380 1563.010 2380.440 ;
        RECT 1603.630 2380.240 1603.950 2380.300 ;
        RECT 1603.435 2380.100 1603.950 2380.240 ;
        RECT 1603.630 2380.040 1603.950 2380.100 ;
        RECT 1603.170 2379.360 1603.490 2379.620 ;
        RECT 1602.250 2379.220 1602.570 2379.280 ;
        RECT 1603.260 2379.220 1603.400 2379.360 ;
        RECT 1602.250 2379.080 1603.400 2379.220 ;
        RECT 1602.250 2379.020 1602.570 2379.080 ;
        RECT 1604.090 2378.880 1604.410 2378.940 ;
        RECT 1603.895 2378.740 1604.410 2378.880 ;
        RECT 1604.090 2378.680 1604.410 2378.740 ;
        RECT 1368.110 2374.120 1368.430 2374.180 ;
        RECT 1548.890 2374.120 1549.210 2374.180 ;
        RECT 1368.110 2373.980 1549.210 2374.120 ;
        RECT 1368.110 2373.920 1368.430 2373.980 ;
        RECT 1548.890 2373.920 1549.210 2373.980 ;
        RECT 1382.370 2373.780 1382.690 2373.840 ;
        RECT 1600.870 2373.780 1601.190 2373.840 ;
        RECT 1382.370 2373.640 1601.190 2373.780 ;
        RECT 1382.370 2373.580 1382.690 2373.640 ;
        RECT 1600.870 2373.580 1601.190 2373.640 ;
        RECT 1367.650 2370.040 1367.970 2370.100 ;
        RECT 1601.790 2370.040 1602.110 2370.100 ;
        RECT 1367.650 2369.900 1602.110 2370.040 ;
        RECT 1367.650 2369.840 1367.970 2369.900 ;
        RECT 1601.790 2369.840 1602.110 2369.900 ;
        RECT 1368.110 2366.980 1368.430 2367.040 ;
        RECT 1541.990 2366.980 1542.310 2367.040 ;
        RECT 1368.110 2366.840 1542.310 2366.980 ;
        RECT 1368.110 2366.780 1368.430 2366.840 ;
        RECT 1541.990 2366.780 1542.310 2366.840 ;
        RECT 1367.190 2360.180 1367.510 2360.240 ;
        RECT 1600.870 2360.180 1601.190 2360.240 ;
        RECT 1367.190 2360.040 1601.190 2360.180 ;
        RECT 1367.190 2359.980 1367.510 2360.040 ;
        RECT 1600.870 2359.980 1601.190 2360.040 ;
        RECT 1367.650 2353.380 1367.970 2353.440 ;
        RECT 1528.190 2353.380 1528.510 2353.440 ;
        RECT 1367.650 2353.240 1528.510 2353.380 ;
        RECT 1367.650 2353.180 1367.970 2353.240 ;
        RECT 1528.190 2353.180 1528.510 2353.240 ;
        RECT 1366.730 2353.040 1367.050 2353.100 ;
        RECT 1601.330 2353.040 1601.650 2353.100 ;
        RECT 1366.730 2352.900 1601.650 2353.040 ;
        RECT 1366.730 2352.840 1367.050 2352.900 ;
        RECT 1601.330 2352.840 1601.650 2352.900 ;
        RECT 1601.330 2352.360 1601.650 2352.420 ;
        RECT 1603.645 2352.360 1603.935 2352.405 ;
        RECT 1601.330 2352.220 1603.935 2352.360 ;
        RECT 1601.330 2352.160 1601.650 2352.220 ;
        RECT 1603.645 2352.175 1603.935 2352.220 ;
        RECT 1367.650 2346.580 1367.970 2346.640 ;
        RECT 1521.290 2346.580 1521.610 2346.640 ;
        RECT 1367.650 2346.440 1521.610 2346.580 ;
        RECT 1367.650 2346.380 1367.970 2346.440 ;
        RECT 1521.290 2346.380 1521.610 2346.440 ;
        RECT 1381.910 2346.240 1382.230 2346.300 ;
        RECT 1601.790 2346.240 1602.110 2346.300 ;
        RECT 1381.910 2346.100 1602.110 2346.240 ;
        RECT 1381.910 2346.040 1382.230 2346.100 ;
        RECT 1601.790 2346.040 1602.110 2346.100 ;
        RECT 1381.450 2339.780 1381.770 2339.840 ;
        RECT 1602.250 2339.780 1602.570 2339.840 ;
        RECT 1381.450 2339.640 1602.570 2339.780 ;
        RECT 1381.450 2339.580 1381.770 2339.640 ;
        RECT 1602.250 2339.580 1602.570 2339.640 ;
        RECT 1380.990 2339.440 1381.310 2339.500 ;
        RECT 1601.330 2339.440 1601.650 2339.500 ;
        RECT 1380.990 2339.300 1601.650 2339.440 ;
        RECT 1380.990 2339.240 1381.310 2339.300 ;
        RECT 1601.330 2339.240 1601.650 2339.300 ;
        RECT 1601.805 2339.100 1602.095 2339.145 ;
        RECT 1602.710 2339.100 1603.030 2339.160 ;
        RECT 1601.805 2338.960 1603.030 2339.100 ;
        RECT 1601.805 2338.915 1602.095 2338.960 ;
        RECT 1602.710 2338.900 1603.030 2338.960 ;
        RECT 1601.330 2338.760 1601.650 2338.820 ;
        RECT 1603.630 2338.760 1603.950 2338.820 ;
        RECT 1601.330 2338.620 1603.950 2338.760 ;
        RECT 1601.330 2338.560 1601.650 2338.620 ;
        RECT 1603.630 2338.560 1603.950 2338.620 ;
        RECT 1600.410 2338.420 1600.730 2338.480 ;
        RECT 1602.710 2338.420 1603.030 2338.480 ;
        RECT 1600.410 2338.280 1603.030 2338.420 ;
        RECT 1600.410 2338.220 1600.730 2338.280 ;
        RECT 1602.710 2338.220 1603.030 2338.280 ;
        RECT 1601.790 2338.080 1602.110 2338.140 ;
        RECT 1601.595 2337.940 1602.110 2338.080 ;
        RECT 1601.790 2337.880 1602.110 2337.940 ;
        RECT 1603.170 2337.740 1603.490 2337.800 ;
        RECT 1603.645 2337.740 1603.935 2337.785 ;
        RECT 1603.170 2337.600 1603.935 2337.740 ;
        RECT 1603.170 2337.540 1603.490 2337.600 ;
        RECT 1603.645 2337.555 1603.935 2337.600 ;
        RECT 1603.630 2337.060 1603.950 2337.120 ;
        RECT 1604.105 2337.060 1604.395 2337.105 ;
        RECT 1603.630 2336.920 1604.395 2337.060 ;
        RECT 1603.630 2336.860 1603.950 2336.920 ;
        RECT 1604.105 2336.875 1604.395 2336.920 ;
        RECT 1367.650 2332.640 1367.970 2332.700 ;
        RECT 1514.850 2332.640 1515.170 2332.700 ;
        RECT 1367.650 2332.500 1515.170 2332.640 ;
        RECT 1367.650 2332.440 1367.970 2332.500 ;
        RECT 1514.850 2332.440 1515.170 2332.500 ;
        RECT 1380.530 2332.300 1380.850 2332.360 ;
        RECT 1600.870 2332.300 1601.190 2332.360 ;
        RECT 1380.530 2332.160 1601.190 2332.300 ;
        RECT 1380.530 2332.100 1380.850 2332.160 ;
        RECT 1600.870 2332.100 1601.190 2332.160 ;
        RECT 1380.070 2325.500 1380.390 2325.560 ;
        RECT 1600.870 2325.500 1601.190 2325.560 ;
        RECT 1380.070 2325.360 1601.190 2325.500 ;
        RECT 1380.070 2325.300 1380.390 2325.360 ;
        RECT 1600.870 2325.300 1601.190 2325.360 ;
        RECT 1366.270 2318.700 1366.590 2318.760 ;
        RECT 1385.590 2318.700 1385.910 2318.760 ;
        RECT 1366.270 2318.560 1385.910 2318.700 ;
        RECT 1366.270 2318.500 1366.590 2318.560 ;
        RECT 1385.590 2318.500 1385.910 2318.560 ;
        RECT 1366.270 2304.760 1366.590 2304.820 ;
        RECT 1393.410 2304.760 1393.730 2304.820 ;
        RECT 1366.270 2304.620 1393.730 2304.760 ;
        RECT 1366.270 2304.560 1366.590 2304.620 ;
        RECT 1393.410 2304.560 1393.730 2304.620 ;
        RECT 1366.270 2300.340 1366.590 2300.400 ;
        RECT 1380.070 2300.340 1380.390 2300.400 ;
        RECT 1366.270 2300.200 1380.390 2300.340 ;
        RECT 1366.270 2300.140 1366.590 2300.200 ;
        RECT 1380.070 2300.140 1380.390 2300.200 ;
        RECT 1366.270 2290.820 1366.590 2290.880 ;
        RECT 1380.530 2290.820 1380.850 2290.880 ;
        RECT 1366.270 2290.680 1380.850 2290.820 ;
        RECT 1366.270 2290.620 1366.590 2290.680 ;
        RECT 1380.530 2290.620 1380.850 2290.680 ;
        RECT 1601.345 2287.420 1601.635 2287.465 ;
        RECT 1602.250 2287.420 1602.570 2287.480 ;
        RECT 1601.345 2287.280 1602.570 2287.420 ;
        RECT 1601.345 2287.235 1601.635 2287.280 ;
        RECT 1602.250 2287.220 1602.570 2287.280 ;
        RECT 1603.170 2287.420 1603.490 2287.480 ;
        RECT 1603.645 2287.420 1603.935 2287.465 ;
        RECT 1603.170 2287.280 1603.935 2287.420 ;
        RECT 1603.170 2287.220 1603.490 2287.280 ;
        RECT 1603.645 2287.235 1603.935 2287.280 ;
        RECT 1603.185 2286.740 1603.475 2286.785 ;
        RECT 1604.090 2286.740 1604.410 2286.800 ;
        RECT 1603.185 2286.600 1604.410 2286.740 ;
        RECT 1603.185 2286.555 1603.475 2286.600 ;
        RECT 1604.090 2286.540 1604.410 2286.600 ;
        RECT 1600.870 2285.520 1601.190 2285.780 ;
        RECT 1600.960 2284.360 1601.100 2285.520 ;
        RECT 1601.790 2284.700 1602.110 2284.760 ;
        RECT 1601.595 2284.560 1602.110 2284.700 ;
        RECT 1601.790 2284.500 1602.110 2284.560 ;
        RECT 1603.630 2284.700 1603.950 2284.760 ;
        RECT 1604.105 2284.700 1604.395 2284.745 ;
        RECT 1603.630 2284.560 1604.395 2284.700 ;
        RECT 1603.630 2284.500 1603.950 2284.560 ;
        RECT 1604.105 2284.515 1604.395 2284.560 ;
        RECT 1600.960 2284.220 1603.860 2284.360 ;
        RECT 1601.790 2283.340 1602.110 2283.400 ;
        RECT 1601.595 2283.200 1602.110 2283.340 ;
        RECT 1601.790 2283.140 1602.110 2283.200 ;
        RECT 1602.250 2283.340 1602.570 2283.400 ;
        RECT 1603.720 2283.340 1603.860 2284.220 ;
        RECT 1602.250 2283.200 1603.860 2283.340 ;
        RECT 1602.250 2283.140 1602.570 2283.200 ;
        RECT 1603.170 2282.660 1603.490 2282.720 ;
        RECT 1604.105 2282.660 1604.395 2282.705 ;
        RECT 1603.170 2282.520 1604.395 2282.660 ;
        RECT 1603.170 2282.460 1603.490 2282.520 ;
        RECT 1604.105 2282.475 1604.395 2282.520 ;
        RECT 1366.270 2281.300 1366.590 2281.360 ;
        RECT 1380.990 2281.300 1381.310 2281.360 ;
        RECT 1366.270 2281.160 1381.310 2281.300 ;
        RECT 1366.270 2281.100 1366.590 2281.160 ;
        RECT 1380.990 2281.100 1381.310 2281.160 ;
        RECT 1366.270 2271.780 1366.590 2271.840 ;
        RECT 1381.450 2271.780 1381.770 2271.840 ;
        RECT 1366.270 2271.640 1381.770 2271.780 ;
        RECT 1366.270 2271.580 1366.590 2271.640 ;
        RECT 1381.450 2271.580 1381.770 2271.640 ;
        RECT 1603.185 2263.280 1603.475 2263.325 ;
        RECT 1604.105 2263.280 1604.395 2263.325 ;
        RECT 1603.185 2263.140 1604.395 2263.280 ;
        RECT 1603.185 2263.095 1603.475 2263.140 ;
        RECT 1604.105 2263.095 1604.395 2263.140 ;
        RECT 1366.270 2262.260 1366.590 2262.320 ;
        RECT 1381.910 2262.260 1382.230 2262.320 ;
        RECT 1366.270 2262.120 1382.230 2262.260 ;
        RECT 1366.270 2262.060 1366.590 2262.120 ;
        RECT 1381.910 2262.060 1382.230 2262.120 ;
        RECT 1600.870 2261.580 1601.190 2261.640 ;
        RECT 1600.675 2261.440 1601.190 2261.580 ;
        RECT 1600.870 2261.380 1601.190 2261.440 ;
        RECT 1603.170 2249.340 1603.490 2249.400 ;
        RECT 1602.975 2249.200 1603.490 2249.340 ;
        RECT 1603.170 2249.140 1603.490 2249.200 ;
        RECT 1601.790 2236.760 1602.110 2236.820 ;
        RECT 1601.595 2236.620 1602.110 2236.760 ;
        RECT 1601.790 2236.560 1602.110 2236.620 ;
        RECT 1602.250 2236.560 1602.570 2236.820 ;
        RECT 1602.710 2236.560 1603.030 2236.820 ;
        RECT 1602.340 2236.140 1602.480 2236.560 ;
        RECT 1602.800 2236.140 1602.940 2236.560 ;
        RECT 1602.250 2235.880 1602.570 2236.140 ;
        RECT 1602.710 2235.880 1603.030 2236.140 ;
        RECT 1603.170 2235.740 1603.490 2235.800 ;
        RECT 1603.645 2235.740 1603.935 2235.785 ;
        RECT 1603.170 2235.600 1603.935 2235.740 ;
        RECT 1603.170 2235.540 1603.490 2235.600 ;
        RECT 1603.645 2235.555 1603.935 2235.600 ;
        RECT 1367.190 2235.400 1367.510 2235.460 ;
        RECT 1604.105 2235.400 1604.395 2235.445 ;
        RECT 1367.190 2235.260 1604.395 2235.400 ;
        RECT 1367.190 2235.200 1367.510 2235.260 ;
        RECT 1604.105 2235.215 1604.395 2235.260 ;
        RECT 1601.790 2235.060 1602.110 2235.120 ;
        RECT 1601.595 2234.920 1602.110 2235.060 ;
        RECT 1601.790 2234.860 1602.110 2234.920 ;
        RECT 1603.185 2234.720 1603.475 2234.765 ;
        RECT 1604.090 2234.720 1604.410 2234.780 ;
        RECT 1603.185 2234.580 1604.410 2234.720 ;
        RECT 1603.185 2234.535 1603.475 2234.580 ;
        RECT 1604.090 2234.520 1604.410 2234.580 ;
        RECT 1601.345 2234.380 1601.635 2234.425 ;
        RECT 1603.630 2234.380 1603.950 2234.440 ;
        RECT 1601.345 2234.240 1603.950 2234.380 ;
        RECT 1601.345 2234.195 1601.635 2234.240 ;
        RECT 1603.630 2234.180 1603.950 2234.240 ;
        RECT 1600.885 2234.040 1601.175 2234.085 ;
        RECT 1604.090 2234.040 1604.410 2234.100 ;
        RECT 1600.885 2233.900 1604.410 2234.040 ;
        RECT 1600.885 2233.855 1601.175 2233.900 ;
        RECT 1604.090 2233.840 1604.410 2233.900 ;
        RECT 1367.190 2224.180 1367.510 2224.240 ;
        RECT 1382.370 2224.180 1382.690 2224.240 ;
        RECT 1367.190 2224.040 1382.690 2224.180 ;
        RECT 1367.190 2223.980 1367.510 2224.040 ;
        RECT 1382.370 2223.980 1382.690 2224.040 ;
        RECT 1367.190 2214.660 1367.510 2214.720 ;
        RECT 1382.830 2214.660 1383.150 2214.720 ;
        RECT 1367.190 2214.520 1383.150 2214.660 ;
        RECT 1367.190 2214.460 1367.510 2214.520 ;
        RECT 1382.830 2214.460 1383.150 2214.520 ;
        RECT 1602.710 2212.080 1603.030 2212.340 ;
        RECT 1603.630 2212.080 1603.950 2212.340 ;
        RECT 1602.800 2210.980 1602.940 2212.080 ;
        RECT 1602.710 2210.720 1603.030 2210.980 ;
        RECT 1602.250 2210.240 1602.570 2210.300 ;
        RECT 1603.720 2210.240 1603.860 2212.080 ;
        RECT 1602.250 2210.100 1603.860 2210.240 ;
        RECT 1602.250 2210.040 1602.570 2210.100 ;
        RECT 1367.190 2206.500 1367.510 2206.560 ;
        RECT 1386.510 2206.500 1386.830 2206.560 ;
        RECT 1367.190 2206.360 1386.830 2206.500 ;
        RECT 1367.190 2206.300 1367.510 2206.360 ;
        RECT 1386.510 2206.300 1386.830 2206.360 ;
      LAYER met1 ;
        RECT 1605.000 2205.000 2051.235 2581.480 ;
      LAYER met1 ;
        RECT 1367.190 2198.680 1367.510 2198.740 ;
        RECT 1386.050 2198.680 1386.370 2198.740 ;
        RECT 1367.190 2198.540 1386.370 2198.680 ;
        RECT 1367.190 2198.480 1367.510 2198.540 ;
        RECT 1386.050 2198.480 1386.370 2198.540 ;
        RECT 1366.270 2167.060 1366.590 2167.120 ;
        RECT 1374.090 2167.060 1374.410 2167.120 ;
        RECT 1366.270 2166.920 1374.410 2167.060 ;
        RECT 1366.270 2166.860 1366.590 2166.920 ;
        RECT 1374.090 2166.860 1374.410 2166.920 ;
        RECT 1601.330 2159.920 1601.650 2159.980 ;
        RECT 1604.090 2159.920 1604.410 2159.980 ;
        RECT 1601.330 2159.780 1604.410 2159.920 ;
        RECT 1601.330 2159.720 1601.650 2159.780 ;
        RECT 1604.090 2159.720 1604.410 2159.780 ;
        RECT 1366.270 2157.540 1366.590 2157.600 ;
        RECT 1374.550 2157.540 1374.870 2157.600 ;
        RECT 1366.270 2157.400 1374.870 2157.540 ;
        RECT 1366.270 2157.340 1366.590 2157.400 ;
        RECT 1374.550 2157.340 1374.870 2157.400 ;
        RECT 1366.270 2148.020 1366.590 2148.080 ;
        RECT 1375.010 2148.020 1375.330 2148.080 ;
        RECT 1366.270 2147.880 1375.330 2148.020 ;
        RECT 1366.270 2147.820 1366.590 2147.880 ;
        RECT 1375.010 2147.820 1375.330 2147.880 ;
        RECT 1601.330 2138.840 1601.650 2138.900 ;
        RECT 1604.090 2138.840 1604.410 2138.900 ;
        RECT 1601.330 2138.700 1604.410 2138.840 ;
        RECT 1601.330 2138.640 1601.650 2138.700 ;
        RECT 1604.090 2138.640 1604.410 2138.700 ;
        RECT 1366.270 2138.500 1366.590 2138.560 ;
        RECT 1375.470 2138.500 1375.790 2138.560 ;
        RECT 1366.270 2138.360 1375.790 2138.500 ;
        RECT 1366.270 2138.300 1366.590 2138.360 ;
        RECT 1375.470 2138.300 1375.790 2138.360 ;
        RECT 1366.270 2128.980 1366.590 2129.040 ;
        RECT 1375.930 2128.980 1376.250 2129.040 ;
        RECT 1366.270 2128.840 1376.250 2128.980 ;
        RECT 1366.270 2128.780 1366.590 2128.840 ;
        RECT 1375.930 2128.780 1376.250 2128.840 ;
        RECT 1367.190 2120.140 1367.510 2120.200 ;
        RECT 1379.610 2120.140 1379.930 2120.200 ;
        RECT 1367.190 2120.000 1379.930 2120.140 ;
        RECT 1367.190 2119.940 1367.510 2120.000 ;
        RECT 1379.610 2119.940 1379.930 2120.000 ;
        RECT 1367.190 2110.280 1367.510 2110.340 ;
        RECT 1379.150 2110.280 1379.470 2110.340 ;
        RECT 1367.190 2110.140 1379.470 2110.280 ;
        RECT 1367.190 2110.080 1367.510 2110.140 ;
        RECT 1379.150 2110.080 1379.470 2110.140 ;
        RECT 1367.190 2100.420 1367.510 2100.480 ;
        RECT 1378.690 2100.420 1379.010 2100.480 ;
        RECT 1367.190 2100.280 1379.010 2100.420 ;
        RECT 1367.190 2100.220 1367.510 2100.280 ;
        RECT 1378.690 2100.220 1379.010 2100.280 ;
        RECT 1367.190 2090.560 1367.510 2090.620 ;
        RECT 1397.550 2090.560 1397.870 2090.620 ;
        RECT 1367.190 2090.420 1397.870 2090.560 ;
        RECT 1367.190 2090.360 1367.510 2090.420 ;
        RECT 1397.550 2090.360 1397.870 2090.420 ;
        RECT 1367.190 2081.380 1367.510 2081.440 ;
        RECT 1392.950 2081.380 1393.270 2081.440 ;
        RECT 1367.190 2081.240 1393.270 2081.380 ;
        RECT 1367.190 2081.180 1367.510 2081.240 ;
        RECT 1392.950 2081.180 1393.270 2081.240 ;
        RECT 1367.190 2071.860 1367.510 2071.920 ;
        RECT 1385.130 2071.860 1385.450 2071.920 ;
        RECT 1367.190 2071.720 1385.450 2071.860 ;
        RECT 1367.190 2071.660 1367.510 2071.720 ;
        RECT 1385.130 2071.660 1385.450 2071.720 ;
        RECT 1367.190 2062.340 1367.510 2062.400 ;
        RECT 1384.670 2062.340 1384.990 2062.400 ;
        RECT 1367.190 2062.200 1384.990 2062.340 ;
        RECT 1367.190 2062.140 1367.510 2062.200 ;
        RECT 1384.670 2062.140 1384.990 2062.200 ;
        RECT 1367.190 2052.820 1367.510 2052.880 ;
        RECT 1384.210 2052.820 1384.530 2052.880 ;
        RECT 1367.190 2052.680 1384.530 2052.820 ;
        RECT 1367.190 2052.620 1367.510 2052.680 ;
        RECT 1384.210 2052.620 1384.530 2052.680 ;
        RECT 1367.190 2043.300 1367.510 2043.360 ;
        RECT 1383.750 2043.300 1384.070 2043.360 ;
        RECT 1367.190 2043.160 1384.070 2043.300 ;
        RECT 1367.190 2043.100 1367.510 2043.160 ;
        RECT 1383.750 2043.100 1384.070 2043.160 ;
        RECT 1367.190 2033.780 1367.510 2033.840 ;
        RECT 1383.290 2033.780 1383.610 2033.840 ;
        RECT 1367.190 2033.640 1383.610 2033.780 ;
        RECT 1367.190 2033.580 1367.510 2033.640 ;
        RECT 1383.290 2033.580 1383.610 2033.640 ;
        RECT 1367.190 2014.740 1367.510 2014.800 ;
        RECT 1378.230 2014.740 1378.550 2014.800 ;
        RECT 1367.190 2014.600 1378.550 2014.740 ;
        RECT 1367.190 2014.540 1367.510 2014.600 ;
        RECT 1378.230 2014.540 1378.550 2014.600 ;
        RECT 1367.190 2005.220 1367.510 2005.280 ;
        RECT 1377.770 2005.220 1378.090 2005.280 ;
        RECT 1367.190 2005.080 1378.090 2005.220 ;
        RECT 1367.190 2005.020 1367.510 2005.080 ;
        RECT 1377.770 2005.020 1378.090 2005.080 ;
        RECT 1367.190 2000.800 1367.510 2000.860 ;
        RECT 1603.630 2000.800 1603.950 2000.860 ;
        RECT 1367.190 2000.660 1603.950 2000.800 ;
        RECT 1367.190 2000.600 1367.510 2000.660 ;
        RECT 1603.630 2000.600 1603.950 2000.660 ;
        RECT 1600.870 1994.340 1601.190 1994.400 ;
        RECT 1604.090 1994.340 1604.410 1994.400 ;
        RECT 1600.870 1994.200 1604.410 1994.340 ;
        RECT 1600.870 1994.140 1601.190 1994.200 ;
        RECT 1604.090 1994.140 1604.410 1994.200 ;
        RECT 1367.190 1987.200 1367.510 1987.260 ;
        RECT 1603.170 1987.200 1603.490 1987.260 ;
        RECT 1367.190 1987.060 1603.490 1987.200 ;
        RECT 1367.190 1987.000 1367.510 1987.060 ;
        RECT 1603.170 1987.000 1603.490 1987.060 ;
        RECT 1366.270 1984.140 1366.590 1984.200 ;
        RECT 1693.330 1984.140 1693.650 1984.200 ;
        RECT 1366.270 1984.000 1693.650 1984.140 ;
        RECT 1366.270 1983.940 1366.590 1984.000 ;
        RECT 1693.330 1983.940 1693.650 1984.000 ;
        RECT 1378.690 1983.800 1379.010 1983.860 ;
        RECT 1987.270 1983.800 1987.590 1983.860 ;
        RECT 1378.690 1983.660 1987.590 1983.800 ;
        RECT 1378.690 1983.600 1379.010 1983.660 ;
        RECT 1987.270 1983.600 1987.590 1983.660 ;
        RECT 1379.610 1983.460 1379.930 1983.520 ;
        RECT 1994.170 1983.460 1994.490 1983.520 ;
        RECT 1379.610 1983.320 1994.490 1983.460 ;
        RECT 1379.610 1983.260 1379.930 1983.320 ;
        RECT 1994.170 1983.260 1994.490 1983.320 ;
        RECT 1375.930 1983.120 1376.250 1983.180 ;
        RECT 2001.070 1983.120 2001.390 1983.180 ;
        RECT 1375.930 1982.980 2001.390 1983.120 ;
        RECT 1375.930 1982.920 1376.250 1982.980 ;
        RECT 2001.070 1982.920 2001.390 1982.980 ;
        RECT 1375.470 1982.780 1375.790 1982.840 ;
        RECT 2007.970 1982.780 2008.290 1982.840 ;
        RECT 1375.470 1982.640 2008.290 1982.780 ;
        RECT 1375.470 1982.580 1375.790 1982.640 ;
        RECT 2007.970 1982.580 2008.290 1982.640 ;
        RECT 1375.010 1982.440 1375.330 1982.500 ;
        RECT 2016.710 1982.440 2017.030 1982.500 ;
        RECT 1375.010 1982.300 2017.030 1982.440 ;
        RECT 1375.010 1982.240 1375.330 1982.300 ;
        RECT 2016.710 1982.240 2017.030 1982.300 ;
        RECT 1374.550 1982.100 1374.870 1982.160 ;
        RECT 2021.770 1982.100 2022.090 1982.160 ;
        RECT 1374.550 1981.960 2022.090 1982.100 ;
        RECT 1374.550 1981.900 1374.870 1981.960 ;
        RECT 2021.770 1981.900 2022.090 1981.960 ;
        RECT 2030.050 1981.900 2030.370 1982.160 ;
        RECT 1374.090 1981.760 1374.410 1981.820 ;
        RECT 2030.140 1981.760 2030.280 1981.900 ;
        RECT 1374.090 1981.620 2030.280 1981.760 ;
        RECT 1374.090 1981.560 1374.410 1981.620 ;
        RECT 1367.190 1980.060 1367.510 1980.120 ;
        RECT 1602.710 1980.060 1603.030 1980.120 ;
        RECT 1367.190 1979.920 1603.030 1980.060 ;
        RECT 1367.190 1979.860 1367.510 1979.920 ;
        RECT 1602.710 1979.860 1603.030 1979.920 ;
        RECT 1367.190 1973.260 1367.510 1973.320 ;
        RECT 1602.250 1973.260 1602.570 1973.320 ;
        RECT 1367.190 1973.120 1602.570 1973.260 ;
        RECT 1367.190 1973.060 1367.510 1973.120 ;
        RECT 1602.250 1973.060 1602.570 1973.120 ;
        RECT 1379.150 1960.340 1379.470 1960.400 ;
        RECT 1600.870 1960.340 1601.190 1960.400 ;
        RECT 1379.150 1960.200 1601.190 1960.340 ;
        RECT 1379.150 1960.140 1379.470 1960.200 ;
        RECT 1600.870 1960.140 1601.190 1960.200 ;
        RECT 1377.770 1960.000 1378.090 1960.060 ;
        RECT 1601.330 1960.000 1601.650 1960.060 ;
        RECT 1377.770 1959.860 1601.650 1960.000 ;
        RECT 1377.770 1959.800 1378.090 1959.860 ;
        RECT 1601.330 1959.800 1601.650 1959.860 ;
        RECT 1367.190 1959.660 1367.510 1959.720 ;
        RECT 1601.790 1959.660 1602.110 1959.720 ;
        RECT 1367.190 1959.520 1602.110 1959.660 ;
        RECT 1367.190 1959.460 1367.510 1959.520 ;
        RECT 1601.790 1959.460 1602.110 1959.520 ;
        RECT 1378.230 1952.860 1378.550 1952.920 ;
        RECT 1600.410 1952.860 1600.730 1952.920 ;
        RECT 1378.230 1952.720 1600.730 1952.860 ;
        RECT 1378.230 1952.660 1378.550 1952.720 ;
        RECT 1600.410 1952.660 1600.730 1952.720 ;
        RECT 1367.650 1952.520 1367.970 1952.580 ;
        RECT 1600.870 1952.520 1601.190 1952.580 ;
        RECT 1367.650 1952.380 1601.190 1952.520 ;
        RECT 1367.650 1952.320 1367.970 1952.380 ;
        RECT 1600.870 1952.320 1601.190 1952.380 ;
        RECT 1367.190 1946.060 1367.510 1946.120 ;
        RECT 1601.330 1946.060 1601.650 1946.120 ;
        RECT 1367.190 1945.920 1601.650 1946.060 ;
        RECT 1367.190 1945.860 1367.510 1945.920 ;
        RECT 1601.330 1945.860 1601.650 1945.920 ;
        RECT 1366.730 1940.280 1367.050 1940.340 ;
        RECT 1367.650 1940.280 1367.970 1940.340 ;
        RECT 1366.730 1940.140 1367.970 1940.280 ;
        RECT 1366.730 1940.080 1367.050 1940.140 ;
        RECT 1367.650 1940.080 1367.970 1940.140 ;
        RECT 1600.870 1939.260 1601.190 1939.320 ;
        RECT 1367.740 1939.120 1601.190 1939.260 ;
        RECT 1367.740 1937.900 1367.880 1939.120 ;
        RECT 1600.870 1939.060 1601.190 1939.120 ;
        RECT 1368.110 1938.920 1368.430 1938.980 ;
        RECT 1604.090 1938.920 1604.410 1938.980 ;
        RECT 1368.110 1938.780 1604.410 1938.920 ;
        RECT 1368.110 1938.720 1368.430 1938.780 ;
        RECT 1604.090 1938.720 1604.410 1938.780 ;
        RECT 1393.410 1938.580 1393.730 1938.640 ;
        RECT 1601.790 1938.580 1602.110 1938.640 ;
        RECT 1393.410 1938.440 1602.110 1938.580 ;
        RECT 1393.410 1938.380 1393.730 1938.440 ;
        RECT 1601.790 1938.380 1602.110 1938.440 ;
        RECT 1368.110 1937.900 1368.430 1937.960 ;
        RECT 1367.740 1937.760 1368.430 1937.900 ;
        RECT 1368.110 1937.700 1368.430 1937.760 ;
        RECT 1385.590 1931.780 1385.910 1931.840 ;
        RECT 1601.330 1931.780 1601.650 1931.840 ;
        RECT 1385.590 1931.640 1601.650 1931.780 ;
        RECT 1385.590 1931.580 1385.910 1931.640 ;
        RECT 1601.330 1931.580 1601.650 1931.640 ;
        RECT 1366.730 1924.980 1367.050 1925.040 ;
        RECT 1600.870 1924.980 1601.190 1925.040 ;
        RECT 1366.730 1924.840 1601.190 1924.980 ;
        RECT 1366.730 1924.780 1367.050 1924.840 ;
        RECT 1600.870 1924.780 1601.190 1924.840 ;
        RECT 1514.850 1924.640 1515.170 1924.700 ;
        RECT 1601.790 1924.640 1602.110 1924.700 ;
        RECT 1514.850 1924.500 1602.110 1924.640 ;
        RECT 1514.850 1924.440 1515.170 1924.500 ;
        RECT 1601.790 1924.440 1602.110 1924.500 ;
        RECT 1521.290 1918.180 1521.610 1918.240 ;
        RECT 1600.870 1918.180 1601.190 1918.240 ;
        RECT 1521.290 1918.040 1601.190 1918.180 ;
        RECT 1521.290 1917.980 1521.610 1918.040 ;
        RECT 1600.870 1917.980 1601.190 1918.040 ;
        RECT 1366.730 1917.640 1367.050 1917.900 ;
        RECT 1366.820 1916.820 1366.960 1917.640 ;
        RECT 1367.190 1916.820 1367.510 1916.880 ;
        RECT 1366.820 1916.680 1367.510 1916.820 ;
        RECT 1367.190 1916.620 1367.510 1916.680 ;
        RECT 1528.190 1911.040 1528.510 1911.100 ;
        RECT 1602.710 1911.040 1603.030 1911.100 ;
        RECT 1528.190 1910.900 1603.030 1911.040 ;
        RECT 1528.190 1910.840 1528.510 1910.900 ;
        RECT 1602.710 1910.840 1603.030 1910.900 ;
        RECT 1603.170 1906.960 1603.490 1907.020 ;
        RECT 1603.645 1906.960 1603.935 1907.005 ;
        RECT 1603.170 1906.820 1603.935 1906.960 ;
        RECT 1603.170 1906.760 1603.490 1906.820 ;
        RECT 1603.645 1906.775 1603.935 1906.820 ;
        RECT 1541.990 1904.240 1542.310 1904.300 ;
        RECT 1600.870 1904.240 1601.190 1904.300 ;
        RECT 1541.990 1904.100 1601.190 1904.240 ;
        RECT 1541.990 1904.040 1542.310 1904.100 ;
        RECT 1600.870 1904.040 1601.190 1904.100 ;
        RECT 1604.090 1901.520 1604.410 1901.580 ;
        RECT 1603.895 1901.380 1604.410 1901.520 ;
        RECT 1604.090 1901.320 1604.410 1901.380 ;
        RECT 1367.650 1901.180 1367.970 1901.240 ;
        RECT 1600.410 1901.180 1600.730 1901.240 ;
        RECT 1367.650 1901.040 1600.730 1901.180 ;
        RECT 1367.650 1900.980 1367.970 1901.040 ;
        RECT 1600.410 1900.980 1600.730 1901.040 ;
        RECT 1368.110 1900.840 1368.430 1900.900 ;
        RECT 1602.250 1900.840 1602.570 1900.900 ;
        RECT 1368.110 1900.700 1602.570 1900.840 ;
        RECT 1368.110 1900.640 1368.430 1900.700 ;
        RECT 1602.250 1900.640 1602.570 1900.700 ;
        RECT 1603.170 1898.800 1603.490 1898.860 ;
        RECT 1602.975 1898.660 1603.490 1898.800 ;
        RECT 1603.170 1898.600 1603.490 1898.660 ;
        RECT 1603.630 1897.780 1603.950 1897.840 ;
        RECT 1603.435 1897.640 1603.950 1897.780 ;
        RECT 1603.630 1897.580 1603.950 1897.640 ;
        RECT 1548.890 1897.440 1549.210 1897.500 ;
        RECT 1601.330 1897.440 1601.650 1897.500 ;
        RECT 1548.890 1897.300 1601.650 1897.440 ;
        RECT 1548.890 1897.240 1549.210 1897.300 ;
        RECT 1601.330 1897.240 1601.650 1897.300 ;
        RECT 1367.650 1894.720 1367.970 1894.780 ;
        RECT 1372.250 1894.720 1372.570 1894.780 ;
        RECT 1367.650 1894.580 1372.570 1894.720 ;
        RECT 1367.650 1894.520 1367.970 1894.580 ;
        RECT 1372.250 1894.520 1372.570 1894.580 ;
        RECT 1373.170 1894.380 1373.490 1894.440 ;
        RECT 1601.790 1894.380 1602.110 1894.440 ;
        RECT 1373.170 1894.240 1602.110 1894.380 ;
        RECT 1373.170 1894.180 1373.490 1894.240 ;
        RECT 1601.790 1894.180 1602.110 1894.240 ;
        RECT 1372.250 1894.040 1372.570 1894.100 ;
        RECT 1604.090 1894.040 1604.410 1894.100 ;
        RECT 1372.250 1893.900 1604.410 1894.040 ;
        RECT 1372.250 1893.840 1372.570 1893.900 ;
        RECT 1604.090 1893.840 1604.410 1893.900 ;
        RECT 1602.710 1891.660 1603.030 1891.720 ;
        RECT 1603.185 1891.660 1603.475 1891.705 ;
        RECT 1602.710 1891.520 1603.475 1891.660 ;
        RECT 1602.710 1891.460 1603.030 1891.520 ;
        RECT 1603.185 1891.475 1603.475 1891.520 ;
        RECT 1576.490 1884.180 1576.810 1884.240 ;
        RECT 1599.950 1884.180 1600.270 1884.240 ;
        RECT 1576.490 1884.040 1600.270 1884.180 ;
        RECT 1576.490 1883.980 1576.810 1884.040 ;
        RECT 1599.950 1883.980 1600.270 1884.040 ;
        RECT 1490.485 1883.840 1490.775 1883.885 ;
        RECT 1514.405 1883.840 1514.695 1883.885 ;
        RECT 1490.485 1883.700 1514.695 1883.840 ;
        RECT 1490.485 1883.655 1490.775 1883.700 ;
        RECT 1514.405 1883.655 1514.695 1883.700 ;
        RECT 1562.690 1883.840 1563.010 1883.900 ;
        RECT 1599.030 1883.840 1599.350 1883.900 ;
        RECT 1562.690 1883.700 1599.350 1883.840 ;
        RECT 1562.690 1883.640 1563.010 1883.700 ;
        RECT 1599.030 1883.640 1599.350 1883.700 ;
        RECT 1392.950 1883.500 1393.270 1883.560 ;
        RECT 1448.625 1883.500 1448.915 1883.545 ;
        RECT 1392.950 1883.360 1448.915 1883.500 ;
        RECT 1392.950 1883.300 1393.270 1883.360 ;
        RECT 1448.625 1883.315 1448.915 1883.360 ;
        RECT 1449.085 1883.500 1449.375 1883.545 ;
        RECT 1449.085 1883.360 1466.320 1883.500 ;
        RECT 1449.085 1883.315 1449.375 1883.360 ;
        RECT 1466.180 1883.160 1466.320 1883.360 ;
        RECT 1490.485 1883.160 1490.775 1883.205 ;
        RECT 1466.180 1883.020 1490.775 1883.160 ;
        RECT 1490.485 1882.975 1490.775 1883.020 ;
        RECT 1514.405 1882.820 1514.695 1882.865 ;
        RECT 1601.790 1882.820 1602.110 1882.880 ;
        RECT 1514.405 1882.680 1602.110 1882.820 ;
        RECT 1514.405 1882.635 1514.695 1882.680 ;
        RECT 1601.790 1882.620 1602.110 1882.680 ;
        RECT 1372.250 1880.100 1372.570 1880.160 ;
        RECT 1602.710 1880.100 1603.030 1880.160 ;
        RECT 1372.250 1879.960 1603.030 1880.100 ;
        RECT 1372.250 1879.900 1372.570 1879.960 ;
        RECT 1602.710 1879.900 1603.030 1879.960 ;
        RECT 1392.030 1876.700 1392.350 1876.760 ;
        RECT 1601.330 1876.700 1601.650 1876.760 ;
        RECT 1392.030 1876.560 1601.650 1876.700 ;
        RECT 1392.030 1876.500 1392.350 1876.560 ;
        RECT 1601.330 1876.500 1601.650 1876.560 ;
        RECT 1368.110 1873.300 1368.430 1873.360 ;
        RECT 1369.030 1873.300 1369.350 1873.360 ;
        RECT 1368.110 1873.160 1369.350 1873.300 ;
        RECT 1368.110 1873.100 1368.430 1873.160 ;
        RECT 1369.030 1873.100 1369.350 1873.160 ;
        RECT 1372.250 1873.300 1372.570 1873.360 ;
        RECT 1600.425 1873.300 1600.715 1873.345 ;
        RECT 1604.105 1873.300 1604.395 1873.345 ;
        RECT 1372.250 1873.160 1604.395 1873.300 ;
        RECT 1372.250 1873.100 1372.570 1873.160 ;
        RECT 1600.425 1873.115 1600.715 1873.160 ;
        RECT 1604.105 1873.115 1604.395 1873.160 ;
        RECT 1367.650 1872.620 1367.970 1872.680 ;
        RECT 1369.030 1872.620 1369.350 1872.680 ;
        RECT 1367.650 1872.480 1369.350 1872.620 ;
        RECT 1367.650 1872.420 1367.970 1872.480 ;
        RECT 1369.030 1872.420 1369.350 1872.480 ;
        RECT 1602.710 1872.080 1603.030 1872.340 ;
        RECT 1602.800 1871.260 1602.940 1872.080 ;
        RECT 1603.170 1871.260 1603.490 1871.320 ;
        RECT 1602.800 1871.120 1603.490 1871.260 ;
        RECT 1603.170 1871.060 1603.490 1871.120 ;
        RECT 1391.570 1869.900 1391.890 1869.960 ;
        RECT 1600.870 1869.900 1601.190 1869.960 ;
        RECT 1391.570 1869.760 1601.190 1869.900 ;
        RECT 1391.570 1869.700 1391.890 1869.760 ;
        RECT 1600.870 1869.700 1601.190 1869.760 ;
        RECT 1600.410 1864.800 1600.730 1864.860 ;
        RECT 1602.265 1864.800 1602.555 1864.845 ;
        RECT 1599.975 1864.660 1602.555 1864.800 ;
        RECT 1600.410 1864.600 1600.730 1864.660 ;
        RECT 1602.265 1864.615 1602.555 1864.660 ;
        RECT 1391.110 1862.760 1391.430 1862.820 ;
        RECT 1391.110 1862.620 1602.020 1862.760 ;
        RECT 1391.110 1862.560 1391.430 1862.620 ;
        RECT 1601.880 1862.480 1602.020 1862.620 ;
        RECT 1601.790 1862.220 1602.110 1862.480 ;
        RECT 1372.250 1859.360 1372.570 1859.420 ;
        RECT 1599.490 1859.360 1599.810 1859.420 ;
        RECT 1602.710 1859.360 1603.030 1859.420 ;
        RECT 1372.250 1859.220 1603.030 1859.360 ;
        RECT 1372.250 1859.160 1372.570 1859.220 ;
        RECT 1599.490 1859.160 1599.810 1859.220 ;
        RECT 1602.710 1859.160 1603.030 1859.220 ;
        RECT 1604.090 1858.000 1604.410 1858.060 ;
        RECT 1603.895 1857.860 1604.410 1858.000 ;
        RECT 1604.090 1857.800 1604.410 1857.860 ;
        RECT 1390.650 1855.960 1390.970 1856.020 ;
        RECT 1601.330 1855.960 1601.650 1856.020 ;
        RECT 1390.650 1855.820 1601.650 1855.960 ;
        RECT 1390.650 1855.760 1390.970 1855.820 ;
        RECT 1601.330 1855.760 1601.650 1855.820 ;
        RECT 1601.345 1855.280 1601.635 1855.325 ;
        RECT 1604.090 1855.280 1604.410 1855.340 ;
        RECT 1601.345 1855.140 1604.410 1855.280 ;
        RECT 1601.345 1855.095 1601.635 1855.140 ;
        RECT 1604.090 1855.080 1604.410 1855.140 ;
        RECT 1372.250 1852.560 1372.570 1852.620 ;
        RECT 1599.950 1852.560 1600.270 1852.620 ;
        RECT 1372.250 1852.420 1600.270 1852.560 ;
        RECT 1372.250 1852.360 1372.570 1852.420 ;
        RECT 1599.950 1852.360 1600.270 1852.420 ;
        RECT 1603.170 1852.360 1603.490 1852.620 ;
        RECT 1604.090 1852.560 1604.410 1852.620 ;
        RECT 1603.895 1852.420 1604.410 1852.560 ;
        RECT 1604.090 1852.360 1604.410 1852.420 ;
        RECT 1603.260 1851.600 1603.400 1852.360 ;
        RECT 1603.170 1851.340 1603.490 1851.600 ;
        RECT 1403.990 1849.160 1404.310 1849.220 ;
        RECT 1600.870 1849.160 1601.190 1849.220 ;
        RECT 1403.990 1849.020 1601.190 1849.160 ;
        RECT 1403.990 1848.960 1404.310 1849.020 ;
        RECT 1600.870 1848.960 1601.190 1849.020 ;
        RECT 1417.790 1848.820 1418.110 1848.880 ;
        RECT 1599.030 1848.820 1599.350 1848.880 ;
        RECT 1417.790 1848.680 1599.350 1848.820 ;
        RECT 1417.790 1848.620 1418.110 1848.680 ;
        RECT 1599.030 1848.620 1599.350 1848.680 ;
        RECT 1599.950 1847.460 1600.270 1847.520 ;
        RECT 1603.170 1847.460 1603.490 1847.520 ;
        RECT 1599.950 1847.320 1603.490 1847.460 ;
        RECT 1599.950 1847.260 1600.270 1847.320 ;
        RECT 1603.170 1847.260 1603.490 1847.320 ;
        RECT 1599.490 1845.420 1599.810 1845.480 ;
        RECT 1601.790 1845.420 1602.110 1845.480 ;
        RECT 1599.490 1845.280 1602.110 1845.420 ;
        RECT 1599.490 1845.220 1599.810 1845.280 ;
        RECT 1601.790 1845.220 1602.110 1845.280 ;
        RECT 1601.805 1843.040 1602.095 1843.085 ;
        RECT 1602.250 1843.040 1602.570 1843.100 ;
        RECT 1601.805 1842.900 1602.570 1843.040 ;
        RECT 1601.805 1842.855 1602.095 1842.900 ;
        RECT 1602.250 1842.840 1602.570 1842.900 ;
        RECT 1390.190 1842.360 1390.510 1842.420 ;
        RECT 1602.250 1842.360 1602.570 1842.420 ;
        RECT 1390.190 1842.220 1602.570 1842.360 ;
        RECT 1390.190 1842.160 1390.510 1842.220 ;
        RECT 1602.250 1842.160 1602.570 1842.220 ;
        RECT 1601.330 1839.300 1601.650 1839.360 ;
        RECT 1601.135 1839.160 1601.650 1839.300 ;
        RECT 1601.330 1839.100 1601.650 1839.160 ;
        RECT 1490.485 1835.220 1490.775 1835.265 ;
        RECT 1463.880 1835.080 1490.775 1835.220 ;
        RECT 1462.885 1834.880 1463.175 1834.925 ;
        RECT 1463.880 1834.880 1464.020 1835.080 ;
        RECT 1490.485 1835.035 1490.775 1835.080 ;
        RECT 1462.885 1834.740 1464.020 1834.880 ;
        RECT 1538.785 1834.880 1539.075 1834.925 ;
        RECT 1587.085 1834.880 1587.375 1834.925 ;
        RECT 1538.785 1834.740 1587.375 1834.880 ;
        RECT 1462.885 1834.695 1463.175 1834.740 ;
        RECT 1538.785 1834.695 1539.075 1834.740 ;
        RECT 1587.085 1834.695 1587.375 1834.740 ;
        RECT 1424.690 1834.540 1425.010 1834.600 ;
        RECT 1462.425 1834.540 1462.715 1834.585 ;
        RECT 1424.690 1834.400 1462.715 1834.540 ;
        RECT 1424.690 1834.340 1425.010 1834.400 ;
        RECT 1462.425 1834.355 1462.715 1834.400 ;
        RECT 1490.485 1834.540 1490.775 1834.585 ;
        RECT 1490.485 1834.400 1538.540 1834.540 ;
        RECT 1490.485 1834.355 1490.775 1834.400 ;
        RECT 1538.400 1834.200 1538.540 1834.400 ;
        RECT 1538.785 1834.200 1539.075 1834.245 ;
        RECT 1538.400 1834.060 1539.075 1834.200 ;
        RECT 1538.785 1834.015 1539.075 1834.060 ;
        RECT 1587.085 1831.480 1587.375 1831.525 ;
        RECT 1593.970 1831.480 1594.290 1831.540 ;
        RECT 1587.085 1831.340 1594.290 1831.480 ;
        RECT 1587.085 1831.295 1587.375 1831.340 ;
        RECT 1593.970 1831.280 1594.290 1831.340 ;
        RECT 1601.790 1829.100 1602.110 1829.160 ;
        RECT 1600.960 1828.960 1602.110 1829.100 ;
        RECT 1600.960 1828.820 1601.100 1828.960 ;
        RECT 1601.790 1828.900 1602.110 1828.960 ;
        RECT 1600.870 1828.560 1601.190 1828.820 ;
        RECT 1431.590 1828.420 1431.910 1828.480 ;
        RECT 1601.790 1828.420 1602.110 1828.480 ;
        RECT 1431.590 1828.280 1602.110 1828.420 ;
        RECT 1431.590 1828.220 1431.910 1828.280 ;
        RECT 1601.790 1828.220 1602.110 1828.280 ;
        RECT 1438.490 1821.620 1438.810 1821.680 ;
        RECT 1601.330 1821.620 1601.650 1821.680 ;
        RECT 1438.490 1821.480 1601.650 1821.620 ;
        RECT 1438.490 1821.420 1438.810 1821.480 ;
        RECT 1601.330 1821.420 1601.650 1821.480 ;
        RECT 1599.950 1818.900 1600.270 1818.960 ;
        RECT 1602.265 1818.900 1602.555 1818.945 ;
        RECT 1599.950 1818.760 1602.555 1818.900 ;
        RECT 1599.950 1818.700 1600.270 1818.760 ;
        RECT 1602.265 1818.715 1602.555 1818.760 ;
        RECT 1368.570 1814.480 1368.890 1814.540 ;
        RECT 1602.250 1814.480 1602.570 1814.540 ;
        RECT 1368.570 1814.340 1602.570 1814.480 ;
        RECT 1368.570 1814.280 1368.890 1814.340 ;
        RECT 1602.250 1814.280 1602.570 1814.340 ;
        RECT 1452.290 1814.140 1452.610 1814.200 ;
        RECT 1599.030 1814.140 1599.350 1814.200 ;
        RECT 1452.290 1814.000 1599.350 1814.140 ;
        RECT 1452.290 1813.940 1452.610 1814.000 ;
        RECT 1599.030 1813.940 1599.350 1814.000 ;
        RECT 1600.410 1813.460 1600.730 1813.520 ;
        RECT 1601.805 1813.460 1602.095 1813.505 ;
        RECT 1600.410 1813.320 1602.095 1813.460 ;
        RECT 1600.410 1813.260 1600.730 1813.320 ;
        RECT 1601.805 1813.275 1602.095 1813.320 ;
        RECT 1367.650 1805.300 1367.970 1805.360 ;
        RECT 1377.310 1805.300 1377.630 1805.360 ;
        RECT 1367.650 1805.160 1377.630 1805.300 ;
        RECT 1367.650 1805.100 1367.970 1805.160 ;
        RECT 1377.310 1805.100 1377.630 1805.160 ;
        RECT 1601.330 1804.620 1601.650 1804.680 ;
        RECT 1603.630 1804.620 1603.950 1804.680 ;
        RECT 1601.330 1804.480 1603.950 1804.620 ;
        RECT 1601.330 1804.420 1601.650 1804.480 ;
        RECT 1603.630 1804.420 1603.950 1804.480 ;
        RECT 1604.090 1801.560 1604.410 1801.620 ;
        RECT 1602.340 1801.420 1604.410 1801.560 ;
        RECT 1602.340 1801.280 1602.480 1801.420 ;
        RECT 1604.090 1801.360 1604.410 1801.420 ;
        RECT 1602.250 1801.020 1602.570 1801.280 ;
        RECT 1601.330 1800.880 1601.650 1800.940 ;
        RECT 1601.330 1800.740 1601.845 1800.880 ;
        RECT 1601.330 1800.680 1601.650 1800.740 ;
        RECT 1601.330 1800.200 1601.650 1800.260 ;
        RECT 1603.630 1800.200 1603.950 1800.260 ;
        RECT 1601.330 1800.060 1603.950 1800.200 ;
        RECT 1601.330 1800.000 1601.650 1800.060 ;
        RECT 1603.630 1800.000 1603.950 1800.060 ;
        RECT 1601.805 1799.520 1602.095 1799.565 ;
        RECT 1603.630 1799.520 1603.950 1799.580 ;
        RECT 1601.805 1799.380 1603.950 1799.520 ;
        RECT 1601.805 1799.335 1602.095 1799.380 ;
        RECT 1603.630 1799.320 1603.950 1799.380 ;
        RECT 1599.950 1799.180 1600.270 1799.240 ;
        RECT 1604.090 1799.180 1604.410 1799.240 ;
        RECT 1599.950 1799.040 1604.410 1799.180 ;
        RECT 1599.950 1798.980 1600.270 1799.040 ;
        RECT 1604.090 1798.980 1604.410 1799.040 ;
        RECT 1369.030 1798.500 1369.350 1798.560 ;
        RECT 1376.850 1798.500 1377.170 1798.560 ;
        RECT 1369.030 1798.360 1377.170 1798.500 ;
        RECT 1369.030 1798.300 1369.350 1798.360 ;
        RECT 1376.850 1798.300 1377.170 1798.360 ;
        RECT 1600.870 1784.560 1601.190 1784.620 ;
        RECT 1601.790 1784.560 1602.110 1784.620 ;
        RECT 1600.870 1784.420 1602.110 1784.560 ;
        RECT 1600.870 1784.360 1601.190 1784.420 ;
        RECT 1601.790 1784.360 1602.110 1784.420 ;
        RECT 1459.190 1780.140 1459.510 1780.200 ;
        RECT 1600.870 1780.140 1601.190 1780.200 ;
        RECT 1459.190 1780.000 1601.190 1780.140 ;
        RECT 1459.190 1779.940 1459.510 1780.000 ;
        RECT 1600.870 1779.940 1601.190 1780.000 ;
        RECT 1371.790 1779.800 1372.110 1779.860 ;
        RECT 1376.390 1779.800 1376.710 1779.860 ;
        RECT 1371.790 1779.660 1376.710 1779.800 ;
        RECT 1371.790 1779.600 1372.110 1779.660 ;
        RECT 1376.390 1779.600 1376.710 1779.660 ;
        RECT 1601.345 1779.460 1601.635 1779.505 ;
        RECT 1603.170 1779.460 1603.490 1779.520 ;
        RECT 1601.345 1779.320 1603.490 1779.460 ;
        RECT 1601.345 1779.275 1601.635 1779.320 ;
        RECT 1603.170 1779.260 1603.490 1779.320 ;
        RECT 1472.990 1773.340 1473.310 1773.400 ;
        RECT 1600.870 1773.340 1601.190 1773.400 ;
        RECT 1472.990 1773.200 1601.190 1773.340 ;
        RECT 1472.990 1773.140 1473.310 1773.200 ;
        RECT 1600.870 1773.140 1601.190 1773.200 ;
        RECT 1369.030 1767.220 1369.350 1767.280 ;
        RECT 1374.090 1767.220 1374.410 1767.280 ;
        RECT 1369.030 1767.080 1374.410 1767.220 ;
        RECT 1369.030 1767.020 1369.350 1767.080 ;
        RECT 1374.090 1767.020 1374.410 1767.080 ;
        RECT 1371.330 1766.200 1371.650 1766.260 ;
        RECT 1600.870 1766.200 1601.190 1766.260 ;
        RECT 1371.330 1766.060 1601.190 1766.200 ;
        RECT 1371.330 1766.000 1371.650 1766.060 ;
        RECT 1600.870 1766.000 1601.190 1766.060 ;
        RECT 1486.790 1759.400 1487.110 1759.460 ;
        RECT 1601.330 1759.400 1601.650 1759.460 ;
        RECT 1486.790 1759.260 1601.650 1759.400 ;
        RECT 1486.790 1759.200 1487.110 1759.260 ;
        RECT 1601.330 1759.200 1601.650 1759.260 ;
        RECT 1370.870 1752.260 1371.190 1752.320 ;
        RECT 1601.330 1752.260 1601.650 1752.320 ;
        RECT 1370.870 1752.120 1601.650 1752.260 ;
        RECT 1370.870 1752.060 1371.190 1752.120 ;
        RECT 1601.330 1752.060 1601.650 1752.120 ;
        RECT 1367.650 1748.180 1367.970 1748.240 ;
        RECT 1375.010 1748.180 1375.330 1748.240 ;
        RECT 1367.650 1748.040 1375.330 1748.180 ;
        RECT 1367.650 1747.980 1367.970 1748.040 ;
        RECT 1375.010 1747.980 1375.330 1748.040 ;
        RECT 1370.410 1745.460 1370.730 1745.520 ;
        RECT 1600.870 1745.460 1601.190 1745.520 ;
        RECT 1370.410 1745.320 1601.190 1745.460 ;
        RECT 1370.410 1745.260 1370.730 1745.320 ;
        RECT 1600.870 1745.260 1601.190 1745.320 ;
        RECT 1493.690 1745.120 1494.010 1745.180 ;
        RECT 1601.790 1745.120 1602.110 1745.180 ;
        RECT 1493.690 1744.980 1602.110 1745.120 ;
        RECT 1493.690 1744.920 1494.010 1744.980 ;
        RECT 1601.790 1744.920 1602.110 1744.980 ;
        RECT 1367.650 1738.660 1367.970 1738.720 ;
        RECT 1375.470 1738.660 1375.790 1738.720 ;
        RECT 1367.650 1738.520 1375.790 1738.660 ;
        RECT 1367.650 1738.460 1367.970 1738.520 ;
        RECT 1375.470 1738.460 1375.790 1738.520 ;
        RECT 1507.490 1738.660 1507.810 1738.720 ;
        RECT 1600.870 1738.660 1601.190 1738.720 ;
        RECT 1507.490 1738.520 1601.190 1738.660 ;
        RECT 1507.490 1738.460 1507.810 1738.520 ;
        RECT 1600.870 1738.460 1601.190 1738.520 ;
        RECT 1369.950 1731.860 1370.270 1731.920 ;
        RECT 1600.870 1731.860 1601.190 1731.920 ;
        RECT 1369.950 1731.720 1601.190 1731.860 ;
        RECT 1369.950 1731.660 1370.270 1731.720 ;
        RECT 1600.870 1731.660 1601.190 1731.720 ;
        RECT 1367.650 1729.480 1367.970 1729.540 ;
        RECT 1375.930 1729.480 1376.250 1729.540 ;
        RECT 1367.650 1729.340 1376.250 1729.480 ;
        RECT 1367.650 1729.280 1367.970 1729.340 ;
        RECT 1375.930 1729.280 1376.250 1729.340 ;
        RECT 1368.110 1719.960 1368.430 1720.020 ;
        RECT 1379.610 1719.960 1379.930 1720.020 ;
        RECT 1368.110 1719.820 1379.930 1719.960 ;
        RECT 1368.110 1719.760 1368.430 1719.820 ;
        RECT 1379.610 1719.760 1379.930 1719.820 ;
        RECT 1367.650 1710.780 1367.970 1710.840 ;
        RECT 1378.690 1710.780 1379.010 1710.840 ;
        RECT 1367.650 1710.640 1379.010 1710.780 ;
        RECT 1367.650 1710.580 1367.970 1710.640 ;
        RECT 1378.690 1710.580 1379.010 1710.640 ;
        RECT 1367.650 1700.580 1367.970 1700.640 ;
        RECT 1379.150 1700.580 1379.470 1700.640 ;
        RECT 1367.650 1700.440 1379.470 1700.580 ;
        RECT 1367.650 1700.380 1367.970 1700.440 ;
        RECT 1379.150 1700.380 1379.470 1700.440 ;
        RECT 1369.030 1676.440 1369.350 1676.500 ;
        RECT 1514.390 1676.440 1514.710 1676.500 ;
        RECT 1369.030 1676.300 1514.710 1676.440 ;
        RECT 1369.030 1676.240 1369.350 1676.300 ;
        RECT 1514.390 1676.240 1514.710 1676.300 ;
        RECT 1371.330 1662.500 1371.650 1662.560 ;
        RECT 1397.090 1662.500 1397.410 1662.560 ;
        RECT 1371.330 1662.360 1397.410 1662.500 ;
        RECT 1371.330 1662.300 1371.650 1662.360 ;
        RECT 1397.090 1662.300 1397.410 1662.360 ;
        RECT 1366.730 1656.720 1367.050 1656.780 ;
        RECT 1367.650 1656.720 1367.970 1656.780 ;
        RECT 1366.730 1656.580 1367.970 1656.720 ;
        RECT 1366.730 1656.520 1367.050 1656.580 ;
        RECT 1367.650 1656.520 1367.970 1656.580 ;
        RECT 1366.730 1656.040 1367.050 1656.100 ;
        RECT 1597.190 1656.040 1597.510 1656.100 ;
        RECT 1366.730 1655.900 1597.510 1656.040 ;
        RECT 1366.730 1655.840 1367.050 1655.900 ;
        RECT 1597.190 1655.840 1597.510 1655.900 ;
        RECT 1369.950 1648.900 1370.270 1648.960 ;
        RECT 1583.390 1648.900 1583.710 1648.960 ;
        RECT 1369.950 1648.760 1583.710 1648.900 ;
        RECT 1369.950 1648.700 1370.270 1648.760 ;
        RECT 1583.390 1648.700 1583.710 1648.760 ;
        RECT 1367.650 1616.600 1367.970 1616.660 ;
        RECT 1378.230 1616.600 1378.550 1616.660 ;
        RECT 1367.650 1616.460 1378.550 1616.600 ;
        RECT 1367.650 1616.400 1367.970 1616.460 ;
        RECT 1378.230 1616.400 1378.550 1616.460 ;
        RECT 1367.190 1606.400 1367.510 1606.460 ;
        RECT 1377.770 1606.400 1378.090 1606.460 ;
        RECT 1367.190 1606.260 1378.090 1606.400 ;
        RECT 1367.190 1606.200 1367.510 1606.260 ;
        RECT 1377.770 1606.200 1378.090 1606.260 ;
      LAYER met1 ;
        RECT 1605.000 1605.000 2051.235 1981.480 ;
      LAYER via ;
        RECT 783.020 3277.640 783.280 3277.900 ;
        RECT 938.500 3277.640 938.760 3277.900 ;
        RECT 597.180 2842.440 597.440 2842.700 ;
        RECT 642.260 2842.440 642.520 2842.700 ;
        RECT 605.000 2841.420 605.260 2841.680 ;
        RECT 700.220 2841.420 700.480 2841.680 ;
        RECT 482.640 2839.720 482.900 2839.980 ;
        RECT 526.340 2839.720 526.600 2839.980 ;
        RECT 573.720 2839.720 573.980 2839.980 ;
        RECT 621.560 2841.080 621.820 2841.340 ;
        RECT 642.260 2840.740 642.520 2841.000 ;
        RECT 745.300 2840.740 745.560 2841.000 ;
        RECT 620.640 2840.400 620.900 2840.660 ;
        RECT 734.720 2840.400 734.980 2840.660 ;
        RECT 1089.380 2840.400 1089.640 2840.660 ;
        RECT 1135.840 2840.400 1136.100 2840.660 ;
        RECT 1180.000 2840.400 1180.260 2840.660 ;
        RECT 600.400 2840.060 600.660 2840.320 ;
        RECT 720.920 2840.060 721.180 2840.320 ;
        RECT 1018.540 2839.720 1018.800 2839.980 ;
        RECT 1065.460 2839.720 1065.720 2839.980 ;
        RECT 1111.920 2839.720 1112.180 2839.980 ;
        RECT 1159.300 2839.720 1159.560 2839.980 ;
        RECT 510.240 2839.380 510.500 2839.640 ;
        RECT 549.340 2839.380 549.600 2839.640 ;
        RECT 627.540 2839.380 627.800 2839.640 ;
        RECT 762.320 2839.380 762.580 2839.640 ;
        RECT 1024.060 2839.380 1024.320 2839.640 ;
        RECT 1070.520 2839.380 1070.780 2839.640 ;
        RECT 1118.360 2839.380 1118.620 2839.640 ;
        RECT 1159.760 2839.380 1160.020 2839.640 ;
        RECT 590.280 2839.040 590.540 2839.300 ;
        RECT 714.020 2839.040 714.280 2839.300 ;
        RECT 427.440 2838.360 427.700 2838.620 ;
        RECT 455.500 2838.360 455.760 2838.620 ;
        RECT 503.340 2838.360 503.600 2838.620 ;
        RECT 783.940 2838.360 784.200 2838.620 ;
        RECT 489.540 2838.020 489.800 2838.280 ;
        RECT 776.120 2838.020 776.380 2838.280 ;
        RECT 475.740 2837.680 476.000 2837.940 ;
        RECT 769.220 2837.680 769.480 2837.940 ;
        RECT 551.640 2837.340 551.900 2837.600 ;
        RECT 693.320 2837.340 693.580 2837.600 ;
        RECT 406.740 2836.660 407.000 2836.920 ;
        RECT 441.700 2836.660 441.960 2836.920 ;
        RECT 627.080 2836.660 627.340 2836.920 ;
        RECT 1024.060 2836.660 1024.320 2836.920 ;
        RECT 1045.220 2836.660 1045.480 2836.920 ;
        RECT 1089.380 2836.660 1089.640 2836.920 ;
        RECT 413.640 2836.320 413.900 2836.580 ;
        RECT 449.980 2836.320 450.240 2836.580 ;
        RECT 390.640 2835.980 390.900 2836.240 ;
        RECT 434.800 2835.980 435.060 2836.240 ;
        RECT 613.280 2835.980 613.540 2836.240 ;
        RECT 1018.540 2835.980 1018.800 2836.240 ;
        RECT 558.540 2628.580 558.800 2628.840 ;
        RECT 907.220 2628.580 907.480 2628.840 ;
        RECT 640.880 2627.900 641.140 2628.160 ;
        RECT 1040.620 2627.900 1040.880 2628.160 ;
        RECT 507.020 2627.560 507.280 2627.820 ;
        RECT 941.720 2627.560 941.980 2627.820 ;
        RECT 497.360 2627.220 497.620 2627.480 ;
        RECT 942.180 2627.220 942.440 2627.480 ;
        RECT 488.160 2626.880 488.420 2627.140 ;
        RECT 942.640 2626.880 942.900 2627.140 ;
        RECT 478.500 2626.540 478.760 2626.800 ;
        RECT 943.100 2626.540 943.360 2626.800 ;
        RECT 468.840 2626.200 469.100 2626.460 ;
        RECT 943.560 2626.200 943.820 2626.460 ;
        RECT 459.180 2625.860 459.440 2626.120 ;
        RECT 944.020 2625.860 944.280 2626.120 ;
        RECT 430.660 2625.520 430.920 2625.780 ;
        RECT 944.480 2625.520 944.740 2625.780 ;
        RECT 449.980 2625.180 450.240 2625.440 ;
        RECT 979.900 2625.180 980.160 2625.440 ;
        RECT 544.740 2624.840 545.000 2625.100 ;
        RECT 878.700 2624.840 878.960 2625.100 ;
        RECT 537.840 2624.500 538.100 2624.760 ;
        RECT 869.040 2624.500 869.300 2624.760 ;
        RECT 524.040 2624.160 524.300 2624.420 ;
        RECT 850.180 2624.160 850.440 2624.420 ;
        RECT 530.940 2623.820 531.200 2624.080 ;
        RECT 859.840 2623.820 860.100 2624.080 ;
        RECT 468.380 2623.480 468.640 2623.740 ;
        RECT 754.960 2623.480 755.220 2623.740 ;
        RECT 373.620 2621.780 373.880 2622.040 ;
        RECT 379.140 2621.780 379.400 2622.040 ;
        RECT 402.140 2621.780 402.400 2622.040 ;
        RECT 406.740 2621.780 407.000 2622.040 ;
        RECT 421.460 2621.780 421.720 2622.040 ;
        RECT 427.440 2621.780 427.700 2622.040 ;
        RECT 475.280 2621.780 475.540 2622.040 ;
        RECT 764.160 2621.780 764.420 2622.040 ;
        RECT 769.220 2621.780 769.480 2622.040 ;
        RECT 773.820 2621.780 774.080 2622.040 ;
        RECT 776.120 2621.780 776.380 2622.040 ;
        RECT 792.680 2621.780 792.940 2622.040 ;
        RECT 495.980 2621.440 496.240 2621.700 ;
        RECT 482.180 2621.100 482.440 2621.360 ;
        RECT 782.100 2621.440 782.360 2621.700 ;
        RECT 783.940 2621.100 784.200 2621.360 ;
        RECT 812.000 2621.780 812.260 2622.040 ;
        RECT 1041.540 2621.780 1041.800 2622.040 ;
        RECT 1097.660 2621.780 1097.920 2622.040 ;
        RECT 1145.040 2621.780 1145.300 2622.040 ;
        RECT 1269.240 2621.780 1269.500 2622.040 ;
        RECT 1138.140 2621.440 1138.400 2621.700 ;
        RECT 1260.040 2621.440 1260.300 2621.700 ;
        RECT 1048.440 2621.100 1048.700 2621.360 ;
        RECT 1107.320 2621.100 1107.580 2621.360 ;
        RECT 1158.840 2621.100 1159.100 2621.360 ;
        RECT 1288.560 2621.100 1288.820 2621.360 ;
        RECT 509.780 2620.760 510.040 2621.020 ;
        RECT 821.660 2620.760 821.920 2621.020 ;
        RECT 1062.240 2620.760 1062.500 2621.020 ;
        RECT 1135.840 2620.760 1136.100 2621.020 ;
        RECT 1151.940 2620.760 1152.200 2621.020 ;
        RECT 1278.900 2620.760 1279.160 2621.020 ;
        RECT 394.320 2620.420 394.580 2620.680 ;
        RECT 440.320 2620.420 440.580 2620.680 ;
        RECT 516.680 2620.420 516.940 2620.680 ;
        RECT 840.520 2620.420 840.780 2620.680 ;
        RECT 1126.640 2620.420 1126.900 2620.680 ;
        RECT 1165.740 2620.420 1166.000 2620.680 ;
        RECT 1297.760 2620.420 1298.020 2620.680 ;
        RECT 393.860 2620.080 394.120 2620.340 ;
        RECT 393.400 2619.740 393.660 2620.000 ;
        RECT 926.540 2620.080 926.800 2620.340 ;
        RECT 1020.840 2620.080 1021.100 2620.340 ;
        RECT 1069.140 2620.080 1069.400 2620.340 ;
        RECT 1069.600 2620.080 1069.860 2620.340 ;
        RECT 1145.500 2620.080 1145.760 2620.340 ;
        RECT 1172.640 2620.080 1172.900 2620.340 ;
        RECT 1317.080 2620.080 1317.340 2620.340 ;
        RECT 391.560 2619.400 391.820 2619.660 ;
        RECT 545.200 2619.740 545.460 2620.000 ;
        RECT 592.580 2619.740 592.840 2620.000 ;
        RECT 955.060 2619.740 955.320 2620.000 ;
        RECT 1027.740 2619.740 1028.000 2620.000 ;
        RECT 1078.800 2619.740 1079.060 2620.000 ;
        RECT 1082.940 2619.740 1083.200 2620.000 ;
        RECT 1164.360 2619.740 1164.620 2620.000 ;
        RECT 1179.540 2619.740 1179.800 2620.000 ;
        RECT 1307.420 2619.740 1307.680 2620.000 ;
        RECT 554.860 2619.400 555.120 2619.660 ;
        RECT 572.340 2619.400 572.600 2619.660 ;
        RECT 613.740 2619.400 614.000 2619.660 ;
        RECT 993.240 2619.400 993.500 2619.660 ;
        RECT 1076.040 2619.400 1076.300 2619.660 ;
        RECT 1155.160 2619.400 1155.420 2619.660 ;
        RECT 1165.280 2619.400 1165.540 2619.660 ;
        RECT 392.020 2619.060 392.280 2619.320 ;
        RECT 573.720 2619.060 573.980 2619.320 ;
        RECT 621.560 2619.060 621.820 2619.320 ;
        RECT 627.080 2619.060 627.340 2619.320 ;
        RECT 1054.880 2619.060 1055.140 2619.320 ;
        RECT 1186.440 2619.400 1186.700 2619.660 ;
        RECT 1335.940 2619.400 1336.200 2619.660 ;
        RECT 392.480 2618.720 392.740 2618.980 ;
        RECT 583.380 2618.720 583.640 2618.980 ;
        RECT 650.080 2618.720 650.340 2618.980 ;
        RECT 1045.220 2618.720 1045.480 2618.980 ;
        RECT 1096.740 2618.720 1097.000 2618.980 ;
        RECT 1191.500 2618.720 1191.760 2618.980 ;
        RECT 392.940 2618.380 393.200 2618.640 ;
        RECT 592.580 2618.380 592.840 2618.640 ;
        RECT 1089.380 2618.380 1089.640 2618.640 ;
        RECT 1183.680 2618.380 1183.940 2618.640 ;
        RECT 1193.340 2619.060 1193.600 2619.320 ;
        RECT 1326.740 2619.060 1327.000 2619.320 ;
        RECT 1345.600 2618.720 1345.860 2618.980 ;
        RECT 391.100 2618.040 391.360 2618.300 ;
        RECT 535.540 2618.040 535.800 2618.300 ;
        RECT 700.220 2618.040 700.480 2618.300 ;
        RECT 983.580 2618.040 983.840 2618.300 ;
        RECT 1131.240 2618.040 1131.500 2618.300 ;
        RECT 1250.380 2618.040 1250.640 2618.300 ;
        RECT 516.680 2617.700 516.940 2617.960 ;
        RECT 779.800 2617.700 780.060 2617.960 ;
        RECT 802.340 2617.700 802.600 2617.960 ;
        RECT 1130.780 2617.700 1131.040 2617.960 ;
        RECT 1240.720 2617.700 1240.980 2617.960 ;
        RECT 433.880 2617.360 434.140 2617.620 ;
        RECT 525.880 2617.360 526.140 2617.620 ;
        RECT 564.060 2617.360 564.320 2617.620 ;
        RECT 734.720 2617.020 734.980 2617.280 ;
        RECT 1002.440 2617.360 1002.700 2617.620 ;
        RECT 1117.440 2617.360 1117.700 2617.620 ;
        RECT 1221.860 2617.360 1222.120 2617.620 ;
        RECT 625.240 2616.680 625.500 2616.940 ;
        RECT 707.120 2616.680 707.380 2616.940 ;
        RECT 720.920 2616.680 721.180 2616.940 ;
        RECT 964.260 2617.020 964.520 2617.280 ;
        RECT 1124.340 2617.020 1124.600 2617.280 ;
        RECT 1231.060 2617.020 1231.320 2617.280 ;
        RECT 1110.540 2616.680 1110.800 2616.940 ;
        RECT 1212.200 2616.680 1212.460 2616.940 ;
        RECT 1103.640 2616.340 1103.900 2616.600 ;
        RECT 1202.540 2616.340 1202.800 2616.600 ;
        RECT 935.740 2616.000 936.000 2616.260 ;
        RECT 693.320 2615.320 693.580 2615.580 ;
        RECT 897.560 2615.320 897.820 2615.580 ;
        RECT 714.020 2614.980 714.280 2615.240 ;
        RECT 1371.360 2594.580 1371.620 2594.840 ;
        RECT 1507.520 2594.580 1507.780 2594.840 ;
        RECT 1369.520 2583.700 1369.780 2583.960 ;
        RECT 1688.760 2583.700 1689.020 2583.960 ;
        RECT 1691.980 2583.700 1692.240 2583.960 ;
        RECT 1704.400 2583.700 1704.660 2583.960 ;
        RECT 1376.880 2583.360 1377.140 2583.620 ;
        RECT 1994.200 2583.360 1994.460 2583.620 ;
        RECT 1377.340 2583.020 1377.600 2583.280 ;
        RECT 2001.100 2583.020 2001.360 2583.280 ;
        RECT 1371.820 2582.680 1372.080 2582.940 ;
        RECT 2008.000 2582.680 2008.260 2582.940 ;
        RECT 1372.280 2582.340 1372.540 2582.600 ;
        RECT 2016.740 2582.340 2017.000 2582.600 ;
        RECT 1372.740 2582.000 1373.000 2582.260 ;
        RECT 2021.800 2582.000 2022.060 2582.260 ;
        RECT 2030.080 2582.000 2030.340 2582.260 ;
        RECT 1369.060 2581.660 1369.320 2581.920 ;
        RECT 1368.140 2573.840 1368.400 2574.100 ;
        RECT 1493.720 2573.840 1493.980 2574.100 ;
        RECT 1376.420 2559.900 1376.680 2560.160 ;
        RECT 1600.900 2559.900 1601.160 2560.160 ;
        RECT 1367.680 2553.100 1367.940 2553.360 ;
        RECT 1486.820 2553.100 1487.080 2553.360 ;
        RECT 1397.120 2546.300 1397.380 2546.560 ;
        RECT 1601.820 2546.300 1602.080 2546.560 ;
        RECT 1514.420 2539.160 1514.680 2539.420 ;
        RECT 1600.900 2539.160 1601.160 2539.420 ;
        RECT 1368.600 2532.700 1368.860 2532.960 ;
        RECT 1473.020 2532.700 1473.280 2532.960 ;
        RECT 1377.800 2532.360 1378.060 2532.620 ;
        RECT 1599.060 2532.360 1599.320 2532.620 ;
        RECT 1367.680 2525.900 1367.940 2526.160 ;
        RECT 1459.220 2525.900 1459.480 2526.160 ;
        RECT 1378.260 2525.560 1378.520 2525.820 ;
        RECT 1600.900 2525.560 1601.160 2525.820 ;
        RECT 1383.320 2518.420 1383.580 2518.680 ;
        RECT 1599.980 2518.420 1600.240 2518.680 ;
        RECT 1601.360 2512.640 1601.620 2512.900 ;
        RECT 1383.780 2512.300 1384.040 2512.560 ;
        RECT 1368.140 2505.160 1368.400 2505.420 ;
        RECT 1452.320 2505.160 1452.580 2505.420 ;
        RECT 1384.240 2504.820 1384.500 2505.080 ;
        RECT 1599.060 2504.820 1599.320 2505.080 ;
        RECT 1368.600 2498.020 1368.860 2498.280 ;
        RECT 1438.520 2498.020 1438.780 2498.280 ;
        RECT 1384.700 2497.680 1384.960 2497.940 ;
        RECT 1600.900 2497.680 1601.160 2497.940 ;
        RECT 1385.160 2490.880 1385.420 2491.140 ;
        RECT 1599.060 2490.880 1599.320 2491.140 ;
        RECT 1368.600 2484.420 1368.860 2484.680 ;
        RECT 1431.620 2484.420 1431.880 2484.680 ;
        RECT 1392.980 2484.080 1393.240 2484.340 ;
        RECT 1600.900 2484.080 1601.160 2484.340 ;
        RECT 1368.600 2477.960 1368.860 2478.220 ;
        RECT 1424.720 2477.960 1424.980 2478.220 ;
        RECT 1397.580 2477.620 1397.840 2477.880 ;
        RECT 1599.060 2477.620 1599.320 2477.880 ;
        RECT 1378.720 2477.280 1378.980 2477.540 ;
        RECT 1599.980 2477.280 1600.240 2477.540 ;
        RECT 1603.200 2477.280 1603.460 2477.540 ;
        RECT 1368.140 2470.480 1368.400 2470.740 ;
        RECT 1390.220 2470.480 1390.480 2470.740 ;
        RECT 1379.180 2470.140 1379.440 2470.400 ;
        RECT 1599.060 2470.140 1599.320 2470.400 ;
        RECT 1379.640 2463.340 1379.900 2463.600 ;
        RECT 1600.900 2463.340 1601.160 2463.600 ;
        RECT 1603.660 2461.640 1603.920 2461.900 ;
        RECT 1604.120 2461.640 1604.380 2461.900 ;
        RECT 1603.660 2460.620 1603.920 2460.880 ;
        RECT 1604.120 2460.620 1604.380 2460.880 ;
        RECT 1368.140 2456.880 1368.400 2457.140 ;
        RECT 1417.820 2456.880 1418.080 2457.140 ;
        RECT 1375.960 2456.540 1376.220 2456.800 ;
        RECT 1599.060 2456.540 1599.320 2456.800 ;
        RECT 1603.200 2454.500 1603.460 2454.760 ;
        RECT 1367.220 2449.740 1367.480 2450.000 ;
        RECT 1404.020 2449.740 1404.280 2450.000 ;
        RECT 1375.500 2449.400 1375.760 2449.660 ;
        RECT 1600.900 2449.400 1601.160 2449.660 ;
        RECT 1603.200 2449.400 1603.460 2449.660 ;
        RECT 1600.440 2449.060 1600.700 2449.320 ;
        RECT 1603.660 2449.060 1603.920 2449.320 ;
        RECT 1604.120 2449.060 1604.380 2449.320 ;
        RECT 1604.120 2447.020 1604.380 2447.280 ;
        RECT 1368.140 2443.280 1368.400 2443.540 ;
        RECT 1390.680 2443.280 1390.940 2443.540 ;
        RECT 1375.040 2442.940 1375.300 2443.200 ;
        RECT 1599.060 2442.940 1599.320 2443.200 ;
        RECT 1374.580 2442.600 1374.840 2442.860 ;
        RECT 1598.600 2442.600 1598.860 2442.860 ;
        RECT 1602.280 2436.140 1602.540 2436.400 ;
        RECT 1374.120 2435.800 1374.380 2436.060 ;
        RECT 1600.900 2435.800 1601.160 2436.060 ;
        RECT 1602.740 2431.040 1603.000 2431.300 ;
        RECT 1603.200 2431.040 1603.460 2431.300 ;
        RECT 1602.740 2430.020 1603.000 2430.280 ;
        RECT 1603.200 2430.020 1603.460 2430.280 ;
        RECT 1367.680 2429.340 1367.940 2429.600 ;
        RECT 1391.140 2429.340 1391.400 2429.600 ;
        RECT 1373.660 2429.000 1373.920 2429.260 ;
        RECT 1599.060 2429.000 1599.320 2429.260 ;
        RECT 1368.140 2422.200 1368.400 2422.460 ;
        RECT 1391.600 2422.200 1391.860 2422.460 ;
        RECT 1373.200 2421.860 1373.460 2422.120 ;
        RECT 1600.900 2421.860 1601.160 2422.120 ;
        RECT 1386.080 2415.060 1386.340 2415.320 ;
        RECT 1599.060 2415.060 1599.320 2415.320 ;
        RECT 1602.280 2414.040 1602.540 2414.300 ;
        RECT 1602.280 2413.360 1602.540 2413.620 ;
        RECT 1603.200 2413.360 1603.460 2413.620 ;
        RECT 1604.120 2413.360 1604.380 2413.620 ;
        RECT 1602.740 2411.660 1603.000 2411.920 ;
        RECT 1368.140 2408.600 1368.400 2408.860 ;
        RECT 1392.060 2408.600 1392.320 2408.860 ;
        RECT 1386.540 2408.260 1386.800 2408.520 ;
        RECT 1600.900 2408.260 1601.160 2408.520 ;
        RECT 1601.360 2402.140 1601.620 2402.400 ;
        RECT 1604.120 2402.140 1604.380 2402.400 ;
        RECT 1368.140 2401.460 1368.400 2401.720 ;
        RECT 1392.520 2401.460 1392.780 2401.720 ;
        RECT 1601.360 2401.460 1601.620 2401.720 ;
        RECT 1382.860 2401.120 1383.120 2401.380 ;
        RECT 1599.060 2401.120 1599.320 2401.380 ;
        RECT 1604.120 2397.040 1604.380 2397.300 ;
        RECT 1600.900 2396.360 1601.160 2396.620 ;
        RECT 1604.120 2396.360 1604.380 2396.620 ;
        RECT 1603.200 2394.660 1603.460 2394.920 ;
        RECT 1368.140 2394.320 1368.400 2394.580 ;
        RECT 1576.520 2394.320 1576.780 2394.580 ;
        RECT 1602.280 2384.800 1602.540 2385.060 ;
        RECT 1603.200 2384.800 1603.460 2385.060 ;
        RECT 1600.900 2384.120 1601.160 2384.380 ;
        RECT 1601.360 2383.100 1601.620 2383.360 ;
        RECT 1368.140 2380.380 1368.400 2380.640 ;
        RECT 1562.720 2380.380 1562.980 2380.640 ;
        RECT 1603.660 2380.040 1603.920 2380.300 ;
        RECT 1603.200 2379.360 1603.460 2379.620 ;
        RECT 1602.280 2379.020 1602.540 2379.280 ;
        RECT 1604.120 2378.680 1604.380 2378.940 ;
        RECT 1368.140 2373.920 1368.400 2374.180 ;
        RECT 1548.920 2373.920 1549.180 2374.180 ;
        RECT 1382.400 2373.580 1382.660 2373.840 ;
        RECT 1600.900 2373.580 1601.160 2373.840 ;
        RECT 1367.680 2369.840 1367.940 2370.100 ;
        RECT 1601.820 2369.840 1602.080 2370.100 ;
        RECT 1368.140 2366.780 1368.400 2367.040 ;
        RECT 1542.020 2366.780 1542.280 2367.040 ;
        RECT 1367.220 2359.980 1367.480 2360.240 ;
        RECT 1600.900 2359.980 1601.160 2360.240 ;
        RECT 1367.680 2353.180 1367.940 2353.440 ;
        RECT 1528.220 2353.180 1528.480 2353.440 ;
        RECT 1366.760 2352.840 1367.020 2353.100 ;
        RECT 1601.360 2352.840 1601.620 2353.100 ;
        RECT 1601.360 2352.160 1601.620 2352.420 ;
        RECT 1367.680 2346.380 1367.940 2346.640 ;
        RECT 1521.320 2346.380 1521.580 2346.640 ;
        RECT 1381.940 2346.040 1382.200 2346.300 ;
        RECT 1601.820 2346.040 1602.080 2346.300 ;
        RECT 1381.480 2339.580 1381.740 2339.840 ;
        RECT 1602.280 2339.580 1602.540 2339.840 ;
        RECT 1381.020 2339.240 1381.280 2339.500 ;
        RECT 1601.360 2339.240 1601.620 2339.500 ;
        RECT 1602.740 2338.900 1603.000 2339.160 ;
        RECT 1601.360 2338.560 1601.620 2338.820 ;
        RECT 1603.660 2338.560 1603.920 2338.820 ;
        RECT 1600.440 2338.220 1600.700 2338.480 ;
        RECT 1602.740 2338.220 1603.000 2338.480 ;
        RECT 1601.820 2337.880 1602.080 2338.140 ;
        RECT 1603.200 2337.540 1603.460 2337.800 ;
        RECT 1603.660 2336.860 1603.920 2337.120 ;
        RECT 1367.680 2332.440 1367.940 2332.700 ;
        RECT 1514.880 2332.440 1515.140 2332.700 ;
        RECT 1380.560 2332.100 1380.820 2332.360 ;
        RECT 1600.900 2332.100 1601.160 2332.360 ;
        RECT 1380.100 2325.300 1380.360 2325.560 ;
        RECT 1600.900 2325.300 1601.160 2325.560 ;
        RECT 1366.300 2318.500 1366.560 2318.760 ;
        RECT 1385.620 2318.500 1385.880 2318.760 ;
        RECT 1366.300 2304.560 1366.560 2304.820 ;
        RECT 1393.440 2304.560 1393.700 2304.820 ;
        RECT 1366.300 2300.140 1366.560 2300.400 ;
        RECT 1380.100 2300.140 1380.360 2300.400 ;
        RECT 1366.300 2290.620 1366.560 2290.880 ;
        RECT 1380.560 2290.620 1380.820 2290.880 ;
        RECT 1602.280 2287.220 1602.540 2287.480 ;
        RECT 1603.200 2287.220 1603.460 2287.480 ;
        RECT 1604.120 2286.540 1604.380 2286.800 ;
        RECT 1600.900 2285.520 1601.160 2285.780 ;
        RECT 1601.820 2284.500 1602.080 2284.760 ;
        RECT 1603.660 2284.500 1603.920 2284.760 ;
        RECT 1601.820 2283.140 1602.080 2283.400 ;
        RECT 1602.280 2283.140 1602.540 2283.400 ;
        RECT 1603.200 2282.460 1603.460 2282.720 ;
        RECT 1366.300 2281.100 1366.560 2281.360 ;
        RECT 1381.020 2281.100 1381.280 2281.360 ;
        RECT 1366.300 2271.580 1366.560 2271.840 ;
        RECT 1381.480 2271.580 1381.740 2271.840 ;
        RECT 1366.300 2262.060 1366.560 2262.320 ;
        RECT 1381.940 2262.060 1382.200 2262.320 ;
        RECT 1600.900 2261.380 1601.160 2261.640 ;
        RECT 1603.200 2249.140 1603.460 2249.400 ;
        RECT 1601.820 2236.560 1602.080 2236.820 ;
        RECT 1602.280 2236.560 1602.540 2236.820 ;
        RECT 1602.740 2236.560 1603.000 2236.820 ;
        RECT 1602.280 2235.880 1602.540 2236.140 ;
        RECT 1602.740 2235.880 1603.000 2236.140 ;
        RECT 1603.200 2235.540 1603.460 2235.800 ;
        RECT 1367.220 2235.200 1367.480 2235.460 ;
        RECT 1601.820 2234.860 1602.080 2235.120 ;
        RECT 1604.120 2234.520 1604.380 2234.780 ;
        RECT 1603.660 2234.180 1603.920 2234.440 ;
        RECT 1604.120 2233.840 1604.380 2234.100 ;
        RECT 1367.220 2223.980 1367.480 2224.240 ;
        RECT 1382.400 2223.980 1382.660 2224.240 ;
        RECT 1367.220 2214.460 1367.480 2214.720 ;
        RECT 1382.860 2214.460 1383.120 2214.720 ;
        RECT 1602.740 2212.080 1603.000 2212.340 ;
        RECT 1603.660 2212.080 1603.920 2212.340 ;
        RECT 1602.740 2210.720 1603.000 2210.980 ;
        RECT 1602.280 2210.040 1602.540 2210.300 ;
        RECT 1367.220 2206.300 1367.480 2206.560 ;
        RECT 1386.540 2206.300 1386.800 2206.560 ;
        RECT 1367.220 2198.480 1367.480 2198.740 ;
        RECT 1386.080 2198.480 1386.340 2198.740 ;
        RECT 1366.300 2166.860 1366.560 2167.120 ;
        RECT 1374.120 2166.860 1374.380 2167.120 ;
        RECT 1601.360 2159.720 1601.620 2159.980 ;
        RECT 1604.120 2159.720 1604.380 2159.980 ;
        RECT 1366.300 2157.340 1366.560 2157.600 ;
        RECT 1374.580 2157.340 1374.840 2157.600 ;
        RECT 1366.300 2147.820 1366.560 2148.080 ;
        RECT 1375.040 2147.820 1375.300 2148.080 ;
        RECT 1601.360 2138.640 1601.620 2138.900 ;
        RECT 1604.120 2138.640 1604.380 2138.900 ;
        RECT 1366.300 2138.300 1366.560 2138.560 ;
        RECT 1375.500 2138.300 1375.760 2138.560 ;
        RECT 1366.300 2128.780 1366.560 2129.040 ;
        RECT 1375.960 2128.780 1376.220 2129.040 ;
        RECT 1367.220 2119.940 1367.480 2120.200 ;
        RECT 1379.640 2119.940 1379.900 2120.200 ;
        RECT 1367.220 2110.080 1367.480 2110.340 ;
        RECT 1379.180 2110.080 1379.440 2110.340 ;
        RECT 1367.220 2100.220 1367.480 2100.480 ;
        RECT 1378.720 2100.220 1378.980 2100.480 ;
        RECT 1367.220 2090.360 1367.480 2090.620 ;
        RECT 1397.580 2090.360 1397.840 2090.620 ;
        RECT 1367.220 2081.180 1367.480 2081.440 ;
        RECT 1392.980 2081.180 1393.240 2081.440 ;
        RECT 1367.220 2071.660 1367.480 2071.920 ;
        RECT 1385.160 2071.660 1385.420 2071.920 ;
        RECT 1367.220 2062.140 1367.480 2062.400 ;
        RECT 1384.700 2062.140 1384.960 2062.400 ;
        RECT 1367.220 2052.620 1367.480 2052.880 ;
        RECT 1384.240 2052.620 1384.500 2052.880 ;
        RECT 1367.220 2043.100 1367.480 2043.360 ;
        RECT 1383.780 2043.100 1384.040 2043.360 ;
        RECT 1367.220 2033.580 1367.480 2033.840 ;
        RECT 1383.320 2033.580 1383.580 2033.840 ;
        RECT 1367.220 2014.540 1367.480 2014.800 ;
        RECT 1378.260 2014.540 1378.520 2014.800 ;
        RECT 1367.220 2005.020 1367.480 2005.280 ;
        RECT 1377.800 2005.020 1378.060 2005.280 ;
        RECT 1367.220 2000.600 1367.480 2000.860 ;
        RECT 1603.660 2000.600 1603.920 2000.860 ;
        RECT 1600.900 1994.140 1601.160 1994.400 ;
        RECT 1604.120 1994.140 1604.380 1994.400 ;
        RECT 1367.220 1987.000 1367.480 1987.260 ;
        RECT 1603.200 1987.000 1603.460 1987.260 ;
        RECT 1366.300 1983.940 1366.560 1984.200 ;
        RECT 1693.360 1983.940 1693.620 1984.200 ;
        RECT 1378.720 1983.600 1378.980 1983.860 ;
        RECT 1987.300 1983.600 1987.560 1983.860 ;
        RECT 1379.640 1983.260 1379.900 1983.520 ;
        RECT 1994.200 1983.260 1994.460 1983.520 ;
        RECT 1375.960 1982.920 1376.220 1983.180 ;
        RECT 2001.100 1982.920 2001.360 1983.180 ;
        RECT 1375.500 1982.580 1375.760 1982.840 ;
        RECT 2008.000 1982.580 2008.260 1982.840 ;
        RECT 1375.040 1982.240 1375.300 1982.500 ;
        RECT 2016.740 1982.240 2017.000 1982.500 ;
        RECT 1374.580 1981.900 1374.840 1982.160 ;
        RECT 2021.800 1981.900 2022.060 1982.160 ;
        RECT 2030.080 1981.900 2030.340 1982.160 ;
        RECT 1374.120 1981.560 1374.380 1981.820 ;
        RECT 1367.220 1979.860 1367.480 1980.120 ;
        RECT 1602.740 1979.860 1603.000 1980.120 ;
        RECT 1367.220 1973.060 1367.480 1973.320 ;
        RECT 1602.280 1973.060 1602.540 1973.320 ;
        RECT 1379.180 1960.140 1379.440 1960.400 ;
        RECT 1600.900 1960.140 1601.160 1960.400 ;
        RECT 1377.800 1959.800 1378.060 1960.060 ;
        RECT 1601.360 1959.800 1601.620 1960.060 ;
        RECT 1367.220 1959.460 1367.480 1959.720 ;
        RECT 1601.820 1959.460 1602.080 1959.720 ;
        RECT 1378.260 1952.660 1378.520 1952.920 ;
        RECT 1600.440 1952.660 1600.700 1952.920 ;
        RECT 1367.680 1952.320 1367.940 1952.580 ;
        RECT 1600.900 1952.320 1601.160 1952.580 ;
        RECT 1367.220 1945.860 1367.480 1946.120 ;
        RECT 1601.360 1945.860 1601.620 1946.120 ;
        RECT 1366.760 1940.080 1367.020 1940.340 ;
        RECT 1367.680 1940.080 1367.940 1940.340 ;
        RECT 1600.900 1939.060 1601.160 1939.320 ;
        RECT 1368.140 1938.720 1368.400 1938.980 ;
        RECT 1604.120 1938.720 1604.380 1938.980 ;
        RECT 1393.440 1938.380 1393.700 1938.640 ;
        RECT 1601.820 1938.380 1602.080 1938.640 ;
        RECT 1368.140 1937.700 1368.400 1937.960 ;
        RECT 1385.620 1931.580 1385.880 1931.840 ;
        RECT 1601.360 1931.580 1601.620 1931.840 ;
        RECT 1366.760 1924.780 1367.020 1925.040 ;
        RECT 1600.900 1924.780 1601.160 1925.040 ;
        RECT 1514.880 1924.440 1515.140 1924.700 ;
        RECT 1601.820 1924.440 1602.080 1924.700 ;
        RECT 1521.320 1917.980 1521.580 1918.240 ;
        RECT 1600.900 1917.980 1601.160 1918.240 ;
        RECT 1366.760 1917.640 1367.020 1917.900 ;
        RECT 1367.220 1916.620 1367.480 1916.880 ;
        RECT 1528.220 1910.840 1528.480 1911.100 ;
        RECT 1602.740 1910.840 1603.000 1911.100 ;
        RECT 1603.200 1906.760 1603.460 1907.020 ;
        RECT 1542.020 1904.040 1542.280 1904.300 ;
        RECT 1600.900 1904.040 1601.160 1904.300 ;
        RECT 1604.120 1901.320 1604.380 1901.580 ;
        RECT 1367.680 1900.980 1367.940 1901.240 ;
        RECT 1600.440 1900.980 1600.700 1901.240 ;
        RECT 1368.140 1900.640 1368.400 1900.900 ;
        RECT 1602.280 1900.640 1602.540 1900.900 ;
        RECT 1603.200 1898.600 1603.460 1898.860 ;
        RECT 1603.660 1897.580 1603.920 1897.840 ;
        RECT 1548.920 1897.240 1549.180 1897.500 ;
        RECT 1601.360 1897.240 1601.620 1897.500 ;
        RECT 1367.680 1894.520 1367.940 1894.780 ;
        RECT 1372.280 1894.520 1372.540 1894.780 ;
        RECT 1373.200 1894.180 1373.460 1894.440 ;
        RECT 1601.820 1894.180 1602.080 1894.440 ;
        RECT 1372.280 1893.840 1372.540 1894.100 ;
        RECT 1604.120 1893.840 1604.380 1894.100 ;
        RECT 1602.740 1891.460 1603.000 1891.720 ;
        RECT 1576.520 1883.980 1576.780 1884.240 ;
        RECT 1599.980 1883.980 1600.240 1884.240 ;
        RECT 1562.720 1883.640 1562.980 1883.900 ;
        RECT 1599.060 1883.640 1599.320 1883.900 ;
        RECT 1392.980 1883.300 1393.240 1883.560 ;
        RECT 1601.820 1882.620 1602.080 1882.880 ;
        RECT 1372.280 1879.900 1372.540 1880.160 ;
        RECT 1602.740 1879.900 1603.000 1880.160 ;
        RECT 1392.060 1876.500 1392.320 1876.760 ;
        RECT 1601.360 1876.500 1601.620 1876.760 ;
        RECT 1368.140 1873.100 1368.400 1873.360 ;
        RECT 1369.060 1873.100 1369.320 1873.360 ;
        RECT 1372.280 1873.100 1372.540 1873.360 ;
        RECT 1367.680 1872.420 1367.940 1872.680 ;
        RECT 1369.060 1872.420 1369.320 1872.680 ;
        RECT 1602.740 1872.080 1603.000 1872.340 ;
        RECT 1603.200 1871.060 1603.460 1871.320 ;
        RECT 1391.600 1869.700 1391.860 1869.960 ;
        RECT 1600.900 1869.700 1601.160 1869.960 ;
        RECT 1600.440 1864.600 1600.700 1864.860 ;
        RECT 1391.140 1862.560 1391.400 1862.820 ;
        RECT 1601.820 1862.220 1602.080 1862.480 ;
        RECT 1372.280 1859.160 1372.540 1859.420 ;
        RECT 1599.520 1859.160 1599.780 1859.420 ;
        RECT 1602.740 1859.160 1603.000 1859.420 ;
        RECT 1604.120 1857.800 1604.380 1858.060 ;
        RECT 1390.680 1855.760 1390.940 1856.020 ;
        RECT 1601.360 1855.760 1601.620 1856.020 ;
        RECT 1604.120 1855.080 1604.380 1855.340 ;
        RECT 1372.280 1852.360 1372.540 1852.620 ;
        RECT 1599.980 1852.360 1600.240 1852.620 ;
        RECT 1603.200 1852.360 1603.460 1852.620 ;
        RECT 1604.120 1852.360 1604.380 1852.620 ;
        RECT 1603.200 1851.340 1603.460 1851.600 ;
        RECT 1404.020 1848.960 1404.280 1849.220 ;
        RECT 1600.900 1848.960 1601.160 1849.220 ;
        RECT 1417.820 1848.620 1418.080 1848.880 ;
        RECT 1599.060 1848.620 1599.320 1848.880 ;
        RECT 1599.980 1847.260 1600.240 1847.520 ;
        RECT 1603.200 1847.260 1603.460 1847.520 ;
        RECT 1599.520 1845.220 1599.780 1845.480 ;
        RECT 1601.820 1845.220 1602.080 1845.480 ;
        RECT 1602.280 1842.840 1602.540 1843.100 ;
        RECT 1390.220 1842.160 1390.480 1842.420 ;
        RECT 1602.280 1842.160 1602.540 1842.420 ;
        RECT 1601.360 1839.100 1601.620 1839.360 ;
        RECT 1424.720 1834.340 1424.980 1834.600 ;
        RECT 1594.000 1831.280 1594.260 1831.540 ;
        RECT 1601.820 1828.900 1602.080 1829.160 ;
        RECT 1600.900 1828.560 1601.160 1828.820 ;
        RECT 1431.620 1828.220 1431.880 1828.480 ;
        RECT 1601.820 1828.220 1602.080 1828.480 ;
        RECT 1438.520 1821.420 1438.780 1821.680 ;
        RECT 1601.360 1821.420 1601.620 1821.680 ;
        RECT 1599.980 1818.700 1600.240 1818.960 ;
        RECT 1368.600 1814.280 1368.860 1814.540 ;
        RECT 1602.280 1814.280 1602.540 1814.540 ;
        RECT 1452.320 1813.940 1452.580 1814.200 ;
        RECT 1599.060 1813.940 1599.320 1814.200 ;
        RECT 1600.440 1813.260 1600.700 1813.520 ;
        RECT 1367.680 1805.100 1367.940 1805.360 ;
        RECT 1377.340 1805.100 1377.600 1805.360 ;
        RECT 1601.360 1804.420 1601.620 1804.680 ;
        RECT 1603.660 1804.420 1603.920 1804.680 ;
        RECT 1604.120 1801.360 1604.380 1801.620 ;
        RECT 1602.280 1801.020 1602.540 1801.280 ;
        RECT 1601.360 1800.680 1601.620 1800.940 ;
        RECT 1601.360 1800.000 1601.620 1800.260 ;
        RECT 1603.660 1800.000 1603.920 1800.260 ;
        RECT 1603.660 1799.320 1603.920 1799.580 ;
        RECT 1599.980 1798.980 1600.240 1799.240 ;
        RECT 1604.120 1798.980 1604.380 1799.240 ;
        RECT 1369.060 1798.300 1369.320 1798.560 ;
        RECT 1376.880 1798.300 1377.140 1798.560 ;
        RECT 1600.900 1784.360 1601.160 1784.620 ;
        RECT 1601.820 1784.360 1602.080 1784.620 ;
        RECT 1459.220 1779.940 1459.480 1780.200 ;
        RECT 1600.900 1779.940 1601.160 1780.200 ;
        RECT 1371.820 1779.600 1372.080 1779.860 ;
        RECT 1376.420 1779.600 1376.680 1779.860 ;
        RECT 1603.200 1779.260 1603.460 1779.520 ;
        RECT 1473.020 1773.140 1473.280 1773.400 ;
        RECT 1600.900 1773.140 1601.160 1773.400 ;
        RECT 1369.060 1767.020 1369.320 1767.280 ;
        RECT 1374.120 1767.020 1374.380 1767.280 ;
        RECT 1371.360 1766.000 1371.620 1766.260 ;
        RECT 1600.900 1766.000 1601.160 1766.260 ;
        RECT 1486.820 1759.200 1487.080 1759.460 ;
        RECT 1601.360 1759.200 1601.620 1759.460 ;
        RECT 1370.900 1752.060 1371.160 1752.320 ;
        RECT 1601.360 1752.060 1601.620 1752.320 ;
        RECT 1367.680 1747.980 1367.940 1748.240 ;
        RECT 1375.040 1747.980 1375.300 1748.240 ;
        RECT 1370.440 1745.260 1370.700 1745.520 ;
        RECT 1600.900 1745.260 1601.160 1745.520 ;
        RECT 1493.720 1744.920 1493.980 1745.180 ;
        RECT 1601.820 1744.920 1602.080 1745.180 ;
        RECT 1367.680 1738.460 1367.940 1738.720 ;
        RECT 1375.500 1738.460 1375.760 1738.720 ;
        RECT 1507.520 1738.460 1507.780 1738.720 ;
        RECT 1600.900 1738.460 1601.160 1738.720 ;
        RECT 1369.980 1731.660 1370.240 1731.920 ;
        RECT 1600.900 1731.660 1601.160 1731.920 ;
        RECT 1367.680 1729.280 1367.940 1729.540 ;
        RECT 1375.960 1729.280 1376.220 1729.540 ;
        RECT 1368.140 1719.760 1368.400 1720.020 ;
        RECT 1379.640 1719.760 1379.900 1720.020 ;
        RECT 1367.680 1710.580 1367.940 1710.840 ;
        RECT 1378.720 1710.580 1378.980 1710.840 ;
        RECT 1367.680 1700.380 1367.940 1700.640 ;
        RECT 1379.180 1700.380 1379.440 1700.640 ;
        RECT 1369.060 1676.240 1369.320 1676.500 ;
        RECT 1514.420 1676.240 1514.680 1676.500 ;
        RECT 1371.360 1662.300 1371.620 1662.560 ;
        RECT 1397.120 1662.300 1397.380 1662.560 ;
        RECT 1366.760 1656.520 1367.020 1656.780 ;
        RECT 1367.680 1656.520 1367.940 1656.780 ;
        RECT 1366.760 1655.840 1367.020 1656.100 ;
        RECT 1597.220 1655.840 1597.480 1656.100 ;
        RECT 1369.980 1648.700 1370.240 1648.960 ;
        RECT 1583.420 1648.700 1583.680 1648.960 ;
        RECT 1367.680 1616.400 1367.940 1616.660 ;
        RECT 1378.260 1616.400 1378.520 1616.660 ;
        RECT 1367.220 1606.200 1367.480 1606.460 ;
        RECT 1377.800 1606.200 1378.060 1606.460 ;
      LAYER met2 ;
        RECT 392.930 3279.795 393.210 3280.165 ;
        RECT 392.470 3274.355 392.750 3274.725 ;
        RECT 392.010 3265.515 392.290 3265.885 ;
        RECT 391.550 3260.075 391.830 3260.445 ;
        RECT 391.090 3237.635 391.370 3238.005 ;
        RECT 379.130 2840.515 379.410 2840.885 ;
        RECT 379.200 2622.070 379.340 2840.515 ;
        RECT 386.030 2839.835 386.310 2840.205 ;
        RECT 373.620 2621.750 373.880 2622.070 ;
        RECT 379.140 2621.750 379.400 2622.070 ;
        RECT 354.750 2618.155 355.030 2618.525 ;
        RECT 354.820 2610.000 354.960 2618.155 ;
        RECT 373.680 2610.000 373.820 2621.750 ;
        RECT 386.100 2610.250 386.240 2839.835 ;
        RECT 390.640 2835.950 390.900 2836.270 ;
        RECT 385.640 2610.110 386.240 2610.250 ;
        RECT 354.620 2609.500 354.960 2610.000 ;
        RECT 373.480 2609.500 373.820 2610.000 ;
        RECT 383.140 2609.570 383.420 2610.000 ;
        RECT 385.640 2609.570 385.780 2610.110 ;
        RECT 354.620 2606.000 354.900 2609.500 ;
        RECT 373.480 2606.000 373.760 2609.500 ;
        RECT 383.140 2609.430 385.780 2609.570 ;
        RECT 390.700 2609.570 390.840 2835.950 ;
        RECT 391.160 2618.330 391.300 3237.635 ;
        RECT 391.620 2619.690 391.760 3260.075 ;
        RECT 391.560 2619.370 391.820 2619.690 ;
        RECT 392.080 2619.350 392.220 3265.515 ;
        RECT 392.020 2619.030 392.280 2619.350 ;
        RECT 392.540 2619.010 392.680 3274.355 ;
        RECT 392.480 2618.690 392.740 2619.010 ;
        RECT 393.000 2618.670 393.140 3279.795 ;
        RECT 393.390 3251.915 393.670 3252.285 ;
        RECT 393.460 2620.030 393.600 3251.915 ;
        RECT 393.850 3245.795 394.130 3246.165 ;
        RECT 393.920 2620.370 394.060 3245.795 ;
        RECT 394.310 2947.955 394.590 2948.325 ;
        RECT 394.380 2620.710 394.520 2947.955 ;
      LAYER met2 ;
        RECT 405.000 2855.000 781.480 3301.235 ;
      LAYER met2 ;
        RECT 938.490 3279.795 938.770 3280.165 ;
        RECT 938.560 3277.930 938.700 3279.795 ;
        RECT 783.020 3277.610 783.280 3277.930 ;
        RECT 938.500 3277.610 938.760 3277.930 ;
        RECT 516.670 2851.395 516.950 2851.765 ;
        RECT 433.870 2842.555 434.150 2842.925 ;
        RECT 509.770 2842.555 510.050 2842.925 ;
        RECT 427.440 2838.330 427.700 2838.650 ;
        RECT 406.740 2836.630 407.000 2836.950 ;
        RECT 406.800 2622.070 406.940 2836.630 ;
        RECT 413.640 2836.290 413.900 2836.610 ;
        RECT 402.140 2621.750 402.400 2622.070 ;
        RECT 406.740 2621.750 407.000 2622.070 ;
        RECT 394.320 2620.390 394.580 2620.710 ;
        RECT 393.860 2620.050 394.120 2620.370 ;
        RECT 393.400 2619.710 393.660 2620.030 ;
        RECT 392.940 2618.350 393.200 2618.670 ;
        RECT 391.100 2618.010 391.360 2618.330 ;
        RECT 402.200 2610.000 402.340 2621.750 ;
        RECT 392.340 2609.570 392.620 2610.000 ;
        RECT 390.700 2609.430 392.620 2609.570 ;
        RECT 383.140 2606.000 383.420 2609.430 ;
        RECT 392.340 2606.000 392.620 2609.430 ;
        RECT 402.000 2609.500 402.340 2610.000 ;
        RECT 411.660 2609.570 411.940 2610.000 ;
        RECT 413.700 2609.570 413.840 2836.290 ;
        RECT 427.500 2622.070 427.640 2838.330 ;
        RECT 430.660 2625.490 430.920 2625.810 ;
        RECT 421.460 2621.750 421.720 2622.070 ;
        RECT 427.440 2621.750 427.700 2622.070 ;
        RECT 421.520 2610.000 421.660 2621.750 ;
        RECT 430.720 2610.000 430.860 2625.490 ;
        RECT 433.940 2617.650 434.080 2842.555 ;
        RECT 475.730 2841.875 476.010 2842.245 ;
        RECT 455.490 2838.475 455.770 2838.845 ;
        RECT 455.500 2838.330 455.760 2838.475 ;
        RECT 475.800 2837.970 475.940 2841.875 ;
        RECT 482.630 2841.195 482.910 2841.565 ;
        RECT 482.700 2840.010 482.840 2841.195 ;
        RECT 482.640 2839.690 482.900 2840.010 ;
        RECT 489.530 2838.475 489.810 2838.845 ;
        RECT 503.330 2838.475 503.610 2838.845 ;
        RECT 489.600 2838.310 489.740 2838.475 ;
        RECT 503.340 2838.330 503.600 2838.475 ;
        RECT 489.540 2837.990 489.800 2838.310 ;
        RECT 475.740 2837.650 476.000 2837.970 ;
        RECT 441.690 2837.115 441.970 2837.485 ;
        RECT 441.760 2836.950 441.900 2837.115 ;
        RECT 434.790 2836.435 435.070 2836.805 ;
        RECT 441.700 2836.630 441.960 2836.950 ;
        RECT 449.970 2836.435 450.250 2836.805 ;
        RECT 434.860 2836.270 435.000 2836.435 ;
        RECT 449.980 2836.290 450.240 2836.435 ;
        RECT 434.800 2835.950 435.060 2836.270 ;
        RECT 468.370 2835.755 468.650 2836.125 ;
        RECT 475.270 2835.755 475.550 2836.125 ;
        RECT 482.170 2835.755 482.450 2836.125 ;
        RECT 495.970 2835.755 496.250 2836.125 ;
        RECT 459.180 2625.830 459.440 2626.150 ;
        RECT 449.980 2625.150 450.240 2625.470 ;
        RECT 440.320 2620.390 440.580 2620.710 ;
        RECT 433.880 2617.330 434.140 2617.650 ;
        RECT 440.380 2610.000 440.520 2620.390 ;
        RECT 450.040 2610.000 450.180 2625.150 ;
        RECT 459.240 2610.000 459.380 2625.830 ;
        RECT 468.440 2623.770 468.580 2835.755 ;
        RECT 468.840 2626.170 469.100 2626.490 ;
        RECT 468.380 2623.450 468.640 2623.770 ;
        RECT 468.900 2610.000 469.040 2626.170 ;
        RECT 475.340 2622.070 475.480 2835.755 ;
        RECT 478.500 2626.510 478.760 2626.830 ;
        RECT 475.280 2621.750 475.540 2622.070 ;
        RECT 478.560 2610.000 478.700 2626.510 ;
        RECT 482.240 2621.390 482.380 2835.755 ;
        RECT 488.160 2626.850 488.420 2627.170 ;
        RECT 482.180 2621.070 482.440 2621.390 ;
        RECT 488.220 2610.000 488.360 2626.850 ;
        RECT 496.040 2621.730 496.180 2835.755 ;
        RECT 507.020 2627.530 507.280 2627.850 ;
        RECT 497.360 2627.190 497.620 2627.510 ;
        RECT 495.980 2621.410 496.240 2621.730 ;
        RECT 497.420 2610.000 497.560 2627.190 ;
        RECT 507.080 2610.000 507.220 2627.530 ;
        RECT 509.840 2621.050 509.980 2842.555 ;
        RECT 510.230 2841.195 510.510 2841.565 ;
        RECT 510.300 2839.670 510.440 2841.195 ;
        RECT 510.240 2839.350 510.500 2839.670 ;
        RECT 509.780 2620.730 510.040 2621.050 ;
        RECT 516.740 2620.710 516.880 2851.395 ;
        RECT 572.330 2847.995 572.610 2848.365 ;
        RECT 600.390 2847.995 600.670 2848.365 ;
        RECT 524.030 2842.555 524.310 2842.925 ;
        RECT 526.330 2842.555 526.610 2842.925 ;
        RECT 530.930 2842.555 531.210 2842.925 ;
        RECT 537.830 2842.555 538.110 2842.925 ;
        RECT 544.730 2842.555 545.010 2842.925 ;
        RECT 558.530 2842.555 558.810 2842.925 ;
        RECT 524.100 2624.450 524.240 2842.555 ;
        RECT 526.400 2840.010 526.540 2842.555 ;
        RECT 526.340 2839.690 526.600 2840.010 ;
        RECT 524.040 2624.130 524.300 2624.450 ;
        RECT 531.000 2624.110 531.140 2842.555 ;
        RECT 537.900 2624.790 538.040 2842.555 ;
        RECT 544.800 2625.130 544.940 2842.555 ;
        RECT 549.330 2841.875 549.610 2842.245 ;
        RECT 549.400 2839.670 549.540 2841.875 ;
        RECT 549.340 2839.350 549.600 2839.670 ;
        RECT 551.630 2838.475 551.910 2838.845 ;
        RECT 551.700 2837.630 551.840 2838.475 ;
        RECT 551.640 2837.310 551.900 2837.630 ;
        RECT 558.600 2628.870 558.740 2842.555 ;
        RECT 558.540 2628.550 558.800 2628.870 ;
        RECT 544.740 2624.810 545.000 2625.130 ;
        RECT 537.840 2624.470 538.100 2624.790 ;
        RECT 530.940 2623.790 531.200 2624.110 ;
        RECT 516.680 2620.390 516.940 2620.710 ;
        RECT 545.200 2619.710 545.460 2620.030 ;
        RECT 535.540 2618.010 535.800 2618.330 ;
        RECT 516.680 2617.670 516.940 2617.990 ;
        RECT 516.740 2610.000 516.880 2617.670 ;
        RECT 525.880 2617.330 526.140 2617.650 ;
        RECT 525.940 2610.000 526.080 2617.330 ;
        RECT 535.600 2610.000 535.740 2618.010 ;
        RECT 545.260 2610.000 545.400 2619.710 ;
        RECT 572.400 2619.690 572.540 2847.995 ;
        RECT 597.170 2845.275 597.450 2845.645 ;
        RECT 573.710 2843.235 573.990 2843.605 ;
        RECT 590.270 2843.235 590.550 2843.605 ;
        RECT 573.780 2840.010 573.920 2843.235 ;
        RECT 573.720 2839.690 573.980 2840.010 ;
        RECT 590.340 2839.330 590.480 2843.235 ;
        RECT 597.240 2842.730 597.380 2845.275 ;
        RECT 597.180 2842.410 597.440 2842.730 ;
        RECT 600.460 2840.350 600.600 2847.995 ;
        RECT 604.990 2845.275 605.270 2845.645 ;
        RECT 605.060 2841.710 605.200 2845.275 ;
        RECT 613.730 2843.915 614.010 2844.285 ;
        RECT 605.000 2841.390 605.260 2841.710 ;
        RECT 600.400 2840.030 600.660 2840.350 ;
        RECT 590.280 2839.010 590.540 2839.330 ;
        RECT 613.280 2835.950 613.540 2836.270 ;
        RECT 592.570 2832.355 592.850 2832.725 ;
        RECT 592.640 2620.030 592.780 2832.355 ;
        RECT 592.580 2619.710 592.840 2620.030 ;
        RECT 554.860 2619.370 555.120 2619.690 ;
        RECT 572.340 2619.370 572.600 2619.690 ;
        RECT 554.920 2610.000 555.060 2619.370 ;
        RECT 573.720 2619.030 573.980 2619.350 ;
        RECT 564.060 2617.330 564.320 2617.650 ;
        RECT 564.120 2610.000 564.260 2617.330 ;
        RECT 573.780 2610.000 573.920 2619.030 ;
        RECT 583.380 2618.690 583.640 2619.010 ;
        RECT 583.440 2610.000 583.580 2618.690 ;
        RECT 592.580 2618.350 592.840 2618.670 ;
        RECT 592.640 2610.000 592.780 2618.350 ;
        RECT 402.000 2606.000 402.280 2609.500 ;
        RECT 411.660 2609.430 413.840 2609.570 ;
        RECT 421.320 2609.500 421.660 2610.000 ;
        RECT 430.520 2609.500 430.860 2610.000 ;
        RECT 440.180 2609.500 440.520 2610.000 ;
        RECT 449.840 2609.500 450.180 2610.000 ;
        RECT 459.040 2609.500 459.380 2610.000 ;
        RECT 468.700 2609.500 469.040 2610.000 ;
        RECT 478.360 2609.500 478.700 2610.000 ;
        RECT 488.020 2609.500 488.360 2610.000 ;
        RECT 497.220 2609.500 497.560 2610.000 ;
        RECT 506.880 2609.500 507.220 2610.000 ;
        RECT 516.540 2609.500 516.880 2610.000 ;
        RECT 525.740 2609.500 526.080 2610.000 ;
        RECT 535.400 2609.500 535.740 2610.000 ;
        RECT 545.060 2609.500 545.400 2610.000 ;
        RECT 554.720 2609.500 555.060 2610.000 ;
        RECT 563.920 2609.500 564.260 2610.000 ;
        RECT 573.580 2609.500 573.920 2610.000 ;
        RECT 583.240 2609.500 583.580 2610.000 ;
        RECT 592.440 2609.500 592.780 2610.000 ;
        RECT 611.760 2609.570 612.040 2610.000 ;
        RECT 613.340 2609.570 613.480 2835.950 ;
        RECT 613.800 2619.690 613.940 2843.915 ;
        RECT 642.250 2842.555 642.530 2842.925 ;
        RECT 642.260 2842.410 642.520 2842.555 ;
        RECT 620.630 2841.195 620.910 2841.565 ;
        RECT 621.550 2841.195 621.830 2841.565 ;
        RECT 627.530 2841.195 627.810 2841.565 ;
        RECT 620.700 2840.690 620.840 2841.195 ;
        RECT 621.560 2841.050 621.820 2841.195 ;
        RECT 620.640 2840.370 620.900 2840.690 ;
        RECT 627.600 2839.670 627.740 2841.195 ;
        RECT 642.320 2841.030 642.460 2842.410 ;
        RECT 700.220 2841.390 700.480 2841.710 ;
        RECT 642.260 2840.710 642.520 2841.030 ;
        RECT 627.540 2839.350 627.800 2839.670 ;
        RECT 693.320 2837.310 693.580 2837.630 ;
        RECT 625.230 2836.435 625.510 2836.805 ;
        RECT 627.080 2836.630 627.340 2836.950 ;
        RECT 613.740 2619.370 614.000 2619.690 ;
        RECT 621.560 2619.030 621.820 2619.350 ;
        RECT 621.620 2610.000 621.760 2619.030 ;
        RECT 625.300 2616.970 625.440 2836.435 ;
        RECT 626.610 2835.755 626.890 2836.125 ;
        RECT 626.680 2619.885 626.820 2835.755 ;
        RECT 626.610 2619.515 626.890 2619.885 ;
        RECT 627.140 2619.350 627.280 2836.630 ;
        RECT 634.430 2835.755 634.710 2836.125 ;
        RECT 640.870 2835.755 641.150 2836.125 ;
        RECT 627.080 2619.030 627.340 2619.350 ;
        RECT 634.500 2619.205 634.640 2835.755 ;
        RECT 640.940 2628.190 641.080 2835.755 ;
        RECT 640.880 2627.870 641.140 2628.190 ;
        RECT 634.430 2618.835 634.710 2619.205 ;
        RECT 650.080 2618.690 650.340 2619.010 ;
        RECT 625.240 2616.650 625.500 2616.970 ;
        RECT 650.140 2610.000 650.280 2618.690 ;
        RECT 693.380 2615.610 693.520 2837.310 ;
        RECT 700.280 2618.330 700.420 2841.390 ;
        RECT 727.810 2841.195 728.090 2841.565 ;
        RECT 720.920 2840.030 721.180 2840.350 ;
        RECT 714.020 2839.010 714.280 2839.330 ;
        RECT 700.220 2618.010 700.480 2618.330 ;
        RECT 707.120 2616.650 707.380 2616.970 ;
        RECT 693.320 2615.290 693.580 2615.610 ;
        RECT 707.180 2610.000 707.320 2616.650 ;
        RECT 714.080 2615.270 714.220 2839.010 ;
        RECT 720.980 2616.970 721.120 2840.030 ;
        RECT 727.880 2620.565 728.020 2841.195 ;
        RECT 745.300 2840.710 745.560 2841.030 ;
        RECT 734.720 2840.370 734.980 2840.690 ;
        RECT 727.810 2620.195 728.090 2620.565 ;
        RECT 734.780 2617.310 734.920 2840.370 ;
        RECT 734.720 2616.990 734.980 2617.310 ;
        RECT 720.920 2616.650 721.180 2616.970 ;
        RECT 714.020 2614.950 714.280 2615.270 ;
        RECT 745.360 2610.000 745.500 2840.710 ;
        RECT 762.320 2839.350 762.580 2839.670 ;
        RECT 754.960 2623.450 755.220 2623.770 ;
        RECT 755.020 2610.000 755.160 2623.450 ;
        RECT 762.380 2621.245 762.520 2839.350 ;
        RECT 776.120 2837.990 776.380 2838.310 ;
        RECT 769.220 2837.650 769.480 2837.970 ;
        RECT 769.280 2622.070 769.420 2837.650 ;
        RECT 776.180 2622.070 776.320 2837.990 ;
        RECT 783.080 2622.490 783.220 3277.610 ;
        RECT 941.710 3274.355 941.990 3274.725 ;
        RECT 783.940 2838.330 784.200 2838.650 ;
        RECT 780.780 2622.350 783.220 2622.490 ;
        RECT 764.160 2621.750 764.420 2622.070 ;
        RECT 769.220 2621.750 769.480 2622.070 ;
        RECT 773.820 2621.750 774.080 2622.070 ;
        RECT 776.120 2621.750 776.380 2622.070 ;
        RECT 762.310 2620.875 762.590 2621.245 ;
        RECT 764.220 2610.000 764.360 2621.750 ;
        RECT 773.880 2610.000 774.020 2621.750 ;
        RECT 779.800 2617.730 780.060 2617.990 ;
        RECT 780.780 2617.730 780.920 2622.350 ;
        RECT 782.100 2621.410 782.360 2621.730 ;
        RECT 779.800 2617.670 780.920 2617.730 ;
        RECT 779.860 2617.590 780.920 2617.670 ;
        RECT 411.660 2606.000 411.940 2609.430 ;
        RECT 421.320 2606.000 421.600 2609.500 ;
        RECT 430.520 2606.000 430.800 2609.500 ;
        RECT 440.180 2606.000 440.460 2609.500 ;
        RECT 449.840 2606.000 450.120 2609.500 ;
        RECT 459.040 2606.000 459.320 2609.500 ;
        RECT 468.700 2606.000 468.980 2609.500 ;
        RECT 478.360 2606.000 478.640 2609.500 ;
        RECT 488.020 2606.000 488.300 2609.500 ;
        RECT 497.220 2606.000 497.500 2609.500 ;
        RECT 506.880 2606.000 507.160 2609.500 ;
        RECT 516.540 2606.000 516.820 2609.500 ;
        RECT 525.740 2606.000 526.020 2609.500 ;
        RECT 535.400 2606.000 535.680 2609.500 ;
        RECT 545.060 2606.000 545.340 2609.500 ;
        RECT 554.720 2606.000 555.000 2609.500 ;
        RECT 563.920 2606.000 564.200 2609.500 ;
        RECT 573.580 2606.000 573.860 2609.500 ;
        RECT 583.240 2606.000 583.520 2609.500 ;
        RECT 592.440 2606.000 592.720 2609.500 ;
        RECT 611.760 2609.430 613.480 2609.570 ;
        RECT 621.420 2609.500 621.760 2610.000 ;
        RECT 649.940 2609.500 650.280 2610.000 ;
        RECT 706.980 2609.500 707.320 2610.000 ;
        RECT 745.160 2609.500 745.500 2610.000 ;
        RECT 754.820 2609.500 755.160 2610.000 ;
        RECT 764.020 2609.500 764.360 2610.000 ;
        RECT 773.680 2609.500 774.020 2610.000 ;
        RECT 782.160 2609.570 782.300 2621.410 ;
        RECT 784.000 2621.390 784.140 2838.330 ;
        RECT 907.220 2628.550 907.480 2628.870 ;
        RECT 878.700 2624.810 878.960 2625.130 ;
        RECT 869.040 2624.470 869.300 2624.790 ;
        RECT 850.180 2624.130 850.440 2624.450 ;
        RECT 792.680 2621.750 792.940 2622.070 ;
        RECT 812.000 2621.750 812.260 2622.070 ;
        RECT 783.940 2621.070 784.200 2621.390 ;
        RECT 792.740 2610.000 792.880 2621.750 ;
        RECT 802.340 2617.670 802.600 2617.990 ;
        RECT 802.400 2610.000 802.540 2617.670 ;
        RECT 812.060 2610.000 812.200 2621.750 ;
        RECT 821.660 2620.730 821.920 2621.050 ;
        RECT 821.720 2610.000 821.860 2620.730 ;
        RECT 840.520 2620.390 840.780 2620.710 ;
        RECT 840.580 2610.000 840.720 2620.390 ;
        RECT 850.240 2610.000 850.380 2624.130 ;
        RECT 859.840 2623.790 860.100 2624.110 ;
        RECT 859.900 2610.000 860.040 2623.790 ;
        RECT 869.100 2610.000 869.240 2624.470 ;
        RECT 878.760 2610.000 878.900 2624.810 ;
        RECT 897.560 2615.290 897.820 2615.610 ;
        RECT 897.620 2610.000 897.760 2615.290 ;
        RECT 907.280 2610.000 907.420 2628.550 ;
        RECT 941.780 2627.850 941.920 3274.355 ;
        RECT 942.170 3265.515 942.450 3265.885 ;
        RECT 941.720 2627.530 941.980 2627.850 ;
        RECT 942.240 2627.510 942.380 3265.515 ;
        RECT 942.630 3260.075 942.910 3260.445 ;
        RECT 942.180 2627.190 942.440 2627.510 ;
        RECT 942.700 2627.170 942.840 3260.075 ;
        RECT 943.090 3251.915 943.370 3252.285 ;
        RECT 942.640 2626.850 942.900 2627.170 ;
        RECT 943.160 2626.830 943.300 3251.915 ;
        RECT 943.550 3245.795 943.830 3246.165 ;
        RECT 943.100 2626.510 943.360 2626.830 ;
        RECT 943.620 2626.490 943.760 3245.795 ;
        RECT 944.010 3237.635 944.290 3238.005 ;
        RECT 943.560 2626.170 943.820 2626.490 ;
        RECT 944.080 2626.150 944.220 3237.635 ;
        RECT 944.470 2947.955 944.750 2948.325 ;
        RECT 944.020 2625.830 944.280 2626.150 ;
        RECT 944.540 2625.810 944.680 2947.955 ;
      LAYER met2 ;
        RECT 955.000 2855.000 1331.480 3301.235 ;
      LAYER met2 ;
        RECT 1103.630 2850.715 1103.910 2851.085 ;
        RECT 1089.370 2847.995 1089.650 2848.365 ;
        RECT 979.890 2842.555 980.170 2842.925 ;
        RECT 987.250 2842.555 987.530 2842.925 ;
        RECT 1020.830 2842.555 1021.110 2842.925 ;
        RECT 1024.050 2842.555 1024.330 2842.925 ;
        RECT 1027.730 2842.555 1028.010 2842.925 ;
        RECT 1065.450 2842.555 1065.730 2842.925 ;
        RECT 1070.510 2842.555 1070.790 2842.925 ;
        RECT 944.480 2625.490 944.740 2625.810 ;
        RECT 979.960 2625.470 980.100 2842.555 ;
        RECT 979.900 2625.150 980.160 2625.470 ;
        RECT 926.540 2620.050 926.800 2620.370 ;
        RECT 926.600 2610.000 926.740 2620.050 ;
        RECT 955.060 2619.710 955.320 2620.030 ;
        RECT 935.740 2615.970 936.000 2616.290 ;
        RECT 935.800 2610.000 935.940 2615.970 ;
        RECT 955.120 2610.000 955.260 2619.710 ;
        RECT 987.320 2618.525 987.460 2842.555 ;
        RECT 1018.530 2841.875 1018.810 2842.245 ;
        RECT 1018.600 2840.010 1018.740 2841.875 ;
        RECT 1018.540 2839.690 1018.800 2840.010 ;
        RECT 1018.600 2836.270 1018.740 2839.690 ;
        RECT 1018.540 2835.950 1018.800 2836.270 ;
        RECT 1020.900 2620.370 1021.040 2842.555 ;
        RECT 1024.120 2839.670 1024.260 2842.555 ;
        RECT 1024.060 2839.350 1024.320 2839.670 ;
        RECT 1024.120 2836.950 1024.260 2839.350 ;
        RECT 1024.060 2836.630 1024.320 2836.950 ;
        RECT 1021.750 2620.875 1022.030 2621.245 ;
        RECT 1020.840 2620.050 1021.100 2620.370 ;
        RECT 993.240 2619.370 993.500 2619.690 ;
        RECT 1012.090 2619.515 1012.370 2619.885 ;
        RECT 983.580 2618.010 983.840 2618.330 ;
        RECT 987.250 2618.155 987.530 2618.525 ;
        RECT 964.260 2616.990 964.520 2617.310 ;
        RECT 964.320 2610.000 964.460 2616.990 ;
        RECT 983.640 2610.000 983.780 2618.010 ;
        RECT 993.300 2610.000 993.440 2619.370 ;
        RECT 1002.440 2617.330 1002.700 2617.650 ;
        RECT 1002.500 2610.000 1002.640 2617.330 ;
        RECT 1012.160 2610.000 1012.300 2619.515 ;
        RECT 1021.820 2610.000 1021.960 2620.875 ;
        RECT 1027.800 2620.030 1027.940 2842.555 ;
        RECT 1065.520 2840.010 1065.660 2842.555 ;
        RECT 1065.460 2839.690 1065.720 2840.010 ;
        RECT 1070.580 2839.670 1070.720 2842.555 ;
        RECT 1089.440 2840.690 1089.580 2847.995 ;
        RECT 1089.380 2840.370 1089.640 2840.690 ;
        RECT 1070.520 2839.350 1070.780 2839.670 ;
        RECT 1045.280 2836.950 1045.420 2837.105 ;
        RECT 1089.440 2836.950 1089.580 2840.370 ;
        RECT 1045.220 2836.805 1045.480 2836.950 ;
        RECT 1045.210 2836.435 1045.490 2836.805 ;
        RECT 1089.380 2836.630 1089.640 2836.950 ;
        RECT 1041.530 2835.755 1041.810 2836.125 ;
        RECT 1040.620 2627.870 1040.880 2628.190 ;
        RECT 1027.740 2619.710 1028.000 2620.030 ;
        RECT 1030.950 2618.835 1031.230 2619.205 ;
        RECT 1031.020 2610.000 1031.160 2618.835 ;
        RECT 1040.680 2610.000 1040.820 2627.870 ;
        RECT 1041.600 2622.070 1041.740 2835.755 ;
        RECT 1041.540 2621.750 1041.800 2622.070 ;
        RECT 1045.280 2619.010 1045.420 2836.435 ;
        RECT 1048.430 2835.755 1048.710 2836.125 ;
        RECT 1054.870 2835.755 1055.150 2836.125 ;
        RECT 1062.230 2835.755 1062.510 2836.125 ;
        RECT 1069.130 2835.755 1069.410 2836.125 ;
        RECT 1076.030 2835.755 1076.310 2836.125 ;
        RECT 1082.930 2835.755 1083.210 2836.125 ;
        RECT 1089.370 2835.755 1089.650 2836.125 ;
        RECT 1096.730 2835.755 1097.010 2836.125 ;
        RECT 1048.500 2621.390 1048.640 2835.755 ;
        RECT 1048.440 2621.070 1048.700 2621.390 ;
        RECT 1050.270 2620.195 1050.550 2620.565 ;
        RECT 1045.220 2618.690 1045.480 2619.010 ;
        RECT 1050.340 2610.000 1050.480 2620.195 ;
        RECT 1054.940 2619.350 1055.080 2835.755 ;
        RECT 1062.300 2621.050 1062.440 2835.755 ;
        RECT 1069.200 2621.130 1069.340 2835.755 ;
        RECT 1062.240 2620.730 1062.500 2621.050 ;
        RECT 1069.200 2620.990 1069.800 2621.130 ;
        RECT 1069.660 2620.370 1069.800 2620.990 ;
        RECT 1069.140 2620.050 1069.400 2620.370 ;
        RECT 1069.600 2620.050 1069.860 2620.370 ;
        RECT 1054.880 2619.030 1055.140 2619.350 ;
        RECT 1069.200 2610.000 1069.340 2620.050 ;
        RECT 1076.100 2619.690 1076.240 2835.755 ;
        RECT 1083.000 2620.030 1083.140 2835.755 ;
        RECT 1078.800 2619.710 1079.060 2620.030 ;
        RECT 1082.940 2619.710 1083.200 2620.030 ;
        RECT 1076.040 2619.370 1076.300 2619.690 ;
        RECT 1078.860 2610.000 1079.000 2619.710 ;
        RECT 1089.440 2618.670 1089.580 2835.755 ;
        RECT 1096.800 2619.010 1096.940 2835.755 ;
        RECT 1097.660 2621.750 1097.920 2622.070 ;
        RECT 1096.740 2618.690 1097.000 2619.010 ;
        RECT 1089.380 2618.350 1089.640 2618.670 ;
        RECT 1097.720 2610.000 1097.860 2621.750 ;
        RECT 1103.700 2616.630 1103.840 2850.715 ;
        RECT 1111.910 2842.555 1112.190 2842.925 ;
        RECT 1118.350 2842.555 1118.630 2842.925 ;
        RECT 1131.230 2842.555 1131.510 2842.925 ;
        RECT 1135.830 2842.555 1136.110 2842.925 ;
        RECT 1138.130 2842.555 1138.410 2842.925 ;
        RECT 1145.030 2842.555 1145.310 2842.925 ;
        RECT 1151.930 2842.555 1152.210 2842.925 ;
        RECT 1158.830 2842.555 1159.110 2842.925 ;
        RECT 1165.270 2842.555 1165.550 2842.925 ;
        RECT 1172.630 2842.555 1172.910 2842.925 ;
        RECT 1179.530 2842.555 1179.810 2842.925 ;
        RECT 1186.430 2842.555 1186.710 2842.925 ;
        RECT 1193.330 2842.555 1193.610 2842.925 ;
        RECT 1111.980 2840.010 1112.120 2842.555 ;
        RECT 1111.920 2839.690 1112.180 2840.010 ;
        RECT 1118.420 2839.670 1118.560 2842.555 ;
        RECT 1130.770 2841.875 1131.050 2842.245 ;
        RECT 1118.360 2839.350 1118.620 2839.670 ;
        RECT 1110.530 2835.755 1110.810 2836.125 ;
        RECT 1117.430 2835.755 1117.710 2836.125 ;
        RECT 1124.330 2835.755 1124.610 2836.125 ;
        RECT 1107.320 2621.070 1107.580 2621.390 ;
        RECT 1103.640 2616.310 1103.900 2616.630 ;
        RECT 1107.380 2610.000 1107.520 2621.070 ;
        RECT 1110.600 2616.970 1110.740 2835.755 ;
        RECT 1117.500 2617.650 1117.640 2835.755 ;
        RECT 1117.440 2617.330 1117.700 2617.650 ;
        RECT 1124.400 2617.310 1124.540 2835.755 ;
        RECT 1126.640 2620.390 1126.900 2620.710 ;
        RECT 1124.340 2616.990 1124.600 2617.310 ;
        RECT 1110.540 2616.650 1110.800 2616.970 ;
        RECT 1126.700 2610.000 1126.840 2620.390 ;
        RECT 1130.840 2617.990 1130.980 2841.875 ;
        RECT 1131.300 2618.330 1131.440 2842.555 ;
        RECT 1135.900 2840.690 1136.040 2842.555 ;
        RECT 1135.840 2840.370 1136.100 2840.690 ;
        RECT 1138.200 2621.730 1138.340 2842.555 ;
        RECT 1145.100 2622.070 1145.240 2842.555 ;
        RECT 1145.040 2621.750 1145.300 2622.070 ;
        RECT 1138.140 2621.410 1138.400 2621.730 ;
        RECT 1152.000 2621.050 1152.140 2842.555 ;
        RECT 1158.900 2621.390 1159.040 2842.555 ;
        RECT 1159.750 2840.515 1160.030 2840.885 ;
        RECT 1159.290 2839.835 1159.570 2840.205 ;
        RECT 1159.300 2839.690 1159.560 2839.835 ;
        RECT 1159.820 2839.670 1159.960 2840.515 ;
        RECT 1159.760 2839.350 1160.020 2839.670 ;
        RECT 1158.840 2621.070 1159.100 2621.390 ;
        RECT 1135.840 2620.730 1136.100 2621.050 ;
        RECT 1151.940 2620.730 1152.200 2621.050 ;
        RECT 1131.240 2618.010 1131.500 2618.330 ;
        RECT 1130.780 2617.670 1131.040 2617.990 ;
        RECT 1135.900 2610.000 1136.040 2620.730 ;
        RECT 1145.500 2620.050 1145.760 2620.370 ;
        RECT 1145.560 2610.000 1145.700 2620.050 ;
        RECT 1164.360 2619.710 1164.620 2620.030 ;
        RECT 1155.160 2619.370 1155.420 2619.690 ;
        RECT 1155.220 2610.000 1155.360 2619.370 ;
        RECT 1164.420 2610.000 1164.560 2619.710 ;
        RECT 1165.340 2619.690 1165.480 2842.555 ;
        RECT 1165.730 2841.875 1166.010 2842.245 ;
        RECT 1165.800 2620.710 1165.940 2841.875 ;
        RECT 1165.740 2620.390 1166.000 2620.710 ;
        RECT 1172.700 2620.370 1172.840 2842.555 ;
        RECT 1172.640 2620.050 1172.900 2620.370 ;
        RECT 1179.600 2620.030 1179.740 2842.555 ;
        RECT 1179.990 2840.515 1180.270 2840.885 ;
        RECT 1180.000 2840.370 1180.260 2840.515 ;
        RECT 1179.540 2619.710 1179.800 2620.030 ;
        RECT 1186.500 2619.690 1186.640 2842.555 ;
        RECT 1165.280 2619.370 1165.540 2619.690 ;
        RECT 1186.440 2619.370 1186.700 2619.690 ;
        RECT 1193.400 2619.350 1193.540 2842.555 ;
        RECT 1269.240 2621.750 1269.500 2622.070 ;
        RECT 1260.040 2621.410 1260.300 2621.730 ;
        RECT 1193.340 2619.030 1193.600 2619.350 ;
        RECT 1191.500 2618.690 1191.760 2619.010 ;
        RECT 1183.680 2618.350 1183.940 2618.670 ;
        RECT 1183.740 2610.000 1183.880 2618.350 ;
        RECT 783.340 2609.570 783.620 2610.000 ;
        RECT 611.760 2606.000 612.040 2609.430 ;
        RECT 621.420 2606.000 621.700 2609.500 ;
        RECT 649.940 2606.000 650.220 2609.500 ;
        RECT 706.980 2606.000 707.260 2609.500 ;
        RECT 745.160 2606.000 745.440 2609.500 ;
        RECT 754.820 2606.000 755.100 2609.500 ;
        RECT 764.020 2606.000 764.300 2609.500 ;
        RECT 773.680 2606.000 773.960 2609.500 ;
        RECT 782.160 2609.430 783.620 2609.570 ;
        RECT 783.340 2606.000 783.620 2609.430 ;
        RECT 792.540 2609.500 792.880 2610.000 ;
        RECT 802.200 2609.500 802.540 2610.000 ;
        RECT 811.860 2609.500 812.200 2610.000 ;
        RECT 821.520 2609.500 821.860 2610.000 ;
        RECT 840.380 2609.500 840.720 2610.000 ;
        RECT 850.040 2609.500 850.380 2610.000 ;
        RECT 859.700 2609.500 860.040 2610.000 ;
        RECT 868.900 2609.500 869.240 2610.000 ;
        RECT 878.560 2609.500 878.900 2610.000 ;
        RECT 897.420 2609.500 897.760 2610.000 ;
        RECT 907.080 2609.500 907.420 2610.000 ;
        RECT 926.400 2609.500 926.740 2610.000 ;
        RECT 935.600 2609.500 935.940 2610.000 ;
        RECT 954.920 2609.500 955.260 2610.000 ;
        RECT 964.120 2609.500 964.460 2610.000 ;
        RECT 983.440 2609.500 983.780 2610.000 ;
        RECT 993.100 2609.500 993.440 2610.000 ;
        RECT 1002.300 2609.500 1002.640 2610.000 ;
        RECT 1011.960 2609.500 1012.300 2610.000 ;
        RECT 1021.620 2609.500 1021.960 2610.000 ;
        RECT 1030.820 2609.500 1031.160 2610.000 ;
        RECT 1040.480 2609.500 1040.820 2610.000 ;
        RECT 1050.140 2609.500 1050.480 2610.000 ;
        RECT 1069.000 2609.500 1069.340 2610.000 ;
        RECT 1078.660 2609.500 1079.000 2610.000 ;
        RECT 1097.520 2609.500 1097.860 2610.000 ;
        RECT 1107.180 2609.500 1107.520 2610.000 ;
        RECT 1126.500 2609.500 1126.840 2610.000 ;
        RECT 1135.700 2609.500 1136.040 2610.000 ;
        RECT 1145.360 2609.500 1145.700 2610.000 ;
        RECT 1155.020 2609.500 1155.360 2610.000 ;
        RECT 1164.220 2609.500 1164.560 2610.000 ;
        RECT 1183.540 2609.500 1183.880 2610.000 ;
        RECT 1191.560 2609.570 1191.700 2618.690 ;
        RECT 1250.380 2618.010 1250.640 2618.330 ;
        RECT 1240.720 2617.670 1240.980 2617.990 ;
        RECT 1221.860 2617.330 1222.120 2617.650 ;
        RECT 1212.200 2616.650 1212.460 2616.970 ;
        RECT 1202.540 2616.310 1202.800 2616.630 ;
        RECT 1202.600 2610.000 1202.740 2616.310 ;
        RECT 1212.260 2610.000 1212.400 2616.650 ;
        RECT 1221.920 2610.000 1222.060 2617.330 ;
        RECT 1231.060 2616.990 1231.320 2617.310 ;
        RECT 1231.120 2610.000 1231.260 2616.990 ;
        RECT 1240.780 2610.000 1240.920 2617.670 ;
        RECT 1250.440 2610.000 1250.580 2618.010 ;
        RECT 1260.100 2610.000 1260.240 2621.410 ;
        RECT 1269.300 2610.000 1269.440 2621.750 ;
        RECT 1288.560 2621.070 1288.820 2621.390 ;
        RECT 1278.900 2620.730 1279.160 2621.050 ;
        RECT 1278.960 2610.000 1279.100 2620.730 ;
        RECT 1288.620 2610.000 1288.760 2621.070 ;
        RECT 1297.760 2620.390 1298.020 2620.710 ;
        RECT 1297.820 2610.000 1297.960 2620.390 ;
        RECT 1317.080 2620.050 1317.340 2620.370 ;
        RECT 1307.420 2619.710 1307.680 2620.030 ;
        RECT 1307.480 2610.000 1307.620 2619.710 ;
        RECT 1317.140 2610.000 1317.280 2620.050 ;
        RECT 1335.940 2619.370 1336.200 2619.690 ;
        RECT 1326.740 2619.030 1327.000 2619.350 ;
        RECT 1326.800 2610.000 1326.940 2619.030 ;
        RECT 1336.000 2610.000 1336.140 2619.370 ;
        RECT 1345.600 2618.690 1345.860 2619.010 ;
        RECT 1345.660 2610.000 1345.800 2618.690 ;
        RECT 1193.200 2609.570 1193.480 2610.000 ;
        RECT 792.540 2606.000 792.820 2609.500 ;
        RECT 802.200 2606.000 802.480 2609.500 ;
        RECT 811.860 2606.000 812.140 2609.500 ;
        RECT 821.520 2606.000 821.800 2609.500 ;
        RECT 840.380 2606.000 840.660 2609.500 ;
        RECT 850.040 2606.000 850.320 2609.500 ;
        RECT 859.700 2606.000 859.980 2609.500 ;
        RECT 868.900 2606.000 869.180 2609.500 ;
        RECT 878.560 2606.000 878.840 2609.500 ;
        RECT 897.420 2606.000 897.700 2609.500 ;
        RECT 907.080 2606.000 907.360 2609.500 ;
        RECT 926.400 2606.000 926.680 2609.500 ;
        RECT 935.600 2606.000 935.880 2609.500 ;
        RECT 954.920 2606.000 955.200 2609.500 ;
        RECT 964.120 2606.000 964.400 2609.500 ;
        RECT 983.440 2606.000 983.720 2609.500 ;
        RECT 993.100 2606.000 993.380 2609.500 ;
        RECT 1002.300 2606.000 1002.580 2609.500 ;
        RECT 1011.960 2606.000 1012.240 2609.500 ;
        RECT 1021.620 2606.000 1021.900 2609.500 ;
        RECT 1030.820 2606.000 1031.100 2609.500 ;
        RECT 1040.480 2606.000 1040.760 2609.500 ;
        RECT 1050.140 2606.000 1050.420 2609.500 ;
        RECT 1069.000 2606.000 1069.280 2609.500 ;
        RECT 1078.660 2606.000 1078.940 2609.500 ;
        RECT 1097.520 2606.000 1097.800 2609.500 ;
        RECT 1107.180 2606.000 1107.460 2609.500 ;
        RECT 1126.500 2606.000 1126.780 2609.500 ;
        RECT 1135.700 2606.000 1135.980 2609.500 ;
        RECT 1145.360 2606.000 1145.640 2609.500 ;
        RECT 1155.020 2606.000 1155.300 2609.500 ;
        RECT 1164.220 2606.000 1164.500 2609.500 ;
        RECT 1183.540 2606.000 1183.820 2609.500 ;
        RECT 1191.560 2609.430 1193.480 2609.570 ;
        RECT 1193.200 2606.000 1193.480 2609.430 ;
        RECT 1202.400 2609.500 1202.740 2610.000 ;
        RECT 1212.060 2609.500 1212.400 2610.000 ;
        RECT 1221.720 2609.500 1222.060 2610.000 ;
        RECT 1230.920 2609.500 1231.260 2610.000 ;
        RECT 1240.580 2609.500 1240.920 2610.000 ;
        RECT 1250.240 2609.500 1250.580 2610.000 ;
        RECT 1259.900 2609.500 1260.240 2610.000 ;
        RECT 1269.100 2609.500 1269.440 2610.000 ;
        RECT 1278.760 2609.500 1279.100 2610.000 ;
        RECT 1288.420 2609.500 1288.760 2610.000 ;
        RECT 1297.620 2609.500 1297.960 2610.000 ;
        RECT 1307.280 2609.500 1307.620 2610.000 ;
        RECT 1316.940 2609.500 1317.280 2610.000 ;
        RECT 1326.600 2609.500 1326.940 2610.000 ;
        RECT 1335.800 2609.500 1336.140 2610.000 ;
        RECT 1345.460 2609.500 1345.800 2610.000 ;
        RECT 1202.400 2606.000 1202.680 2609.500 ;
        RECT 1212.060 2606.000 1212.340 2609.500 ;
        RECT 1221.720 2606.000 1222.000 2609.500 ;
        RECT 1230.920 2606.000 1231.200 2609.500 ;
        RECT 1240.580 2606.000 1240.860 2609.500 ;
        RECT 1250.240 2606.000 1250.520 2609.500 ;
        RECT 1259.900 2606.000 1260.180 2609.500 ;
        RECT 1269.100 2606.000 1269.380 2609.500 ;
        RECT 1278.760 2606.000 1279.040 2609.500 ;
        RECT 1288.420 2606.000 1288.700 2609.500 ;
        RECT 1297.620 2606.000 1297.900 2609.500 ;
        RECT 1307.280 2606.000 1307.560 2609.500 ;
        RECT 1316.940 2606.000 1317.220 2609.500 ;
        RECT 1326.600 2606.000 1326.880 2609.500 ;
        RECT 1335.800 2606.000 1336.080 2609.500 ;
        RECT 1345.460 2606.000 1345.740 2609.500 ;
      LAYER met2 ;
        RECT 350.030 2605.720 354.340 2606.000 ;
        RECT 355.180 2605.720 363.540 2606.000 ;
        RECT 364.380 2605.720 373.200 2606.000 ;
        RECT 374.040 2605.720 382.860 2606.000 ;
        RECT 383.700 2605.720 392.060 2606.000 ;
        RECT 392.900 2605.720 401.720 2606.000 ;
        RECT 402.560 2605.720 411.380 2606.000 ;
        RECT 412.220 2605.720 421.040 2606.000 ;
        RECT 421.880 2605.720 430.240 2606.000 ;
        RECT 431.080 2605.720 439.900 2606.000 ;
        RECT 440.740 2605.720 449.560 2606.000 ;
        RECT 450.400 2605.720 458.760 2606.000 ;
        RECT 459.600 2605.720 468.420 2606.000 ;
        RECT 469.260 2605.720 478.080 2606.000 ;
        RECT 478.920 2605.720 487.740 2606.000 ;
        RECT 488.580 2605.720 496.940 2606.000 ;
        RECT 497.780 2605.720 506.600 2606.000 ;
        RECT 507.440 2605.720 516.260 2606.000 ;
        RECT 517.100 2605.720 525.460 2606.000 ;
        RECT 526.300 2605.720 535.120 2606.000 ;
        RECT 535.960 2605.720 544.780 2606.000 ;
        RECT 545.620 2605.720 554.440 2606.000 ;
        RECT 555.280 2605.720 563.640 2606.000 ;
        RECT 564.480 2605.720 573.300 2606.000 ;
        RECT 574.140 2605.720 582.960 2606.000 ;
        RECT 583.800 2605.720 592.160 2606.000 ;
        RECT 593.000 2605.720 601.820 2606.000 ;
        RECT 602.660 2605.720 611.480 2606.000 ;
        RECT 612.320 2605.720 621.140 2606.000 ;
        RECT 621.980 2605.720 630.340 2606.000 ;
        RECT 631.180 2605.720 640.000 2606.000 ;
        RECT 640.840 2605.720 649.660 2606.000 ;
        RECT 650.500 2605.720 658.860 2606.000 ;
        RECT 659.700 2605.720 668.520 2606.000 ;
        RECT 669.360 2605.720 678.180 2606.000 ;
        RECT 679.020 2605.720 687.840 2606.000 ;
        RECT 688.680 2605.720 697.040 2606.000 ;
        RECT 697.880 2605.720 706.700 2606.000 ;
        RECT 707.540 2605.720 716.360 2606.000 ;
        RECT 717.200 2605.720 725.560 2606.000 ;
        RECT 726.400 2605.720 735.220 2606.000 ;
        RECT 736.060 2605.720 744.880 2606.000 ;
        RECT 745.720 2605.720 754.540 2606.000 ;
        RECT 755.380 2605.720 763.740 2606.000 ;
        RECT 764.580 2605.720 773.400 2606.000 ;
        RECT 774.240 2605.720 783.060 2606.000 ;
        RECT 783.900 2605.720 792.260 2606.000 ;
        RECT 793.100 2605.720 801.920 2606.000 ;
        RECT 802.760 2605.720 811.580 2606.000 ;
        RECT 812.420 2605.720 821.240 2606.000 ;
        RECT 822.080 2605.720 830.440 2606.000 ;
        RECT 831.280 2605.720 840.100 2606.000 ;
        RECT 840.940 2605.720 849.760 2606.000 ;
        RECT 850.600 2605.720 859.420 2606.000 ;
        RECT 860.260 2605.720 868.620 2606.000 ;
        RECT 869.460 2605.720 878.280 2606.000 ;
        RECT 879.120 2605.720 887.940 2606.000 ;
        RECT 888.780 2605.720 897.140 2606.000 ;
        RECT 897.980 2605.720 906.800 2606.000 ;
        RECT 907.640 2605.720 916.460 2606.000 ;
        RECT 917.300 2605.720 926.120 2606.000 ;
        RECT 926.960 2605.720 935.320 2606.000 ;
        RECT 936.160 2605.720 944.980 2606.000 ;
        RECT 945.820 2605.720 954.640 2606.000 ;
        RECT 955.480 2605.720 963.840 2606.000 ;
        RECT 964.680 2605.720 973.500 2606.000 ;
        RECT 974.340 2605.720 983.160 2606.000 ;
        RECT 984.000 2605.720 992.820 2606.000 ;
        RECT 993.660 2605.720 1002.020 2606.000 ;
        RECT 1002.860 2605.720 1011.680 2606.000 ;
        RECT 1012.520 2605.720 1021.340 2606.000 ;
        RECT 1022.180 2605.720 1030.540 2606.000 ;
        RECT 1031.380 2605.720 1040.200 2606.000 ;
        RECT 1041.040 2605.720 1049.860 2606.000 ;
        RECT 1050.700 2605.720 1059.520 2606.000 ;
        RECT 1060.360 2605.720 1068.720 2606.000 ;
        RECT 1069.560 2605.720 1078.380 2606.000 ;
        RECT 1079.220 2605.720 1088.040 2606.000 ;
        RECT 1088.880 2605.720 1097.240 2606.000 ;
        RECT 1098.080 2605.720 1106.900 2606.000 ;
        RECT 1107.740 2605.720 1116.560 2606.000 ;
        RECT 1117.400 2605.720 1126.220 2606.000 ;
        RECT 1127.060 2605.720 1135.420 2606.000 ;
        RECT 1136.260 2605.720 1145.080 2606.000 ;
        RECT 1145.920 2605.720 1154.740 2606.000 ;
        RECT 1155.580 2605.720 1163.940 2606.000 ;
        RECT 1164.780 2605.720 1173.600 2606.000 ;
        RECT 1174.440 2605.720 1183.260 2606.000 ;
        RECT 1184.100 2605.720 1192.920 2606.000 ;
        RECT 1193.760 2605.720 1202.120 2606.000 ;
        RECT 1202.960 2605.720 1211.780 2606.000 ;
        RECT 1212.620 2605.720 1221.440 2606.000 ;
        RECT 1222.280 2605.720 1230.640 2606.000 ;
        RECT 1231.480 2605.720 1240.300 2606.000 ;
        RECT 1241.140 2605.720 1249.960 2606.000 ;
        RECT 1250.800 2605.720 1259.620 2606.000 ;
        RECT 1260.460 2605.720 1268.820 2606.000 ;
        RECT 1269.660 2605.720 1278.480 2606.000 ;
        RECT 1279.320 2605.720 1288.140 2606.000 ;
        RECT 1288.980 2605.720 1297.340 2606.000 ;
        RECT 1298.180 2605.720 1307.000 2606.000 ;
        RECT 1307.840 2605.720 1316.660 2606.000 ;
        RECT 1317.500 2605.720 1326.320 2606.000 ;
        RECT 1327.160 2605.720 1335.520 2606.000 ;
        RECT 1336.360 2605.720 1345.180 2606.000 ;
        RECT 1346.020 2605.720 1354.840 2606.000 ;
        RECT 1355.680 2605.720 1357.230 2606.000 ;
        RECT 350.030 1604.280 1357.230 2605.720 ;
      LAYER met2 ;
        RECT 1369.970 2604.555 1370.250 2604.925 ;
        RECT 1369.520 2583.670 1369.780 2583.990 ;
        RECT 1369.060 2581.630 1369.320 2581.950 ;
        RECT 1368.130 2575.995 1368.410 2576.365 ;
        RECT 1368.200 2574.130 1368.340 2575.995 ;
        RECT 1368.140 2573.810 1368.400 2574.130 ;
        RECT 1367.670 2556.955 1367.950 2557.325 ;
        RECT 1367.740 2553.390 1367.880 2556.955 ;
        RECT 1367.680 2553.070 1367.940 2553.390 ;
        RECT 1368.590 2537.915 1368.870 2538.285 ;
        RECT 1368.660 2532.990 1368.800 2537.915 ;
        RECT 1368.600 2532.670 1368.860 2532.990 ;
        RECT 1367.670 2528.395 1367.950 2528.765 ;
        RECT 1367.740 2526.190 1367.880 2528.395 ;
        RECT 1367.680 2525.870 1367.940 2526.190 ;
        RECT 1367.670 2518.875 1367.950 2519.245 ;
        RECT 1367.740 2477.650 1367.880 2518.875 ;
        RECT 1368.130 2509.355 1368.410 2509.725 ;
        RECT 1368.200 2505.450 1368.340 2509.355 ;
        RECT 1368.140 2505.130 1368.400 2505.450 ;
        RECT 1368.590 2499.835 1368.870 2500.205 ;
        RECT 1368.660 2498.310 1368.800 2499.835 ;
        RECT 1368.600 2497.990 1368.860 2498.310 ;
        RECT 1368.590 2490.315 1368.870 2490.685 ;
        RECT 1368.660 2484.710 1368.800 2490.315 ;
        RECT 1368.600 2484.390 1368.860 2484.710 ;
        RECT 1368.590 2480.795 1368.870 2481.165 ;
        RECT 1368.660 2478.250 1368.800 2480.795 ;
        RECT 1368.600 2477.930 1368.860 2478.250 ;
        RECT 1367.740 2477.510 1368.800 2477.650 ;
        RECT 1368.130 2471.275 1368.410 2471.645 ;
        RECT 1368.200 2470.770 1368.340 2471.275 ;
        RECT 1368.140 2470.450 1368.400 2470.770 ;
        RECT 1368.130 2461.755 1368.410 2462.125 ;
        RECT 1368.200 2457.170 1368.340 2461.755 ;
        RECT 1368.140 2456.850 1368.400 2457.170 ;
        RECT 1367.210 2452.235 1367.490 2452.605 ;
        RECT 1367.280 2450.030 1367.420 2452.235 ;
        RECT 1367.220 2449.710 1367.480 2450.030 ;
        RECT 1368.140 2443.250 1368.400 2443.570 ;
        RECT 1368.200 2443.085 1368.340 2443.250 ;
        RECT 1368.130 2442.715 1368.410 2443.085 ;
        RECT 1367.670 2433.195 1367.950 2433.565 ;
        RECT 1367.740 2429.630 1367.880 2433.195 ;
        RECT 1367.680 2429.310 1367.940 2429.630 ;
        RECT 1368.130 2423.675 1368.410 2424.045 ;
        RECT 1368.200 2422.490 1368.340 2423.675 ;
        RECT 1368.140 2422.170 1368.400 2422.490 ;
        RECT 1368.130 2414.155 1368.410 2414.525 ;
        RECT 1368.200 2408.890 1368.340 2414.155 ;
        RECT 1368.140 2408.570 1368.400 2408.890 ;
        RECT 1368.130 2404.635 1368.410 2405.005 ;
        RECT 1368.200 2401.750 1368.340 2404.635 ;
        RECT 1368.140 2401.430 1368.400 2401.750 ;
        RECT 1368.130 2395.115 1368.410 2395.485 ;
        RECT 1368.200 2394.610 1368.340 2395.115 ;
        RECT 1368.140 2394.290 1368.400 2394.610 ;
        RECT 1368.130 2385.595 1368.410 2385.965 ;
        RECT 1368.200 2380.670 1368.340 2385.595 ;
        RECT 1368.140 2380.350 1368.400 2380.670 ;
        RECT 1368.130 2376.075 1368.410 2376.445 ;
        RECT 1368.200 2374.210 1368.340 2376.075 ;
        RECT 1368.140 2373.890 1368.400 2374.210 ;
        RECT 1367.680 2369.810 1367.940 2370.130 ;
        RECT 1367.740 2361.370 1367.880 2369.810 ;
        RECT 1368.140 2366.925 1368.400 2367.070 ;
        RECT 1368.130 2366.555 1368.410 2366.925 ;
        RECT 1367.740 2361.230 1368.340 2361.370 ;
        RECT 1367.220 2359.950 1367.480 2360.270 ;
        RECT 1366.760 2352.810 1367.020 2353.130 ;
        RECT 1366.290 2318.955 1366.570 2319.325 ;
        RECT 1366.360 2318.790 1366.500 2318.955 ;
        RECT 1366.300 2318.470 1366.560 2318.790 ;
        RECT 1366.290 2309.435 1366.570 2309.805 ;
        RECT 1366.360 2304.850 1366.500 2309.435 ;
        RECT 1366.300 2304.530 1366.560 2304.850 ;
        RECT 1366.300 2300.285 1366.560 2300.430 ;
        RECT 1366.290 2299.915 1366.570 2300.285 ;
        RECT 1366.300 2290.765 1366.560 2290.910 ;
        RECT 1366.290 2290.395 1366.570 2290.765 ;
        RECT 1366.300 2281.245 1366.560 2281.390 ;
        RECT 1366.290 2280.875 1366.570 2281.245 ;
        RECT 1366.300 2271.725 1366.560 2271.870 ;
        RECT 1366.290 2271.355 1366.570 2271.725 ;
        RECT 1366.300 2262.205 1366.560 2262.350 ;
        RECT 1366.290 2261.835 1366.570 2262.205 ;
        RECT 1366.820 2252.685 1366.960 2352.810 ;
        RECT 1366.750 2252.315 1367.030 2252.685 ;
        RECT 1367.280 2243.165 1367.420 2359.950 ;
        RECT 1367.670 2357.035 1367.950 2357.405 ;
        RECT 1367.740 2353.470 1367.880 2357.035 ;
        RECT 1367.680 2353.150 1367.940 2353.470 ;
        RECT 1367.670 2347.515 1367.950 2347.885 ;
        RECT 1367.740 2346.670 1367.880 2347.515 ;
        RECT 1367.680 2346.350 1367.940 2346.670 ;
        RECT 1367.670 2337.995 1367.950 2338.365 ;
        RECT 1367.740 2332.730 1367.880 2337.995 ;
        RECT 1367.680 2332.410 1367.940 2332.730 ;
        RECT 1367.670 2328.475 1367.950 2328.845 ;
        RECT 1367.210 2242.795 1367.490 2243.165 ;
        RECT 1367.220 2235.170 1367.480 2235.490 ;
        RECT 1367.280 2233.645 1367.420 2235.170 ;
        RECT 1367.210 2233.275 1367.490 2233.645 ;
        RECT 1367.220 2224.125 1367.480 2224.270 ;
        RECT 1367.210 2223.755 1367.490 2224.125 ;
        RECT 1367.220 2214.605 1367.480 2214.750 ;
        RECT 1367.210 2214.235 1367.490 2214.605 ;
        RECT 1367.220 2206.270 1367.480 2206.590 ;
        RECT 1367.280 2205.085 1367.420 2206.270 ;
        RECT 1367.210 2204.715 1367.490 2205.085 ;
        RECT 1367.220 2198.450 1367.480 2198.770 ;
        RECT 1367.280 2195.565 1367.420 2198.450 ;
        RECT 1367.210 2195.195 1367.490 2195.565 ;
        RECT 1366.300 2167.005 1366.560 2167.150 ;
        RECT 1366.290 2166.635 1366.570 2167.005 ;
        RECT 1366.300 2157.485 1366.560 2157.630 ;
        RECT 1366.290 2157.115 1366.570 2157.485 ;
        RECT 1366.300 2147.965 1366.560 2148.110 ;
        RECT 1366.290 2147.595 1366.570 2147.965 ;
        RECT 1366.300 2138.445 1366.560 2138.590 ;
        RECT 1366.290 2138.075 1366.570 2138.445 ;
        RECT 1366.300 2128.925 1366.560 2129.070 ;
        RECT 1366.290 2128.555 1366.570 2128.925 ;
        RECT 1367.220 2119.910 1367.480 2120.230 ;
        RECT 1367.280 2119.405 1367.420 2119.910 ;
        RECT 1367.210 2119.035 1367.490 2119.405 ;
        RECT 1367.220 2110.050 1367.480 2110.370 ;
        RECT 1367.280 2109.885 1367.420 2110.050 ;
        RECT 1367.210 2109.515 1367.490 2109.885 ;
        RECT 1367.220 2100.365 1367.480 2100.510 ;
        RECT 1367.210 2099.995 1367.490 2100.365 ;
        RECT 1367.210 2090.475 1367.490 2090.845 ;
        RECT 1367.220 2090.330 1367.480 2090.475 ;
        RECT 1367.220 2081.325 1367.480 2081.470 ;
        RECT 1367.210 2080.955 1367.490 2081.325 ;
        RECT 1367.220 2071.805 1367.480 2071.950 ;
        RECT 1367.210 2071.435 1367.490 2071.805 ;
        RECT 1367.220 2062.285 1367.480 2062.430 ;
        RECT 1367.210 2061.915 1367.490 2062.285 ;
        RECT 1367.220 2052.765 1367.480 2052.910 ;
        RECT 1367.210 2052.395 1367.490 2052.765 ;
        RECT 1367.220 2043.245 1367.480 2043.390 ;
        RECT 1367.210 2042.875 1367.490 2043.245 ;
        RECT 1367.220 2033.725 1367.480 2033.870 ;
        RECT 1367.210 2033.355 1367.490 2033.725 ;
        RECT 1367.220 2014.685 1367.480 2014.830 ;
        RECT 1367.210 2014.315 1367.490 2014.685 ;
        RECT 1367.220 2005.165 1367.480 2005.310 ;
        RECT 1367.210 2004.795 1367.490 2005.165 ;
        RECT 1367.220 2000.570 1367.480 2000.890 ;
        RECT 1367.280 1995.645 1367.420 2000.570 ;
        RECT 1367.210 1995.275 1367.490 1995.645 ;
        RECT 1367.220 1986.970 1367.480 1987.290 ;
        RECT 1367.280 1986.125 1367.420 1986.970 ;
        RECT 1367.210 1985.755 1367.490 1986.125 ;
        RECT 1366.300 1983.910 1366.560 1984.230 ;
        RECT 1366.360 1681.485 1366.500 1983.910 ;
        RECT 1367.220 1979.830 1367.480 1980.150 ;
        RECT 1367.280 1976.605 1367.420 1979.830 ;
        RECT 1367.210 1976.235 1367.490 1976.605 ;
        RECT 1367.220 1973.030 1367.480 1973.350 ;
        RECT 1367.280 1967.085 1367.420 1973.030 ;
        RECT 1367.210 1966.715 1367.490 1967.085 ;
        RECT 1367.220 1959.430 1367.480 1959.750 ;
        RECT 1367.280 1957.565 1367.420 1959.430 ;
        RECT 1367.210 1957.195 1367.490 1957.565 ;
        RECT 1367.740 1953.370 1367.880 2328.475 ;
        RECT 1367.280 1953.230 1367.880 1953.370 ;
        RECT 1367.280 1947.250 1367.420 1953.230 ;
        RECT 1367.680 1952.290 1367.940 1952.610 ;
        RECT 1367.740 1948.045 1367.880 1952.290 ;
        RECT 1367.670 1947.675 1367.950 1948.045 ;
        RECT 1367.280 1947.110 1367.880 1947.250 ;
        RECT 1367.220 1945.830 1367.480 1946.150 ;
        RECT 1366.760 1940.050 1367.020 1940.370 ;
        RECT 1366.820 1925.070 1366.960 1940.050 ;
        RECT 1366.760 1924.750 1367.020 1925.070 ;
        RECT 1367.280 1919.370 1367.420 1945.830 ;
        RECT 1367.740 1940.370 1367.880 1947.110 ;
        RECT 1367.680 1940.050 1367.940 1940.370 ;
        RECT 1368.200 1939.770 1368.340 2361.230 ;
        RECT 1367.740 1939.630 1368.340 1939.770 ;
        RECT 1367.740 1929.005 1367.880 1939.630 ;
        RECT 1368.140 1938.690 1368.400 1939.010 ;
        RECT 1368.200 1938.525 1368.340 1938.690 ;
        RECT 1368.130 1938.155 1368.410 1938.525 ;
        RECT 1368.140 1937.670 1368.400 1937.990 ;
        RECT 1367.670 1928.635 1367.950 1929.005 ;
        RECT 1366.820 1919.230 1367.420 1919.370 ;
        RECT 1366.820 1917.930 1366.960 1919.230 ;
        RECT 1366.760 1917.610 1367.020 1917.930 ;
        RECT 1368.200 1917.330 1368.340 1937.670 ;
        RECT 1366.820 1917.190 1368.340 1917.330 ;
        RECT 1366.290 1681.115 1366.570 1681.485 ;
        RECT 1366.820 1656.810 1366.960 1917.190 ;
        RECT 1367.220 1916.590 1367.480 1916.910 ;
        RECT 1366.760 1656.490 1367.020 1656.810 ;
        RECT 1366.760 1655.810 1367.020 1656.130 ;
        RECT 1366.820 1652.925 1366.960 1655.810 ;
        RECT 1366.750 1652.555 1367.030 1652.925 ;
        RECT 1367.280 1624.365 1367.420 1916.590 ;
        RECT 1367.670 1909.595 1367.950 1909.965 ;
        RECT 1367.740 1901.270 1367.880 1909.595 ;
        RECT 1368.130 1901.435 1368.410 1901.805 ;
        RECT 1367.680 1900.950 1367.940 1901.270 ;
        RECT 1368.200 1900.930 1368.340 1901.435 ;
        RECT 1368.140 1900.610 1368.400 1900.930 ;
        RECT 1367.680 1894.490 1367.940 1894.810 ;
        RECT 1367.740 1872.710 1367.880 1894.490 ;
        RECT 1368.140 1873.070 1368.400 1873.390 ;
        RECT 1367.680 1872.390 1367.940 1872.710 ;
        RECT 1368.200 1843.325 1368.340 1873.070 ;
        RECT 1368.130 1842.955 1368.410 1843.325 ;
        RECT 1368.660 1814.570 1368.800 2477.510 ;
        RECT 1369.120 1873.390 1369.260 2581.630 ;
        RECT 1369.060 1873.070 1369.320 1873.390 ;
        RECT 1369.060 1872.390 1369.320 1872.710 ;
        RECT 1369.120 1824.285 1369.260 1872.390 ;
        RECT 1369.050 1823.915 1369.330 1824.285 ;
        RECT 1368.600 1814.250 1368.860 1814.570 ;
        RECT 1367.680 1805.245 1367.940 1805.390 ;
        RECT 1367.670 1804.875 1367.950 1805.245 ;
        RECT 1369.060 1798.270 1369.320 1798.590 ;
        RECT 1369.120 1795.725 1369.260 1798.270 ;
        RECT 1369.050 1795.355 1369.330 1795.725 ;
        RECT 1369.060 1767.165 1369.320 1767.310 ;
        RECT 1369.050 1766.795 1369.330 1767.165 ;
        RECT 1367.680 1748.125 1367.940 1748.270 ;
        RECT 1367.670 1747.755 1367.950 1748.125 ;
        RECT 1367.680 1738.605 1367.940 1738.750 ;
        RECT 1367.670 1738.235 1367.950 1738.605 ;
        RECT 1367.680 1729.250 1367.940 1729.570 ;
        RECT 1367.740 1729.085 1367.880 1729.250 ;
        RECT 1367.670 1728.715 1367.950 1729.085 ;
        RECT 1368.140 1719.730 1368.400 1720.050 ;
        RECT 1368.200 1719.565 1368.340 1719.730 ;
        RECT 1368.130 1719.195 1368.410 1719.565 ;
        RECT 1367.680 1710.550 1367.940 1710.870 ;
        RECT 1367.740 1710.045 1367.880 1710.550 ;
        RECT 1367.670 1709.675 1367.950 1710.045 ;
        RECT 1367.680 1700.525 1367.940 1700.670 ;
        RECT 1367.670 1700.155 1367.950 1700.525 ;
        RECT 1369.580 1691.005 1369.720 2583.670 ;
        RECT 1370.040 1731.950 1370.180 2604.555 ;
        RECT 1371.350 2595.035 1371.630 2595.405 ;
        RECT 1371.420 2594.870 1371.560 2595.035 ;
        RECT 1371.360 2594.550 1371.620 2594.870 ;
        RECT 1507.520 2594.550 1507.780 2594.870 ;
        RECT 1370.430 2585.515 1370.710 2585.885 ;
        RECT 1370.500 1745.550 1370.640 2585.515 ;
        RECT 1376.880 2583.330 1377.140 2583.650 ;
        RECT 1371.820 2582.650 1372.080 2582.970 ;
        RECT 1370.890 2566.475 1371.170 2566.845 ;
        RECT 1370.960 1752.350 1371.100 2566.475 ;
        RECT 1371.350 2547.435 1371.630 2547.805 ;
        RECT 1371.420 1766.290 1371.560 2547.435 ;
        RECT 1371.880 1814.765 1372.020 2582.650 ;
        RECT 1372.280 2582.310 1372.540 2582.630 ;
        RECT 1372.340 1894.810 1372.480 2582.310 ;
        RECT 1372.740 2581.970 1373.000 2582.290 ;
        RECT 1372.280 1894.490 1372.540 1894.810 ;
        RECT 1372.280 1893.810 1372.540 1894.130 ;
        RECT 1372.340 1890.925 1372.480 1893.810 ;
        RECT 1372.270 1890.555 1372.550 1890.925 ;
        RECT 1372.270 1881.035 1372.550 1881.405 ;
        RECT 1372.340 1880.190 1372.480 1881.035 ;
        RECT 1372.280 1879.870 1372.540 1880.190 ;
        RECT 1372.280 1873.070 1372.540 1873.390 ;
        RECT 1372.340 1871.885 1372.480 1873.070 ;
        RECT 1372.270 1871.515 1372.550 1871.885 ;
        RECT 1372.270 1861.995 1372.550 1862.365 ;
        RECT 1372.340 1859.450 1372.480 1861.995 ;
        RECT 1372.280 1859.130 1372.540 1859.450 ;
        RECT 1372.270 1852.475 1372.550 1852.845 ;
        RECT 1372.280 1852.330 1372.540 1852.475 ;
        RECT 1372.800 1833.805 1372.940 2581.970 ;
        RECT 1376.420 2559.870 1376.680 2560.190 ;
        RECT 1375.960 2456.510 1376.220 2456.830 ;
        RECT 1375.500 2449.370 1375.760 2449.690 ;
        RECT 1375.040 2442.910 1375.300 2443.230 ;
        RECT 1374.580 2442.570 1374.840 2442.890 ;
        RECT 1374.120 2435.770 1374.380 2436.090 ;
        RECT 1373.660 2428.970 1373.920 2429.290 ;
        RECT 1373.200 2421.830 1373.460 2422.150 ;
        RECT 1373.260 2186.045 1373.400 2421.830 ;
        RECT 1373.190 2185.675 1373.470 2186.045 ;
        RECT 1373.720 2176.525 1373.860 2428.970 ;
        RECT 1373.650 2176.155 1373.930 2176.525 ;
        RECT 1374.180 2167.150 1374.320 2435.770 ;
        RECT 1374.120 2166.830 1374.380 2167.150 ;
        RECT 1374.640 2157.630 1374.780 2442.570 ;
        RECT 1374.580 2157.310 1374.840 2157.630 ;
        RECT 1375.100 2148.110 1375.240 2442.910 ;
        RECT 1375.040 2147.790 1375.300 2148.110 ;
        RECT 1375.560 2138.590 1375.700 2449.370 ;
        RECT 1375.500 2138.270 1375.760 2138.590 ;
        RECT 1376.020 2129.070 1376.160 2456.510 ;
        RECT 1375.960 2128.750 1376.220 2129.070 ;
        RECT 1375.960 1982.890 1376.220 1983.210 ;
        RECT 1375.500 1982.550 1375.760 1982.870 ;
        RECT 1375.040 1982.210 1375.300 1982.530 ;
        RECT 1374.580 1981.870 1374.840 1982.190 ;
        RECT 1374.120 1981.530 1374.380 1981.850 ;
        RECT 1373.190 1919.115 1373.470 1919.485 ;
        RECT 1373.260 1894.470 1373.400 1919.115 ;
        RECT 1373.200 1894.150 1373.460 1894.470 ;
        RECT 1372.730 1833.435 1373.010 1833.805 ;
        RECT 1371.810 1814.395 1372.090 1814.765 ;
        RECT 1371.820 1779.570 1372.080 1779.890 ;
        RECT 1371.880 1776.685 1372.020 1779.570 ;
        RECT 1371.810 1776.315 1372.090 1776.685 ;
        RECT 1374.180 1767.310 1374.320 1981.530 ;
        RECT 1374.120 1766.990 1374.380 1767.310 ;
        RECT 1371.360 1765.970 1371.620 1766.290 ;
        RECT 1374.640 1758.210 1374.780 1981.870 ;
        RECT 1372.800 1758.070 1374.780 1758.210 ;
        RECT 1372.800 1757.645 1372.940 1758.070 ;
        RECT 1372.730 1757.275 1373.010 1757.645 ;
        RECT 1370.900 1752.030 1371.160 1752.350 ;
        RECT 1375.100 1748.270 1375.240 1982.210 ;
        RECT 1375.040 1747.950 1375.300 1748.270 ;
        RECT 1370.440 1745.230 1370.700 1745.550 ;
        RECT 1375.560 1738.750 1375.700 1982.550 ;
        RECT 1375.500 1738.430 1375.760 1738.750 ;
        RECT 1369.980 1731.630 1370.240 1731.950 ;
        RECT 1376.020 1729.570 1376.160 1982.890 ;
        RECT 1376.480 1779.890 1376.620 2559.870 ;
        RECT 1376.940 1798.590 1377.080 2583.330 ;
        RECT 1377.340 2582.990 1377.600 2583.310 ;
        RECT 1377.400 1805.390 1377.540 2582.990 ;
        RECT 1493.720 2573.810 1493.980 2574.130 ;
        RECT 1486.820 2553.070 1487.080 2553.390 ;
        RECT 1397.120 2546.270 1397.380 2546.590 ;
        RECT 1377.800 2532.330 1378.060 2532.650 ;
        RECT 1377.860 2005.310 1378.000 2532.330 ;
        RECT 1378.260 2525.530 1378.520 2525.850 ;
        RECT 1378.320 2014.830 1378.460 2525.530 ;
        RECT 1383.320 2518.390 1383.580 2518.710 ;
        RECT 1378.720 2477.250 1378.980 2477.570 ;
        RECT 1378.780 2100.510 1378.920 2477.250 ;
        RECT 1379.180 2470.110 1379.440 2470.430 ;
        RECT 1379.240 2110.370 1379.380 2470.110 ;
        RECT 1379.640 2463.310 1379.900 2463.630 ;
        RECT 1379.700 2120.230 1379.840 2463.310 ;
        RECT 1382.860 2401.090 1383.120 2401.410 ;
        RECT 1382.400 2373.550 1382.660 2373.870 ;
        RECT 1381.940 2346.010 1382.200 2346.330 ;
        RECT 1381.480 2339.550 1381.740 2339.870 ;
        RECT 1381.020 2339.210 1381.280 2339.530 ;
        RECT 1380.560 2332.070 1380.820 2332.390 ;
        RECT 1380.100 2325.270 1380.360 2325.590 ;
        RECT 1380.160 2300.430 1380.300 2325.270 ;
        RECT 1380.100 2300.110 1380.360 2300.430 ;
        RECT 1380.620 2290.910 1380.760 2332.070 ;
        RECT 1380.560 2290.590 1380.820 2290.910 ;
        RECT 1381.080 2281.390 1381.220 2339.210 ;
        RECT 1381.020 2281.070 1381.280 2281.390 ;
        RECT 1381.540 2271.870 1381.680 2339.550 ;
        RECT 1381.480 2271.550 1381.740 2271.870 ;
        RECT 1382.000 2262.350 1382.140 2346.010 ;
        RECT 1381.940 2262.030 1382.200 2262.350 ;
        RECT 1382.460 2224.270 1382.600 2373.550 ;
        RECT 1382.400 2223.950 1382.660 2224.270 ;
        RECT 1382.920 2214.750 1383.060 2401.090 ;
        RECT 1382.860 2214.430 1383.120 2214.750 ;
        RECT 1379.640 2119.910 1379.900 2120.230 ;
        RECT 1379.180 2110.050 1379.440 2110.370 ;
        RECT 1378.720 2100.190 1378.980 2100.510 ;
        RECT 1383.380 2033.870 1383.520 2518.390 ;
        RECT 1383.780 2512.270 1384.040 2512.590 ;
        RECT 1383.840 2043.390 1383.980 2512.270 ;
        RECT 1384.240 2504.790 1384.500 2505.110 ;
        RECT 1384.300 2052.910 1384.440 2504.790 ;
        RECT 1384.700 2497.650 1384.960 2497.970 ;
        RECT 1384.760 2062.430 1384.900 2497.650 ;
        RECT 1385.160 2490.850 1385.420 2491.170 ;
        RECT 1385.220 2071.950 1385.360 2490.850 ;
        RECT 1392.980 2484.050 1393.240 2484.370 ;
        RECT 1390.220 2470.450 1390.480 2470.770 ;
        RECT 1386.080 2415.030 1386.340 2415.350 ;
        RECT 1385.620 2318.470 1385.880 2318.790 ;
        RECT 1385.160 2071.630 1385.420 2071.950 ;
        RECT 1384.700 2062.110 1384.960 2062.430 ;
        RECT 1384.240 2052.590 1384.500 2052.910 ;
        RECT 1383.780 2043.070 1384.040 2043.390 ;
        RECT 1383.320 2033.550 1383.580 2033.870 ;
        RECT 1378.260 2014.510 1378.520 2014.830 ;
        RECT 1377.800 2004.990 1378.060 2005.310 ;
        RECT 1378.720 1983.570 1378.980 1983.890 ;
        RECT 1377.800 1959.770 1378.060 1960.090 ;
        RECT 1377.340 1805.070 1377.600 1805.390 ;
        RECT 1376.880 1798.270 1377.140 1798.590 ;
        RECT 1376.420 1779.570 1376.680 1779.890 ;
        RECT 1375.960 1729.250 1376.220 1729.570 ;
        RECT 1369.510 1690.635 1369.790 1691.005 ;
        RECT 1369.060 1676.210 1369.320 1676.530 ;
        RECT 1369.120 1671.965 1369.260 1676.210 ;
        RECT 1369.050 1671.595 1369.330 1671.965 ;
        RECT 1371.360 1662.445 1371.620 1662.590 ;
        RECT 1371.350 1662.075 1371.630 1662.445 ;
        RECT 1367.680 1656.490 1367.940 1656.810 ;
        RECT 1367.740 1633.885 1367.880 1656.490 ;
        RECT 1369.980 1648.670 1370.240 1648.990 ;
        RECT 1370.040 1643.405 1370.180 1648.670 ;
        RECT 1369.970 1643.035 1370.250 1643.405 ;
        RECT 1367.670 1633.515 1367.950 1633.885 ;
        RECT 1367.210 1623.995 1367.490 1624.365 ;
        RECT 1367.680 1616.370 1367.940 1616.690 ;
        RECT 1367.740 1614.845 1367.880 1616.370 ;
        RECT 1367.670 1614.475 1367.950 1614.845 ;
        RECT 1377.860 1606.490 1378.000 1959.770 ;
        RECT 1378.260 1952.630 1378.520 1952.950 ;
        RECT 1378.320 1616.690 1378.460 1952.630 ;
        RECT 1378.780 1710.870 1378.920 1983.570 ;
        RECT 1379.640 1983.230 1379.900 1983.550 ;
        RECT 1379.180 1960.110 1379.440 1960.430 ;
        RECT 1378.720 1710.550 1378.980 1710.870 ;
        RECT 1379.240 1700.670 1379.380 1960.110 ;
        RECT 1379.700 1720.050 1379.840 1983.230 ;
        RECT 1385.680 1931.870 1385.820 2318.470 ;
        RECT 1386.140 2198.770 1386.280 2415.030 ;
        RECT 1386.540 2408.230 1386.800 2408.550 ;
        RECT 1386.600 2206.590 1386.740 2408.230 ;
        RECT 1386.540 2206.270 1386.800 2206.590 ;
        RECT 1386.080 2198.450 1386.340 2198.770 ;
        RECT 1385.620 1931.550 1385.880 1931.870 ;
        RECT 1390.280 1842.450 1390.420 2470.450 ;
        RECT 1390.680 2443.250 1390.940 2443.570 ;
        RECT 1390.740 1856.050 1390.880 2443.250 ;
        RECT 1391.140 2429.310 1391.400 2429.630 ;
        RECT 1391.200 1862.850 1391.340 2429.310 ;
        RECT 1391.600 2422.170 1391.860 2422.490 ;
        RECT 1391.660 1869.990 1391.800 2422.170 ;
        RECT 1392.060 2408.570 1392.320 2408.890 ;
        RECT 1392.120 1876.790 1392.260 2408.570 ;
        RECT 1392.520 2401.430 1392.780 2401.750 ;
        RECT 1392.580 1905.770 1392.720 2401.430 ;
        RECT 1393.040 2081.470 1393.180 2484.050 ;
        RECT 1393.440 2304.530 1393.700 2304.850 ;
        RECT 1392.980 2081.150 1393.240 2081.470 ;
        RECT 1393.500 1938.670 1393.640 2304.530 ;
        RECT 1393.440 1938.350 1393.700 1938.670 ;
        RECT 1392.580 1905.630 1393.180 1905.770 ;
        RECT 1393.040 1883.590 1393.180 1905.630 ;
        RECT 1392.980 1883.270 1393.240 1883.590 ;
        RECT 1392.060 1876.470 1392.320 1876.790 ;
        RECT 1391.600 1869.670 1391.860 1869.990 ;
        RECT 1391.140 1862.530 1391.400 1862.850 ;
        RECT 1390.680 1855.730 1390.940 1856.050 ;
        RECT 1390.220 1842.130 1390.480 1842.450 ;
        RECT 1379.640 1719.730 1379.900 1720.050 ;
        RECT 1379.180 1700.350 1379.440 1700.670 ;
        RECT 1397.180 1662.590 1397.320 2546.270 ;
        RECT 1473.020 2532.670 1473.280 2532.990 ;
        RECT 1459.220 2525.870 1459.480 2526.190 ;
        RECT 1452.320 2505.130 1452.580 2505.450 ;
        RECT 1438.520 2497.990 1438.780 2498.310 ;
        RECT 1431.620 2484.390 1431.880 2484.710 ;
        RECT 1424.720 2477.930 1424.980 2478.250 ;
        RECT 1397.580 2477.590 1397.840 2477.910 ;
        RECT 1397.640 2090.650 1397.780 2477.590 ;
        RECT 1417.820 2456.850 1418.080 2457.170 ;
        RECT 1404.020 2449.710 1404.280 2450.030 ;
        RECT 1397.580 2090.330 1397.840 2090.650 ;
        RECT 1404.080 1849.250 1404.220 2449.710 ;
        RECT 1404.020 1848.930 1404.280 1849.250 ;
        RECT 1417.880 1848.910 1418.020 2456.850 ;
        RECT 1417.820 1848.590 1418.080 1848.910 ;
        RECT 1424.780 1834.630 1424.920 2477.930 ;
        RECT 1424.720 1834.310 1424.980 1834.630 ;
        RECT 1431.680 1828.510 1431.820 2484.390 ;
        RECT 1431.620 1828.190 1431.880 1828.510 ;
        RECT 1438.580 1821.710 1438.720 2497.990 ;
        RECT 1438.520 1821.390 1438.780 1821.710 ;
        RECT 1452.380 1814.230 1452.520 2505.130 ;
        RECT 1452.320 1813.910 1452.580 1814.230 ;
        RECT 1459.280 1780.230 1459.420 2525.870 ;
        RECT 1459.220 1779.910 1459.480 1780.230 ;
        RECT 1473.080 1773.430 1473.220 2532.670 ;
        RECT 1473.020 1773.110 1473.280 1773.430 ;
        RECT 1486.880 1759.490 1487.020 2553.070 ;
        RECT 1486.820 1759.170 1487.080 1759.490 ;
        RECT 1493.780 1745.210 1493.920 2573.810 ;
        RECT 1493.720 1744.890 1493.980 1745.210 ;
        RECT 1507.580 1738.750 1507.720 2594.550 ;
        RECT 1688.750 2586.875 1689.030 2587.245 ;
        RECT 1688.820 2583.990 1688.960 2586.875 ;
        RECT 1688.760 2583.670 1689.020 2583.990 ;
        RECT 1691.980 2583.670 1692.240 2583.990 ;
        RECT 1704.400 2583.670 1704.660 2583.990 ;
        RECT 1692.040 2582.485 1692.180 2583.670 ;
        RECT 1704.460 2582.485 1704.600 2583.670 ;
        RECT 1994.190 2583.475 1994.470 2583.845 ;
        RECT 1994.200 2583.330 1994.460 2583.475 ;
        RECT 2001.100 2583.165 2001.360 2583.310 ;
        RECT 2001.090 2582.795 2001.370 2583.165 ;
        RECT 2007.990 2582.795 2008.270 2583.165 ;
        RECT 2008.000 2582.650 2008.260 2582.795 ;
        RECT 2016.740 2582.485 2017.000 2582.630 ;
        RECT 1691.970 2582.115 1692.250 2582.485 ;
        RECT 1704.390 2582.115 1704.670 2582.485 ;
        RECT 2016.730 2582.115 2017.010 2582.485 ;
        RECT 2021.790 2582.115 2022.070 2582.485 ;
        RECT 2030.070 2582.115 2030.350 2582.485 ;
        RECT 2021.800 2581.970 2022.060 2582.115 ;
        RECT 2030.080 2581.970 2030.340 2582.115 ;
        RECT 1600.890 2560.355 1601.170 2560.725 ;
        RECT 1600.960 2560.190 1601.100 2560.355 ;
        RECT 1600.900 2559.870 1601.160 2560.190 ;
        RECT 1601.820 2546.270 1602.080 2546.590 ;
        RECT 1583.410 2545.395 1583.690 2545.765 ;
        RECT 1514.420 2539.130 1514.680 2539.450 ;
        RECT 1507.520 1738.430 1507.780 1738.750 ;
        RECT 1514.480 1676.530 1514.620 2539.130 ;
        RECT 1576.520 2394.290 1576.780 2394.610 ;
        RECT 1562.720 2380.350 1562.980 2380.670 ;
        RECT 1548.920 2373.890 1549.180 2374.210 ;
        RECT 1542.020 2366.750 1542.280 2367.070 ;
        RECT 1528.220 2353.150 1528.480 2353.470 ;
        RECT 1521.320 2346.350 1521.580 2346.670 ;
        RECT 1514.880 2332.410 1515.140 2332.730 ;
        RECT 1514.940 1924.730 1515.080 2332.410 ;
        RECT 1514.880 1924.410 1515.140 1924.730 ;
        RECT 1521.380 1918.270 1521.520 2346.350 ;
        RECT 1521.320 1917.950 1521.580 1918.270 ;
        RECT 1528.280 1911.130 1528.420 2353.150 ;
        RECT 1528.220 1910.810 1528.480 1911.130 ;
        RECT 1542.080 1904.330 1542.220 2366.750 ;
        RECT 1542.020 1904.010 1542.280 1904.330 ;
        RECT 1548.980 1897.530 1549.120 2373.890 ;
        RECT 1548.920 1897.210 1549.180 1897.530 ;
        RECT 1562.780 1883.930 1562.920 2380.350 ;
        RECT 1576.580 1884.270 1576.720 2394.290 ;
        RECT 1576.520 1883.950 1576.780 1884.270 ;
        RECT 1562.720 1883.610 1562.980 1883.930 ;
        RECT 1514.420 1676.210 1514.680 1676.530 ;
        RECT 1397.120 1662.270 1397.380 1662.590 ;
        RECT 1583.480 1648.990 1583.620 2545.395 ;
        RECT 1597.210 2539.275 1597.490 2539.645 ;
        RECT 1594.000 1831.250 1594.260 1831.570 ;
        RECT 1594.060 1817.485 1594.200 1831.250 ;
        RECT 1593.990 1817.115 1594.270 1817.485 ;
        RECT 1597.280 1656.130 1597.420 2539.275 ;
        RECT 1600.900 2539.130 1601.160 2539.450 ;
        RECT 1599.060 2532.330 1599.320 2532.650 ;
        RECT 1599.120 2531.485 1599.260 2532.330 ;
        RECT 1600.960 2531.485 1601.100 2539.130 ;
        RECT 1601.880 2537.605 1602.020 2546.270 ;
        RECT 1601.810 2537.235 1602.090 2537.605 ;
        RECT 1599.050 2531.115 1599.330 2531.485 ;
        RECT 1600.890 2531.115 1601.170 2531.485 ;
        RECT 1600.900 2525.530 1601.160 2525.850 ;
        RECT 1599.980 2518.390 1600.240 2518.710 ;
        RECT 1599.060 2504.965 1599.320 2505.110 ;
        RECT 1599.050 2504.595 1599.330 2504.965 ;
        RECT 1600.040 2504.285 1600.180 2518.390 ;
        RECT 1600.960 2515.845 1601.100 2525.530 ;
        RECT 1603.650 2523.635 1603.930 2524.005 ;
        RECT 1602.730 2518.195 1603.010 2518.565 ;
        RECT 1600.890 2515.475 1601.170 2515.845 ;
        RECT 1601.360 2512.610 1601.620 2512.930 ;
        RECT 1599.970 2503.915 1600.250 2504.285 ;
        RECT 1601.420 2498.165 1601.560 2512.610 ;
        RECT 1601.810 2512.075 1602.090 2512.445 ;
        RECT 1600.900 2497.650 1601.160 2497.970 ;
        RECT 1601.350 2497.795 1601.630 2498.165 ;
        RECT 1599.060 2490.850 1599.320 2491.170 ;
        RECT 1599.120 2490.005 1599.260 2490.850 ;
        RECT 1599.050 2489.635 1599.330 2490.005 ;
        RECT 1600.960 2486.605 1601.100 2497.650 ;
        RECT 1601.350 2488.955 1601.630 2489.325 ;
        RECT 1600.890 2486.235 1601.170 2486.605 ;
        RECT 1600.900 2484.050 1601.160 2484.370 ;
        RECT 1599.060 2477.590 1599.320 2477.910 ;
        RECT 1599.120 2476.405 1599.260 2477.590 ;
        RECT 1599.980 2477.250 1600.240 2477.570 ;
        RECT 1599.050 2476.035 1599.330 2476.405 ;
        RECT 1599.060 2470.110 1599.320 2470.430 ;
        RECT 1599.120 2468.925 1599.260 2470.110 ;
        RECT 1599.050 2468.555 1599.330 2468.925 ;
        RECT 1600.040 2463.485 1600.180 2477.250 ;
        RECT 1600.960 2475.045 1601.100 2484.050 ;
        RECT 1600.890 2474.675 1601.170 2475.045 ;
        RECT 1599.970 2463.115 1600.250 2463.485 ;
        RECT 1600.900 2463.310 1601.160 2463.630 ;
        RECT 1599.060 2456.510 1599.320 2456.830 ;
        RECT 1599.120 2456.005 1599.260 2456.510 ;
        RECT 1599.050 2455.635 1599.330 2456.005 ;
        RECT 1600.960 2451.925 1601.100 2463.310 ;
        RECT 1600.890 2451.555 1601.170 2451.925 ;
        RECT 1600.900 2449.370 1601.160 2449.690 ;
        RECT 1600.440 2449.205 1600.700 2449.350 ;
        RECT 1600.430 2448.835 1600.710 2449.205 ;
        RECT 1599.060 2442.910 1599.320 2443.230 ;
        RECT 1598.600 2442.570 1598.860 2442.890 ;
        RECT 1598.660 2433.565 1598.800 2442.570 ;
        RECT 1599.120 2439.685 1599.260 2442.910 ;
        RECT 1600.960 2439.685 1601.100 2449.370 ;
        RECT 1601.420 2442.405 1601.560 2488.955 ;
        RECT 1601.880 2467.565 1602.020 2512.075 ;
        RECT 1602.270 2482.835 1602.550 2483.205 ;
        RECT 1601.810 2467.195 1602.090 2467.565 ;
        RECT 1601.350 2442.035 1601.630 2442.405 ;
        RECT 1599.050 2439.315 1599.330 2439.685 ;
        RECT 1600.890 2439.315 1601.170 2439.685 ;
        RECT 1601.350 2436.595 1601.630 2436.965 ;
        RECT 1600.900 2435.770 1601.160 2436.090 ;
        RECT 1598.590 2433.195 1598.870 2433.565 ;
        RECT 1599.060 2428.970 1599.320 2429.290 ;
        RECT 1599.120 2428.125 1599.260 2428.970 ;
        RECT 1599.050 2427.755 1599.330 2428.125 ;
        RECT 1600.960 2422.685 1601.100 2435.770 ;
        RECT 1600.890 2422.315 1601.170 2422.685 ;
        RECT 1600.900 2421.830 1601.160 2422.150 ;
        RECT 1599.060 2415.205 1599.320 2415.350 ;
        RECT 1599.050 2414.835 1599.330 2415.205 ;
        RECT 1600.960 2410.445 1601.100 2421.830 ;
        RECT 1600.890 2410.075 1601.170 2410.445 ;
        RECT 1600.900 2408.230 1601.160 2408.550 ;
        RECT 1599.060 2401.090 1599.320 2401.410 ;
        RECT 1599.120 2398.885 1599.260 2401.090 ;
        RECT 1600.960 2398.885 1601.100 2408.230 ;
        RECT 1601.420 2402.430 1601.560 2436.595 ;
        RECT 1601.880 2420.645 1602.020 2467.195 ;
        RECT 1602.340 2436.965 1602.480 2482.835 ;
        RECT 1602.800 2473.005 1602.940 2518.195 ;
        RECT 1603.190 2500.515 1603.470 2500.885 ;
        RECT 1603.260 2477.570 1603.400 2500.515 ;
        RECT 1603.720 2495.330 1603.860 2523.635 ;
        RECT 1604.110 2506.890 1604.390 2507.005 ;
        RECT 1604.110 2506.750 1604.780 2506.890 ;
        RECT 1604.110 2506.635 1604.390 2506.750 ;
        RECT 1603.720 2495.190 1604.320 2495.330 ;
        RECT 1603.650 2494.395 1603.930 2494.765 ;
        RECT 1603.200 2477.250 1603.460 2477.570 ;
        RECT 1602.730 2472.635 1603.010 2473.005 ;
        RECT 1602.270 2436.595 1602.550 2436.965 ;
        RECT 1602.280 2436.110 1602.540 2436.430 ;
        RECT 1602.340 2430.845 1602.480 2436.110 ;
        RECT 1602.800 2431.330 1602.940 2472.635 ;
        RECT 1603.720 2461.930 1603.860 2494.395 ;
        RECT 1604.180 2477.765 1604.320 2495.190 ;
        RECT 1604.110 2477.395 1604.390 2477.765 ;
        RECT 1604.180 2461.930 1604.320 2477.395 ;
        RECT 1603.660 2461.610 1603.920 2461.930 ;
        RECT 1604.120 2461.610 1604.380 2461.930 ;
        RECT 1603.190 2461.330 1603.470 2461.445 ;
        RECT 1604.640 2461.330 1604.780 2506.750 ;
        RECT 1603.190 2461.190 1604.780 2461.330 ;
        RECT 1603.190 2461.075 1603.470 2461.190 ;
        RECT 1603.660 2460.590 1603.920 2460.910 ;
        RECT 1604.120 2460.590 1604.380 2460.910 ;
        RECT 1603.200 2454.645 1603.460 2454.790 ;
        RECT 1603.190 2454.275 1603.470 2454.645 ;
        RECT 1603.200 2449.370 1603.460 2449.690 ;
        RECT 1603.260 2431.330 1603.400 2449.370 ;
        RECT 1603.720 2449.350 1603.860 2460.590 ;
        RECT 1604.180 2449.350 1604.320 2460.590 ;
        RECT 1603.660 2449.030 1603.920 2449.350 ;
        RECT 1604.120 2449.030 1604.380 2449.350 ;
        RECT 1604.120 2446.990 1604.380 2447.310 ;
        RECT 1603.650 2442.035 1603.930 2442.405 ;
        RECT 1602.740 2431.010 1603.000 2431.330 ;
        RECT 1603.200 2431.010 1603.460 2431.330 ;
        RECT 1602.270 2430.475 1602.550 2430.845 ;
        RECT 1601.810 2420.275 1602.090 2420.645 ;
        RECT 1601.360 2402.110 1601.620 2402.430 ;
        RECT 1601.360 2401.430 1601.620 2401.750 ;
        RECT 1599.050 2398.515 1599.330 2398.885 ;
        RECT 1600.890 2398.515 1601.170 2398.885 ;
        RECT 1600.900 2396.330 1601.160 2396.650 ;
        RECT 1600.960 2384.410 1601.100 2396.330 ;
        RECT 1600.900 2384.090 1601.160 2384.410 ;
        RECT 1600.890 2383.555 1601.170 2383.925 ;
        RECT 1601.420 2383.810 1601.560 2401.430 ;
        RECT 1601.880 2384.490 1602.020 2420.275 ;
        RECT 1602.340 2414.330 1602.480 2430.475 ;
        RECT 1602.740 2429.990 1603.000 2430.310 ;
        RECT 1603.200 2429.990 1603.460 2430.310 ;
        RECT 1602.800 2424.725 1602.940 2429.990 ;
        RECT 1602.730 2424.355 1603.010 2424.725 ;
        RECT 1602.280 2414.010 1602.540 2414.330 ;
        RECT 1602.280 2413.330 1602.540 2413.650 ;
        RECT 1602.340 2407.725 1602.480 2413.330 ;
        RECT 1602.800 2412.370 1602.940 2424.355 ;
        RECT 1603.260 2413.650 1603.400 2429.990 ;
        RECT 1603.720 2413.845 1603.860 2442.035 ;
        RECT 1603.200 2413.330 1603.460 2413.650 ;
        RECT 1603.650 2413.475 1603.930 2413.845 ;
        RECT 1604.180 2413.650 1604.320 2446.990 ;
        RECT 1604.120 2413.330 1604.380 2413.650 ;
        RECT 1603.190 2413.050 1603.470 2413.165 ;
        RECT 1604.640 2413.050 1604.780 2461.190 ;
        RECT 1603.190 2412.910 1604.780 2413.050 ;
        RECT 1603.190 2412.795 1603.470 2412.910 ;
        RECT 1602.800 2412.230 1603.860 2412.370 ;
        RECT 1602.740 2411.630 1603.000 2411.950 ;
        RECT 1602.270 2407.355 1602.550 2407.725 ;
        RECT 1602.340 2385.090 1602.480 2407.355 ;
        RECT 1602.800 2401.605 1602.940 2411.630 ;
        RECT 1603.190 2411.435 1603.470 2411.805 ;
        RECT 1602.730 2401.235 1603.010 2401.605 ;
        RECT 1602.280 2384.770 1602.540 2385.090 ;
        RECT 1601.880 2384.350 1602.480 2384.490 ;
        RECT 1601.810 2383.810 1602.090 2383.925 ;
        RECT 1601.420 2383.670 1602.090 2383.810 ;
        RECT 1601.810 2383.555 1602.090 2383.670 ;
        RECT 1600.960 2373.870 1601.100 2383.555 ;
        RECT 1601.360 2383.070 1601.620 2383.390 ;
        RECT 1600.900 2373.550 1601.160 2373.870 ;
        RECT 1600.890 2371.995 1601.170 2372.365 ;
        RECT 1600.960 2360.270 1601.100 2371.995 ;
        RECT 1601.420 2366.925 1601.560 2383.070 ;
        RECT 1601.880 2370.130 1602.020 2383.555 ;
        RECT 1602.340 2379.845 1602.480 2384.350 ;
        RECT 1602.270 2379.475 1602.550 2379.845 ;
        RECT 1602.280 2378.990 1602.540 2379.310 ;
        RECT 1601.820 2369.810 1602.080 2370.130 ;
        RECT 1602.340 2369.530 1602.480 2378.990 ;
        RECT 1601.880 2369.390 1602.480 2369.530 ;
        RECT 1601.350 2366.555 1601.630 2366.925 ;
        RECT 1601.350 2365.875 1601.630 2366.245 ;
        RECT 1600.900 2359.950 1601.160 2360.270 ;
        RECT 1600.890 2354.995 1601.170 2355.365 ;
        RECT 1600.960 2343.690 1601.100 2354.995 ;
        RECT 1601.420 2353.130 1601.560 2365.875 ;
        RECT 1601.880 2361.485 1602.020 2369.390 ;
        RECT 1602.800 2366.810 1602.940 2401.235 ;
        RECT 1603.260 2395.485 1603.400 2411.435 ;
        RECT 1603.720 2396.050 1603.860 2412.230 ;
        RECT 1604.120 2402.110 1604.380 2402.430 ;
        RECT 1604.180 2397.330 1604.320 2402.110 ;
        RECT 1604.120 2397.010 1604.380 2397.330 ;
        RECT 1604.640 2396.730 1604.780 2412.910 ;
        RECT 1604.180 2396.650 1604.780 2396.730 ;
        RECT 1604.120 2396.590 1604.780 2396.650 ;
        RECT 1604.120 2396.330 1604.380 2396.590 ;
        RECT 1603.720 2395.910 1604.320 2396.050 ;
        RECT 1603.190 2395.370 1603.470 2395.485 ;
        RECT 1603.190 2395.230 1603.860 2395.370 ;
        RECT 1603.190 2395.115 1603.470 2395.230 ;
        RECT 1603.200 2394.630 1603.460 2394.950 ;
        RECT 1603.260 2390.045 1603.400 2394.630 ;
        RECT 1603.190 2389.675 1603.470 2390.045 ;
        RECT 1603.200 2384.770 1603.460 2385.090 ;
        RECT 1603.260 2379.650 1603.400 2384.770 ;
        RECT 1603.720 2380.330 1603.860 2395.230 ;
        RECT 1603.660 2380.010 1603.920 2380.330 ;
        RECT 1603.200 2379.330 1603.460 2379.650 ;
        RECT 1603.650 2379.475 1603.930 2379.845 ;
        RECT 1603.190 2378.795 1603.470 2379.165 ;
        RECT 1602.340 2366.670 1602.940 2366.810 ;
        RECT 1601.810 2361.115 1602.090 2361.485 ;
        RECT 1601.810 2360.435 1602.090 2360.805 ;
        RECT 1601.360 2352.810 1601.620 2353.130 ;
        RECT 1601.360 2352.130 1601.620 2352.450 ;
        RECT 1601.420 2350.605 1601.560 2352.130 ;
        RECT 1601.350 2350.235 1601.630 2350.605 ;
        RECT 1601.350 2348.875 1601.630 2349.245 ;
        RECT 1600.500 2343.550 1601.100 2343.690 ;
        RECT 1600.500 2338.510 1600.640 2343.550 ;
        RECT 1600.890 2342.755 1601.170 2343.125 ;
        RECT 1600.440 2338.190 1600.700 2338.510 ;
        RECT 1600.960 2332.390 1601.100 2342.755 ;
        RECT 1601.420 2339.530 1601.560 2348.875 ;
        RECT 1601.880 2346.330 1602.020 2360.435 ;
        RECT 1602.340 2355.365 1602.480 2366.670 ;
        RECT 1602.730 2365.875 1603.010 2366.245 ;
        RECT 1602.270 2354.995 1602.550 2355.365 ;
        RECT 1602.270 2354.315 1602.550 2354.685 ;
        RECT 1601.820 2346.010 1602.080 2346.330 ;
        RECT 1601.810 2345.475 1602.090 2345.845 ;
        RECT 1601.360 2339.210 1601.620 2339.530 ;
        RECT 1601.880 2338.930 1602.020 2345.475 ;
        RECT 1602.340 2339.870 1602.480 2354.315 ;
        RECT 1602.280 2339.550 1602.540 2339.870 ;
        RECT 1602.800 2339.190 1602.940 2365.875 ;
        RECT 1603.260 2344.485 1603.400 2378.795 ;
        RECT 1603.720 2372.365 1603.860 2379.475 ;
        RECT 1604.180 2379.165 1604.320 2395.910 ;
        RECT 1604.110 2378.795 1604.390 2379.165 ;
        RECT 1604.120 2378.650 1604.380 2378.795 ;
        RECT 1604.180 2378.495 1604.320 2378.650 ;
        RECT 1604.110 2377.435 1604.390 2377.805 ;
        RECT 1603.650 2371.995 1603.930 2372.365 ;
        RECT 1603.190 2344.115 1603.470 2344.485 ;
        RECT 1601.360 2338.530 1601.620 2338.850 ;
        RECT 1601.880 2338.790 1602.480 2338.930 ;
        RECT 1602.740 2338.870 1603.000 2339.190 ;
        RECT 1600.900 2332.070 1601.160 2332.390 ;
        RECT 1600.890 2325.755 1601.170 2326.125 ;
        RECT 1600.960 2325.590 1601.100 2325.755 ;
        RECT 1600.900 2325.270 1601.160 2325.590 ;
        RECT 1600.890 2324.395 1601.170 2324.765 ;
        RECT 1600.960 2285.810 1601.100 2324.395 ;
        RECT 1600.900 2285.490 1601.160 2285.810 ;
        RECT 1601.420 2285.210 1601.560 2338.530 ;
        RECT 1601.820 2337.850 1602.080 2338.170 ;
        RECT 1600.960 2285.070 1601.560 2285.210 ;
        RECT 1600.960 2261.670 1601.100 2285.070 ;
        RECT 1601.880 2284.790 1602.020 2337.850 ;
        RECT 1602.340 2287.510 1602.480 2338.790 ;
        RECT 1602.740 2338.190 1603.000 2338.510 ;
        RECT 1603.260 2338.365 1603.400 2344.115 ;
        RECT 1603.720 2338.850 1603.860 2371.995 ;
        RECT 1603.660 2338.530 1603.920 2338.850 ;
        RECT 1602.280 2287.190 1602.540 2287.510 ;
        RECT 1601.820 2284.470 1602.080 2284.790 ;
        RECT 1601.820 2283.110 1602.080 2283.430 ;
        RECT 1602.280 2283.110 1602.540 2283.430 ;
        RECT 1600.900 2261.350 1601.160 2261.670 ;
        RECT 1601.880 2236.850 1602.020 2283.110 ;
        RECT 1602.340 2236.850 1602.480 2283.110 ;
        RECT 1602.800 2236.850 1602.940 2338.190 ;
        RECT 1603.190 2337.995 1603.470 2338.365 ;
        RECT 1603.200 2337.510 1603.460 2337.830 ;
        RECT 1603.260 2287.510 1603.400 2337.510 ;
        RECT 1603.660 2336.830 1603.920 2337.150 ;
        RECT 1603.200 2287.190 1603.460 2287.510 ;
        RECT 1603.720 2284.790 1603.860 2336.830 ;
        RECT 1604.180 2286.830 1604.320 2377.435 ;
        RECT 1604.120 2286.510 1604.380 2286.830 ;
        RECT 1603.660 2284.470 1603.920 2284.790 ;
        RECT 1603.200 2282.430 1603.460 2282.750 ;
        RECT 1603.260 2249.430 1603.400 2282.430 ;
        RECT 1603.200 2249.110 1603.460 2249.430 ;
        RECT 1601.820 2236.530 1602.080 2236.850 ;
        RECT 1602.280 2236.530 1602.540 2236.850 ;
        RECT 1602.740 2236.530 1603.000 2236.850 ;
        RECT 1602.280 2235.850 1602.540 2236.170 ;
        RECT 1602.740 2235.850 1603.000 2236.170 ;
        RECT 1601.820 2234.830 1602.080 2235.150 ;
        RECT 1601.360 2159.690 1601.620 2160.010 ;
        RECT 1601.420 2138.930 1601.560 2159.690 ;
        RECT 1601.360 2138.610 1601.620 2138.930 ;
        RECT 1600.900 1994.110 1601.160 1994.430 ;
        RECT 1600.960 1960.850 1601.100 1994.110 ;
        RECT 1600.500 1960.710 1601.100 1960.850 ;
        RECT 1600.500 1959.490 1600.640 1960.710 ;
        RECT 1600.900 1960.285 1601.160 1960.430 ;
        RECT 1600.890 1959.915 1601.170 1960.285 ;
        RECT 1601.360 1959.770 1601.620 1960.090 ;
        RECT 1600.500 1959.350 1601.100 1959.490 ;
        RECT 1600.440 1952.630 1600.700 1952.950 ;
        RECT 1600.500 1945.325 1600.640 1952.630 ;
        RECT 1600.960 1952.610 1601.100 1959.350 ;
        RECT 1600.900 1952.290 1601.160 1952.610 ;
        RECT 1601.420 1949.405 1601.560 1959.770 ;
        RECT 1601.880 1959.750 1602.020 2234.830 ;
        RECT 1602.340 2211.885 1602.480 2235.850 ;
        RECT 1602.800 2212.370 1602.940 2235.850 ;
        RECT 1603.200 2235.510 1603.460 2235.830 ;
        RECT 1602.740 2212.050 1603.000 2212.370 ;
        RECT 1602.270 2211.515 1602.550 2211.885 ;
        RECT 1602.740 2210.690 1603.000 2211.010 ;
        RECT 1602.280 2210.010 1602.540 2210.330 ;
        RECT 1602.340 1973.350 1602.480 2210.010 ;
        RECT 1602.800 1980.150 1602.940 2210.690 ;
        RECT 1603.260 1987.290 1603.400 2235.510 ;
        RECT 1604.180 2234.810 1604.780 2234.890 ;
        RECT 1604.120 2234.750 1604.780 2234.810 ;
        RECT 1604.120 2234.490 1604.380 2234.750 ;
        RECT 1603.660 2234.150 1603.920 2234.470 ;
        RECT 1603.720 2212.370 1603.860 2234.150 ;
        RECT 1604.120 2233.810 1604.380 2234.130 ;
        RECT 1603.660 2212.050 1603.920 2212.370 ;
        RECT 1603.650 2211.515 1603.930 2211.885 ;
        RECT 1603.720 2000.890 1603.860 2211.515 ;
        RECT 1604.180 2160.010 1604.320 2233.810 ;
        RECT 1604.120 2159.690 1604.380 2160.010 ;
        RECT 1604.120 2138.610 1604.380 2138.930 ;
        RECT 1603.660 2000.570 1603.920 2000.890 ;
        RECT 1604.180 1994.430 1604.320 2138.610 ;
        RECT 1604.120 1994.110 1604.380 1994.430 ;
        RECT 1603.200 1986.970 1603.460 1987.290 ;
        RECT 1602.740 1979.830 1603.000 1980.150 ;
        RECT 1602.280 1973.030 1602.540 1973.350 ;
        RECT 1601.820 1959.430 1602.080 1959.750 ;
        RECT 1601.350 1949.035 1601.630 1949.405 ;
        RECT 1601.360 1945.830 1601.620 1946.150 ;
        RECT 1600.430 1944.955 1600.710 1945.325 ;
        RECT 1600.900 1939.030 1601.160 1939.350 ;
        RECT 1600.960 1931.725 1601.100 1939.030 ;
        RECT 1601.420 1937.845 1601.560 1945.830 ;
        RECT 1604.640 1939.090 1604.780 2234.750 ;
      LAYER met2 ;
        RECT 1605.000 2205.000 2051.235 2581.480 ;
      LAYER met2 ;
        RECT 1693.360 1984.085 1693.620 1984.230 ;
        RECT 1693.350 1983.715 1693.630 1984.085 ;
        RECT 1987.290 1983.715 1987.570 1984.085 ;
        RECT 1987.300 1983.570 1987.560 1983.715 ;
        RECT 1994.200 1983.405 1994.460 1983.550 ;
        RECT 1994.190 1983.035 1994.470 1983.405 ;
        RECT 2001.090 1983.035 2001.370 1983.405 ;
        RECT 2001.100 1982.890 2001.360 1983.035 ;
        RECT 2008.000 1982.725 2008.260 1982.870 ;
        RECT 2007.990 1982.355 2008.270 1982.725 ;
        RECT 2016.730 1982.355 2017.010 1982.725 ;
        RECT 2021.790 1982.355 2022.070 1982.725 ;
        RECT 2030.070 1982.355 2030.350 1982.725 ;
        RECT 2016.740 1982.210 2017.000 1982.355 ;
        RECT 2021.860 1982.190 2022.000 1982.355 ;
        RECT 2030.140 1982.190 2030.280 1982.355 ;
        RECT 2021.800 1981.870 2022.060 1982.190 ;
        RECT 2030.080 1981.870 2030.340 1982.190 ;
        RECT 1604.180 1939.010 1604.780 1939.090 ;
        RECT 1604.120 1938.950 1604.780 1939.010 ;
        RECT 1604.120 1938.690 1604.380 1938.950 ;
        RECT 1601.820 1938.350 1602.080 1938.670 ;
        RECT 1601.350 1937.475 1601.630 1937.845 ;
        RECT 1601.880 1932.405 1602.020 1938.350 ;
        RECT 1601.810 1932.035 1602.090 1932.405 ;
        RECT 1600.890 1931.355 1601.170 1931.725 ;
        RECT 1601.360 1931.550 1601.620 1931.870 ;
        RECT 1600.900 1924.750 1601.160 1925.070 ;
        RECT 1600.960 1918.805 1601.100 1924.750 ;
        RECT 1600.890 1918.435 1601.170 1918.805 ;
        RECT 1600.900 1917.950 1601.160 1918.270 ;
        RECT 1600.960 1915.290 1601.100 1917.950 ;
        RECT 1601.420 1916.085 1601.560 1931.550 ;
        RECT 1601.820 1924.410 1602.080 1924.730 ;
        RECT 1601.350 1915.715 1601.630 1916.085 ;
        RECT 1600.960 1915.150 1601.560 1915.290 ;
        RECT 1600.900 1904.010 1601.160 1904.330 ;
        RECT 1600.440 1900.950 1600.700 1901.270 ;
        RECT 1600.500 1896.930 1600.640 1900.950 ;
        RECT 1600.960 1897.725 1601.100 1904.010 ;
        RECT 1601.420 1898.405 1601.560 1915.150 ;
        RECT 1601.880 1904.525 1602.020 1924.410 ;
        RECT 1603.190 1923.875 1603.470 1924.245 ;
        RECT 1602.740 1910.810 1603.000 1911.130 ;
        RECT 1601.810 1904.155 1602.090 1904.525 ;
        RECT 1602.280 1900.610 1602.540 1900.930 ;
        RECT 1601.350 1898.035 1601.630 1898.405 ;
        RECT 1600.890 1897.355 1601.170 1897.725 ;
        RECT 1601.360 1897.210 1601.620 1897.530 ;
        RECT 1600.500 1896.790 1601.100 1896.930 ;
        RECT 1600.960 1888.885 1601.100 1896.790 ;
        RECT 1600.890 1888.515 1601.170 1888.885 ;
        RECT 1599.980 1883.950 1600.240 1884.270 ;
        RECT 1599.060 1883.610 1599.320 1883.930 ;
        RECT 1599.120 1875.965 1599.260 1883.610 ;
        RECT 1599.050 1875.595 1599.330 1875.965 ;
        RECT 1600.040 1869.165 1600.180 1883.950 ;
        RECT 1600.890 1883.755 1601.170 1884.125 ;
        RECT 1600.960 1877.325 1601.100 1883.755 ;
        RECT 1601.420 1880.725 1601.560 1897.210 ;
        RECT 1602.340 1895.005 1602.480 1900.610 ;
        RECT 1602.270 1894.635 1602.550 1895.005 ;
        RECT 1601.820 1894.150 1602.080 1894.470 ;
        RECT 1601.880 1883.445 1602.020 1894.150 ;
        RECT 1601.810 1883.075 1602.090 1883.445 ;
        RECT 1601.820 1882.590 1602.080 1882.910 ;
        RECT 1601.350 1880.355 1601.630 1880.725 ;
        RECT 1600.890 1876.955 1601.170 1877.325 ;
        RECT 1600.960 1870.410 1601.100 1876.955 ;
        RECT 1601.360 1876.470 1601.620 1876.790 ;
        RECT 1600.500 1870.270 1601.100 1870.410 ;
        RECT 1599.970 1868.795 1600.250 1869.165 ;
        RECT 1600.500 1867.690 1600.640 1870.270 ;
        RECT 1600.900 1869.670 1601.160 1869.990 ;
        RECT 1600.040 1867.550 1600.640 1867.690 ;
        RECT 1599.520 1859.130 1599.780 1859.450 ;
        RECT 1599.060 1848.590 1599.320 1848.910 ;
        RECT 1599.120 1828.365 1599.260 1848.590 ;
        RECT 1599.580 1845.510 1599.720 1859.130 ;
        RECT 1600.040 1852.650 1600.180 1867.550 ;
        RECT 1600.430 1865.395 1600.710 1865.765 ;
        RECT 1600.500 1864.890 1600.640 1865.395 ;
        RECT 1600.440 1864.570 1600.700 1864.890 ;
        RECT 1600.960 1863.725 1601.100 1869.670 ;
        RECT 1600.890 1863.355 1601.170 1863.725 ;
        RECT 1601.420 1857.605 1601.560 1876.470 ;
        RECT 1601.880 1863.045 1602.020 1882.590 ;
        RECT 1601.810 1862.675 1602.090 1863.045 ;
        RECT 1601.820 1862.190 1602.080 1862.510 ;
        RECT 1601.350 1857.235 1601.630 1857.605 ;
        RECT 1601.360 1855.730 1601.620 1856.050 ;
        RECT 1599.980 1852.330 1600.240 1852.650 ;
        RECT 1600.040 1847.550 1600.180 1852.330 ;
        RECT 1600.900 1848.930 1601.160 1849.250 ;
        RECT 1599.980 1847.230 1600.240 1847.550 ;
        RECT 1599.520 1845.190 1599.780 1845.510 ;
        RECT 1600.960 1842.645 1601.100 1848.930 ;
        RECT 1600.890 1842.275 1601.170 1842.645 ;
        RECT 1601.420 1839.925 1601.560 1855.730 ;
        RECT 1601.880 1846.045 1602.020 1862.190 ;
        RECT 1602.340 1848.765 1602.480 1894.635 ;
        RECT 1602.800 1892.285 1602.940 1910.810 ;
        RECT 1603.260 1907.050 1603.400 1923.875 ;
        RECT 1603.650 1917.755 1603.930 1918.125 ;
        RECT 1603.200 1906.730 1603.460 1907.050 ;
        RECT 1603.190 1906.195 1603.470 1906.565 ;
        RECT 1603.260 1898.890 1603.400 1906.195 ;
        RECT 1603.200 1898.570 1603.460 1898.890 ;
        RECT 1603.720 1898.290 1603.860 1917.755 ;
        RECT 1604.110 1912.315 1604.390 1912.685 ;
        RECT 1604.180 1901.610 1604.320 1912.315 ;
        RECT 1604.120 1901.290 1604.380 1901.610 ;
        RECT 1604.110 1900.755 1604.390 1901.125 ;
        RECT 1603.260 1898.150 1603.860 1898.290 ;
        RECT 1602.730 1891.915 1603.010 1892.285 ;
        RECT 1602.740 1891.430 1603.000 1891.750 ;
        RECT 1602.800 1880.190 1602.940 1891.430 ;
        RECT 1602.740 1879.870 1603.000 1880.190 ;
        RECT 1602.800 1872.370 1602.940 1879.870 ;
        RECT 1602.740 1872.050 1603.000 1872.370 ;
        RECT 1602.730 1871.770 1603.010 1871.885 ;
        RECT 1603.260 1871.770 1603.400 1898.150 ;
        RECT 1603.660 1897.550 1603.920 1897.870 ;
        RECT 1603.720 1884.125 1603.860 1897.550 ;
        RECT 1604.180 1894.130 1604.320 1900.755 ;
        RECT 1604.120 1893.810 1604.380 1894.130 ;
        RECT 1604.180 1889.450 1604.320 1893.810 ;
        RECT 1604.180 1889.310 1604.780 1889.450 ;
        RECT 1604.110 1888.515 1604.390 1888.885 ;
        RECT 1603.650 1883.755 1603.930 1884.125 ;
        RECT 1602.730 1871.630 1603.400 1871.770 ;
        RECT 1602.730 1871.515 1603.010 1871.630 ;
        RECT 1602.800 1859.450 1602.940 1871.515 ;
        RECT 1603.200 1871.030 1603.460 1871.350 ;
        RECT 1603.260 1861.685 1603.400 1871.030 ;
        RECT 1603.190 1861.315 1603.470 1861.685 ;
        RECT 1602.740 1859.130 1603.000 1859.450 ;
        RECT 1603.260 1852.650 1603.400 1861.315 ;
        RECT 1604.180 1858.090 1604.320 1888.515 ;
        RECT 1604.120 1857.770 1604.380 1858.090 ;
        RECT 1604.110 1856.130 1604.390 1856.245 ;
        RECT 1604.640 1856.130 1604.780 1889.310 ;
        RECT 1604.110 1855.990 1604.780 1856.130 ;
        RECT 1604.110 1855.875 1604.390 1855.990 ;
        RECT 1604.180 1855.370 1604.320 1855.875 ;
        RECT 1604.120 1855.050 1604.380 1855.370 ;
        RECT 1603.200 1852.330 1603.460 1852.650 ;
        RECT 1604.120 1852.560 1604.380 1852.650 ;
        RECT 1604.120 1852.420 1604.780 1852.560 ;
        RECT 1604.120 1852.330 1604.380 1852.420 ;
        RECT 1603.200 1851.310 1603.460 1851.630 ;
        RECT 1602.270 1848.395 1602.550 1848.765 ;
        RECT 1603.260 1847.970 1603.400 1851.310 ;
        RECT 1602.340 1847.830 1603.400 1847.970 ;
        RECT 1601.810 1845.675 1602.090 1846.045 ;
        RECT 1601.820 1845.190 1602.080 1845.510 ;
        RECT 1601.350 1839.555 1601.630 1839.925 ;
        RECT 1601.360 1839.070 1601.620 1839.390 ;
        RECT 1600.900 1828.530 1601.160 1828.850 ;
        RECT 1599.050 1827.995 1599.330 1828.365 ;
        RECT 1600.960 1824.965 1601.100 1828.530 ;
        RECT 1600.890 1824.595 1601.170 1824.965 ;
        RECT 1601.420 1822.130 1601.560 1839.070 ;
        RECT 1601.880 1829.190 1602.020 1845.190 ;
        RECT 1602.340 1843.130 1602.480 1847.830 ;
        RECT 1603.200 1847.230 1603.460 1847.550 ;
        RECT 1602.280 1842.810 1602.540 1843.130 ;
        RECT 1602.280 1842.130 1602.540 1842.450 ;
        RECT 1601.820 1828.870 1602.080 1829.190 ;
        RECT 1601.820 1828.190 1602.080 1828.510 ;
        RECT 1600.960 1821.990 1601.560 1822.130 ;
        RECT 1600.040 1818.990 1600.180 1819.145 ;
        RECT 1599.980 1818.845 1600.240 1818.990 ;
        RECT 1599.970 1818.475 1600.250 1818.845 ;
        RECT 1599.060 1813.910 1599.320 1814.230 ;
        RECT 1599.120 1807.285 1599.260 1813.910 ;
        RECT 1599.050 1806.915 1599.330 1807.285 ;
        RECT 1600.040 1799.270 1600.180 1818.475 ;
        RECT 1600.440 1813.405 1600.700 1813.550 ;
        RECT 1600.430 1813.035 1600.710 1813.405 ;
        RECT 1600.960 1807.285 1601.100 1821.990 ;
        RECT 1601.360 1821.390 1601.620 1821.710 ;
        RECT 1600.890 1806.915 1601.170 1807.285 ;
        RECT 1600.960 1801.730 1601.100 1806.915 ;
        RECT 1601.420 1805.245 1601.560 1821.390 ;
        RECT 1601.880 1810.685 1602.020 1828.190 ;
        RECT 1602.340 1822.245 1602.480 1842.130 ;
        RECT 1603.260 1831.085 1603.400 1847.230 ;
        RECT 1603.650 1847.035 1603.930 1847.405 ;
        RECT 1603.190 1830.715 1603.470 1831.085 ;
        RECT 1603.260 1826.890 1603.400 1830.715 ;
        RECT 1602.800 1826.750 1603.400 1826.890 ;
        RECT 1602.270 1821.875 1602.550 1822.245 ;
        RECT 1602.280 1814.250 1602.540 1814.570 ;
        RECT 1601.810 1810.315 1602.090 1810.685 ;
        RECT 1602.340 1809.890 1602.480 1814.250 ;
        RECT 1601.880 1809.750 1602.480 1809.890 ;
        RECT 1601.350 1804.875 1601.630 1805.245 ;
        RECT 1601.360 1804.390 1601.620 1804.710 ;
        RECT 1601.420 1801.845 1601.560 1804.390 ;
        RECT 1600.500 1801.590 1601.100 1801.730 ;
        RECT 1600.500 1800.370 1600.640 1801.590 ;
        RECT 1601.350 1801.475 1601.630 1801.845 ;
        RECT 1601.420 1800.970 1601.560 1801.475 ;
        RECT 1601.360 1800.650 1601.620 1800.970 ;
        RECT 1600.500 1800.230 1601.100 1800.370 ;
        RECT 1599.980 1798.950 1600.240 1799.270 ;
        RECT 1600.960 1784.650 1601.100 1800.230 ;
        RECT 1601.360 1799.970 1601.620 1800.290 ;
        RECT 1601.420 1789.605 1601.560 1799.970 ;
        RECT 1601.880 1793.005 1602.020 1809.750 ;
        RECT 1602.280 1800.990 1602.540 1801.310 ;
        RECT 1602.340 1799.125 1602.480 1800.990 ;
        RECT 1602.270 1798.755 1602.550 1799.125 ;
        RECT 1601.810 1792.635 1602.090 1793.005 ;
        RECT 1601.350 1789.235 1601.630 1789.605 ;
        RECT 1600.900 1784.330 1601.160 1784.650 ;
        RECT 1600.890 1783.795 1601.170 1784.165 ;
        RECT 1600.960 1780.230 1601.100 1783.795 ;
        RECT 1600.900 1779.910 1601.160 1780.230 ;
        RECT 1600.890 1777.675 1601.170 1778.045 ;
        RECT 1600.960 1773.430 1601.100 1777.675 ;
        RECT 1600.900 1773.110 1601.160 1773.430 ;
        RECT 1600.890 1772.235 1601.170 1772.605 ;
        RECT 1600.960 1766.290 1601.100 1772.235 ;
        RECT 1601.420 1767.165 1601.560 1789.235 ;
        RECT 1602.800 1785.525 1602.940 1826.750 ;
        RECT 1603.190 1824.595 1603.470 1824.965 ;
        RECT 1602.730 1785.155 1603.010 1785.525 ;
        RECT 1601.820 1784.330 1602.080 1784.650 ;
        RECT 1601.350 1766.795 1601.630 1767.165 ;
        RECT 1600.900 1765.970 1601.160 1766.290 ;
        RECT 1601.350 1766.115 1601.630 1766.485 ;
        RECT 1600.890 1762.715 1601.170 1763.085 ;
        RECT 1600.960 1756.170 1601.100 1762.715 ;
        RECT 1601.420 1759.490 1601.560 1766.115 ;
        RECT 1601.880 1762.405 1602.020 1784.330 ;
        RECT 1603.260 1780.085 1603.400 1824.595 ;
        RECT 1603.720 1804.710 1603.860 1847.035 ;
        RECT 1604.110 1842.530 1604.390 1842.645 ;
        RECT 1604.640 1842.530 1604.780 1852.420 ;
        RECT 1604.110 1842.390 1604.780 1842.530 ;
        RECT 1604.110 1842.275 1604.390 1842.390 ;
        RECT 1604.110 1836.155 1604.390 1836.525 ;
        RECT 1603.660 1804.390 1603.920 1804.710 ;
        RECT 1604.180 1803.770 1604.320 1836.155 ;
        RECT 1603.720 1803.630 1604.320 1803.770 ;
        RECT 1603.720 1800.290 1603.860 1803.630 ;
        RECT 1604.640 1803.090 1604.780 1842.390 ;
        RECT 1604.180 1802.950 1604.780 1803.090 ;
        RECT 1604.180 1801.650 1604.320 1802.950 ;
        RECT 1604.120 1801.330 1604.380 1801.650 ;
        RECT 1603.660 1799.970 1603.920 1800.290 ;
        RECT 1603.720 1799.610 1604.780 1799.690 ;
        RECT 1603.660 1799.550 1604.780 1799.610 ;
        RECT 1603.660 1799.290 1603.920 1799.550 ;
        RECT 1603.650 1798.755 1603.930 1799.125 ;
        RECT 1604.120 1798.950 1604.380 1799.270 ;
        RECT 1603.190 1779.715 1603.470 1780.085 ;
        RECT 1603.200 1779.230 1603.460 1779.550 ;
        RECT 1601.810 1762.035 1602.090 1762.405 ;
        RECT 1601.360 1759.170 1601.620 1759.490 ;
        RECT 1603.260 1756.285 1603.400 1779.230 ;
        RECT 1600.960 1756.030 1601.560 1756.170 ;
        RECT 1601.420 1752.350 1601.560 1756.030 ;
        RECT 1603.190 1755.915 1603.470 1756.285 ;
        RECT 1601.810 1754.555 1602.090 1754.925 ;
        RECT 1601.360 1752.030 1601.620 1752.350 ;
        RECT 1600.890 1748.435 1601.170 1748.805 ;
        RECT 1600.960 1745.550 1601.100 1748.435 ;
        RECT 1600.900 1745.230 1601.160 1745.550 ;
        RECT 1601.880 1745.210 1602.020 1754.555 ;
        RECT 1603.720 1750.845 1603.860 1798.755 ;
        RECT 1604.180 1773.285 1604.320 1798.950 ;
        RECT 1604.110 1772.915 1604.390 1773.285 ;
        RECT 1604.110 1766.370 1604.390 1766.485 ;
        RECT 1604.640 1766.370 1604.780 1799.550 ;
        RECT 1604.110 1766.230 1604.780 1766.370 ;
        RECT 1604.110 1766.115 1604.390 1766.230 ;
        RECT 1603.650 1750.475 1603.930 1750.845 ;
        RECT 1601.820 1744.890 1602.080 1745.210 ;
        RECT 1600.890 1742.995 1601.170 1743.365 ;
        RECT 1600.960 1738.750 1601.100 1742.995 ;
        RECT 1600.900 1738.430 1601.160 1738.750 ;
        RECT 1600.900 1731.805 1601.160 1731.950 ;
        RECT 1600.890 1731.435 1601.170 1731.805 ;
        RECT 1597.220 1655.810 1597.480 1656.130 ;
        RECT 1583.420 1648.670 1583.680 1648.990 ;
        RECT 1378.260 1616.370 1378.520 1616.690 ;
        RECT 1367.220 1606.170 1367.480 1606.490 ;
        RECT 1377.800 1606.170 1378.060 1606.490 ;
        RECT 1367.280 1605.325 1367.420 1606.170 ;
        RECT 1367.210 1604.955 1367.490 1605.325 ;
      LAYER met2 ;
        RECT 1605.000 1605.000 2051.235 1981.480 ;
        RECT 350.030 1604.000 350.660 1604.280 ;
        RECT 351.500 1604.000 352.500 1604.280 ;
        RECT 353.340 1604.000 354.340 1604.280 ;
        RECT 355.180 1604.000 356.640 1604.280 ;
        RECT 357.480 1604.000 358.480 1604.280 ;
        RECT 359.320 1604.000 360.780 1604.280 ;
        RECT 361.620 1604.000 362.620 1604.280 ;
        RECT 363.460 1604.000 364.920 1604.280 ;
        RECT 365.760 1604.000 366.760 1604.280 ;
        RECT 367.600 1604.000 369.060 1604.280 ;
        RECT 369.900 1604.000 370.900 1604.280 ;
        RECT 371.740 1604.000 373.200 1604.280 ;
        RECT 374.040 1604.000 375.040 1604.280 ;
        RECT 375.880 1604.000 377.340 1604.280 ;
        RECT 378.180 1604.000 379.180 1604.280 ;
        RECT 380.020 1604.000 381.480 1604.280 ;
        RECT 382.320 1604.000 383.320 1604.280 ;
        RECT 384.160 1604.000 385.620 1604.280 ;
        RECT 386.460 1604.000 387.460 1604.280 ;
        RECT 388.300 1604.000 389.760 1604.280 ;
        RECT 390.600 1604.000 391.600 1604.280 ;
        RECT 392.440 1604.000 393.900 1604.280 ;
        RECT 394.740 1604.000 395.740 1604.280 ;
        RECT 396.580 1604.000 398.040 1604.280 ;
        RECT 398.880 1604.000 399.880 1604.280 ;
        RECT 400.720 1604.000 402.180 1604.280 ;
        RECT 403.020 1604.000 404.020 1604.280 ;
        RECT 404.860 1604.000 406.320 1604.280 ;
        RECT 407.160 1604.000 408.160 1604.280 ;
        RECT 409.000 1604.000 410.000 1604.280 ;
        RECT 410.840 1604.000 412.300 1604.280 ;
        RECT 413.140 1604.000 414.140 1604.280 ;
        RECT 414.980 1604.000 416.440 1604.280 ;
        RECT 417.280 1604.000 418.280 1604.280 ;
        RECT 419.120 1604.000 420.580 1604.280 ;
        RECT 421.420 1604.000 422.420 1604.280 ;
        RECT 423.260 1604.000 424.720 1604.280 ;
        RECT 425.560 1604.000 426.560 1604.280 ;
        RECT 427.400 1604.000 428.860 1604.280 ;
        RECT 429.700 1604.000 430.700 1604.280 ;
        RECT 431.540 1604.000 433.000 1604.280 ;
        RECT 433.840 1604.000 434.840 1604.280 ;
        RECT 435.680 1604.000 437.140 1604.280 ;
        RECT 437.980 1604.000 438.980 1604.280 ;
        RECT 439.820 1604.000 441.280 1604.280 ;
        RECT 442.120 1604.000 443.120 1604.280 ;
        RECT 443.960 1604.000 445.420 1604.280 ;
        RECT 446.260 1604.000 447.260 1604.280 ;
        RECT 448.100 1604.000 449.560 1604.280 ;
        RECT 450.400 1604.000 451.400 1604.280 ;
        RECT 452.240 1604.000 453.700 1604.280 ;
        RECT 454.540 1604.000 455.540 1604.280 ;
        RECT 456.380 1604.000 457.840 1604.280 ;
        RECT 458.680 1604.000 459.680 1604.280 ;
        RECT 460.520 1604.000 461.980 1604.280 ;
        RECT 462.820 1604.000 463.820 1604.280 ;
        RECT 464.660 1604.000 465.660 1604.280 ;
        RECT 466.500 1604.000 467.960 1604.280 ;
        RECT 468.800 1604.000 469.800 1604.280 ;
        RECT 470.640 1604.000 472.100 1604.280 ;
        RECT 472.940 1604.000 473.940 1604.280 ;
        RECT 474.780 1604.000 476.240 1604.280 ;
        RECT 477.080 1604.000 478.080 1604.280 ;
        RECT 478.920 1604.000 480.380 1604.280 ;
        RECT 481.220 1604.000 482.220 1604.280 ;
        RECT 483.060 1604.000 484.520 1604.280 ;
        RECT 485.360 1604.000 486.360 1604.280 ;
        RECT 487.200 1604.000 488.660 1604.280 ;
        RECT 489.500 1604.000 490.500 1604.280 ;
        RECT 491.340 1604.000 492.800 1604.280 ;
        RECT 493.640 1604.000 494.640 1604.280 ;
        RECT 495.480 1604.000 496.940 1604.280 ;
        RECT 497.780 1604.000 498.780 1604.280 ;
        RECT 499.620 1604.000 501.080 1604.280 ;
        RECT 501.920 1604.000 502.920 1604.280 ;
        RECT 503.760 1604.000 505.220 1604.280 ;
        RECT 506.060 1604.000 507.060 1604.280 ;
        RECT 507.900 1604.000 509.360 1604.280 ;
        RECT 510.200 1604.000 511.200 1604.280 ;
        RECT 512.040 1604.000 513.500 1604.280 ;
        RECT 514.340 1604.000 515.340 1604.280 ;
        RECT 516.180 1604.000 517.640 1604.280 ;
        RECT 518.480 1604.000 519.480 1604.280 ;
        RECT 520.320 1604.000 521.320 1604.280 ;
        RECT 522.160 1604.000 523.620 1604.280 ;
        RECT 524.460 1604.000 525.460 1604.280 ;
        RECT 526.300 1604.000 527.760 1604.280 ;
        RECT 528.600 1604.000 529.600 1604.280 ;
        RECT 530.440 1604.000 531.900 1604.280 ;
        RECT 532.740 1604.000 533.740 1604.280 ;
        RECT 534.580 1604.000 536.040 1604.280 ;
        RECT 536.880 1604.000 537.880 1604.280 ;
        RECT 538.720 1604.000 540.180 1604.280 ;
        RECT 541.020 1604.000 542.020 1604.280 ;
        RECT 542.860 1604.000 544.320 1604.280 ;
        RECT 545.160 1604.000 546.160 1604.280 ;
        RECT 547.000 1604.000 548.460 1604.280 ;
        RECT 549.300 1604.000 550.300 1604.280 ;
        RECT 551.140 1604.000 552.600 1604.280 ;
        RECT 553.440 1604.000 554.440 1604.280 ;
        RECT 555.280 1604.000 556.740 1604.280 ;
        RECT 557.580 1604.000 558.580 1604.280 ;
        RECT 559.420 1604.000 560.880 1604.280 ;
        RECT 561.720 1604.000 562.720 1604.280 ;
        RECT 563.560 1604.000 565.020 1604.280 ;
        RECT 565.860 1604.000 566.860 1604.280 ;
        RECT 567.700 1604.000 569.160 1604.280 ;
        RECT 570.000 1604.000 571.000 1604.280 ;
        RECT 571.840 1604.000 573.300 1604.280 ;
        RECT 574.140 1604.000 575.140 1604.280 ;
        RECT 575.980 1604.000 576.980 1604.280 ;
        RECT 577.820 1604.000 579.280 1604.280 ;
        RECT 580.120 1604.000 581.120 1604.280 ;
        RECT 581.960 1604.000 583.420 1604.280 ;
        RECT 584.260 1604.000 585.260 1604.280 ;
        RECT 586.100 1604.000 587.560 1604.280 ;
        RECT 588.400 1604.000 589.400 1604.280 ;
        RECT 590.240 1604.000 591.700 1604.280 ;
        RECT 592.540 1604.000 593.540 1604.280 ;
        RECT 594.380 1604.000 595.840 1604.280 ;
        RECT 596.680 1604.000 597.680 1604.280 ;
        RECT 598.520 1604.000 599.980 1604.280 ;
        RECT 600.820 1604.000 601.820 1604.280 ;
        RECT 602.660 1604.000 604.120 1604.280 ;
        RECT 604.960 1604.000 605.960 1604.280 ;
        RECT 606.800 1604.000 608.260 1604.280 ;
        RECT 609.100 1604.000 610.100 1604.280 ;
        RECT 610.940 1604.000 612.400 1604.280 ;
        RECT 613.240 1604.000 614.240 1604.280 ;
        RECT 615.080 1604.000 616.540 1604.280 ;
        RECT 617.380 1604.000 618.380 1604.280 ;
        RECT 619.220 1604.000 620.680 1604.280 ;
        RECT 621.520 1604.000 622.520 1604.280 ;
        RECT 623.360 1604.000 624.820 1604.280 ;
        RECT 625.660 1604.000 626.660 1604.280 ;
        RECT 627.500 1604.000 628.960 1604.280 ;
        RECT 629.800 1604.000 630.800 1604.280 ;
        RECT 631.640 1604.000 632.640 1604.280 ;
        RECT 633.480 1604.000 634.940 1604.280 ;
        RECT 635.780 1604.000 636.780 1604.280 ;
        RECT 637.620 1604.000 639.080 1604.280 ;
        RECT 639.920 1604.000 640.920 1604.280 ;
        RECT 641.760 1604.000 643.220 1604.280 ;
        RECT 644.060 1604.000 645.060 1604.280 ;
        RECT 645.900 1604.000 647.360 1604.280 ;
        RECT 648.200 1604.000 649.200 1604.280 ;
        RECT 650.040 1604.000 651.500 1604.280 ;
        RECT 652.340 1604.000 653.340 1604.280 ;
        RECT 654.180 1604.000 655.640 1604.280 ;
        RECT 656.480 1604.000 657.480 1604.280 ;
        RECT 658.320 1604.000 659.780 1604.280 ;
        RECT 660.620 1604.000 661.620 1604.280 ;
        RECT 662.460 1604.000 663.920 1604.280 ;
        RECT 664.760 1604.000 665.760 1604.280 ;
        RECT 666.600 1604.000 668.060 1604.280 ;
        RECT 668.900 1604.000 669.900 1604.280 ;
        RECT 670.740 1604.000 672.200 1604.280 ;
        RECT 673.040 1604.000 674.040 1604.280 ;
        RECT 674.880 1604.000 676.340 1604.280 ;
        RECT 677.180 1604.000 678.180 1604.280 ;
        RECT 679.020 1604.000 680.480 1604.280 ;
        RECT 681.320 1604.000 682.320 1604.280 ;
        RECT 683.160 1604.000 684.620 1604.280 ;
        RECT 685.460 1604.000 686.460 1604.280 ;
        RECT 687.300 1604.000 688.300 1604.280 ;
        RECT 689.140 1604.000 690.600 1604.280 ;
        RECT 691.440 1604.000 692.440 1604.280 ;
        RECT 693.280 1604.000 694.740 1604.280 ;
        RECT 695.580 1604.000 696.580 1604.280 ;
        RECT 697.420 1604.000 698.880 1604.280 ;
        RECT 699.720 1604.000 700.720 1604.280 ;
        RECT 701.560 1604.000 703.020 1604.280 ;
        RECT 703.860 1604.000 704.860 1604.280 ;
        RECT 705.700 1604.000 707.160 1604.280 ;
        RECT 708.000 1604.000 709.000 1604.280 ;
        RECT 709.840 1604.000 711.300 1604.280 ;
        RECT 712.140 1604.000 713.140 1604.280 ;
        RECT 713.980 1604.000 715.440 1604.280 ;
        RECT 716.280 1604.000 717.280 1604.280 ;
        RECT 718.120 1604.000 719.580 1604.280 ;
        RECT 720.420 1604.000 721.420 1604.280 ;
        RECT 722.260 1604.000 723.720 1604.280 ;
        RECT 724.560 1604.000 725.560 1604.280 ;
        RECT 726.400 1604.000 727.860 1604.280 ;
        RECT 728.700 1604.000 729.700 1604.280 ;
        RECT 730.540 1604.000 732.000 1604.280 ;
        RECT 732.840 1604.000 733.840 1604.280 ;
        RECT 734.680 1604.000 736.140 1604.280 ;
        RECT 736.980 1604.000 737.980 1604.280 ;
        RECT 738.820 1604.000 740.280 1604.280 ;
        RECT 741.120 1604.000 742.120 1604.280 ;
        RECT 742.960 1604.000 743.960 1604.280 ;
        RECT 744.800 1604.000 746.260 1604.280 ;
        RECT 747.100 1604.000 748.100 1604.280 ;
        RECT 748.940 1604.000 750.400 1604.280 ;
        RECT 751.240 1604.000 752.240 1604.280 ;
        RECT 753.080 1604.000 754.540 1604.280 ;
        RECT 755.380 1604.000 756.380 1604.280 ;
        RECT 757.220 1604.000 758.680 1604.280 ;
        RECT 759.520 1604.000 760.520 1604.280 ;
        RECT 761.360 1604.000 762.820 1604.280 ;
        RECT 763.660 1604.000 764.660 1604.280 ;
        RECT 765.500 1604.000 766.960 1604.280 ;
        RECT 767.800 1604.000 768.800 1604.280 ;
        RECT 769.640 1604.000 771.100 1604.280 ;
        RECT 771.940 1604.000 772.940 1604.280 ;
        RECT 773.780 1604.000 775.240 1604.280 ;
        RECT 776.080 1604.000 777.080 1604.280 ;
        RECT 777.920 1604.000 779.380 1604.280 ;
        RECT 780.220 1604.000 781.220 1604.280 ;
        RECT 782.060 1604.000 783.520 1604.280 ;
        RECT 784.360 1604.000 785.360 1604.280 ;
        RECT 786.200 1604.000 787.660 1604.280 ;
        RECT 788.500 1604.000 789.500 1604.280 ;
        RECT 790.340 1604.000 791.800 1604.280 ;
        RECT 792.640 1604.000 793.640 1604.280 ;
        RECT 794.480 1604.000 795.940 1604.280 ;
        RECT 796.780 1604.000 797.780 1604.280 ;
        RECT 798.620 1604.000 799.620 1604.280 ;
        RECT 800.460 1604.000 801.920 1604.280 ;
        RECT 802.760 1604.000 803.760 1604.280 ;
        RECT 804.600 1604.000 806.060 1604.280 ;
        RECT 806.900 1604.000 807.900 1604.280 ;
        RECT 808.740 1604.000 810.200 1604.280 ;
        RECT 811.040 1604.000 812.040 1604.280 ;
        RECT 812.880 1604.000 814.340 1604.280 ;
        RECT 815.180 1604.000 816.180 1604.280 ;
        RECT 817.020 1604.000 818.480 1604.280 ;
        RECT 819.320 1604.000 820.320 1604.280 ;
        RECT 821.160 1604.000 822.620 1604.280 ;
        RECT 823.460 1604.000 824.460 1604.280 ;
        RECT 825.300 1604.000 826.760 1604.280 ;
        RECT 827.600 1604.000 828.600 1604.280 ;
        RECT 829.440 1604.000 830.900 1604.280 ;
        RECT 831.740 1604.000 832.740 1604.280 ;
        RECT 833.580 1604.000 835.040 1604.280 ;
        RECT 835.880 1604.000 836.880 1604.280 ;
        RECT 837.720 1604.000 839.180 1604.280 ;
        RECT 840.020 1604.000 841.020 1604.280 ;
        RECT 841.860 1604.000 843.320 1604.280 ;
        RECT 844.160 1604.000 845.160 1604.280 ;
        RECT 846.000 1604.000 847.460 1604.280 ;
        RECT 848.300 1604.000 849.300 1604.280 ;
        RECT 850.140 1604.000 851.600 1604.280 ;
        RECT 852.440 1604.000 853.440 1604.280 ;
        RECT 854.280 1604.000 855.740 1604.280 ;
        RECT 856.580 1604.000 857.580 1604.280 ;
        RECT 858.420 1604.000 859.420 1604.280 ;
        RECT 860.260 1604.000 861.720 1604.280 ;
        RECT 862.560 1604.000 863.560 1604.280 ;
        RECT 864.400 1604.000 865.860 1604.280 ;
        RECT 866.700 1604.000 867.700 1604.280 ;
        RECT 868.540 1604.000 870.000 1604.280 ;
        RECT 870.840 1604.000 871.840 1604.280 ;
        RECT 872.680 1604.000 874.140 1604.280 ;
        RECT 874.980 1604.000 875.980 1604.280 ;
        RECT 876.820 1604.000 878.280 1604.280 ;
        RECT 879.120 1604.000 880.120 1604.280 ;
        RECT 880.960 1604.000 882.420 1604.280 ;
        RECT 883.260 1604.000 884.260 1604.280 ;
        RECT 885.100 1604.000 886.560 1604.280 ;
        RECT 887.400 1604.000 888.400 1604.280 ;
        RECT 889.240 1604.000 890.700 1604.280 ;
        RECT 891.540 1604.000 892.540 1604.280 ;
        RECT 893.380 1604.000 894.840 1604.280 ;
        RECT 895.680 1604.000 896.680 1604.280 ;
        RECT 897.520 1604.000 898.980 1604.280 ;
        RECT 899.820 1604.000 900.820 1604.280 ;
        RECT 901.660 1604.000 903.120 1604.280 ;
        RECT 903.960 1604.000 904.960 1604.280 ;
        RECT 905.800 1604.000 907.260 1604.280 ;
        RECT 908.100 1604.000 909.100 1604.280 ;
        RECT 909.940 1604.000 911.400 1604.280 ;
        RECT 912.240 1604.000 913.240 1604.280 ;
        RECT 914.080 1604.000 915.080 1604.280 ;
        RECT 915.920 1604.000 917.380 1604.280 ;
        RECT 918.220 1604.000 919.220 1604.280 ;
        RECT 920.060 1604.000 921.520 1604.280 ;
        RECT 922.360 1604.000 923.360 1604.280 ;
        RECT 924.200 1604.000 925.660 1604.280 ;
        RECT 926.500 1604.000 927.500 1604.280 ;
        RECT 928.340 1604.000 929.800 1604.280 ;
        RECT 930.640 1604.000 931.640 1604.280 ;
        RECT 932.480 1604.000 933.940 1604.280 ;
        RECT 934.780 1604.000 935.780 1604.280 ;
        RECT 936.620 1604.000 938.080 1604.280 ;
        RECT 938.920 1604.000 939.920 1604.280 ;
        RECT 940.760 1604.000 942.220 1604.280 ;
        RECT 943.060 1604.000 944.060 1604.280 ;
        RECT 944.900 1604.000 946.360 1604.280 ;
        RECT 947.200 1604.000 948.200 1604.280 ;
        RECT 949.040 1604.000 950.500 1604.280 ;
        RECT 951.340 1604.000 952.340 1604.280 ;
        RECT 953.180 1604.000 954.640 1604.280 ;
        RECT 955.480 1604.000 956.480 1604.280 ;
        RECT 957.320 1604.000 958.780 1604.280 ;
        RECT 959.620 1604.000 960.620 1604.280 ;
        RECT 961.460 1604.000 962.920 1604.280 ;
        RECT 963.760 1604.000 964.760 1604.280 ;
        RECT 965.600 1604.000 967.060 1604.280 ;
        RECT 967.900 1604.000 968.900 1604.280 ;
        RECT 969.740 1604.000 970.740 1604.280 ;
        RECT 971.580 1604.000 973.040 1604.280 ;
        RECT 973.880 1604.000 974.880 1604.280 ;
        RECT 975.720 1604.000 977.180 1604.280 ;
        RECT 978.020 1604.000 979.020 1604.280 ;
        RECT 979.860 1604.000 981.320 1604.280 ;
        RECT 982.160 1604.000 983.160 1604.280 ;
        RECT 984.000 1604.000 985.460 1604.280 ;
        RECT 986.300 1604.000 987.300 1604.280 ;
        RECT 988.140 1604.000 989.600 1604.280 ;
        RECT 990.440 1604.000 991.440 1604.280 ;
        RECT 992.280 1604.000 993.740 1604.280 ;
        RECT 994.580 1604.000 995.580 1604.280 ;
        RECT 996.420 1604.000 997.880 1604.280 ;
        RECT 998.720 1604.000 999.720 1604.280 ;
        RECT 1000.560 1604.000 1002.020 1604.280 ;
        RECT 1002.860 1604.000 1003.860 1604.280 ;
        RECT 1004.700 1604.000 1006.160 1604.280 ;
        RECT 1007.000 1604.000 1008.000 1604.280 ;
        RECT 1008.840 1604.000 1010.300 1604.280 ;
        RECT 1011.140 1604.000 1012.140 1604.280 ;
        RECT 1012.980 1604.000 1014.440 1604.280 ;
        RECT 1015.280 1604.000 1016.280 1604.280 ;
        RECT 1017.120 1604.000 1018.580 1604.280 ;
        RECT 1019.420 1604.000 1020.420 1604.280 ;
        RECT 1021.260 1604.000 1022.720 1604.280 ;
        RECT 1023.560 1604.000 1024.560 1604.280 ;
        RECT 1025.400 1604.000 1026.400 1604.280 ;
        RECT 1027.240 1604.000 1028.700 1604.280 ;
        RECT 1029.540 1604.000 1030.540 1604.280 ;
        RECT 1031.380 1604.000 1032.840 1604.280 ;
        RECT 1033.680 1604.000 1034.680 1604.280 ;
        RECT 1035.520 1604.000 1036.980 1604.280 ;
        RECT 1037.820 1604.000 1038.820 1604.280 ;
        RECT 1039.660 1604.000 1041.120 1604.280 ;
        RECT 1041.960 1604.000 1042.960 1604.280 ;
        RECT 1043.800 1604.000 1045.260 1604.280 ;
        RECT 1046.100 1604.000 1047.100 1604.280 ;
        RECT 1047.940 1604.000 1049.400 1604.280 ;
        RECT 1050.240 1604.000 1051.240 1604.280 ;
        RECT 1052.080 1604.000 1053.540 1604.280 ;
        RECT 1054.380 1604.000 1055.380 1604.280 ;
        RECT 1056.220 1604.000 1057.680 1604.280 ;
        RECT 1058.520 1604.000 1059.520 1604.280 ;
        RECT 1060.360 1604.000 1061.820 1604.280 ;
        RECT 1062.660 1604.000 1063.660 1604.280 ;
        RECT 1064.500 1604.000 1065.960 1604.280 ;
        RECT 1066.800 1604.000 1067.800 1604.280 ;
        RECT 1068.640 1604.000 1070.100 1604.280 ;
        RECT 1070.940 1604.000 1071.940 1604.280 ;
        RECT 1072.780 1604.000 1074.240 1604.280 ;
        RECT 1075.080 1604.000 1076.080 1604.280 ;
        RECT 1076.920 1604.000 1078.380 1604.280 ;
        RECT 1079.220 1604.000 1080.220 1604.280 ;
        RECT 1081.060 1604.000 1082.060 1604.280 ;
        RECT 1082.900 1604.000 1084.360 1604.280 ;
        RECT 1085.200 1604.000 1086.200 1604.280 ;
        RECT 1087.040 1604.000 1088.500 1604.280 ;
        RECT 1089.340 1604.000 1090.340 1604.280 ;
        RECT 1091.180 1604.000 1092.640 1604.280 ;
        RECT 1093.480 1604.000 1094.480 1604.280 ;
        RECT 1095.320 1604.000 1096.780 1604.280 ;
        RECT 1097.620 1604.000 1098.620 1604.280 ;
        RECT 1099.460 1604.000 1100.920 1604.280 ;
        RECT 1101.760 1604.000 1102.760 1604.280 ;
        RECT 1103.600 1604.000 1105.060 1604.280 ;
        RECT 1105.900 1604.000 1106.900 1604.280 ;
        RECT 1107.740 1604.000 1109.200 1604.280 ;
        RECT 1110.040 1604.000 1111.040 1604.280 ;
        RECT 1111.880 1604.000 1113.340 1604.280 ;
        RECT 1114.180 1604.000 1115.180 1604.280 ;
        RECT 1116.020 1604.000 1117.480 1604.280 ;
        RECT 1118.320 1604.000 1119.320 1604.280 ;
        RECT 1120.160 1604.000 1121.620 1604.280 ;
        RECT 1122.460 1604.000 1123.460 1604.280 ;
        RECT 1124.300 1604.000 1125.760 1604.280 ;
        RECT 1126.600 1604.000 1127.600 1604.280 ;
        RECT 1128.440 1604.000 1129.900 1604.280 ;
        RECT 1130.740 1604.000 1131.740 1604.280 ;
        RECT 1132.580 1604.000 1134.040 1604.280 ;
        RECT 1134.880 1604.000 1135.880 1604.280 ;
        RECT 1136.720 1604.000 1137.720 1604.280 ;
        RECT 1138.560 1604.000 1140.020 1604.280 ;
        RECT 1140.860 1604.000 1141.860 1604.280 ;
        RECT 1142.700 1604.000 1144.160 1604.280 ;
        RECT 1145.000 1604.000 1146.000 1604.280 ;
        RECT 1146.840 1604.000 1148.300 1604.280 ;
        RECT 1149.140 1604.000 1150.140 1604.280 ;
        RECT 1150.980 1604.000 1152.440 1604.280 ;
        RECT 1153.280 1604.000 1154.280 1604.280 ;
        RECT 1155.120 1604.000 1156.580 1604.280 ;
        RECT 1157.420 1604.000 1158.420 1604.280 ;
        RECT 1159.260 1604.000 1160.720 1604.280 ;
        RECT 1161.560 1604.000 1162.560 1604.280 ;
        RECT 1163.400 1604.000 1164.860 1604.280 ;
        RECT 1165.700 1604.000 1166.700 1604.280 ;
        RECT 1167.540 1604.000 1169.000 1604.280 ;
        RECT 1169.840 1604.000 1170.840 1604.280 ;
        RECT 1171.680 1604.000 1173.140 1604.280 ;
        RECT 1173.980 1604.000 1174.980 1604.280 ;
        RECT 1175.820 1604.000 1177.280 1604.280 ;
        RECT 1178.120 1604.000 1179.120 1604.280 ;
        RECT 1179.960 1604.000 1181.420 1604.280 ;
        RECT 1182.260 1604.000 1183.260 1604.280 ;
        RECT 1184.100 1604.000 1185.560 1604.280 ;
        RECT 1186.400 1604.000 1187.400 1604.280 ;
        RECT 1188.240 1604.000 1189.700 1604.280 ;
        RECT 1190.540 1604.000 1191.540 1604.280 ;
        RECT 1192.380 1604.000 1193.380 1604.280 ;
        RECT 1194.220 1604.000 1195.680 1604.280 ;
        RECT 1196.520 1604.000 1197.520 1604.280 ;
        RECT 1198.360 1604.000 1199.820 1604.280 ;
        RECT 1200.660 1604.000 1201.660 1604.280 ;
        RECT 1202.500 1604.000 1203.960 1604.280 ;
        RECT 1204.800 1604.000 1205.800 1604.280 ;
        RECT 1206.640 1604.000 1208.100 1604.280 ;
        RECT 1208.940 1604.000 1209.940 1604.280 ;
        RECT 1210.780 1604.000 1212.240 1604.280 ;
        RECT 1213.080 1604.000 1214.080 1604.280 ;
        RECT 1214.920 1604.000 1216.380 1604.280 ;
        RECT 1217.220 1604.000 1218.220 1604.280 ;
        RECT 1219.060 1604.000 1220.520 1604.280 ;
        RECT 1221.360 1604.000 1222.360 1604.280 ;
        RECT 1223.200 1604.000 1224.660 1604.280 ;
        RECT 1225.500 1604.000 1226.500 1604.280 ;
        RECT 1227.340 1604.000 1228.800 1604.280 ;
        RECT 1229.640 1604.000 1230.640 1604.280 ;
        RECT 1231.480 1604.000 1232.940 1604.280 ;
        RECT 1233.780 1604.000 1234.780 1604.280 ;
        RECT 1235.620 1604.000 1237.080 1604.280 ;
        RECT 1237.920 1604.000 1238.920 1604.280 ;
        RECT 1239.760 1604.000 1241.220 1604.280 ;
        RECT 1242.060 1604.000 1243.060 1604.280 ;
        RECT 1243.900 1604.000 1245.360 1604.280 ;
        RECT 1246.200 1604.000 1247.200 1604.280 ;
        RECT 1248.040 1604.000 1249.040 1604.280 ;
        RECT 1249.880 1604.000 1251.340 1604.280 ;
        RECT 1252.180 1604.000 1253.180 1604.280 ;
        RECT 1254.020 1604.000 1255.480 1604.280 ;
        RECT 1256.320 1604.000 1257.320 1604.280 ;
        RECT 1258.160 1604.000 1259.620 1604.280 ;
        RECT 1260.460 1604.000 1261.460 1604.280 ;
        RECT 1262.300 1604.000 1263.760 1604.280 ;
        RECT 1264.600 1604.000 1265.600 1604.280 ;
        RECT 1266.440 1604.000 1267.900 1604.280 ;
        RECT 1268.740 1604.000 1269.740 1604.280 ;
        RECT 1270.580 1604.000 1272.040 1604.280 ;
        RECT 1272.880 1604.000 1273.880 1604.280 ;
        RECT 1274.720 1604.000 1276.180 1604.280 ;
        RECT 1277.020 1604.000 1278.020 1604.280 ;
        RECT 1278.860 1604.000 1280.320 1604.280 ;
        RECT 1281.160 1604.000 1282.160 1604.280 ;
        RECT 1283.000 1604.000 1284.460 1604.280 ;
        RECT 1285.300 1604.000 1286.300 1604.280 ;
        RECT 1287.140 1604.000 1288.600 1604.280 ;
        RECT 1289.440 1604.000 1290.440 1604.280 ;
        RECT 1291.280 1604.000 1292.740 1604.280 ;
        RECT 1293.580 1604.000 1294.580 1604.280 ;
        RECT 1295.420 1604.000 1296.880 1604.280 ;
        RECT 1297.720 1604.000 1298.720 1604.280 ;
        RECT 1299.560 1604.000 1301.020 1604.280 ;
        RECT 1301.860 1604.000 1302.860 1604.280 ;
        RECT 1303.700 1604.000 1304.700 1604.280 ;
        RECT 1305.540 1604.000 1307.000 1604.280 ;
        RECT 1307.840 1604.000 1308.840 1604.280 ;
        RECT 1309.680 1604.000 1311.140 1604.280 ;
        RECT 1311.980 1604.000 1312.980 1604.280 ;
        RECT 1313.820 1604.000 1315.280 1604.280 ;
        RECT 1316.120 1604.000 1317.120 1604.280 ;
        RECT 1317.960 1604.000 1319.420 1604.280 ;
        RECT 1320.260 1604.000 1321.260 1604.280 ;
        RECT 1322.100 1604.000 1323.560 1604.280 ;
        RECT 1324.400 1604.000 1325.400 1604.280 ;
        RECT 1326.240 1604.000 1327.700 1604.280 ;
        RECT 1328.540 1604.000 1329.540 1604.280 ;
        RECT 1330.380 1604.000 1331.840 1604.280 ;
        RECT 1332.680 1604.000 1333.680 1604.280 ;
        RECT 1334.520 1604.000 1335.980 1604.280 ;
        RECT 1336.820 1604.000 1337.820 1604.280 ;
        RECT 1338.660 1604.000 1340.120 1604.280 ;
        RECT 1340.960 1604.000 1341.960 1604.280 ;
        RECT 1342.800 1604.000 1344.260 1604.280 ;
        RECT 1345.100 1604.000 1346.100 1604.280 ;
        RECT 1346.940 1604.000 1348.400 1604.280 ;
        RECT 1349.240 1604.000 1350.240 1604.280 ;
        RECT 1351.080 1604.000 1352.540 1604.280 ;
        RECT 1353.380 1604.000 1354.380 1604.280 ;
        RECT 1355.220 1604.000 1356.680 1604.280 ;
      LAYER via2 ;
        RECT 392.930 3279.840 393.210 3280.120 ;
        RECT 392.470 3274.400 392.750 3274.680 ;
        RECT 392.010 3265.560 392.290 3265.840 ;
        RECT 391.550 3260.120 391.830 3260.400 ;
        RECT 391.090 3237.680 391.370 3237.960 ;
        RECT 379.130 2840.560 379.410 2840.840 ;
        RECT 386.030 2839.880 386.310 2840.160 ;
        RECT 354.750 2618.200 355.030 2618.480 ;
        RECT 393.390 3251.960 393.670 3252.240 ;
        RECT 393.850 3245.840 394.130 3246.120 ;
        RECT 394.310 2948.000 394.590 2948.280 ;
        RECT 938.490 3279.840 938.770 3280.120 ;
        RECT 516.670 2851.440 516.950 2851.720 ;
        RECT 433.870 2842.600 434.150 2842.880 ;
        RECT 509.770 2842.600 510.050 2842.880 ;
        RECT 475.730 2841.920 476.010 2842.200 ;
        RECT 455.490 2838.520 455.770 2838.800 ;
        RECT 482.630 2841.240 482.910 2841.520 ;
        RECT 489.530 2838.520 489.810 2838.800 ;
        RECT 503.330 2838.520 503.610 2838.800 ;
        RECT 441.690 2837.160 441.970 2837.440 ;
        RECT 434.790 2836.480 435.070 2836.760 ;
        RECT 449.970 2836.480 450.250 2836.760 ;
        RECT 468.370 2835.800 468.650 2836.080 ;
        RECT 475.270 2835.800 475.550 2836.080 ;
        RECT 482.170 2835.800 482.450 2836.080 ;
        RECT 495.970 2835.800 496.250 2836.080 ;
        RECT 510.230 2841.240 510.510 2841.520 ;
        RECT 572.330 2848.040 572.610 2848.320 ;
        RECT 600.390 2848.040 600.670 2848.320 ;
        RECT 524.030 2842.600 524.310 2842.880 ;
        RECT 526.330 2842.600 526.610 2842.880 ;
        RECT 530.930 2842.600 531.210 2842.880 ;
        RECT 537.830 2842.600 538.110 2842.880 ;
        RECT 544.730 2842.600 545.010 2842.880 ;
        RECT 558.530 2842.600 558.810 2842.880 ;
        RECT 549.330 2841.920 549.610 2842.200 ;
        RECT 551.630 2838.520 551.910 2838.800 ;
        RECT 597.170 2845.320 597.450 2845.600 ;
        RECT 573.710 2843.280 573.990 2843.560 ;
        RECT 590.270 2843.280 590.550 2843.560 ;
        RECT 604.990 2845.320 605.270 2845.600 ;
        RECT 613.730 2843.960 614.010 2844.240 ;
        RECT 592.570 2832.400 592.850 2832.680 ;
        RECT 642.250 2842.600 642.530 2842.880 ;
        RECT 620.630 2841.240 620.910 2841.520 ;
        RECT 621.550 2841.240 621.830 2841.520 ;
        RECT 627.530 2841.240 627.810 2841.520 ;
        RECT 625.230 2836.480 625.510 2836.760 ;
        RECT 626.610 2835.800 626.890 2836.080 ;
        RECT 626.610 2619.560 626.890 2619.840 ;
        RECT 634.430 2835.800 634.710 2836.080 ;
        RECT 640.870 2835.800 641.150 2836.080 ;
        RECT 634.430 2618.880 634.710 2619.160 ;
        RECT 727.810 2841.240 728.090 2841.520 ;
        RECT 727.810 2620.240 728.090 2620.520 ;
        RECT 941.710 3274.400 941.990 3274.680 ;
        RECT 762.310 2620.920 762.590 2621.200 ;
        RECT 942.170 3265.560 942.450 3265.840 ;
        RECT 942.630 3260.120 942.910 3260.400 ;
        RECT 943.090 3251.960 943.370 3252.240 ;
        RECT 943.550 3245.840 943.830 3246.120 ;
        RECT 944.010 3237.680 944.290 3237.960 ;
        RECT 944.470 2948.000 944.750 2948.280 ;
        RECT 1103.630 2850.760 1103.910 2851.040 ;
        RECT 1089.370 2848.040 1089.650 2848.320 ;
        RECT 979.890 2842.600 980.170 2842.880 ;
        RECT 987.250 2842.600 987.530 2842.880 ;
        RECT 1020.830 2842.600 1021.110 2842.880 ;
        RECT 1024.050 2842.600 1024.330 2842.880 ;
        RECT 1027.730 2842.600 1028.010 2842.880 ;
        RECT 1065.450 2842.600 1065.730 2842.880 ;
        RECT 1070.510 2842.600 1070.790 2842.880 ;
        RECT 1018.530 2841.920 1018.810 2842.200 ;
        RECT 1021.750 2620.920 1022.030 2621.200 ;
        RECT 1012.090 2619.560 1012.370 2619.840 ;
        RECT 987.250 2618.200 987.530 2618.480 ;
        RECT 1045.210 2836.480 1045.490 2836.760 ;
        RECT 1041.530 2835.800 1041.810 2836.080 ;
        RECT 1030.950 2618.880 1031.230 2619.160 ;
        RECT 1048.430 2835.800 1048.710 2836.080 ;
        RECT 1054.870 2835.800 1055.150 2836.080 ;
        RECT 1062.230 2835.800 1062.510 2836.080 ;
        RECT 1069.130 2835.800 1069.410 2836.080 ;
        RECT 1076.030 2835.800 1076.310 2836.080 ;
        RECT 1082.930 2835.800 1083.210 2836.080 ;
        RECT 1089.370 2835.800 1089.650 2836.080 ;
        RECT 1096.730 2835.800 1097.010 2836.080 ;
        RECT 1050.270 2620.240 1050.550 2620.520 ;
        RECT 1111.910 2842.600 1112.190 2842.880 ;
        RECT 1118.350 2842.600 1118.630 2842.880 ;
        RECT 1131.230 2842.600 1131.510 2842.880 ;
        RECT 1135.830 2842.600 1136.110 2842.880 ;
        RECT 1138.130 2842.600 1138.410 2842.880 ;
        RECT 1145.030 2842.600 1145.310 2842.880 ;
        RECT 1151.930 2842.600 1152.210 2842.880 ;
        RECT 1158.830 2842.600 1159.110 2842.880 ;
        RECT 1165.270 2842.600 1165.550 2842.880 ;
        RECT 1172.630 2842.600 1172.910 2842.880 ;
        RECT 1179.530 2842.600 1179.810 2842.880 ;
        RECT 1186.430 2842.600 1186.710 2842.880 ;
        RECT 1193.330 2842.600 1193.610 2842.880 ;
        RECT 1130.770 2841.920 1131.050 2842.200 ;
        RECT 1110.530 2835.800 1110.810 2836.080 ;
        RECT 1117.430 2835.800 1117.710 2836.080 ;
        RECT 1124.330 2835.800 1124.610 2836.080 ;
        RECT 1159.750 2840.560 1160.030 2840.840 ;
        RECT 1159.290 2839.880 1159.570 2840.160 ;
        RECT 1165.730 2841.920 1166.010 2842.200 ;
        RECT 1179.990 2840.560 1180.270 2840.840 ;
        RECT 1369.970 2604.600 1370.250 2604.880 ;
        RECT 1368.130 2576.040 1368.410 2576.320 ;
        RECT 1367.670 2557.000 1367.950 2557.280 ;
        RECT 1368.590 2537.960 1368.870 2538.240 ;
        RECT 1367.670 2528.440 1367.950 2528.720 ;
        RECT 1367.670 2518.920 1367.950 2519.200 ;
        RECT 1368.130 2509.400 1368.410 2509.680 ;
        RECT 1368.590 2499.880 1368.870 2500.160 ;
        RECT 1368.590 2490.360 1368.870 2490.640 ;
        RECT 1368.590 2480.840 1368.870 2481.120 ;
        RECT 1368.130 2471.320 1368.410 2471.600 ;
        RECT 1368.130 2461.800 1368.410 2462.080 ;
        RECT 1367.210 2452.280 1367.490 2452.560 ;
        RECT 1368.130 2442.760 1368.410 2443.040 ;
        RECT 1367.670 2433.240 1367.950 2433.520 ;
        RECT 1368.130 2423.720 1368.410 2424.000 ;
        RECT 1368.130 2414.200 1368.410 2414.480 ;
        RECT 1368.130 2404.680 1368.410 2404.960 ;
        RECT 1368.130 2395.160 1368.410 2395.440 ;
        RECT 1368.130 2385.640 1368.410 2385.920 ;
        RECT 1368.130 2376.120 1368.410 2376.400 ;
        RECT 1368.130 2366.600 1368.410 2366.880 ;
        RECT 1366.290 2319.000 1366.570 2319.280 ;
        RECT 1366.290 2309.480 1366.570 2309.760 ;
        RECT 1366.290 2299.960 1366.570 2300.240 ;
        RECT 1366.290 2290.440 1366.570 2290.720 ;
        RECT 1366.290 2280.920 1366.570 2281.200 ;
        RECT 1366.290 2271.400 1366.570 2271.680 ;
        RECT 1366.290 2261.880 1366.570 2262.160 ;
        RECT 1366.750 2252.360 1367.030 2252.640 ;
        RECT 1367.670 2357.080 1367.950 2357.360 ;
        RECT 1367.670 2347.560 1367.950 2347.840 ;
        RECT 1367.670 2338.040 1367.950 2338.320 ;
        RECT 1367.670 2328.520 1367.950 2328.800 ;
        RECT 1367.210 2242.840 1367.490 2243.120 ;
        RECT 1367.210 2233.320 1367.490 2233.600 ;
        RECT 1367.210 2223.800 1367.490 2224.080 ;
        RECT 1367.210 2214.280 1367.490 2214.560 ;
        RECT 1367.210 2204.760 1367.490 2205.040 ;
        RECT 1367.210 2195.240 1367.490 2195.520 ;
        RECT 1366.290 2166.680 1366.570 2166.960 ;
        RECT 1366.290 2157.160 1366.570 2157.440 ;
        RECT 1366.290 2147.640 1366.570 2147.920 ;
        RECT 1366.290 2138.120 1366.570 2138.400 ;
        RECT 1366.290 2128.600 1366.570 2128.880 ;
        RECT 1367.210 2119.080 1367.490 2119.360 ;
        RECT 1367.210 2109.560 1367.490 2109.840 ;
        RECT 1367.210 2100.040 1367.490 2100.320 ;
        RECT 1367.210 2090.520 1367.490 2090.800 ;
        RECT 1367.210 2081.000 1367.490 2081.280 ;
        RECT 1367.210 2071.480 1367.490 2071.760 ;
        RECT 1367.210 2061.960 1367.490 2062.240 ;
        RECT 1367.210 2052.440 1367.490 2052.720 ;
        RECT 1367.210 2042.920 1367.490 2043.200 ;
        RECT 1367.210 2033.400 1367.490 2033.680 ;
        RECT 1367.210 2014.360 1367.490 2014.640 ;
        RECT 1367.210 2004.840 1367.490 2005.120 ;
        RECT 1367.210 1995.320 1367.490 1995.600 ;
        RECT 1367.210 1985.800 1367.490 1986.080 ;
        RECT 1367.210 1976.280 1367.490 1976.560 ;
        RECT 1367.210 1966.760 1367.490 1967.040 ;
        RECT 1367.210 1957.240 1367.490 1957.520 ;
        RECT 1367.670 1947.720 1367.950 1948.000 ;
        RECT 1368.130 1938.200 1368.410 1938.480 ;
        RECT 1367.670 1928.680 1367.950 1928.960 ;
        RECT 1366.290 1681.160 1366.570 1681.440 ;
        RECT 1366.750 1652.600 1367.030 1652.880 ;
        RECT 1367.670 1909.640 1367.950 1909.920 ;
        RECT 1368.130 1901.480 1368.410 1901.760 ;
        RECT 1368.130 1843.000 1368.410 1843.280 ;
        RECT 1369.050 1823.960 1369.330 1824.240 ;
        RECT 1367.670 1804.920 1367.950 1805.200 ;
        RECT 1369.050 1795.400 1369.330 1795.680 ;
        RECT 1369.050 1766.840 1369.330 1767.120 ;
        RECT 1367.670 1747.800 1367.950 1748.080 ;
        RECT 1367.670 1738.280 1367.950 1738.560 ;
        RECT 1367.670 1728.760 1367.950 1729.040 ;
        RECT 1368.130 1719.240 1368.410 1719.520 ;
        RECT 1367.670 1709.720 1367.950 1710.000 ;
        RECT 1367.670 1700.200 1367.950 1700.480 ;
        RECT 1371.350 2595.080 1371.630 2595.360 ;
        RECT 1370.430 2585.560 1370.710 2585.840 ;
        RECT 1370.890 2566.520 1371.170 2566.800 ;
        RECT 1371.350 2547.480 1371.630 2547.760 ;
        RECT 1372.270 1890.600 1372.550 1890.880 ;
        RECT 1372.270 1881.080 1372.550 1881.360 ;
        RECT 1372.270 1871.560 1372.550 1871.840 ;
        RECT 1372.270 1862.040 1372.550 1862.320 ;
        RECT 1372.270 1852.520 1372.550 1852.800 ;
        RECT 1373.190 2185.720 1373.470 2186.000 ;
        RECT 1373.650 2176.200 1373.930 2176.480 ;
        RECT 1373.190 1919.160 1373.470 1919.440 ;
        RECT 1372.730 1833.480 1373.010 1833.760 ;
        RECT 1371.810 1814.440 1372.090 1814.720 ;
        RECT 1371.810 1776.360 1372.090 1776.640 ;
        RECT 1372.730 1757.320 1373.010 1757.600 ;
        RECT 1369.510 1690.680 1369.790 1690.960 ;
        RECT 1369.050 1671.640 1369.330 1671.920 ;
        RECT 1371.350 1662.120 1371.630 1662.400 ;
        RECT 1369.970 1643.080 1370.250 1643.360 ;
        RECT 1367.670 1633.560 1367.950 1633.840 ;
        RECT 1367.210 1624.040 1367.490 1624.320 ;
        RECT 1367.670 1614.520 1367.950 1614.800 ;
        RECT 1688.750 2586.920 1689.030 2587.200 ;
        RECT 1994.190 2583.520 1994.470 2583.800 ;
        RECT 2001.090 2582.840 2001.370 2583.120 ;
        RECT 2007.990 2582.840 2008.270 2583.120 ;
        RECT 1691.970 2582.160 1692.250 2582.440 ;
        RECT 1704.390 2582.160 1704.670 2582.440 ;
        RECT 2016.730 2582.160 2017.010 2582.440 ;
        RECT 2021.790 2582.160 2022.070 2582.440 ;
        RECT 2030.070 2582.160 2030.350 2582.440 ;
        RECT 1600.890 2560.400 1601.170 2560.680 ;
        RECT 1583.410 2545.440 1583.690 2545.720 ;
        RECT 1597.210 2539.320 1597.490 2539.600 ;
        RECT 1593.990 1817.160 1594.270 1817.440 ;
        RECT 1601.810 2537.280 1602.090 2537.560 ;
        RECT 1599.050 2531.160 1599.330 2531.440 ;
        RECT 1600.890 2531.160 1601.170 2531.440 ;
        RECT 1599.050 2504.640 1599.330 2504.920 ;
        RECT 1603.650 2523.680 1603.930 2523.960 ;
        RECT 1602.730 2518.240 1603.010 2518.520 ;
        RECT 1600.890 2515.520 1601.170 2515.800 ;
        RECT 1599.970 2503.960 1600.250 2504.240 ;
        RECT 1601.810 2512.120 1602.090 2512.400 ;
        RECT 1601.350 2497.840 1601.630 2498.120 ;
        RECT 1599.050 2489.680 1599.330 2489.960 ;
        RECT 1601.350 2489.000 1601.630 2489.280 ;
        RECT 1600.890 2486.280 1601.170 2486.560 ;
        RECT 1599.050 2476.080 1599.330 2476.360 ;
        RECT 1599.050 2468.600 1599.330 2468.880 ;
        RECT 1600.890 2474.720 1601.170 2475.000 ;
        RECT 1599.970 2463.160 1600.250 2463.440 ;
        RECT 1599.050 2455.680 1599.330 2455.960 ;
        RECT 1600.890 2451.600 1601.170 2451.880 ;
        RECT 1600.430 2448.880 1600.710 2449.160 ;
        RECT 1602.270 2482.880 1602.550 2483.160 ;
        RECT 1601.810 2467.240 1602.090 2467.520 ;
        RECT 1601.350 2442.080 1601.630 2442.360 ;
        RECT 1599.050 2439.360 1599.330 2439.640 ;
        RECT 1600.890 2439.360 1601.170 2439.640 ;
        RECT 1601.350 2436.640 1601.630 2436.920 ;
        RECT 1598.590 2433.240 1598.870 2433.520 ;
        RECT 1599.050 2427.800 1599.330 2428.080 ;
        RECT 1600.890 2422.360 1601.170 2422.640 ;
        RECT 1599.050 2414.880 1599.330 2415.160 ;
        RECT 1600.890 2410.120 1601.170 2410.400 ;
        RECT 1603.190 2500.560 1603.470 2500.840 ;
        RECT 1604.110 2506.680 1604.390 2506.960 ;
        RECT 1603.650 2494.440 1603.930 2494.720 ;
        RECT 1602.730 2472.680 1603.010 2472.960 ;
        RECT 1602.270 2436.640 1602.550 2436.920 ;
        RECT 1604.110 2477.440 1604.390 2477.720 ;
        RECT 1603.190 2461.120 1603.470 2461.400 ;
        RECT 1603.190 2454.320 1603.470 2454.600 ;
        RECT 1603.650 2442.080 1603.930 2442.360 ;
        RECT 1602.270 2430.520 1602.550 2430.800 ;
        RECT 1601.810 2420.320 1602.090 2420.600 ;
        RECT 1599.050 2398.560 1599.330 2398.840 ;
        RECT 1600.890 2398.560 1601.170 2398.840 ;
        RECT 1600.890 2383.600 1601.170 2383.880 ;
        RECT 1602.730 2424.400 1603.010 2424.680 ;
        RECT 1603.650 2413.520 1603.930 2413.800 ;
        RECT 1603.190 2412.840 1603.470 2413.120 ;
        RECT 1602.270 2407.400 1602.550 2407.680 ;
        RECT 1603.190 2411.480 1603.470 2411.760 ;
        RECT 1602.730 2401.280 1603.010 2401.560 ;
        RECT 1601.810 2383.600 1602.090 2383.880 ;
        RECT 1600.890 2372.040 1601.170 2372.320 ;
        RECT 1602.270 2379.520 1602.550 2379.800 ;
        RECT 1601.350 2366.600 1601.630 2366.880 ;
        RECT 1601.350 2365.920 1601.630 2366.200 ;
        RECT 1600.890 2355.040 1601.170 2355.320 ;
        RECT 1603.190 2395.160 1603.470 2395.440 ;
        RECT 1603.190 2389.720 1603.470 2390.000 ;
        RECT 1603.650 2379.520 1603.930 2379.800 ;
        RECT 1603.190 2378.840 1603.470 2379.120 ;
        RECT 1601.810 2361.160 1602.090 2361.440 ;
        RECT 1601.810 2360.480 1602.090 2360.760 ;
        RECT 1601.350 2350.280 1601.630 2350.560 ;
        RECT 1601.350 2348.920 1601.630 2349.200 ;
        RECT 1600.890 2342.800 1601.170 2343.080 ;
        RECT 1602.730 2365.920 1603.010 2366.200 ;
        RECT 1602.270 2355.040 1602.550 2355.320 ;
        RECT 1602.270 2354.360 1602.550 2354.640 ;
        RECT 1601.810 2345.520 1602.090 2345.800 ;
        RECT 1604.110 2378.840 1604.390 2379.120 ;
        RECT 1604.110 2377.480 1604.390 2377.760 ;
        RECT 1603.650 2372.040 1603.930 2372.320 ;
        RECT 1603.190 2344.160 1603.470 2344.440 ;
        RECT 1600.890 2325.800 1601.170 2326.080 ;
        RECT 1600.890 2324.440 1601.170 2324.720 ;
        RECT 1603.190 2338.040 1603.470 2338.320 ;
        RECT 1600.890 1959.960 1601.170 1960.240 ;
        RECT 1602.270 2211.560 1602.550 2211.840 ;
        RECT 1603.650 2211.560 1603.930 2211.840 ;
        RECT 1601.350 1949.080 1601.630 1949.360 ;
        RECT 1600.430 1945.000 1600.710 1945.280 ;
        RECT 1693.350 1983.760 1693.630 1984.040 ;
        RECT 1987.290 1983.760 1987.570 1984.040 ;
        RECT 1994.190 1983.080 1994.470 1983.360 ;
        RECT 2001.090 1983.080 2001.370 1983.360 ;
        RECT 2007.990 1982.400 2008.270 1982.680 ;
        RECT 2016.730 1982.400 2017.010 1982.680 ;
        RECT 2021.790 1982.400 2022.070 1982.680 ;
        RECT 2030.070 1982.400 2030.350 1982.680 ;
        RECT 1601.350 1937.520 1601.630 1937.800 ;
        RECT 1601.810 1932.080 1602.090 1932.360 ;
        RECT 1600.890 1931.400 1601.170 1931.680 ;
        RECT 1600.890 1918.480 1601.170 1918.760 ;
        RECT 1601.350 1915.760 1601.630 1916.040 ;
        RECT 1603.190 1923.920 1603.470 1924.200 ;
        RECT 1601.810 1904.200 1602.090 1904.480 ;
        RECT 1601.350 1898.080 1601.630 1898.360 ;
        RECT 1600.890 1897.400 1601.170 1897.680 ;
        RECT 1600.890 1888.560 1601.170 1888.840 ;
        RECT 1599.050 1875.640 1599.330 1875.920 ;
        RECT 1600.890 1883.800 1601.170 1884.080 ;
        RECT 1602.270 1894.680 1602.550 1894.960 ;
        RECT 1601.810 1883.120 1602.090 1883.400 ;
        RECT 1601.350 1880.400 1601.630 1880.680 ;
        RECT 1600.890 1877.000 1601.170 1877.280 ;
        RECT 1599.970 1868.840 1600.250 1869.120 ;
        RECT 1600.430 1865.440 1600.710 1865.720 ;
        RECT 1600.890 1863.400 1601.170 1863.680 ;
        RECT 1601.810 1862.720 1602.090 1863.000 ;
        RECT 1601.350 1857.280 1601.630 1857.560 ;
        RECT 1600.890 1842.320 1601.170 1842.600 ;
        RECT 1603.650 1917.800 1603.930 1918.080 ;
        RECT 1603.190 1906.240 1603.470 1906.520 ;
        RECT 1604.110 1912.360 1604.390 1912.640 ;
        RECT 1604.110 1900.800 1604.390 1901.080 ;
        RECT 1602.730 1891.960 1603.010 1892.240 ;
        RECT 1602.730 1871.560 1603.010 1871.840 ;
        RECT 1604.110 1888.560 1604.390 1888.840 ;
        RECT 1603.650 1883.800 1603.930 1884.080 ;
        RECT 1603.190 1861.360 1603.470 1861.640 ;
        RECT 1604.110 1855.920 1604.390 1856.200 ;
        RECT 1602.270 1848.440 1602.550 1848.720 ;
        RECT 1601.810 1845.720 1602.090 1846.000 ;
        RECT 1601.350 1839.600 1601.630 1839.880 ;
        RECT 1599.050 1828.040 1599.330 1828.320 ;
        RECT 1600.890 1824.640 1601.170 1824.920 ;
        RECT 1599.970 1818.520 1600.250 1818.800 ;
        RECT 1599.050 1806.960 1599.330 1807.240 ;
        RECT 1600.430 1813.080 1600.710 1813.360 ;
        RECT 1600.890 1806.960 1601.170 1807.240 ;
        RECT 1603.650 1847.080 1603.930 1847.360 ;
        RECT 1603.190 1830.760 1603.470 1831.040 ;
        RECT 1602.270 1821.920 1602.550 1822.200 ;
        RECT 1601.810 1810.360 1602.090 1810.640 ;
        RECT 1601.350 1804.920 1601.630 1805.200 ;
        RECT 1601.350 1801.520 1601.630 1801.800 ;
        RECT 1602.270 1798.800 1602.550 1799.080 ;
        RECT 1601.810 1792.680 1602.090 1792.960 ;
        RECT 1601.350 1789.280 1601.630 1789.560 ;
        RECT 1600.890 1783.840 1601.170 1784.120 ;
        RECT 1600.890 1777.720 1601.170 1778.000 ;
        RECT 1600.890 1772.280 1601.170 1772.560 ;
        RECT 1603.190 1824.640 1603.470 1824.920 ;
        RECT 1602.730 1785.200 1603.010 1785.480 ;
        RECT 1601.350 1766.840 1601.630 1767.120 ;
        RECT 1601.350 1766.160 1601.630 1766.440 ;
        RECT 1600.890 1762.760 1601.170 1763.040 ;
        RECT 1604.110 1842.320 1604.390 1842.600 ;
        RECT 1604.110 1836.200 1604.390 1836.480 ;
        RECT 1603.650 1798.800 1603.930 1799.080 ;
        RECT 1603.190 1779.760 1603.470 1780.040 ;
        RECT 1601.810 1762.080 1602.090 1762.360 ;
        RECT 1603.190 1755.960 1603.470 1756.240 ;
        RECT 1601.810 1754.600 1602.090 1754.880 ;
        RECT 1600.890 1748.480 1601.170 1748.760 ;
        RECT 1604.110 1772.960 1604.390 1773.240 ;
        RECT 1604.110 1766.160 1604.390 1766.440 ;
        RECT 1603.650 1750.520 1603.930 1750.800 ;
        RECT 1600.890 1743.040 1601.170 1743.320 ;
        RECT 1600.890 1731.480 1601.170 1731.760 ;
        RECT 1367.210 1605.000 1367.490 1605.280 ;
      LAYER met3 ;
        RECT 759.280 3301.235 761.020 3302.140 ;
        RECT 781.040 3301.235 786.300 3302.140 ;
        RECT 1309.280 3301.235 1311.020 3302.140 ;
        RECT 1331.040 3301.235 1336.300 3302.140 ;
        RECT 400.000 3282.785 404.600 3283.085 ;
        RECT 392.905 3280.130 393.235 3280.145 ;
        RECT 400.510 3280.130 400.810 3282.785 ;
        RECT 392.905 3279.830 400.810 3280.130 ;
        RECT 392.905 3279.815 393.235 3279.830 ;
        RECT 400.000 3277.145 404.600 3277.445 ;
        RECT 392.445 3274.690 392.775 3274.705 ;
        RECT 400.510 3274.690 400.810 3277.145 ;
        RECT 392.445 3274.390 400.810 3274.690 ;
        RECT 392.445 3274.375 392.775 3274.390 ;
        RECT 400.000 3268.645 404.600 3268.945 ;
        RECT 391.985 3265.850 392.315 3265.865 ;
        RECT 400.510 3265.850 400.810 3268.645 ;
        RECT 391.985 3265.550 400.810 3265.850 ;
        RECT 391.985 3265.535 392.315 3265.550 ;
        RECT 400.000 3263.005 404.600 3263.305 ;
        RECT 391.525 3260.410 391.855 3260.425 ;
        RECT 400.510 3260.410 400.810 3263.005 ;
        RECT 391.525 3260.110 400.810 3260.410 ;
        RECT 391.525 3260.095 391.855 3260.110 ;
        RECT 400.000 3254.505 404.600 3254.805 ;
        RECT 393.365 3252.250 393.695 3252.265 ;
        RECT 400.510 3252.250 400.810 3254.505 ;
        RECT 393.365 3251.950 400.810 3252.250 ;
        RECT 393.365 3251.935 393.695 3251.950 ;
        RECT 400.000 3248.865 404.600 3249.165 ;
        RECT 393.825 3246.130 394.155 3246.145 ;
        RECT 400.510 3246.130 400.810 3248.865 ;
        RECT 393.825 3245.830 400.810 3246.130 ;
        RECT 393.825 3245.815 394.155 3245.830 ;
        RECT 400.000 3240.365 404.600 3240.665 ;
        RECT 391.065 3237.970 391.395 3237.985 ;
        RECT 400.510 3237.970 400.810 3240.365 ;
        RECT 391.065 3237.670 400.810 3237.970 ;
        RECT 391.065 3237.655 391.395 3237.670 ;
        RECT 400.000 2951.125 404.600 2951.425 ;
        RECT 394.285 2948.290 394.615 2948.305 ;
        RECT 400.510 2948.290 400.810 2951.125 ;
        RECT 394.285 2947.990 400.810 2948.290 ;
        RECT 394.285 2947.975 394.615 2947.990 ;
        RECT 400.000 2942.625 404.600 2942.925 ;
      LAYER met3 ;
        RECT 405.000 2855.000 781.480 3301.235 ;
      LAYER met3 ;
        RECT 781.480 3300.400 786.300 3301.235 ;
        RECT 781.880 3298.265 786.480 3298.565 ;
        RECT 781.480 3293.600 784.050 3294.660 ;
        RECT 950.000 3282.785 954.600 3283.085 ;
        RECT 938.465 3280.130 938.795 3280.145 ;
        RECT 950.670 3280.130 950.970 3282.785 ;
        RECT 938.465 3279.830 950.970 3280.130 ;
        RECT 938.465 3279.815 938.795 3279.830 ;
        RECT 950.000 3277.145 954.600 3277.445 ;
        RECT 941.685 3274.690 942.015 3274.705 ;
        RECT 950.670 3274.690 950.970 3277.145 ;
        RECT 941.685 3274.390 950.970 3274.690 ;
        RECT 941.685 3274.375 942.015 3274.390 ;
        RECT 950.000 3268.645 954.600 3268.945 ;
        RECT 942.145 3265.850 942.475 3265.865 ;
        RECT 950.670 3265.850 950.970 3268.645 ;
        RECT 942.145 3265.550 950.970 3265.850 ;
        RECT 942.145 3265.535 942.475 3265.550 ;
        RECT 950.000 3263.005 954.600 3263.305 ;
        RECT 942.605 3260.410 942.935 3260.425 ;
        RECT 950.670 3260.410 950.970 3263.005 ;
        RECT 942.605 3260.110 950.970 3260.410 ;
        RECT 942.605 3260.095 942.935 3260.110 ;
        RECT 950.000 3254.505 954.600 3254.805 ;
        RECT 943.065 3252.250 943.395 3252.265 ;
        RECT 950.670 3252.250 950.970 3254.505 ;
        RECT 943.065 3251.950 950.970 3252.250 ;
        RECT 943.065 3251.935 943.395 3251.950 ;
        RECT 950.000 3248.865 954.600 3249.165 ;
        RECT 943.525 3246.130 943.855 3246.145 ;
        RECT 950.670 3246.130 950.970 3248.865 ;
        RECT 943.525 3245.830 950.970 3246.130 ;
        RECT 943.525 3245.815 943.855 3245.830 ;
        RECT 950.000 3240.365 954.600 3240.665 ;
        RECT 943.985 3237.970 944.315 3237.985 ;
        RECT 950.670 3237.970 950.970 3240.365 ;
        RECT 943.985 3237.670 950.970 3237.970 ;
        RECT 943.985 3237.655 944.315 3237.670 ;
        RECT 781.880 2996.910 786.480 2997.210 ;
        RECT 781.880 2988.410 786.480 2988.710 ;
        RECT 781.880 2982.770 786.480 2983.070 ;
        RECT 781.880 2974.270 786.480 2974.570 ;
        RECT 781.880 2968.630 786.480 2968.930 ;
        RECT 781.880 2960.130 786.480 2960.430 ;
        RECT 781.880 2954.490 786.480 2954.790 ;
        RECT 950.000 2951.125 954.600 2951.425 ;
        RECT 944.445 2948.290 944.775 2948.305 ;
        RECT 950.670 2948.290 950.970 2951.125 ;
        RECT 944.445 2947.990 950.970 2948.290 ;
        RECT 944.445 2947.975 944.775 2947.990 ;
        RECT 950.000 2942.625 954.600 2942.925 ;
      LAYER met3 ;
        RECT 955.000 2855.000 1331.480 3301.235 ;
      LAYER met3 ;
        RECT 1331.480 3300.400 1336.300 3301.235 ;
        RECT 1331.880 3298.265 1336.480 3298.565 ;
        RECT 1331.480 3293.600 1334.050 3294.660 ;
        RECT 1331.880 2996.910 1336.480 2997.210 ;
        RECT 1331.880 2988.410 1336.480 2988.710 ;
        RECT 1331.880 2982.770 1336.480 2983.070 ;
        RECT 1331.880 2974.270 1336.480 2974.570 ;
        RECT 1331.880 2968.630 1336.480 2968.930 ;
        RECT 1331.880 2960.130 1336.480 2960.430 ;
        RECT 1331.880 2954.490 1336.480 2954.790 ;
        RECT 516.645 2851.730 516.975 2851.745 ;
        RECT 517.310 2851.730 517.690 2851.740 ;
        RECT 516.645 2851.430 517.690 2851.730 ;
        RECT 516.645 2851.415 516.975 2851.430 ;
        RECT 517.310 2851.420 517.690 2851.430 ;
        RECT 1103.605 2851.060 1103.935 2851.065 ;
        RECT 1103.350 2851.050 1103.935 2851.060 ;
        RECT 1103.350 2850.750 1104.160 2851.050 ;
        RECT 1103.350 2850.740 1103.935 2850.750 ;
        RECT 1103.605 2850.735 1103.935 2850.740 ;
        RECT 568.910 2848.330 569.290 2848.340 ;
        RECT 572.305 2848.330 572.635 2848.345 ;
        RECT 568.910 2848.030 572.635 2848.330 ;
        RECT 568.910 2848.020 569.290 2848.030 ;
        RECT 572.305 2848.015 572.635 2848.030 ;
        RECT 592.270 2848.330 592.650 2848.340 ;
        RECT 600.365 2848.330 600.695 2848.345 ;
        RECT 1089.345 2848.340 1089.675 2848.345 ;
        RECT 1089.090 2848.330 1089.675 2848.340 ;
        RECT 592.270 2848.030 600.695 2848.330 ;
        RECT 1088.890 2848.030 1089.675 2848.330 ;
        RECT 592.270 2848.020 592.650 2848.030 ;
        RECT 600.365 2848.015 600.695 2848.030 ;
        RECT 1089.090 2848.020 1089.675 2848.030 ;
        RECT 1089.345 2848.015 1089.675 2848.020 ;
        RECT 597.145 2845.620 597.475 2845.625 ;
        RECT 604.965 2845.620 605.295 2845.625 ;
        RECT 597.145 2845.610 597.730 2845.620 ;
        RECT 604.710 2845.610 605.295 2845.620 ;
        RECT 597.145 2845.310 597.930 2845.610 ;
        RECT 604.510 2845.310 605.295 2845.610 ;
        RECT 597.145 2845.300 597.730 2845.310 ;
        RECT 604.710 2845.300 605.295 2845.310 ;
        RECT 597.145 2845.295 597.475 2845.300 ;
        RECT 604.965 2845.295 605.295 2845.300 ;
        RECT 612.990 2844.250 613.370 2844.260 ;
        RECT 613.705 2844.250 614.035 2844.265 ;
        RECT 612.990 2843.950 614.035 2844.250 ;
        RECT 612.990 2843.940 613.370 2843.950 ;
        RECT 613.705 2843.935 614.035 2843.950 ;
        RECT 573.685 2843.580 574.015 2843.585 ;
        RECT 573.430 2843.570 574.015 2843.580 ;
        RECT 573.230 2843.270 574.015 2843.570 ;
        RECT 573.430 2843.260 574.015 2843.270 ;
        RECT 575.270 2843.570 575.650 2843.580 ;
        RECT 590.245 2843.570 590.575 2843.585 ;
        RECT 575.270 2843.270 590.575 2843.570 ;
        RECT 575.270 2843.260 575.650 2843.270 ;
        RECT 573.685 2843.255 574.015 2843.260 ;
        RECT 590.245 2843.255 590.575 2843.270 ;
        RECT 432.670 2842.890 433.050 2842.900 ;
        RECT 433.845 2842.890 434.175 2842.905 ;
        RECT 432.670 2842.590 434.175 2842.890 ;
        RECT 432.670 2842.580 433.050 2842.590 ;
        RECT 433.845 2842.575 434.175 2842.590 ;
        RECT 507.190 2842.890 507.570 2842.900 ;
        RECT 509.745 2842.890 510.075 2842.905 ;
        RECT 524.005 2842.900 524.335 2842.905 ;
        RECT 507.190 2842.590 510.075 2842.890 ;
        RECT 507.190 2842.580 507.570 2842.590 ;
        RECT 509.745 2842.575 510.075 2842.590 ;
        RECT 523.750 2842.890 524.335 2842.900 ;
        RECT 526.305 2842.900 526.635 2842.905 ;
        RECT 526.305 2842.890 526.890 2842.900 ;
        RECT 529.270 2842.890 529.650 2842.900 ;
        RECT 530.905 2842.890 531.235 2842.905 ;
        RECT 523.750 2842.590 524.560 2842.890 ;
        RECT 526.305 2842.590 527.090 2842.890 ;
        RECT 529.270 2842.590 531.235 2842.890 ;
        RECT 523.750 2842.580 524.335 2842.590 ;
        RECT 524.005 2842.575 524.335 2842.580 ;
        RECT 526.305 2842.580 526.890 2842.590 ;
        RECT 529.270 2842.580 529.650 2842.590 ;
        RECT 526.305 2842.575 526.635 2842.580 ;
        RECT 530.905 2842.575 531.235 2842.590 ;
        RECT 533.870 2842.890 534.250 2842.900 ;
        RECT 537.805 2842.890 538.135 2842.905 ;
        RECT 533.870 2842.590 538.135 2842.890 ;
        RECT 533.870 2842.580 534.250 2842.590 ;
        RECT 537.805 2842.575 538.135 2842.590 ;
        RECT 543.070 2842.890 543.450 2842.900 ;
        RECT 544.705 2842.890 545.035 2842.905 ;
        RECT 543.070 2842.590 545.035 2842.890 ;
        RECT 543.070 2842.580 543.450 2842.590 ;
        RECT 544.705 2842.575 545.035 2842.590 ;
        RECT 557.790 2842.890 558.170 2842.900 ;
        RECT 558.505 2842.890 558.835 2842.905 ;
        RECT 557.790 2842.590 558.835 2842.890 ;
        RECT 557.790 2842.580 558.170 2842.590 ;
        RECT 558.505 2842.575 558.835 2842.590 ;
        RECT 642.225 2842.900 642.555 2842.905 ;
        RECT 642.225 2842.890 642.810 2842.900 ;
        RECT 979.865 2842.890 980.195 2842.905 ;
        RECT 980.990 2842.890 981.370 2842.900 ;
        RECT 642.225 2842.590 643.010 2842.890 ;
        RECT 979.865 2842.590 981.370 2842.890 ;
        RECT 642.225 2842.580 642.810 2842.590 ;
        RECT 642.225 2842.575 642.555 2842.580 ;
        RECT 979.865 2842.575 980.195 2842.590 ;
        RECT 980.990 2842.580 981.370 2842.590 ;
        RECT 987.225 2842.890 987.555 2842.905 ;
        RECT 988.350 2842.890 988.730 2842.900 ;
        RECT 987.225 2842.590 988.730 2842.890 ;
        RECT 987.225 2842.575 987.555 2842.590 ;
        RECT 988.350 2842.580 988.730 2842.590 ;
        RECT 1019.630 2842.890 1020.010 2842.900 ;
        RECT 1020.805 2842.890 1021.135 2842.905 ;
        RECT 1019.630 2842.590 1021.135 2842.890 ;
        RECT 1019.630 2842.580 1020.010 2842.590 ;
        RECT 1020.805 2842.575 1021.135 2842.590 ;
        RECT 1024.025 2842.900 1024.355 2842.905 ;
        RECT 1024.025 2842.890 1024.610 2842.900 ;
        RECT 1026.990 2842.890 1027.370 2842.900 ;
        RECT 1027.705 2842.890 1028.035 2842.905 ;
        RECT 1024.025 2842.590 1024.810 2842.890 ;
        RECT 1026.990 2842.590 1028.035 2842.890 ;
        RECT 1024.025 2842.580 1024.610 2842.590 ;
        RECT 1026.990 2842.580 1027.370 2842.590 ;
        RECT 1024.025 2842.575 1024.355 2842.580 ;
        RECT 1027.705 2842.575 1028.035 2842.590 ;
        RECT 1065.425 2842.900 1065.755 2842.905 ;
        RECT 1070.485 2842.900 1070.815 2842.905 ;
        RECT 1111.885 2842.900 1112.215 2842.905 ;
        RECT 1118.325 2842.900 1118.655 2842.905 ;
        RECT 1131.205 2842.900 1131.535 2842.905 ;
        RECT 1135.805 2842.900 1136.135 2842.905 ;
        RECT 1065.425 2842.890 1066.010 2842.900 ;
        RECT 1070.230 2842.890 1070.815 2842.900 ;
        RECT 1111.630 2842.890 1112.215 2842.900 ;
        RECT 1118.070 2842.890 1118.655 2842.900 ;
        RECT 1065.425 2842.590 1066.210 2842.890 ;
        RECT 1070.030 2842.590 1070.815 2842.890 ;
        RECT 1111.430 2842.590 1112.215 2842.890 ;
        RECT 1117.870 2842.590 1118.655 2842.890 ;
        RECT 1065.425 2842.580 1066.010 2842.590 ;
        RECT 1070.230 2842.580 1070.815 2842.590 ;
        RECT 1111.630 2842.580 1112.215 2842.590 ;
        RECT 1118.070 2842.580 1118.655 2842.590 ;
        RECT 1130.950 2842.890 1131.535 2842.900 ;
        RECT 1135.550 2842.890 1136.135 2842.900 ;
        RECT 1130.950 2842.590 1131.760 2842.890 ;
        RECT 1135.350 2842.590 1136.135 2842.890 ;
        RECT 1130.950 2842.580 1131.535 2842.590 ;
        RECT 1135.550 2842.580 1136.135 2842.590 ;
        RECT 1136.470 2842.890 1136.850 2842.900 ;
        RECT 1138.105 2842.890 1138.435 2842.905 ;
        RECT 1136.470 2842.590 1138.435 2842.890 ;
        RECT 1136.470 2842.580 1136.850 2842.590 ;
        RECT 1065.425 2842.575 1065.755 2842.580 ;
        RECT 1070.485 2842.575 1070.815 2842.580 ;
        RECT 1111.885 2842.575 1112.215 2842.580 ;
        RECT 1118.325 2842.575 1118.655 2842.580 ;
        RECT 1131.205 2842.575 1131.535 2842.580 ;
        RECT 1135.805 2842.575 1136.135 2842.580 ;
        RECT 1138.105 2842.575 1138.435 2842.590 ;
        RECT 1143.830 2842.890 1144.210 2842.900 ;
        RECT 1145.005 2842.890 1145.335 2842.905 ;
        RECT 1143.830 2842.590 1145.335 2842.890 ;
        RECT 1143.830 2842.580 1144.210 2842.590 ;
        RECT 1145.005 2842.575 1145.335 2842.590 ;
        RECT 1151.190 2842.890 1151.570 2842.900 ;
        RECT 1151.905 2842.890 1152.235 2842.905 ;
        RECT 1151.190 2842.590 1152.235 2842.890 ;
        RECT 1151.190 2842.580 1151.570 2842.590 ;
        RECT 1151.905 2842.575 1152.235 2842.590 ;
        RECT 1153.950 2842.890 1154.330 2842.900 ;
        RECT 1158.805 2842.890 1159.135 2842.905 ;
        RECT 1165.245 2842.900 1165.575 2842.905 ;
        RECT 1172.605 2842.900 1172.935 2842.905 ;
        RECT 1153.950 2842.590 1159.135 2842.890 ;
        RECT 1153.950 2842.580 1154.330 2842.590 ;
        RECT 1158.805 2842.575 1159.135 2842.590 ;
        RECT 1164.990 2842.890 1165.575 2842.900 ;
        RECT 1172.350 2842.890 1172.935 2842.900 ;
        RECT 1178.790 2842.890 1179.170 2842.900 ;
        RECT 1179.505 2842.890 1179.835 2842.905 ;
        RECT 1186.405 2842.900 1186.735 2842.905 ;
        RECT 1164.990 2842.590 1165.800 2842.890 ;
        RECT 1172.350 2842.590 1173.160 2842.890 ;
        RECT 1178.790 2842.590 1179.835 2842.890 ;
        RECT 1164.990 2842.580 1165.575 2842.590 ;
        RECT 1172.350 2842.580 1172.935 2842.590 ;
        RECT 1178.790 2842.580 1179.170 2842.590 ;
        RECT 1165.245 2842.575 1165.575 2842.580 ;
        RECT 1172.605 2842.575 1172.935 2842.580 ;
        RECT 1179.505 2842.575 1179.835 2842.590 ;
        RECT 1186.150 2842.890 1186.735 2842.900 ;
        RECT 1190.750 2842.890 1191.130 2842.900 ;
        RECT 1193.305 2842.890 1193.635 2842.905 ;
        RECT 1186.150 2842.590 1186.960 2842.890 ;
        RECT 1190.750 2842.590 1193.635 2842.890 ;
        RECT 1186.150 2842.580 1186.735 2842.590 ;
        RECT 1190.750 2842.580 1191.130 2842.590 ;
        RECT 1186.405 2842.575 1186.735 2842.580 ;
        RECT 1193.305 2842.575 1193.635 2842.590 ;
        RECT 475.705 2842.220 476.035 2842.225 ;
        RECT 549.305 2842.220 549.635 2842.225 ;
        RECT 1018.505 2842.220 1018.835 2842.225 ;
        RECT 475.705 2842.210 476.290 2842.220 ;
        RECT 475.480 2841.910 476.290 2842.210 ;
        RECT 475.705 2841.900 476.290 2841.910 ;
        RECT 549.305 2842.210 549.890 2842.220 ;
        RECT 1018.505 2842.210 1019.090 2842.220 ;
        RECT 1128.190 2842.210 1128.570 2842.220 ;
        RECT 1130.745 2842.210 1131.075 2842.225 ;
        RECT 549.305 2841.910 550.090 2842.210 ;
        RECT 1018.505 2841.910 1019.290 2842.210 ;
        RECT 1128.190 2841.910 1131.075 2842.210 ;
        RECT 549.305 2841.900 549.890 2841.910 ;
        RECT 1018.505 2841.900 1019.090 2841.910 ;
        RECT 1128.190 2841.900 1128.570 2841.910 ;
        RECT 475.705 2841.895 476.035 2841.900 ;
        RECT 549.305 2841.895 549.635 2841.900 ;
        RECT 1018.505 2841.895 1018.835 2841.900 ;
        RECT 1130.745 2841.895 1131.075 2841.910 ;
        RECT 1163.150 2842.210 1163.530 2842.220 ;
        RECT 1165.705 2842.210 1166.035 2842.225 ;
        RECT 1163.150 2841.910 1166.035 2842.210 ;
        RECT 1163.150 2841.900 1163.530 2841.910 ;
        RECT 1165.705 2841.895 1166.035 2841.910 ;
        RECT 480.510 2841.530 480.890 2841.540 ;
        RECT 482.605 2841.530 482.935 2841.545 ;
        RECT 480.510 2841.230 482.935 2841.530 ;
        RECT 480.510 2841.220 480.890 2841.230 ;
        RECT 482.605 2841.215 482.935 2841.230 ;
        RECT 504.430 2841.530 504.810 2841.540 ;
        RECT 510.205 2841.530 510.535 2841.545 ;
        RECT 504.430 2841.230 510.535 2841.530 ;
        RECT 504.430 2841.220 504.810 2841.230 ;
        RECT 510.205 2841.215 510.535 2841.230 ;
        RECT 618.510 2841.530 618.890 2841.540 ;
        RECT 620.605 2841.530 620.935 2841.545 ;
        RECT 621.525 2841.540 621.855 2841.545 ;
        RECT 618.510 2841.230 620.935 2841.530 ;
        RECT 618.510 2841.220 618.890 2841.230 ;
        RECT 620.605 2841.215 620.935 2841.230 ;
        RECT 621.270 2841.530 621.855 2841.540 ;
        RECT 626.790 2841.530 627.170 2841.540 ;
        RECT 627.505 2841.530 627.835 2841.545 ;
        RECT 621.270 2841.230 622.080 2841.530 ;
        RECT 626.790 2841.230 627.835 2841.530 ;
        RECT 621.270 2841.220 621.855 2841.230 ;
        RECT 626.790 2841.220 627.170 2841.230 ;
        RECT 621.525 2841.215 621.855 2841.220 ;
        RECT 627.505 2841.215 627.835 2841.230 ;
        RECT 647.950 2841.530 648.330 2841.540 ;
        RECT 727.785 2841.530 728.115 2841.545 ;
        RECT 647.950 2841.230 728.115 2841.530 ;
        RECT 647.950 2841.220 648.330 2841.230 ;
        RECT 727.785 2841.215 728.115 2841.230 ;
        RECT 379.105 2840.850 379.435 2840.865 ;
        RECT 1001.230 2840.850 1001.610 2840.860 ;
        RECT 379.105 2840.550 1001.610 2840.850 ;
        RECT 379.105 2840.535 379.435 2840.550 ;
        RECT 1001.230 2840.540 1001.610 2840.550 ;
        RECT 1159.725 2840.850 1160.055 2840.865 ;
        RECT 1164.070 2840.850 1164.450 2840.860 ;
        RECT 1159.725 2840.550 1164.450 2840.850 ;
        RECT 1159.725 2840.535 1160.055 2840.550 ;
        RECT 1164.070 2840.540 1164.450 2840.550 ;
        RECT 1179.965 2840.850 1180.295 2840.865 ;
        RECT 1180.630 2840.850 1181.010 2840.860 ;
        RECT 1179.965 2840.550 1181.010 2840.850 ;
        RECT 1179.965 2840.535 1180.295 2840.550 ;
        RECT 1180.630 2840.540 1181.010 2840.550 ;
        RECT 386.005 2840.170 386.335 2840.185 ;
        RECT 1159.265 2840.180 1159.595 2840.185 ;
        RECT 1007.670 2840.170 1008.050 2840.180 ;
        RECT 1159.265 2840.170 1159.850 2840.180 ;
        RECT 386.005 2839.870 1008.050 2840.170 ;
        RECT 1159.040 2839.870 1159.850 2840.170 ;
        RECT 386.005 2839.855 386.335 2839.870 ;
        RECT 1007.670 2839.860 1008.050 2839.870 ;
        RECT 1159.265 2839.860 1159.850 2839.870 ;
        RECT 1159.265 2839.855 1159.595 2839.860 ;
        RECT 455.465 2838.810 455.795 2838.825 ;
        RECT 457.510 2838.810 457.890 2838.820 ;
        RECT 455.465 2838.510 457.890 2838.810 ;
        RECT 455.465 2838.495 455.795 2838.510 ;
        RECT 457.510 2838.500 457.890 2838.510 ;
        RECT 488.790 2838.810 489.170 2838.820 ;
        RECT 489.505 2838.810 489.835 2838.825 ;
        RECT 488.790 2838.510 489.835 2838.810 ;
        RECT 488.790 2838.500 489.170 2838.510 ;
        RECT 489.505 2838.495 489.835 2838.510 ;
        RECT 501.670 2838.810 502.050 2838.820 ;
        RECT 503.305 2838.810 503.635 2838.825 ;
        RECT 551.605 2838.820 551.935 2838.825 ;
        RECT 501.670 2838.510 503.635 2838.810 ;
        RECT 501.670 2838.500 502.050 2838.510 ;
        RECT 503.305 2838.495 503.635 2838.510 ;
        RECT 551.350 2838.810 551.935 2838.820 ;
        RECT 551.350 2838.510 552.160 2838.810 ;
        RECT 551.350 2838.500 551.935 2838.510 ;
        RECT 551.605 2838.495 551.935 2838.500 ;
        RECT 441.665 2837.450 441.995 2837.465 ;
        RECT 442.790 2837.450 443.170 2837.460 ;
        RECT 441.665 2837.150 443.170 2837.450 ;
        RECT 441.665 2837.135 441.995 2837.150 ;
        RECT 442.790 2837.140 443.170 2837.150 ;
        RECT 434.765 2836.770 435.095 2836.785 ;
        RECT 449.945 2836.780 450.275 2836.785 ;
        RECT 437.270 2836.770 437.650 2836.780 ;
        RECT 449.945 2836.770 450.530 2836.780 ;
        RECT 434.765 2836.470 437.650 2836.770 ;
        RECT 449.720 2836.470 450.530 2836.770 ;
        RECT 434.765 2836.455 435.095 2836.470 ;
        RECT 437.270 2836.460 437.650 2836.470 ;
        RECT 449.945 2836.460 450.530 2836.470 ;
        RECT 621.270 2836.770 621.650 2836.780 ;
        RECT 625.205 2836.770 625.535 2836.785 ;
        RECT 621.270 2836.470 625.535 2836.770 ;
        RECT 621.270 2836.460 621.650 2836.470 ;
        RECT 449.945 2836.455 450.275 2836.460 ;
        RECT 625.205 2836.455 625.535 2836.470 ;
        RECT 1041.710 2836.770 1042.090 2836.780 ;
        RECT 1045.185 2836.770 1045.515 2836.785 ;
        RECT 1041.710 2836.470 1045.515 2836.770 ;
        RECT 1041.710 2836.460 1042.090 2836.470 ;
        RECT 1045.185 2836.455 1045.515 2836.470 ;
        RECT 466.710 2836.090 467.090 2836.100 ;
        RECT 468.345 2836.090 468.675 2836.105 ;
        RECT 466.710 2835.790 468.675 2836.090 ;
        RECT 466.710 2835.780 467.090 2835.790 ;
        RECT 468.345 2835.775 468.675 2835.790 ;
        RECT 471.310 2836.090 471.690 2836.100 ;
        RECT 475.245 2836.090 475.575 2836.105 ;
        RECT 471.310 2835.790 475.575 2836.090 ;
        RECT 471.310 2835.780 471.690 2835.790 ;
        RECT 475.245 2835.775 475.575 2835.790 ;
        RECT 481.430 2836.090 481.810 2836.100 ;
        RECT 482.145 2836.090 482.475 2836.105 ;
        RECT 481.430 2835.790 482.475 2836.090 ;
        RECT 481.430 2835.780 481.810 2835.790 ;
        RECT 482.145 2835.775 482.475 2835.790 ;
        RECT 494.310 2836.090 494.690 2836.100 ;
        RECT 495.945 2836.090 496.275 2836.105 ;
        RECT 494.310 2835.790 496.275 2836.090 ;
        RECT 494.310 2835.780 494.690 2835.790 ;
        RECT 495.945 2835.775 496.275 2835.790 ;
        RECT 624.030 2836.090 624.410 2836.100 ;
        RECT 626.585 2836.090 626.915 2836.105 ;
        RECT 624.030 2835.790 626.915 2836.090 ;
        RECT 624.030 2835.780 624.410 2835.790 ;
        RECT 626.585 2835.775 626.915 2835.790 ;
        RECT 633.230 2836.090 633.610 2836.100 ;
        RECT 634.405 2836.090 634.735 2836.105 ;
        RECT 640.845 2836.100 641.175 2836.105 ;
        RECT 633.230 2835.790 634.735 2836.090 ;
        RECT 633.230 2835.780 633.610 2835.790 ;
        RECT 634.405 2835.775 634.735 2835.790 ;
        RECT 640.590 2836.090 641.175 2836.100 ;
        RECT 1039.870 2836.090 1040.250 2836.100 ;
        RECT 1041.505 2836.090 1041.835 2836.105 ;
        RECT 640.590 2835.790 641.400 2836.090 ;
        RECT 1039.870 2835.790 1041.835 2836.090 ;
        RECT 640.590 2835.780 641.175 2835.790 ;
        RECT 1039.870 2835.780 1040.250 2835.790 ;
        RECT 640.845 2835.775 641.175 2835.780 ;
        RECT 1041.505 2835.775 1041.835 2835.790 ;
        RECT 1046.310 2836.090 1046.690 2836.100 ;
        RECT 1048.405 2836.090 1048.735 2836.105 ;
        RECT 1054.845 2836.100 1055.175 2836.105 ;
        RECT 1062.205 2836.100 1062.535 2836.105 ;
        RECT 1046.310 2835.790 1048.735 2836.090 ;
        RECT 1046.310 2835.780 1046.690 2835.790 ;
        RECT 1048.405 2835.775 1048.735 2835.790 ;
        RECT 1054.590 2836.090 1055.175 2836.100 ;
        RECT 1061.950 2836.090 1062.535 2836.100 ;
        RECT 1067.470 2836.090 1067.850 2836.100 ;
        RECT 1069.105 2836.090 1069.435 2836.105 ;
        RECT 1054.590 2835.790 1055.400 2836.090 ;
        RECT 1061.950 2835.790 1062.760 2836.090 ;
        RECT 1067.470 2835.790 1069.435 2836.090 ;
        RECT 1054.590 2835.780 1055.175 2835.790 ;
        RECT 1061.950 2835.780 1062.535 2835.790 ;
        RECT 1067.470 2835.780 1067.850 2835.790 ;
        RECT 1054.845 2835.775 1055.175 2835.780 ;
        RECT 1062.205 2835.775 1062.535 2835.780 ;
        RECT 1069.105 2835.775 1069.435 2835.790 ;
        RECT 1073.910 2836.090 1074.290 2836.100 ;
        RECT 1076.005 2836.090 1076.335 2836.105 ;
        RECT 1073.910 2835.790 1076.335 2836.090 ;
        RECT 1073.910 2835.780 1074.290 2835.790 ;
        RECT 1076.005 2835.775 1076.335 2835.790 ;
        RECT 1081.270 2836.090 1081.650 2836.100 ;
        RECT 1082.905 2836.090 1083.235 2836.105 ;
        RECT 1089.345 2836.100 1089.675 2836.105 ;
        RECT 1089.345 2836.090 1089.930 2836.100 ;
        RECT 1081.270 2835.790 1083.235 2836.090 ;
        RECT 1089.120 2835.790 1089.930 2836.090 ;
        RECT 1081.270 2835.780 1081.650 2835.790 ;
        RECT 1082.905 2835.775 1083.235 2835.790 ;
        RECT 1089.345 2835.780 1089.930 2835.790 ;
        RECT 1095.990 2836.090 1096.370 2836.100 ;
        RECT 1096.705 2836.090 1097.035 2836.105 ;
        RECT 1095.990 2835.790 1097.035 2836.090 ;
        RECT 1095.990 2835.780 1096.370 2835.790 ;
        RECT 1089.345 2835.775 1089.675 2835.780 ;
        RECT 1096.705 2835.775 1097.035 2835.790 ;
        RECT 1109.790 2836.090 1110.170 2836.100 ;
        RECT 1110.505 2836.090 1110.835 2836.105 ;
        RECT 1109.790 2835.790 1110.835 2836.090 ;
        RECT 1109.790 2835.780 1110.170 2835.790 ;
        RECT 1110.505 2835.775 1110.835 2835.790 ;
        RECT 1116.230 2836.090 1116.610 2836.100 ;
        RECT 1117.405 2836.090 1117.735 2836.105 ;
        RECT 1116.230 2835.790 1117.735 2836.090 ;
        RECT 1116.230 2835.780 1116.610 2835.790 ;
        RECT 1117.405 2835.775 1117.735 2835.790 ;
        RECT 1118.990 2836.090 1119.370 2836.100 ;
        RECT 1124.305 2836.090 1124.635 2836.105 ;
        RECT 1118.990 2835.790 1124.635 2836.090 ;
        RECT 1118.990 2835.780 1119.370 2835.790 ;
        RECT 1124.305 2835.775 1124.635 2835.790 ;
        RECT 586.310 2832.690 586.690 2832.700 ;
        RECT 592.545 2832.690 592.875 2832.705 ;
        RECT 586.310 2832.390 592.875 2832.690 ;
        RECT 586.310 2832.380 586.690 2832.390 ;
        RECT 592.545 2832.375 592.875 2832.390 ;
        RECT 762.285 2621.210 762.615 2621.225 ;
        RECT 1021.725 2621.210 1022.055 2621.225 ;
        RECT 762.285 2620.910 1022.055 2621.210 ;
        RECT 762.285 2620.895 762.615 2620.910 ;
        RECT 1021.725 2620.895 1022.055 2620.910 ;
        RECT 727.785 2620.530 728.115 2620.545 ;
        RECT 1050.245 2620.530 1050.575 2620.545 ;
        RECT 727.785 2620.230 1050.575 2620.530 ;
        RECT 727.785 2620.215 728.115 2620.230 ;
        RECT 1050.245 2620.215 1050.575 2620.230 ;
        RECT 626.585 2619.850 626.915 2619.865 ;
        RECT 1012.065 2619.850 1012.395 2619.865 ;
        RECT 626.585 2619.550 1012.395 2619.850 ;
        RECT 626.585 2619.535 626.915 2619.550 ;
        RECT 1012.065 2619.535 1012.395 2619.550 ;
        RECT 634.405 2619.170 634.735 2619.185 ;
        RECT 1030.925 2619.170 1031.255 2619.185 ;
        RECT 634.405 2618.870 1031.255 2619.170 ;
        RECT 634.405 2618.855 634.735 2618.870 ;
        RECT 1030.925 2618.855 1031.255 2618.870 ;
        RECT 354.725 2618.490 355.055 2618.505 ;
        RECT 987.225 2618.490 987.555 2618.505 ;
        RECT 354.725 2618.190 987.555 2618.490 ;
        RECT 354.725 2618.175 355.055 2618.190 ;
        RECT 987.225 2618.175 987.555 2618.190 ;
        RECT 1355.930 2604.890 1359.930 2605.000 ;
        RECT 1369.945 2604.890 1370.275 2604.905 ;
      LAYER met3 ;
        RECT 357.355 2604.000 1355.530 2604.865 ;
      LAYER met3 ;
        RECT 1355.930 2604.590 1370.275 2604.890 ;
        RECT 1355.930 2604.400 1359.930 2604.590 ;
        RECT 1369.945 2604.575 1370.275 2604.590 ;
      LAYER met3 ;
        RECT 357.355 2595.880 1355.930 2604.000 ;
        RECT 357.355 2594.480 1355.530 2595.880 ;
      LAYER met3 ;
        RECT 1355.930 2595.370 1359.930 2595.480 ;
        RECT 1371.325 2595.370 1371.655 2595.385 ;
        RECT 1355.930 2595.070 1371.655 2595.370 ;
        RECT 1355.930 2594.880 1359.930 2595.070 ;
        RECT 1371.325 2595.055 1371.655 2595.070 ;
      LAYER met3 ;
        RECT 357.355 2586.360 1355.930 2594.480 ;
      LAYER met3 ;
        RECT 1688.725 2587.210 1689.055 2587.225 ;
        RECT 1688.725 2586.910 1701.425 2587.210 ;
        RECT 1688.725 2586.895 1689.055 2586.910 ;
      LAYER met3 ;
        RECT 357.355 2584.960 1355.530 2586.360 ;
      LAYER met3 ;
        RECT 1355.930 2585.850 1359.930 2585.960 ;
        RECT 1370.405 2585.850 1370.735 2585.865 ;
        RECT 1355.930 2585.550 1370.735 2585.850 ;
        RECT 1355.930 2585.360 1359.930 2585.550 ;
        RECT 1370.405 2585.535 1370.735 2585.550 ;
      LAYER met3 ;
        RECT 357.355 2576.840 1355.930 2584.960 ;
      LAYER met3 ;
        RECT 1369.230 2582.450 1369.610 2582.460 ;
        RECT 1691.945 2582.450 1692.275 2582.465 ;
        RECT 1369.230 2582.150 1692.275 2582.450 ;
        RECT 1369.230 2582.140 1369.610 2582.150 ;
        RECT 1691.945 2582.135 1692.275 2582.150 ;
        RECT 1692.625 2581.880 1692.925 2586.480 ;
        RECT 1701.125 2581.880 1701.425 2586.910 ;
        RECT 1704.365 2582.450 1704.695 2582.465 ;
        RECT 1990.365 2582.450 1990.665 2586.480 ;
        RECT 1994.165 2583.810 1994.495 2583.825 ;
        RECT 1998.865 2583.810 1999.165 2586.480 ;
        RECT 1994.165 2583.510 1999.165 2583.810 ;
        RECT 1994.165 2583.495 1994.495 2583.510 ;
        RECT 1704.365 2582.150 1990.665 2582.450 ;
        RECT 1704.365 2582.135 1704.695 2582.150 ;
        RECT 1990.365 2581.880 1990.665 2582.150 ;
        RECT 1998.865 2581.880 1999.165 2583.510 ;
        RECT 2001.065 2583.130 2001.395 2583.145 ;
        RECT 2004.505 2583.130 2004.805 2586.480 ;
        RECT 2001.065 2582.830 2004.805 2583.130 ;
        RECT 2001.065 2582.815 2001.395 2582.830 ;
        RECT 2004.505 2581.880 2004.805 2582.830 ;
        RECT 2007.965 2583.130 2008.295 2583.145 ;
        RECT 2013.005 2583.130 2013.305 2586.480 ;
        RECT 2007.965 2582.830 2013.305 2583.130 ;
        RECT 2007.965 2582.815 2008.295 2582.830 ;
        RECT 2013.005 2581.880 2013.305 2582.830 ;
        RECT 2016.705 2582.450 2017.035 2582.465 ;
        RECT 2018.645 2582.450 2018.945 2586.480 ;
        RECT 2016.705 2582.150 2018.945 2582.450 ;
        RECT 2016.705 2582.135 2017.035 2582.150 ;
        RECT 2018.645 2581.880 2018.945 2582.150 ;
        RECT 2021.765 2582.450 2022.095 2582.465 ;
        RECT 2027.145 2582.450 2027.445 2586.480 ;
        RECT 2021.765 2582.150 2027.445 2582.450 ;
        RECT 2021.765 2582.135 2022.095 2582.150 ;
        RECT 2027.145 2581.880 2027.445 2582.150 ;
        RECT 2030.045 2582.450 2030.375 2582.465 ;
        RECT 2032.785 2582.450 2033.085 2586.480 ;
        RECT 2030.045 2582.150 2033.085 2582.450 ;
        RECT 2030.045 2582.135 2030.375 2582.150 ;
        RECT 2032.785 2581.880 2033.085 2582.150 ;
      LAYER met3 ;
        RECT 357.355 2575.440 1355.530 2576.840 ;
      LAYER met3 ;
        RECT 1355.930 2576.330 1359.930 2576.440 ;
        RECT 1368.105 2576.330 1368.435 2576.345 ;
        RECT 1355.930 2576.030 1368.435 2576.330 ;
        RECT 1355.930 2575.840 1359.930 2576.030 ;
        RECT 1368.105 2576.015 1368.435 2576.030 ;
      LAYER met3 ;
        RECT 357.355 2567.320 1355.930 2575.440 ;
        RECT 357.355 2565.920 1355.530 2567.320 ;
      LAYER met3 ;
        RECT 1355.930 2566.810 1359.930 2566.920 ;
        RECT 1370.865 2566.810 1371.195 2566.825 ;
        RECT 1355.930 2566.510 1371.195 2566.810 ;
        RECT 1355.930 2566.320 1359.930 2566.510 ;
        RECT 1370.865 2566.495 1371.195 2566.510 ;
      LAYER met3 ;
        RECT 357.355 2557.800 1355.930 2565.920 ;
      LAYER met3 ;
        RECT 1600.865 2560.700 1601.195 2560.705 ;
        RECT 1600.865 2560.690 1601.450 2560.700 ;
        RECT 1600.640 2560.390 1601.450 2560.690 ;
        RECT 1600.865 2560.380 1601.450 2560.390 ;
        RECT 1600.865 2560.375 1601.195 2560.380 ;
      LAYER met3 ;
        RECT 357.355 2556.400 1355.530 2557.800 ;
      LAYER met3 ;
        RECT 1355.930 2557.290 1359.930 2557.400 ;
        RECT 1367.645 2557.290 1367.975 2557.305 ;
        RECT 1355.930 2556.990 1367.975 2557.290 ;
        RECT 1355.930 2556.800 1359.930 2556.990 ;
        RECT 1367.645 2556.975 1367.975 2556.990 ;
      LAYER met3 ;
        RECT 357.355 2548.280 1355.930 2556.400 ;
        RECT 357.355 2546.880 1355.530 2548.280 ;
      LAYER met3 ;
        RECT 1355.930 2547.770 1359.930 2547.880 ;
        RECT 1371.325 2547.770 1371.655 2547.785 ;
        RECT 1355.930 2547.470 1371.655 2547.770 ;
        RECT 1355.930 2547.280 1359.930 2547.470 ;
        RECT 1371.325 2547.455 1371.655 2547.470 ;
      LAYER met3 ;
        RECT 357.355 2538.760 1355.930 2546.880 ;
      LAYER met3 ;
        RECT 1583.385 2545.730 1583.715 2545.745 ;
        RECT 1600.150 2545.730 1600.530 2545.740 ;
        RECT 1583.385 2545.430 1600.530 2545.730 ;
        RECT 1583.385 2545.415 1583.715 2545.430 ;
        RECT 1600.150 2545.420 1600.530 2545.430 ;
        RECT 1597.185 2539.610 1597.515 2539.625 ;
        RECT 1600.150 2539.610 1600.530 2539.620 ;
        RECT 1597.185 2539.310 1600.530 2539.610 ;
        RECT 1597.185 2539.295 1597.515 2539.310 ;
        RECT 1600.150 2539.300 1600.530 2539.310 ;
      LAYER met3 ;
        RECT 357.355 2537.360 1355.530 2538.760 ;
      LAYER met3 ;
        RECT 1355.930 2538.250 1359.930 2538.360 ;
        RECT 1368.565 2538.250 1368.895 2538.265 ;
        RECT 1355.930 2537.950 1368.895 2538.250 ;
        RECT 1355.930 2537.760 1359.930 2537.950 ;
        RECT 1368.565 2537.935 1368.895 2537.950 ;
        RECT 1601.785 2537.580 1602.115 2537.585 ;
        RECT 1601.785 2537.570 1602.370 2537.580 ;
      LAYER met3 ;
        RECT 357.355 2529.240 1355.930 2537.360 ;
      LAYER met3 ;
        RECT 1601.560 2537.270 1602.370 2537.570 ;
        RECT 1601.785 2537.260 1602.370 2537.270 ;
        RECT 1601.785 2537.255 1602.115 2537.260 ;
        RECT 1599.025 2531.460 1599.355 2531.465 ;
        RECT 1600.865 2531.460 1601.195 2531.465 ;
        RECT 1599.025 2531.450 1599.610 2531.460 ;
        RECT 1600.865 2531.450 1601.450 2531.460 ;
        RECT 1598.800 2531.150 1599.610 2531.450 ;
        RECT 1600.640 2531.150 1601.450 2531.450 ;
        RECT 1599.025 2531.140 1599.610 2531.150 ;
        RECT 1600.865 2531.140 1601.450 2531.150 ;
        RECT 1599.025 2531.135 1599.355 2531.140 ;
        RECT 1600.865 2531.135 1601.195 2531.140 ;
      LAYER met3 ;
        RECT 357.355 2527.840 1355.530 2529.240 ;
      LAYER met3 ;
        RECT 1355.930 2528.730 1359.930 2528.840 ;
        RECT 1367.645 2528.730 1367.975 2528.745 ;
        RECT 1355.930 2528.430 1367.975 2528.730 ;
        RECT 1355.930 2528.240 1359.930 2528.430 ;
        RECT 1367.645 2528.415 1367.975 2528.430 ;
      LAYER met3 ;
        RECT 357.355 2519.720 1355.930 2527.840 ;
      LAYER met3 ;
        RECT 1603.625 2523.980 1603.955 2523.985 ;
        RECT 1603.625 2523.970 1604.210 2523.980 ;
        RECT 1603.400 2523.670 1604.210 2523.970 ;
        RECT 1603.625 2523.660 1604.210 2523.670 ;
        RECT 1603.625 2523.655 1603.955 2523.660 ;
      LAYER met3 ;
        RECT 357.355 2518.320 1355.530 2519.720 ;
      LAYER met3 ;
        RECT 1355.930 2519.210 1359.930 2519.320 ;
        RECT 1367.645 2519.210 1367.975 2519.225 ;
        RECT 1355.930 2518.910 1367.975 2519.210 ;
        RECT 1355.930 2518.720 1359.930 2518.910 ;
        RECT 1367.645 2518.895 1367.975 2518.910 ;
        RECT 1383.030 2519.210 1383.410 2519.220 ;
        RECT 1599.230 2519.210 1599.610 2519.220 ;
        RECT 1383.030 2518.910 1599.610 2519.210 ;
        RECT 1383.030 2518.900 1383.410 2518.910 ;
        RECT 1599.230 2518.900 1599.610 2518.910 ;
        RECT 1602.705 2518.540 1603.035 2518.545 ;
        RECT 1602.705 2518.530 1603.290 2518.540 ;
      LAYER met3 ;
        RECT 357.355 2510.200 1355.930 2518.320 ;
      LAYER met3 ;
        RECT 1602.480 2518.230 1603.290 2518.530 ;
        RECT 1602.705 2518.220 1603.290 2518.230 ;
        RECT 1602.705 2518.215 1603.035 2518.220 ;
        RECT 1600.865 2515.820 1601.195 2515.825 ;
        RECT 1600.865 2515.810 1601.450 2515.820 ;
        RECT 1600.640 2515.510 1601.450 2515.810 ;
        RECT 1600.865 2515.500 1601.450 2515.510 ;
        RECT 1600.865 2515.495 1601.195 2515.500 ;
        RECT 1601.785 2512.420 1602.115 2512.425 ;
        RECT 1601.785 2512.410 1602.370 2512.420 ;
        RECT 1601.560 2512.110 1602.370 2512.410 ;
        RECT 1601.785 2512.100 1602.370 2512.110 ;
        RECT 1601.785 2512.095 1602.115 2512.100 ;
      LAYER met3 ;
        RECT 357.355 2508.800 1355.530 2510.200 ;
      LAYER met3 ;
        RECT 1355.930 2509.690 1359.930 2509.800 ;
        RECT 1368.105 2509.690 1368.435 2509.705 ;
        RECT 1355.930 2509.390 1368.435 2509.690 ;
        RECT 1355.930 2509.200 1359.930 2509.390 ;
        RECT 1368.105 2509.375 1368.435 2509.390 ;
      LAYER met3 ;
        RECT 357.355 2500.680 1355.930 2508.800 ;
      LAYER met3 ;
        RECT 1604.085 2506.980 1604.415 2506.985 ;
        RECT 1603.830 2506.970 1604.415 2506.980 ;
        RECT 1603.830 2506.670 1604.640 2506.970 ;
        RECT 1603.830 2506.660 1604.415 2506.670 ;
        RECT 1604.085 2506.655 1604.415 2506.660 ;
        RECT 1599.025 2504.940 1599.355 2504.945 ;
        RECT 1599.025 2504.930 1599.610 2504.940 ;
        RECT 1598.800 2504.630 1599.610 2504.930 ;
        RECT 1599.025 2504.620 1599.610 2504.630 ;
        RECT 1599.025 2504.615 1599.355 2504.620 ;
        RECT 1599.945 2504.260 1600.275 2504.265 ;
        RECT 1599.945 2504.250 1600.530 2504.260 ;
        RECT 1599.720 2503.950 1600.530 2504.250 ;
        RECT 1599.945 2503.940 1600.530 2503.950 ;
        RECT 1599.945 2503.935 1600.275 2503.940 ;
        RECT 1603.165 2500.860 1603.495 2500.865 ;
        RECT 1602.910 2500.850 1603.495 2500.860 ;
      LAYER met3 ;
        RECT 357.355 2499.280 1355.530 2500.680 ;
      LAYER met3 ;
        RECT 1602.910 2500.550 1603.720 2500.850 ;
        RECT 1602.910 2500.540 1603.495 2500.550 ;
        RECT 1603.165 2500.535 1603.495 2500.540 ;
        RECT 1355.930 2500.170 1359.930 2500.280 ;
        RECT 1368.565 2500.170 1368.895 2500.185 ;
        RECT 1355.930 2499.870 1368.895 2500.170 ;
        RECT 1355.930 2499.680 1359.930 2499.870 ;
        RECT 1368.565 2499.855 1368.895 2499.870 ;
      LAYER met3 ;
        RECT 357.355 2491.160 1355.930 2499.280 ;
      LAYER met3 ;
        RECT 1601.325 2498.140 1601.655 2498.145 ;
        RECT 1601.070 2498.130 1601.655 2498.140 ;
        RECT 1601.070 2497.830 1601.880 2498.130 ;
        RECT 1601.070 2497.820 1601.655 2497.830 ;
        RECT 1601.325 2497.815 1601.655 2497.820 ;
        RECT 1603.625 2494.740 1603.955 2494.745 ;
        RECT 1603.625 2494.730 1604.210 2494.740 ;
        RECT 1603.400 2494.430 1604.210 2494.730 ;
        RECT 1603.625 2494.420 1604.210 2494.430 ;
        RECT 1603.625 2494.415 1603.955 2494.420 ;
      LAYER met3 ;
        RECT 357.355 2489.760 1355.530 2491.160 ;
      LAYER met3 ;
        RECT 1355.930 2490.650 1359.930 2490.760 ;
        RECT 1368.565 2490.650 1368.895 2490.665 ;
        RECT 1355.930 2490.350 1368.895 2490.650 ;
        RECT 1355.930 2490.160 1359.930 2490.350 ;
        RECT 1368.565 2490.335 1368.895 2490.350 ;
        RECT 1599.025 2489.980 1599.355 2489.985 ;
        RECT 1599.025 2489.970 1599.610 2489.980 ;
      LAYER met3 ;
        RECT 357.355 2481.640 1355.930 2489.760 ;
      LAYER met3 ;
        RECT 1598.800 2489.670 1599.610 2489.970 ;
        RECT 1599.025 2489.660 1599.610 2489.670 ;
        RECT 1599.025 2489.655 1599.355 2489.660 ;
        RECT 1601.325 2489.300 1601.655 2489.305 ;
        RECT 1601.070 2489.290 1601.655 2489.300 ;
        RECT 1601.070 2488.990 1601.880 2489.290 ;
        RECT 1601.070 2488.980 1601.655 2488.990 ;
        RECT 1601.325 2488.975 1601.655 2488.980 ;
        RECT 1600.865 2486.580 1601.195 2486.585 ;
        RECT 1600.865 2486.570 1601.450 2486.580 ;
        RECT 1600.640 2486.270 1601.450 2486.570 ;
        RECT 1600.865 2486.260 1601.450 2486.270 ;
        RECT 1600.865 2486.255 1601.195 2486.260 ;
        RECT 1602.245 2483.180 1602.575 2483.185 ;
        RECT 1601.990 2483.170 1602.575 2483.180 ;
        RECT 1601.990 2482.870 1602.800 2483.170 ;
        RECT 1601.990 2482.860 1602.575 2482.870 ;
        RECT 1602.245 2482.855 1602.575 2482.860 ;
      LAYER met3 ;
        RECT 357.355 2480.240 1355.530 2481.640 ;
      LAYER met3 ;
        RECT 1355.930 2481.130 1359.930 2481.240 ;
        RECT 1368.565 2481.130 1368.895 2481.145 ;
        RECT 1355.930 2480.830 1368.895 2481.130 ;
        RECT 1355.930 2480.640 1359.930 2480.830 ;
        RECT 1368.565 2480.815 1368.895 2480.830 ;
      LAYER met3 ;
        RECT 357.355 2472.120 1355.930 2480.240 ;
      LAYER met3 ;
        RECT 1604.085 2477.740 1604.415 2477.745 ;
        RECT 1603.830 2477.730 1604.415 2477.740 ;
        RECT 1603.630 2477.430 1604.415 2477.730 ;
        RECT 1603.830 2477.420 1604.415 2477.430 ;
        RECT 1604.085 2477.415 1604.415 2477.420 ;
        RECT 1599.025 2476.380 1599.355 2476.385 ;
        RECT 1599.025 2476.370 1599.610 2476.380 ;
        RECT 1598.800 2476.070 1599.610 2476.370 ;
        RECT 1599.025 2476.060 1599.610 2476.070 ;
        RECT 1599.025 2476.055 1599.355 2476.060 ;
        RECT 1600.865 2475.020 1601.195 2475.025 ;
        RECT 1600.865 2475.010 1601.450 2475.020 ;
        RECT 1600.640 2474.710 1601.450 2475.010 ;
        RECT 1600.865 2474.700 1601.450 2474.710 ;
        RECT 1600.865 2474.695 1601.195 2474.700 ;
        RECT 1602.705 2472.980 1603.035 2472.985 ;
        RECT 1602.705 2472.970 1603.290 2472.980 ;
        RECT 1602.705 2472.670 1603.490 2472.970 ;
        RECT 1602.705 2472.660 1603.290 2472.670 ;
        RECT 1602.705 2472.655 1603.035 2472.660 ;
      LAYER met3 ;
        RECT 357.355 2470.720 1355.530 2472.120 ;
      LAYER met3 ;
        RECT 1355.930 2471.610 1359.930 2471.720 ;
        RECT 1368.105 2471.610 1368.435 2471.625 ;
        RECT 1355.930 2471.310 1368.435 2471.610 ;
        RECT 1355.930 2471.120 1359.930 2471.310 ;
        RECT 1368.105 2471.295 1368.435 2471.310 ;
      LAYER met3 ;
        RECT 357.355 2462.600 1355.930 2470.720 ;
      LAYER met3 ;
        RECT 1599.025 2468.900 1599.355 2468.905 ;
        RECT 1599.025 2468.890 1599.610 2468.900 ;
        RECT 1598.800 2468.590 1599.610 2468.890 ;
        RECT 1599.025 2468.580 1599.610 2468.590 ;
        RECT 1599.025 2468.575 1599.355 2468.580 ;
        RECT 1601.785 2467.540 1602.115 2467.545 ;
        RECT 1601.785 2467.530 1602.370 2467.540 ;
        RECT 1601.785 2467.230 1602.570 2467.530 ;
        RECT 1601.785 2467.220 1602.370 2467.230 ;
        RECT 1601.785 2467.215 1602.115 2467.220 ;
        RECT 1599.945 2463.460 1600.275 2463.465 ;
        RECT 1599.945 2463.450 1600.530 2463.460 ;
        RECT 1599.720 2463.150 1600.530 2463.450 ;
        RECT 1599.945 2463.140 1600.530 2463.150 ;
        RECT 1599.945 2463.135 1600.275 2463.140 ;
      LAYER met3 ;
        RECT 357.355 2461.200 1355.530 2462.600 ;
      LAYER met3 ;
        RECT 1355.930 2462.090 1359.930 2462.200 ;
        RECT 1368.105 2462.090 1368.435 2462.105 ;
        RECT 1355.930 2461.790 1368.435 2462.090 ;
        RECT 1355.930 2461.600 1359.930 2461.790 ;
        RECT 1368.105 2461.775 1368.435 2461.790 ;
        RECT 1603.165 2461.420 1603.495 2461.425 ;
        RECT 1602.910 2461.410 1603.495 2461.420 ;
      LAYER met3 ;
        RECT 357.355 2453.080 1355.930 2461.200 ;
      LAYER met3 ;
        RECT 1602.710 2461.110 1603.495 2461.410 ;
        RECT 1602.910 2461.100 1603.495 2461.110 ;
        RECT 1603.165 2461.095 1603.495 2461.100 ;
        RECT 1599.025 2455.980 1599.355 2455.985 ;
        RECT 1599.025 2455.970 1599.610 2455.980 ;
        RECT 1598.800 2455.670 1599.610 2455.970 ;
        RECT 1599.025 2455.660 1599.610 2455.670 ;
        RECT 1599.025 2455.655 1599.355 2455.660 ;
        RECT 1603.165 2454.620 1603.495 2454.625 ;
        RECT 1602.910 2454.610 1603.495 2454.620 ;
        RECT 1602.710 2454.310 1603.495 2454.610 ;
        RECT 1602.910 2454.300 1603.495 2454.310 ;
        RECT 1603.165 2454.295 1603.495 2454.300 ;
      LAYER met3 ;
        RECT 357.355 2451.680 1355.530 2453.080 ;
      LAYER met3 ;
        RECT 1355.930 2452.570 1359.930 2452.680 ;
        RECT 1367.185 2452.570 1367.515 2452.585 ;
        RECT 1355.930 2452.270 1367.515 2452.570 ;
        RECT 1355.930 2452.080 1359.930 2452.270 ;
        RECT 1367.185 2452.255 1367.515 2452.270 ;
        RECT 1600.865 2451.900 1601.195 2451.905 ;
        RECT 1600.865 2451.890 1601.450 2451.900 ;
      LAYER met3 ;
        RECT 357.355 2443.560 1355.930 2451.680 ;
      LAYER met3 ;
        RECT 1600.640 2451.590 1601.450 2451.890 ;
        RECT 1600.865 2451.580 1601.450 2451.590 ;
        RECT 1600.865 2451.575 1601.195 2451.580 ;
        RECT 1600.405 2449.170 1600.735 2449.185 ;
        RECT 1601.070 2449.170 1601.450 2449.180 ;
        RECT 1600.405 2448.870 1601.450 2449.170 ;
        RECT 1600.405 2448.855 1600.735 2448.870 ;
        RECT 1601.070 2448.860 1601.450 2448.870 ;
      LAYER met3 ;
        RECT 357.355 2442.160 1355.530 2443.560 ;
      LAYER met3 ;
        RECT 1355.930 2443.050 1359.930 2443.160 ;
        RECT 1368.105 2443.050 1368.435 2443.065 ;
        RECT 1355.930 2442.750 1368.435 2443.050 ;
        RECT 1355.930 2442.560 1359.930 2442.750 ;
        RECT 1368.105 2442.735 1368.435 2442.750 ;
        RECT 1601.325 2442.370 1601.655 2442.385 ;
        RECT 1603.625 2442.380 1603.955 2442.385 ;
        RECT 1603.625 2442.370 1604.210 2442.380 ;
      LAYER met3 ;
        RECT 357.355 2434.040 1355.930 2442.160 ;
      LAYER met3 ;
        RECT 1601.325 2442.070 1604.410 2442.370 ;
        RECT 1601.325 2442.055 1601.655 2442.070 ;
        RECT 1603.625 2442.060 1604.210 2442.070 ;
        RECT 1603.625 2442.055 1603.955 2442.060 ;
        RECT 1599.025 2439.660 1599.355 2439.665 ;
        RECT 1600.865 2439.660 1601.195 2439.665 ;
        RECT 1599.025 2439.650 1599.610 2439.660 ;
        RECT 1600.865 2439.650 1601.450 2439.660 ;
        RECT 1598.800 2439.350 1599.610 2439.650 ;
        RECT 1600.640 2439.350 1601.450 2439.650 ;
        RECT 1599.025 2439.340 1599.610 2439.350 ;
        RECT 1600.865 2439.340 1601.450 2439.350 ;
        RECT 1599.025 2439.335 1599.355 2439.340 ;
        RECT 1600.865 2439.335 1601.195 2439.340 ;
        RECT 1601.325 2436.940 1601.655 2436.945 ;
        RECT 1601.070 2436.930 1601.655 2436.940 ;
        RECT 1602.245 2436.930 1602.575 2436.945 ;
        RECT 1600.870 2436.630 1602.575 2436.930 ;
        RECT 1601.070 2436.620 1601.655 2436.630 ;
        RECT 1601.325 2436.615 1601.655 2436.620 ;
        RECT 1602.245 2436.615 1602.575 2436.630 ;
      LAYER met3 ;
        RECT 357.355 2432.640 1355.530 2434.040 ;
      LAYER met3 ;
        RECT 1355.930 2433.530 1359.930 2433.640 ;
        RECT 1367.645 2433.530 1367.975 2433.545 ;
        RECT 1355.930 2433.230 1367.975 2433.530 ;
        RECT 1355.930 2433.040 1359.930 2433.230 ;
        RECT 1367.645 2433.215 1367.975 2433.230 ;
        RECT 1598.565 2433.530 1598.895 2433.545 ;
        RECT 1599.230 2433.530 1599.610 2433.540 ;
        RECT 1598.565 2433.230 1599.610 2433.530 ;
        RECT 1598.565 2433.215 1598.895 2433.230 ;
        RECT 1599.230 2433.220 1599.610 2433.230 ;
      LAYER met3 ;
        RECT 357.355 2424.520 1355.930 2432.640 ;
      LAYER met3 ;
        RECT 1602.245 2430.820 1602.575 2430.825 ;
        RECT 1601.990 2430.810 1602.575 2430.820 ;
        RECT 1601.790 2430.510 1602.575 2430.810 ;
        RECT 1601.990 2430.500 1602.575 2430.510 ;
        RECT 1602.245 2430.495 1602.575 2430.500 ;
        RECT 1599.025 2428.100 1599.355 2428.105 ;
        RECT 1599.025 2428.090 1599.610 2428.100 ;
        RECT 1598.800 2427.790 1599.610 2428.090 ;
        RECT 1599.025 2427.780 1599.610 2427.790 ;
        RECT 1599.025 2427.775 1599.355 2427.780 ;
        RECT 1602.705 2424.700 1603.035 2424.705 ;
        RECT 1602.705 2424.690 1603.290 2424.700 ;
      LAYER met3 ;
        RECT 357.355 2423.120 1355.530 2424.520 ;
      LAYER met3 ;
        RECT 1602.705 2424.390 1603.490 2424.690 ;
        RECT 1602.705 2424.380 1603.290 2424.390 ;
        RECT 1602.705 2424.375 1603.035 2424.380 ;
        RECT 1355.930 2424.010 1359.930 2424.120 ;
        RECT 1368.105 2424.010 1368.435 2424.025 ;
        RECT 1355.930 2423.710 1368.435 2424.010 ;
        RECT 1355.930 2423.520 1359.930 2423.710 ;
        RECT 1368.105 2423.695 1368.435 2423.710 ;
      LAYER met3 ;
        RECT 357.355 2415.000 1355.930 2423.120 ;
      LAYER met3 ;
        RECT 1600.865 2422.660 1601.195 2422.665 ;
        RECT 1600.865 2422.650 1601.450 2422.660 ;
        RECT 1600.640 2422.350 1601.450 2422.650 ;
        RECT 1600.865 2422.340 1601.450 2422.350 ;
        RECT 1600.865 2422.335 1601.195 2422.340 ;
        RECT 1601.785 2420.620 1602.115 2420.625 ;
        RECT 1601.785 2420.610 1602.370 2420.620 ;
        RECT 1601.785 2420.310 1602.570 2420.610 ;
        RECT 1601.785 2420.300 1602.370 2420.310 ;
        RECT 1601.785 2420.295 1602.115 2420.300 ;
        RECT 1599.025 2415.180 1599.355 2415.185 ;
        RECT 1599.025 2415.170 1599.610 2415.180 ;
      LAYER met3 ;
        RECT 357.355 2413.600 1355.530 2415.000 ;
      LAYER met3 ;
        RECT 1598.800 2414.870 1599.610 2415.170 ;
        RECT 1599.025 2414.860 1599.610 2414.870 ;
        RECT 1599.025 2414.855 1599.355 2414.860 ;
        RECT 1355.930 2414.490 1359.930 2414.600 ;
        RECT 1368.105 2414.490 1368.435 2414.505 ;
        RECT 1355.930 2414.190 1368.435 2414.490 ;
        RECT 1355.930 2414.000 1359.930 2414.190 ;
        RECT 1368.105 2414.175 1368.435 2414.190 ;
        RECT 1603.625 2413.810 1603.955 2413.825 ;
      LAYER met3 ;
        RECT 357.355 2405.480 1355.930 2413.600 ;
      LAYER met3 ;
        RECT 1603.625 2413.495 1604.170 2413.810 ;
        RECT 1603.165 2413.140 1603.495 2413.145 ;
        RECT 1602.910 2413.130 1603.495 2413.140 ;
        RECT 1602.710 2412.830 1603.495 2413.130 ;
        RECT 1602.910 2412.820 1603.495 2412.830 ;
        RECT 1603.165 2412.815 1603.495 2412.820 ;
        RECT 1603.165 2411.770 1603.495 2411.785 ;
        RECT 1603.870 2411.770 1604.170 2413.495 ;
        RECT 1603.165 2411.470 1604.170 2411.770 ;
        RECT 1603.165 2411.455 1603.495 2411.470 ;
        RECT 1600.865 2410.420 1601.195 2410.425 ;
        RECT 1600.865 2410.410 1601.450 2410.420 ;
        RECT 1600.640 2410.110 1601.450 2410.410 ;
        RECT 1600.865 2410.100 1601.450 2410.110 ;
        RECT 1600.865 2410.095 1601.195 2410.100 ;
        RECT 1602.245 2407.700 1602.575 2407.705 ;
        RECT 1601.990 2407.690 1602.575 2407.700 ;
        RECT 1601.790 2407.390 1602.575 2407.690 ;
        RECT 1601.990 2407.380 1602.575 2407.390 ;
        RECT 1602.245 2407.375 1602.575 2407.380 ;
      LAYER met3 ;
        RECT 357.355 2404.080 1355.530 2405.480 ;
      LAYER met3 ;
        RECT 1355.930 2404.970 1359.930 2405.080 ;
        RECT 1368.105 2404.970 1368.435 2404.985 ;
        RECT 1355.930 2404.670 1368.435 2404.970 ;
        RECT 1355.930 2404.480 1359.930 2404.670 ;
        RECT 1368.105 2404.655 1368.435 2404.670 ;
      LAYER met3 ;
        RECT 357.355 2395.960 1355.930 2404.080 ;
      LAYER met3 ;
        RECT 1602.705 2401.580 1603.035 2401.585 ;
        RECT 1602.705 2401.570 1603.290 2401.580 ;
        RECT 1602.705 2401.270 1603.490 2401.570 ;
        RECT 1602.705 2401.260 1603.290 2401.270 ;
        RECT 1602.705 2401.255 1603.035 2401.260 ;
        RECT 1599.025 2398.860 1599.355 2398.865 ;
        RECT 1600.865 2398.860 1601.195 2398.865 ;
        RECT 1599.025 2398.850 1599.610 2398.860 ;
        RECT 1600.865 2398.850 1601.450 2398.860 ;
        RECT 1598.800 2398.550 1599.610 2398.850 ;
        RECT 1600.640 2398.550 1601.450 2398.850 ;
        RECT 1599.025 2398.540 1599.610 2398.550 ;
        RECT 1600.865 2398.540 1601.450 2398.550 ;
        RECT 1599.025 2398.535 1599.355 2398.540 ;
        RECT 1600.865 2398.535 1601.195 2398.540 ;
      LAYER met3 ;
        RECT 357.355 2394.560 1355.530 2395.960 ;
      LAYER met3 ;
        RECT 1355.930 2395.450 1359.930 2395.560 ;
        RECT 1368.105 2395.450 1368.435 2395.465 ;
        RECT 1603.165 2395.460 1603.495 2395.465 ;
        RECT 1602.910 2395.450 1603.495 2395.460 ;
        RECT 1355.930 2395.150 1368.435 2395.450 ;
        RECT 1602.710 2395.150 1603.495 2395.450 ;
        RECT 1355.930 2394.960 1359.930 2395.150 ;
        RECT 1368.105 2395.135 1368.435 2395.150 ;
        RECT 1602.910 2395.140 1603.495 2395.150 ;
        RECT 1603.165 2395.135 1603.495 2395.140 ;
      LAYER met3 ;
        RECT 357.355 2386.440 1355.930 2394.560 ;
      LAYER met3 ;
        RECT 1603.165 2390.020 1603.495 2390.025 ;
        RECT 1602.910 2390.010 1603.495 2390.020 ;
        RECT 1602.910 2389.710 1603.720 2390.010 ;
        RECT 1602.910 2389.700 1603.495 2389.710 ;
        RECT 1603.165 2389.695 1603.495 2389.700 ;
      LAYER met3 ;
        RECT 357.355 2385.040 1355.530 2386.440 ;
      LAYER met3 ;
        RECT 1355.930 2385.930 1359.930 2386.040 ;
        RECT 1368.105 2385.930 1368.435 2385.945 ;
        RECT 1355.930 2385.630 1368.435 2385.930 ;
        RECT 1355.930 2385.440 1359.930 2385.630 ;
        RECT 1368.105 2385.615 1368.435 2385.630 ;
      LAYER met3 ;
        RECT 357.355 2376.920 1355.930 2385.040 ;
      LAYER met3 ;
        RECT 1600.865 2383.900 1601.195 2383.905 ;
        RECT 1601.785 2383.900 1602.115 2383.905 ;
        RECT 1600.865 2383.890 1601.450 2383.900 ;
        RECT 1600.640 2383.590 1601.450 2383.890 ;
        RECT 1600.865 2383.580 1601.450 2383.590 ;
        RECT 1601.785 2383.890 1602.370 2383.900 ;
        RECT 1601.785 2383.590 1602.570 2383.890 ;
        RECT 1601.785 2383.580 1602.370 2383.590 ;
        RECT 1600.865 2383.575 1601.195 2383.580 ;
        RECT 1601.785 2383.575 1602.115 2383.580 ;
        RECT 1602.245 2379.810 1602.575 2379.825 ;
        RECT 1603.625 2379.810 1603.955 2379.825 ;
        RECT 1602.245 2379.510 1603.955 2379.810 ;
        RECT 1602.245 2379.495 1602.575 2379.510 ;
        RECT 1603.625 2379.495 1603.955 2379.510 ;
        RECT 1599.230 2379.130 1599.610 2379.140 ;
        RECT 1603.165 2379.130 1603.495 2379.145 ;
        RECT 1604.085 2379.140 1604.415 2379.145 ;
        RECT 1599.230 2378.830 1603.495 2379.130 ;
        RECT 1599.230 2378.820 1599.610 2378.830 ;
        RECT 1603.165 2378.815 1603.495 2378.830 ;
        RECT 1603.830 2379.130 1604.415 2379.140 ;
        RECT 1603.830 2378.830 1604.640 2379.130 ;
        RECT 1603.830 2378.820 1604.415 2378.830 ;
        RECT 1604.085 2378.815 1604.415 2378.820 ;
        RECT 1602.910 2378.450 1603.290 2378.460 ;
        RECT 1602.910 2378.150 1604.170 2378.450 ;
        RECT 1602.910 2378.140 1603.290 2378.150 ;
        RECT 1603.870 2377.785 1604.170 2378.150 ;
        RECT 1603.870 2377.470 1604.415 2377.785 ;
        RECT 1604.085 2377.455 1604.415 2377.470 ;
      LAYER met3 ;
        RECT 357.355 2375.520 1355.530 2376.920 ;
      LAYER met3 ;
        RECT 1355.930 2376.410 1359.930 2376.520 ;
        RECT 1368.105 2376.410 1368.435 2376.425 ;
        RECT 1355.930 2376.110 1368.435 2376.410 ;
        RECT 1355.930 2375.920 1359.930 2376.110 ;
        RECT 1368.105 2376.095 1368.435 2376.110 ;
      LAYER met3 ;
        RECT 357.355 2367.400 1355.930 2375.520 ;
      LAYER met3 ;
        RECT 1600.865 2372.340 1601.195 2372.345 ;
        RECT 1603.625 2372.340 1603.955 2372.345 ;
        RECT 1600.865 2372.330 1601.450 2372.340 ;
        RECT 1600.640 2372.030 1601.450 2372.330 ;
        RECT 1600.865 2372.020 1601.450 2372.030 ;
        RECT 1603.625 2372.330 1604.210 2372.340 ;
        RECT 1603.625 2372.030 1604.410 2372.330 ;
        RECT 1603.625 2372.020 1604.210 2372.030 ;
        RECT 1600.865 2372.015 1601.195 2372.020 ;
        RECT 1603.625 2372.015 1603.955 2372.020 ;
      LAYER met3 ;
        RECT 357.355 2366.000 1355.530 2367.400 ;
      LAYER met3 ;
        RECT 1355.930 2366.890 1359.930 2367.000 ;
        RECT 1368.105 2366.890 1368.435 2366.905 ;
        RECT 1355.930 2366.590 1368.435 2366.890 ;
        RECT 1355.930 2366.400 1359.930 2366.590 ;
        RECT 1368.105 2366.575 1368.435 2366.590 ;
        RECT 1601.325 2366.890 1601.655 2366.905 ;
        RECT 1601.325 2366.590 1603.250 2366.890 ;
        RECT 1601.325 2366.575 1601.655 2366.590 ;
        RECT 1602.950 2366.225 1603.250 2366.590 ;
        RECT 1601.325 2366.220 1601.655 2366.225 ;
        RECT 1601.070 2366.210 1601.655 2366.220 ;
        RECT 1602.705 2366.220 1603.250 2366.225 ;
        RECT 1602.705 2366.210 1603.290 2366.220 ;
      LAYER met3 ;
        RECT 357.355 2357.880 1355.930 2366.000 ;
      LAYER met3 ;
        RECT 1601.070 2365.910 1601.880 2366.210 ;
        RECT 1602.705 2365.910 1603.490 2366.210 ;
        RECT 1601.070 2365.900 1601.655 2365.910 ;
        RECT 1601.325 2365.895 1601.655 2365.900 ;
        RECT 1602.705 2365.900 1603.290 2365.910 ;
        RECT 1602.705 2365.895 1603.035 2365.900 ;
        RECT 1601.070 2361.450 1601.450 2361.460 ;
        RECT 1601.785 2361.450 1602.115 2361.465 ;
        RECT 1601.070 2361.150 1602.115 2361.450 ;
        RECT 1601.070 2361.140 1601.450 2361.150 ;
        RECT 1601.785 2361.135 1602.115 2361.150 ;
        RECT 1601.785 2360.780 1602.115 2360.785 ;
        RECT 1601.785 2360.770 1602.370 2360.780 ;
        RECT 1601.560 2360.470 1602.370 2360.770 ;
        RECT 1601.785 2360.460 1602.370 2360.470 ;
        RECT 1601.785 2360.455 1602.115 2360.460 ;
      LAYER met3 ;
        RECT 357.355 2356.480 1355.530 2357.880 ;
      LAYER met3 ;
        RECT 1355.930 2357.370 1359.930 2357.480 ;
        RECT 1367.645 2357.370 1367.975 2357.385 ;
        RECT 1355.930 2357.070 1367.975 2357.370 ;
        RECT 1355.930 2356.880 1359.930 2357.070 ;
        RECT 1367.645 2357.055 1367.975 2357.070 ;
      LAYER met3 ;
        RECT 357.355 2348.360 1355.930 2356.480 ;
      LAYER met3 ;
        RECT 1600.865 2355.330 1601.195 2355.345 ;
        RECT 1602.245 2355.330 1602.575 2355.345 ;
        RECT 1602.910 2355.330 1603.290 2355.340 ;
        RECT 1600.865 2355.030 1603.290 2355.330 ;
        RECT 1600.865 2355.015 1601.195 2355.030 ;
        RECT 1602.245 2355.015 1602.575 2355.030 ;
        RECT 1602.910 2355.020 1603.290 2355.030 ;
        RECT 1602.245 2354.660 1602.575 2354.665 ;
        RECT 1601.990 2354.650 1602.575 2354.660 ;
        RECT 1601.990 2354.350 1602.800 2354.650 ;
        RECT 1601.990 2354.340 1602.575 2354.350 ;
        RECT 1602.245 2354.335 1602.575 2354.340 ;
        RECT 1601.325 2350.570 1601.655 2350.585 ;
        RECT 1601.990 2350.570 1602.370 2350.580 ;
        RECT 1601.325 2350.270 1602.370 2350.570 ;
        RECT 1601.325 2350.255 1601.655 2350.270 ;
        RECT 1601.990 2350.260 1602.370 2350.270 ;
        RECT 1601.325 2349.220 1601.655 2349.225 ;
        RECT 1601.070 2349.210 1601.655 2349.220 ;
        RECT 1601.070 2348.910 1601.880 2349.210 ;
        RECT 1601.070 2348.900 1601.655 2348.910 ;
        RECT 1601.325 2348.895 1601.655 2348.900 ;
      LAYER met3 ;
        RECT 357.355 2346.960 1355.530 2348.360 ;
      LAYER met3 ;
        RECT 1355.930 2347.850 1359.930 2347.960 ;
        RECT 1367.645 2347.850 1367.975 2347.865 ;
        RECT 1355.930 2347.550 1367.975 2347.850 ;
        RECT 1355.930 2347.360 1359.930 2347.550 ;
        RECT 1367.645 2347.535 1367.975 2347.550 ;
      LAYER met3 ;
        RECT 357.355 2338.840 1355.930 2346.960 ;
      LAYER met3 ;
        RECT 1599.230 2345.810 1599.610 2345.820 ;
        RECT 1601.785 2345.810 1602.115 2345.825 ;
        RECT 1599.230 2345.510 1602.115 2345.810 ;
        RECT 1599.230 2345.500 1599.610 2345.510 ;
        RECT 1601.785 2345.495 1602.115 2345.510 ;
        RECT 1603.165 2344.460 1603.495 2344.465 ;
        RECT 1602.910 2344.450 1603.495 2344.460 ;
        RECT 1602.710 2344.150 1603.495 2344.450 ;
        RECT 1602.910 2344.140 1603.495 2344.150 ;
        RECT 1603.165 2344.135 1603.495 2344.140 ;
        RECT 1600.865 2343.100 1601.195 2343.105 ;
        RECT 1600.865 2343.090 1601.450 2343.100 ;
        RECT 1600.640 2342.790 1601.450 2343.090 ;
        RECT 1600.865 2342.780 1601.450 2342.790 ;
        RECT 1600.865 2342.775 1601.195 2342.780 ;
      LAYER met3 ;
        RECT 357.355 2337.440 1355.530 2338.840 ;
      LAYER met3 ;
        RECT 1355.930 2338.330 1359.930 2338.440 ;
        RECT 1367.645 2338.330 1367.975 2338.345 ;
        RECT 1355.930 2338.030 1367.975 2338.330 ;
        RECT 1355.930 2337.840 1359.930 2338.030 ;
        RECT 1367.645 2338.015 1367.975 2338.030 ;
        RECT 1601.990 2338.330 1602.370 2338.340 ;
        RECT 1603.165 2338.330 1603.495 2338.345 ;
        RECT 1601.990 2338.030 1603.495 2338.330 ;
        RECT 1601.990 2338.020 1602.370 2338.030 ;
        RECT 1603.165 2338.015 1603.495 2338.030 ;
      LAYER met3 ;
        RECT 357.355 2329.320 1355.930 2337.440 ;
        RECT 357.355 2327.920 1355.530 2329.320 ;
      LAYER met3 ;
        RECT 1355.930 2328.810 1359.930 2328.920 ;
        RECT 1367.645 2328.810 1367.975 2328.825 ;
        RECT 1355.930 2328.510 1367.975 2328.810 ;
        RECT 1355.930 2328.320 1359.930 2328.510 ;
        RECT 1367.645 2328.495 1367.975 2328.510 ;
      LAYER met3 ;
        RECT 357.355 2319.800 1355.930 2327.920 ;
      LAYER met3 ;
        RECT 1600.865 2326.100 1601.195 2326.105 ;
        RECT 1600.865 2326.090 1601.450 2326.100 ;
        RECT 1600.640 2325.790 1601.450 2326.090 ;
        RECT 1600.865 2325.780 1601.450 2325.790 ;
        RECT 1601.990 2325.780 1602.370 2326.100 ;
        RECT 1600.865 2325.775 1601.195 2325.780 ;
        RECT 1600.865 2324.730 1601.195 2324.745 ;
        RECT 1602.030 2324.730 1602.330 2325.780 ;
        RECT 1600.865 2324.430 1602.330 2324.730 ;
        RECT 1600.865 2324.415 1601.195 2324.430 ;
      LAYER met3 ;
        RECT 357.355 2318.400 1355.530 2319.800 ;
      LAYER met3 ;
        RECT 1355.930 2319.290 1359.930 2319.400 ;
        RECT 1366.265 2319.290 1366.595 2319.305 ;
        RECT 1355.930 2318.990 1366.595 2319.290 ;
        RECT 1355.930 2318.800 1359.930 2318.990 ;
        RECT 1366.265 2318.975 1366.595 2318.990 ;
      LAYER met3 ;
        RECT 357.355 2310.280 1355.930 2318.400 ;
        RECT 357.355 2308.880 1355.530 2310.280 ;
      LAYER met3 ;
        RECT 1355.930 2309.770 1359.930 2309.880 ;
        RECT 1366.265 2309.770 1366.595 2309.785 ;
        RECT 1355.930 2309.470 1366.595 2309.770 ;
        RECT 1355.930 2309.280 1359.930 2309.470 ;
        RECT 1366.265 2309.455 1366.595 2309.470 ;
      LAYER met3 ;
        RECT 357.355 2300.760 1355.930 2308.880 ;
        RECT 357.355 2299.360 1355.530 2300.760 ;
      LAYER met3 ;
        RECT 1355.930 2300.250 1359.930 2300.360 ;
        RECT 1366.265 2300.250 1366.595 2300.265 ;
        RECT 1355.930 2299.950 1366.595 2300.250 ;
        RECT 1355.930 2299.760 1359.930 2299.950 ;
        RECT 1366.265 2299.935 1366.595 2299.950 ;
      LAYER met3 ;
        RECT 357.355 2291.240 1355.930 2299.360 ;
        RECT 357.355 2289.840 1355.530 2291.240 ;
      LAYER met3 ;
        RECT 1355.930 2290.730 1359.930 2290.840 ;
        RECT 1366.265 2290.730 1366.595 2290.745 ;
        RECT 1355.930 2290.430 1366.595 2290.730 ;
        RECT 1355.930 2290.240 1359.930 2290.430 ;
        RECT 1366.265 2290.415 1366.595 2290.430 ;
      LAYER met3 ;
        RECT 357.355 2281.720 1355.930 2289.840 ;
        RECT 357.355 2280.320 1355.530 2281.720 ;
      LAYER met3 ;
        RECT 1355.930 2281.210 1359.930 2281.320 ;
        RECT 1366.265 2281.210 1366.595 2281.225 ;
        RECT 1355.930 2280.910 1366.595 2281.210 ;
        RECT 1355.930 2280.720 1359.930 2280.910 ;
        RECT 1366.265 2280.895 1366.595 2280.910 ;
      LAYER met3 ;
        RECT 357.355 2272.200 1355.930 2280.320 ;
        RECT 357.355 2270.800 1355.530 2272.200 ;
      LAYER met3 ;
        RECT 1355.930 2271.690 1359.930 2271.800 ;
        RECT 1366.265 2271.690 1366.595 2271.705 ;
        RECT 1355.930 2271.390 1366.595 2271.690 ;
        RECT 1355.930 2271.200 1359.930 2271.390 ;
        RECT 1366.265 2271.375 1366.595 2271.390 ;
      LAYER met3 ;
        RECT 357.355 2262.680 1355.930 2270.800 ;
        RECT 357.355 2261.280 1355.530 2262.680 ;
      LAYER met3 ;
        RECT 1355.930 2262.170 1359.930 2262.280 ;
        RECT 1366.265 2262.170 1366.595 2262.185 ;
        RECT 1355.930 2261.870 1366.595 2262.170 ;
        RECT 1355.930 2261.680 1359.930 2261.870 ;
        RECT 1366.265 2261.855 1366.595 2261.870 ;
      LAYER met3 ;
        RECT 357.355 2253.160 1355.930 2261.280 ;
        RECT 357.355 2251.760 1355.530 2253.160 ;
      LAYER met3 ;
        RECT 1355.930 2252.650 1359.930 2252.760 ;
        RECT 1366.725 2252.650 1367.055 2252.665 ;
        RECT 1355.930 2252.350 1367.055 2252.650 ;
        RECT 1355.930 2252.160 1359.930 2252.350 ;
        RECT 1366.725 2252.335 1367.055 2252.350 ;
      LAYER met3 ;
        RECT 357.355 2243.640 1355.930 2251.760 ;
        RECT 357.355 2242.240 1355.530 2243.640 ;
      LAYER met3 ;
        RECT 1355.930 2243.130 1359.930 2243.240 ;
        RECT 1367.185 2243.130 1367.515 2243.145 ;
        RECT 1355.930 2242.830 1367.515 2243.130 ;
        RECT 1355.930 2242.640 1359.930 2242.830 ;
        RECT 1367.185 2242.815 1367.515 2242.830 ;
      LAYER met3 ;
        RECT 357.355 2234.120 1355.930 2242.240 ;
        RECT 357.355 2232.720 1355.530 2234.120 ;
      LAYER met3 ;
        RECT 1355.930 2233.610 1359.930 2233.720 ;
        RECT 1367.185 2233.610 1367.515 2233.625 ;
        RECT 1355.930 2233.310 1367.515 2233.610 ;
        RECT 1355.930 2233.120 1359.930 2233.310 ;
        RECT 1367.185 2233.295 1367.515 2233.310 ;
      LAYER met3 ;
        RECT 357.355 2224.600 1355.930 2232.720 ;
        RECT 357.355 2223.200 1355.530 2224.600 ;
      LAYER met3 ;
        RECT 1355.930 2224.090 1359.930 2224.200 ;
        RECT 1367.185 2224.090 1367.515 2224.105 ;
        RECT 1355.930 2223.790 1367.515 2224.090 ;
        RECT 1355.930 2223.600 1359.930 2223.790 ;
        RECT 1367.185 2223.775 1367.515 2223.790 ;
      LAYER met3 ;
        RECT 357.355 2215.080 1355.930 2223.200 ;
        RECT 357.355 2213.680 1355.530 2215.080 ;
      LAYER met3 ;
        RECT 1355.930 2214.570 1359.930 2214.680 ;
        RECT 1367.185 2214.570 1367.515 2214.585 ;
        RECT 1355.930 2214.270 1367.515 2214.570 ;
        RECT 1355.930 2214.080 1359.930 2214.270 ;
        RECT 1367.185 2214.255 1367.515 2214.270 ;
      LAYER met3 ;
        RECT 357.355 2205.560 1355.930 2213.680 ;
      LAYER met3 ;
        RECT 1602.245 2211.850 1602.575 2211.865 ;
        RECT 1603.625 2211.850 1603.955 2211.865 ;
        RECT 1602.245 2211.550 1603.955 2211.850 ;
        RECT 1602.245 2211.535 1602.575 2211.550 ;
        RECT 1603.625 2211.535 1603.955 2211.550 ;
      LAYER met3 ;
        RECT 357.355 2204.160 1355.530 2205.560 ;
      LAYER met3 ;
        RECT 1355.930 2205.050 1359.930 2205.160 ;
        RECT 1367.185 2205.050 1367.515 2205.065 ;
        RECT 1355.930 2204.750 1367.515 2205.050 ;
      LAYER met3 ;
        RECT 1605.000 2205.000 2051.235 2581.480 ;
      LAYER met3 ;
        RECT 2051.235 2225.460 2052.140 2227.200 ;
        RECT 2051.235 2205.000 2052.140 2205.440 ;
        RECT 1355.930 2204.560 1359.930 2204.750 ;
        RECT 1367.185 2204.735 1367.515 2204.750 ;
      LAYER met3 ;
        RECT 357.355 2196.040 1355.930 2204.160 ;
      LAYER met3 ;
        RECT 1704.490 2200.000 1704.790 2204.600 ;
        RECT 1710.130 2200.000 1710.430 2204.600 ;
        RECT 1718.630 2200.000 1718.930 2204.600 ;
        RECT 1724.270 2200.000 1724.570 2204.600 ;
        RECT 1732.770 2200.000 1733.070 2204.600 ;
        RECT 1738.410 2200.000 1738.710 2204.600 ;
        RECT 1746.910 2200.000 1747.210 2204.600 ;
        RECT 2043.600 2202.430 2044.660 2205.000 ;
        RECT 2048.265 2200.000 2048.565 2204.600 ;
        RECT 2050.400 2200.180 2052.140 2205.000 ;
      LAYER met3 ;
        RECT 357.355 2194.640 1355.530 2196.040 ;
      LAYER met3 ;
        RECT 1355.930 2195.530 1359.930 2195.640 ;
        RECT 1367.185 2195.530 1367.515 2195.545 ;
        RECT 1355.930 2195.230 1367.515 2195.530 ;
        RECT 1355.930 2195.040 1359.930 2195.230 ;
        RECT 1367.185 2195.215 1367.515 2195.230 ;
      LAYER met3 ;
        RECT 357.355 2186.520 1355.930 2194.640 ;
        RECT 357.355 2185.120 1355.530 2186.520 ;
      LAYER met3 ;
        RECT 1355.930 2186.010 1359.930 2186.120 ;
        RECT 1373.165 2186.010 1373.495 2186.025 ;
        RECT 1355.930 2185.710 1373.495 2186.010 ;
        RECT 1355.930 2185.520 1359.930 2185.710 ;
        RECT 1373.165 2185.695 1373.495 2185.710 ;
      LAYER met3 ;
        RECT 357.355 2177.000 1355.930 2185.120 ;
        RECT 357.355 2175.600 1355.530 2177.000 ;
      LAYER met3 ;
        RECT 1355.930 2176.490 1359.930 2176.600 ;
        RECT 1373.625 2176.490 1373.955 2176.505 ;
        RECT 1355.930 2176.190 1373.955 2176.490 ;
        RECT 1355.930 2176.000 1359.930 2176.190 ;
        RECT 1373.625 2176.175 1373.955 2176.190 ;
      LAYER met3 ;
        RECT 357.355 2167.480 1355.930 2175.600 ;
        RECT 357.355 2166.080 1355.530 2167.480 ;
      LAYER met3 ;
        RECT 1355.930 2166.970 1359.930 2167.080 ;
        RECT 1366.265 2166.970 1366.595 2166.985 ;
        RECT 1355.930 2166.670 1366.595 2166.970 ;
        RECT 1355.930 2166.480 1359.930 2166.670 ;
        RECT 1366.265 2166.655 1366.595 2166.670 ;
      LAYER met3 ;
        RECT 357.355 2157.960 1355.930 2166.080 ;
        RECT 357.355 2156.560 1355.530 2157.960 ;
      LAYER met3 ;
        RECT 1355.930 2157.450 1359.930 2157.560 ;
        RECT 1366.265 2157.450 1366.595 2157.465 ;
        RECT 1355.930 2157.150 1366.595 2157.450 ;
        RECT 1355.930 2156.960 1359.930 2157.150 ;
        RECT 1366.265 2157.135 1366.595 2157.150 ;
      LAYER met3 ;
        RECT 357.355 2148.440 1355.930 2156.560 ;
        RECT 357.355 2147.040 1355.530 2148.440 ;
      LAYER met3 ;
        RECT 1355.930 2147.930 1359.930 2148.040 ;
        RECT 1366.265 2147.930 1366.595 2147.945 ;
        RECT 1355.930 2147.630 1366.595 2147.930 ;
        RECT 1355.930 2147.440 1359.930 2147.630 ;
        RECT 1366.265 2147.615 1366.595 2147.630 ;
      LAYER met3 ;
        RECT 357.355 2138.920 1355.930 2147.040 ;
        RECT 357.355 2137.520 1355.530 2138.920 ;
      LAYER met3 ;
        RECT 1355.930 2138.410 1359.930 2138.520 ;
        RECT 1366.265 2138.410 1366.595 2138.425 ;
        RECT 1355.930 2138.110 1366.595 2138.410 ;
        RECT 1355.930 2137.920 1359.930 2138.110 ;
        RECT 1366.265 2138.095 1366.595 2138.110 ;
      LAYER met3 ;
        RECT 357.355 2129.400 1355.930 2137.520 ;
        RECT 357.355 2128.000 1355.530 2129.400 ;
      LAYER met3 ;
        RECT 1355.930 2128.890 1359.930 2129.000 ;
        RECT 1366.265 2128.890 1366.595 2128.905 ;
        RECT 1355.930 2128.590 1366.595 2128.890 ;
        RECT 1355.930 2128.400 1359.930 2128.590 ;
        RECT 1366.265 2128.575 1366.595 2128.590 ;
      LAYER met3 ;
        RECT 357.355 2119.880 1355.930 2128.000 ;
        RECT 357.355 2118.480 1355.530 2119.880 ;
      LAYER met3 ;
        RECT 1355.930 2119.370 1359.930 2119.480 ;
        RECT 1367.185 2119.370 1367.515 2119.385 ;
        RECT 1355.930 2119.070 1367.515 2119.370 ;
        RECT 1355.930 2118.880 1359.930 2119.070 ;
        RECT 1367.185 2119.055 1367.515 2119.070 ;
      LAYER met3 ;
        RECT 357.355 2110.360 1355.930 2118.480 ;
        RECT 357.355 2108.960 1355.530 2110.360 ;
      LAYER met3 ;
        RECT 1355.930 2109.850 1359.930 2109.960 ;
        RECT 1367.185 2109.850 1367.515 2109.865 ;
        RECT 1355.930 2109.550 1367.515 2109.850 ;
        RECT 1355.930 2109.360 1359.930 2109.550 ;
        RECT 1367.185 2109.535 1367.515 2109.550 ;
      LAYER met3 ;
        RECT 357.355 2100.840 1355.930 2108.960 ;
        RECT 357.355 2099.440 1355.530 2100.840 ;
      LAYER met3 ;
        RECT 1355.930 2100.330 1359.930 2100.440 ;
        RECT 1367.185 2100.330 1367.515 2100.345 ;
        RECT 1355.930 2100.030 1367.515 2100.330 ;
        RECT 1355.930 2099.840 1359.930 2100.030 ;
        RECT 1367.185 2100.015 1367.515 2100.030 ;
      LAYER met3 ;
        RECT 357.355 2091.320 1355.930 2099.440 ;
        RECT 357.355 2089.920 1355.530 2091.320 ;
      LAYER met3 ;
        RECT 1355.930 2090.810 1359.930 2090.920 ;
        RECT 1367.185 2090.810 1367.515 2090.825 ;
        RECT 1355.930 2090.510 1367.515 2090.810 ;
        RECT 1355.930 2090.320 1359.930 2090.510 ;
        RECT 1367.185 2090.495 1367.515 2090.510 ;
      LAYER met3 ;
        RECT 357.355 2081.800 1355.930 2089.920 ;
        RECT 357.355 2080.400 1355.530 2081.800 ;
      LAYER met3 ;
        RECT 1355.930 2081.290 1359.930 2081.400 ;
        RECT 1367.185 2081.290 1367.515 2081.305 ;
        RECT 1355.930 2080.990 1367.515 2081.290 ;
        RECT 1355.930 2080.800 1359.930 2080.990 ;
        RECT 1367.185 2080.975 1367.515 2080.990 ;
      LAYER met3 ;
        RECT 357.355 2072.280 1355.930 2080.400 ;
        RECT 357.355 2070.880 1355.530 2072.280 ;
      LAYER met3 ;
        RECT 1355.930 2071.770 1359.930 2071.880 ;
        RECT 1367.185 2071.770 1367.515 2071.785 ;
        RECT 1355.930 2071.470 1367.515 2071.770 ;
        RECT 1355.930 2071.280 1359.930 2071.470 ;
        RECT 1367.185 2071.455 1367.515 2071.470 ;
      LAYER met3 ;
        RECT 357.355 2062.760 1355.930 2070.880 ;
        RECT 357.355 2061.360 1355.530 2062.760 ;
      LAYER met3 ;
        RECT 1355.930 2062.250 1359.930 2062.360 ;
        RECT 1367.185 2062.250 1367.515 2062.265 ;
        RECT 1355.930 2061.950 1367.515 2062.250 ;
        RECT 1355.930 2061.760 1359.930 2061.950 ;
        RECT 1367.185 2061.935 1367.515 2061.950 ;
      LAYER met3 ;
        RECT 357.355 2053.240 1355.930 2061.360 ;
        RECT 357.355 2051.840 1355.530 2053.240 ;
      LAYER met3 ;
        RECT 1355.930 2052.730 1359.930 2052.840 ;
        RECT 1367.185 2052.730 1367.515 2052.745 ;
        RECT 1355.930 2052.430 1367.515 2052.730 ;
        RECT 1355.930 2052.240 1359.930 2052.430 ;
        RECT 1367.185 2052.415 1367.515 2052.430 ;
      LAYER met3 ;
        RECT 357.355 2043.720 1355.930 2051.840 ;
        RECT 357.355 2042.320 1355.530 2043.720 ;
      LAYER met3 ;
        RECT 1355.930 2043.210 1359.930 2043.320 ;
        RECT 1367.185 2043.210 1367.515 2043.225 ;
        RECT 1355.930 2042.910 1367.515 2043.210 ;
        RECT 1355.930 2042.720 1359.930 2042.910 ;
        RECT 1367.185 2042.895 1367.515 2042.910 ;
      LAYER met3 ;
        RECT 357.355 2034.200 1355.930 2042.320 ;
        RECT 357.355 2032.800 1355.530 2034.200 ;
      LAYER met3 ;
        RECT 1355.930 2033.690 1359.930 2033.800 ;
        RECT 1367.185 2033.690 1367.515 2033.705 ;
        RECT 1355.930 2033.390 1367.515 2033.690 ;
        RECT 1355.930 2033.200 1359.930 2033.390 ;
        RECT 1367.185 2033.375 1367.515 2033.390 ;
      LAYER met3 ;
        RECT 357.355 2024.680 1355.930 2032.800 ;
        RECT 357.355 2023.280 1355.530 2024.680 ;
      LAYER met3 ;
        RECT 1355.930 2024.170 1359.930 2024.280 ;
        RECT 1383.030 2024.170 1383.410 2024.180 ;
        RECT 1355.930 2023.870 1383.410 2024.170 ;
        RECT 1355.930 2023.680 1359.930 2023.870 ;
        RECT 1383.030 2023.860 1383.410 2023.870 ;
      LAYER met3 ;
        RECT 357.355 2015.160 1355.930 2023.280 ;
        RECT 357.355 2013.760 1355.530 2015.160 ;
      LAYER met3 ;
        RECT 1355.930 2014.650 1359.930 2014.760 ;
        RECT 1367.185 2014.650 1367.515 2014.665 ;
        RECT 1355.930 2014.350 1367.515 2014.650 ;
        RECT 1355.930 2014.160 1359.930 2014.350 ;
        RECT 1367.185 2014.335 1367.515 2014.350 ;
      LAYER met3 ;
        RECT 357.355 2005.640 1355.930 2013.760 ;
        RECT 357.355 2004.240 1355.530 2005.640 ;
      LAYER met3 ;
        RECT 1355.930 2005.130 1359.930 2005.240 ;
        RECT 1367.185 2005.130 1367.515 2005.145 ;
        RECT 1355.930 2004.830 1367.515 2005.130 ;
        RECT 1355.930 2004.640 1359.930 2004.830 ;
        RECT 1367.185 2004.815 1367.515 2004.830 ;
      LAYER met3 ;
        RECT 357.355 1996.120 1355.930 2004.240 ;
        RECT 357.355 1994.720 1355.530 1996.120 ;
      LAYER met3 ;
        RECT 1355.930 1995.610 1359.930 1995.720 ;
        RECT 1367.185 1995.610 1367.515 1995.625 ;
        RECT 1355.930 1995.310 1367.515 1995.610 ;
        RECT 1355.930 1995.120 1359.930 1995.310 ;
        RECT 1367.185 1995.295 1367.515 1995.310 ;
      LAYER met3 ;
        RECT 357.355 1986.600 1355.930 1994.720 ;
        RECT 357.355 1985.200 1355.530 1986.600 ;
      LAYER met3 ;
        RECT 1355.930 1986.090 1359.930 1986.200 ;
        RECT 1367.185 1986.090 1367.515 1986.105 ;
        RECT 1355.930 1985.790 1367.515 1986.090 ;
        RECT 1355.930 1985.600 1359.930 1985.790 ;
        RECT 1367.185 1985.775 1367.515 1985.790 ;
      LAYER met3 ;
        RECT 357.355 1977.080 1355.930 1985.200 ;
      LAYER met3 ;
        RECT 1692.625 1981.880 1692.925 1986.480 ;
        RECT 1693.325 1984.050 1693.655 1984.065 ;
        RECT 1701.125 1984.050 1701.425 1986.480 ;
        RECT 1693.325 1983.750 1701.425 1984.050 ;
        RECT 1693.325 1983.735 1693.655 1983.750 ;
        RECT 1701.125 1981.880 1701.425 1983.750 ;
        RECT 1987.265 1984.050 1987.595 1984.065 ;
        RECT 1990.365 1984.050 1990.665 1986.480 ;
        RECT 1987.265 1983.750 1990.665 1984.050 ;
        RECT 1987.265 1983.735 1987.595 1983.750 ;
        RECT 1990.365 1981.880 1990.665 1983.750 ;
        RECT 1994.165 1983.370 1994.495 1983.385 ;
        RECT 1998.865 1983.370 1999.165 1986.480 ;
        RECT 1994.165 1983.070 1999.165 1983.370 ;
        RECT 1994.165 1983.055 1994.495 1983.070 ;
        RECT 1998.865 1981.880 1999.165 1983.070 ;
        RECT 2001.065 1983.370 2001.395 1983.385 ;
        RECT 2004.505 1983.370 2004.805 1986.480 ;
        RECT 2001.065 1983.070 2004.805 1983.370 ;
        RECT 2001.065 1983.055 2001.395 1983.070 ;
        RECT 2004.505 1981.880 2004.805 1983.070 ;
        RECT 2007.965 1982.690 2008.295 1982.705 ;
        RECT 2013.005 1982.690 2013.305 1986.480 ;
        RECT 2007.965 1982.390 2013.305 1982.690 ;
        RECT 2007.965 1982.375 2008.295 1982.390 ;
        RECT 2013.005 1981.880 2013.305 1982.390 ;
        RECT 2016.705 1982.690 2017.035 1982.705 ;
        RECT 2018.645 1982.690 2018.945 1986.480 ;
        RECT 2016.705 1982.390 2018.945 1982.690 ;
        RECT 2016.705 1982.375 2017.035 1982.390 ;
        RECT 2018.645 1981.880 2018.945 1982.390 ;
        RECT 2021.765 1982.690 2022.095 1982.705 ;
        RECT 2027.145 1982.690 2027.445 1986.480 ;
        RECT 2021.765 1982.390 2027.445 1982.690 ;
        RECT 2021.765 1982.375 2022.095 1982.390 ;
        RECT 2027.145 1981.880 2027.445 1982.390 ;
        RECT 2030.045 1982.690 2030.375 1982.705 ;
        RECT 2032.785 1982.690 2033.085 1986.480 ;
        RECT 2030.045 1982.390 2033.085 1982.690 ;
        RECT 2030.045 1982.375 2030.375 1982.390 ;
        RECT 2032.785 1981.880 2033.085 1982.390 ;
      LAYER met3 ;
        RECT 357.355 1975.680 1355.530 1977.080 ;
      LAYER met3 ;
        RECT 1355.930 1976.570 1359.930 1976.680 ;
        RECT 1367.185 1976.570 1367.515 1976.585 ;
        RECT 1355.930 1976.270 1367.515 1976.570 ;
        RECT 1355.930 1976.080 1359.930 1976.270 ;
        RECT 1367.185 1976.255 1367.515 1976.270 ;
      LAYER met3 ;
        RECT 357.355 1967.560 1355.930 1975.680 ;
        RECT 357.355 1966.160 1355.530 1967.560 ;
      LAYER met3 ;
        RECT 1355.930 1967.050 1359.930 1967.160 ;
        RECT 1367.185 1967.050 1367.515 1967.065 ;
        RECT 1355.930 1966.750 1367.515 1967.050 ;
        RECT 1355.930 1966.560 1359.930 1966.750 ;
        RECT 1367.185 1966.735 1367.515 1966.750 ;
      LAYER met3 ;
        RECT 357.355 1958.040 1355.930 1966.160 ;
      LAYER met3 ;
        RECT 1600.865 1960.260 1601.195 1960.265 ;
        RECT 1600.865 1960.250 1601.450 1960.260 ;
        RECT 1600.640 1959.950 1601.450 1960.250 ;
        RECT 1600.865 1959.940 1601.450 1959.950 ;
        RECT 1600.865 1959.935 1601.195 1959.940 ;
      LAYER met3 ;
        RECT 357.355 1956.640 1355.530 1958.040 ;
      LAYER met3 ;
        RECT 1355.930 1957.530 1359.930 1957.640 ;
        RECT 1367.185 1957.530 1367.515 1957.545 ;
        RECT 1355.930 1957.230 1367.515 1957.530 ;
        RECT 1355.930 1957.040 1359.930 1957.230 ;
        RECT 1367.185 1957.215 1367.515 1957.230 ;
      LAYER met3 ;
        RECT 357.355 1948.520 1355.930 1956.640 ;
      LAYER met3 ;
        RECT 1601.325 1949.380 1601.655 1949.385 ;
        RECT 1601.070 1949.370 1601.655 1949.380 ;
        RECT 1601.070 1949.070 1601.880 1949.370 ;
        RECT 1601.070 1949.060 1601.655 1949.070 ;
        RECT 1601.325 1949.055 1601.655 1949.060 ;
      LAYER met3 ;
        RECT 357.355 1947.120 1355.530 1948.520 ;
      LAYER met3 ;
        RECT 1355.930 1948.010 1359.930 1948.120 ;
        RECT 1367.645 1948.010 1367.975 1948.025 ;
        RECT 1355.930 1947.710 1367.975 1948.010 ;
        RECT 1355.930 1947.520 1359.930 1947.710 ;
        RECT 1367.645 1947.695 1367.975 1947.710 ;
      LAYER met3 ;
        RECT 357.355 1939.000 1355.930 1947.120 ;
      LAYER met3 ;
        RECT 1600.405 1945.290 1600.735 1945.305 ;
        RECT 1601.070 1945.290 1601.450 1945.300 ;
        RECT 1600.405 1944.990 1601.450 1945.290 ;
        RECT 1600.405 1944.975 1600.735 1944.990 ;
        RECT 1601.070 1944.980 1601.450 1944.990 ;
      LAYER met3 ;
        RECT 357.355 1937.600 1355.530 1939.000 ;
      LAYER met3 ;
        RECT 1355.930 1938.490 1359.930 1938.600 ;
        RECT 1368.105 1938.490 1368.435 1938.505 ;
        RECT 1355.930 1938.190 1368.435 1938.490 ;
        RECT 1355.930 1938.000 1359.930 1938.190 ;
        RECT 1368.105 1938.175 1368.435 1938.190 ;
        RECT 1601.325 1937.820 1601.655 1937.825 ;
        RECT 1601.070 1937.810 1601.655 1937.820 ;
      LAYER met3 ;
        RECT 357.355 1929.480 1355.930 1937.600 ;
      LAYER met3 ;
        RECT 1601.070 1937.510 1601.880 1937.810 ;
        RECT 1601.070 1937.500 1601.655 1937.510 ;
        RECT 1601.325 1937.495 1601.655 1937.500 ;
        RECT 1599.230 1932.370 1599.610 1932.380 ;
        RECT 1601.785 1932.370 1602.115 1932.385 ;
        RECT 1599.230 1932.070 1602.115 1932.370 ;
        RECT 1599.230 1932.060 1599.610 1932.070 ;
        RECT 1601.785 1932.055 1602.115 1932.070 ;
        RECT 1600.865 1931.700 1601.195 1931.705 ;
        RECT 1600.865 1931.690 1601.450 1931.700 ;
        RECT 1600.640 1931.390 1601.450 1931.690 ;
        RECT 1600.865 1931.380 1601.450 1931.390 ;
        RECT 1600.865 1931.375 1601.195 1931.380 ;
      LAYER met3 ;
        RECT 357.355 1928.080 1355.530 1929.480 ;
      LAYER met3 ;
        RECT 1355.930 1928.970 1359.930 1929.080 ;
        RECT 1367.645 1928.970 1367.975 1928.985 ;
        RECT 1355.930 1928.670 1367.975 1928.970 ;
        RECT 1355.930 1928.480 1359.930 1928.670 ;
        RECT 1367.645 1928.655 1367.975 1928.670 ;
      LAYER met3 ;
        RECT 357.355 1919.960 1355.930 1928.080 ;
      LAYER met3 ;
        RECT 1603.165 1924.220 1603.495 1924.225 ;
        RECT 1602.910 1924.210 1603.495 1924.220 ;
        RECT 1602.910 1923.910 1603.720 1924.210 ;
        RECT 1602.910 1923.900 1603.495 1923.910 ;
        RECT 1603.165 1923.895 1603.495 1923.900 ;
      LAYER met3 ;
        RECT 357.355 1918.560 1355.530 1919.960 ;
      LAYER met3 ;
        RECT 1355.930 1919.450 1359.930 1919.560 ;
        RECT 1373.165 1919.450 1373.495 1919.465 ;
        RECT 1355.930 1919.150 1373.495 1919.450 ;
        RECT 1355.930 1918.960 1359.930 1919.150 ;
        RECT 1373.165 1919.135 1373.495 1919.150 ;
        RECT 1599.230 1918.770 1599.610 1918.780 ;
        RECT 1600.865 1918.770 1601.195 1918.785 ;
      LAYER met3 ;
        RECT 357.355 1910.440 1355.930 1918.560 ;
      LAYER met3 ;
        RECT 1599.230 1918.470 1601.195 1918.770 ;
        RECT 1599.230 1918.460 1599.610 1918.470 ;
        RECT 1600.865 1918.455 1601.195 1918.470 ;
        RECT 1603.625 1918.100 1603.955 1918.105 ;
        RECT 1603.625 1918.090 1604.210 1918.100 ;
        RECT 1603.400 1917.790 1604.210 1918.090 ;
        RECT 1603.625 1917.780 1604.210 1917.790 ;
        RECT 1603.625 1917.775 1603.955 1917.780 ;
        RECT 1601.325 1916.060 1601.655 1916.065 ;
        RECT 1601.070 1916.050 1601.655 1916.060 ;
        RECT 1601.070 1915.750 1601.880 1916.050 ;
        RECT 1601.070 1915.740 1601.655 1915.750 ;
        RECT 1601.325 1915.735 1601.655 1915.740 ;
        RECT 1604.085 1912.660 1604.415 1912.665 ;
        RECT 1603.830 1912.650 1604.415 1912.660 ;
        RECT 1603.830 1912.350 1604.640 1912.650 ;
        RECT 1603.830 1912.340 1604.415 1912.350 ;
        RECT 1604.085 1912.335 1604.415 1912.340 ;
      LAYER met3 ;
        RECT 357.355 1909.040 1355.530 1910.440 ;
      LAYER met3 ;
        RECT 1355.930 1909.930 1359.930 1910.040 ;
        RECT 1367.645 1909.930 1367.975 1909.945 ;
        RECT 1355.930 1909.630 1367.975 1909.930 ;
        RECT 1355.930 1909.440 1359.930 1909.630 ;
        RECT 1367.645 1909.615 1367.975 1909.630 ;
      LAYER met3 ;
        RECT 357.355 1900.920 1355.930 1909.040 ;
      LAYER met3 ;
        RECT 1603.165 1906.540 1603.495 1906.545 ;
        RECT 1602.910 1906.530 1603.495 1906.540 ;
        RECT 1602.910 1906.230 1603.720 1906.530 ;
        RECT 1602.910 1906.220 1603.495 1906.230 ;
        RECT 1603.165 1906.215 1603.495 1906.220 ;
        RECT 1601.785 1904.500 1602.115 1904.505 ;
        RECT 1601.785 1904.490 1602.370 1904.500 ;
        RECT 1601.560 1904.190 1602.370 1904.490 ;
        RECT 1601.785 1904.180 1602.370 1904.190 ;
        RECT 1601.785 1904.175 1602.115 1904.180 ;
        RECT 1368.105 1901.770 1368.435 1901.785 ;
        RECT 1358.230 1901.470 1368.435 1901.770 ;
      LAYER met3 ;
        RECT 357.355 1899.520 1355.530 1900.920 ;
      LAYER met3 ;
        RECT 1358.230 1900.520 1358.530 1901.470 ;
        RECT 1368.105 1901.455 1368.435 1901.470 ;
        RECT 1604.085 1901.100 1604.415 1901.105 ;
        RECT 1603.830 1901.090 1604.415 1901.100 ;
        RECT 1603.830 1900.790 1604.640 1901.090 ;
        RECT 1603.830 1900.780 1604.415 1900.790 ;
        RECT 1604.085 1900.775 1604.415 1900.780 ;
        RECT 1355.930 1899.920 1359.930 1900.520 ;
      LAYER met3 ;
        RECT 357.355 1891.400 1355.930 1899.520 ;
      LAYER met3 ;
        RECT 1601.325 1898.380 1601.655 1898.385 ;
        RECT 1601.070 1898.370 1601.655 1898.380 ;
        RECT 1601.070 1898.070 1601.880 1898.370 ;
        RECT 1601.070 1898.060 1601.655 1898.070 ;
        RECT 1601.325 1898.055 1601.655 1898.060 ;
        RECT 1599.230 1897.690 1599.610 1897.700 ;
        RECT 1600.865 1897.690 1601.195 1897.705 ;
        RECT 1599.230 1897.390 1601.195 1897.690 ;
        RECT 1599.230 1897.380 1599.610 1897.390 ;
        RECT 1600.865 1897.375 1601.195 1897.390 ;
        RECT 1602.245 1894.980 1602.575 1894.985 ;
        RECT 1601.990 1894.970 1602.575 1894.980 ;
        RECT 1601.790 1894.670 1602.575 1894.970 ;
        RECT 1601.990 1894.660 1602.575 1894.670 ;
        RECT 1602.245 1894.655 1602.575 1894.660 ;
        RECT 1602.705 1892.260 1603.035 1892.265 ;
        RECT 1602.705 1892.250 1603.290 1892.260 ;
        RECT 1602.480 1891.950 1603.290 1892.250 ;
        RECT 1602.705 1891.940 1603.290 1891.950 ;
        RECT 1602.705 1891.935 1603.035 1891.940 ;
      LAYER met3 ;
        RECT 357.355 1890.000 1355.530 1891.400 ;
      LAYER met3 ;
        RECT 1355.930 1890.890 1359.930 1891.000 ;
        RECT 1372.245 1890.890 1372.575 1890.905 ;
        RECT 1355.930 1890.590 1372.575 1890.890 ;
        RECT 1355.930 1890.400 1359.930 1890.590 ;
        RECT 1372.245 1890.575 1372.575 1890.590 ;
      LAYER met3 ;
        RECT 357.355 1881.880 1355.930 1890.000 ;
      LAYER met3 ;
        RECT 1600.865 1888.850 1601.195 1888.865 ;
        RECT 1604.085 1888.860 1604.415 1888.865 ;
        RECT 1603.830 1888.850 1604.415 1888.860 ;
        RECT 1600.865 1888.550 1604.415 1888.850 ;
        RECT 1600.865 1888.535 1601.195 1888.550 ;
        RECT 1603.830 1888.540 1604.415 1888.550 ;
        RECT 1604.085 1888.535 1604.415 1888.540 ;
        RECT 1600.865 1884.090 1601.195 1884.105 ;
        RECT 1603.625 1884.090 1603.955 1884.105 ;
        RECT 1600.865 1883.790 1603.955 1884.090 ;
        RECT 1600.865 1883.775 1601.195 1883.790 ;
        RECT 1603.625 1883.775 1603.955 1883.790 ;
        RECT 1600.150 1883.410 1600.530 1883.420 ;
        RECT 1601.785 1883.410 1602.115 1883.425 ;
        RECT 1600.150 1883.110 1602.115 1883.410 ;
        RECT 1600.150 1883.100 1600.530 1883.110 ;
        RECT 1601.785 1883.095 1602.115 1883.110 ;
      LAYER met3 ;
        RECT 357.355 1880.480 1355.530 1881.880 ;
      LAYER met3 ;
        RECT 1355.930 1881.370 1359.930 1881.480 ;
        RECT 1372.245 1881.370 1372.575 1881.385 ;
        RECT 1355.930 1881.070 1372.575 1881.370 ;
        RECT 1355.930 1880.880 1359.930 1881.070 ;
        RECT 1372.245 1881.055 1372.575 1881.070 ;
        RECT 1601.325 1880.700 1601.655 1880.705 ;
        RECT 1601.070 1880.690 1601.655 1880.700 ;
      LAYER met3 ;
        RECT 357.355 1872.360 1355.930 1880.480 ;
      LAYER met3 ;
        RECT 1601.070 1880.390 1601.880 1880.690 ;
        RECT 1601.070 1880.380 1601.655 1880.390 ;
        RECT 1601.325 1880.375 1601.655 1880.380 ;
        RECT 1600.865 1877.300 1601.195 1877.305 ;
        RECT 1600.865 1877.290 1601.450 1877.300 ;
        RECT 1600.865 1876.990 1601.650 1877.290 ;
        RECT 1600.865 1876.980 1601.450 1876.990 ;
        RECT 1600.865 1876.975 1601.195 1876.980 ;
        RECT 1599.025 1875.940 1599.355 1875.945 ;
        RECT 1599.025 1875.930 1599.610 1875.940 ;
        RECT 1598.800 1875.630 1599.610 1875.930 ;
        RECT 1599.025 1875.620 1599.610 1875.630 ;
        RECT 1599.025 1875.615 1599.355 1875.620 ;
      LAYER met3 ;
        RECT 357.355 1870.960 1355.530 1872.360 ;
      LAYER met3 ;
        RECT 1355.930 1871.850 1359.930 1871.960 ;
        RECT 1372.245 1871.850 1372.575 1871.865 ;
        RECT 1355.930 1871.550 1372.575 1871.850 ;
        RECT 1355.930 1871.360 1359.930 1871.550 ;
        RECT 1372.245 1871.535 1372.575 1871.550 ;
        RECT 1602.705 1871.860 1603.035 1871.865 ;
        RECT 1602.705 1871.850 1603.290 1871.860 ;
        RECT 1602.705 1871.550 1603.490 1871.850 ;
        RECT 1602.705 1871.540 1603.290 1871.550 ;
        RECT 1602.705 1871.535 1603.035 1871.540 ;
      LAYER met3 ;
        RECT 357.355 1862.840 1355.930 1870.960 ;
      LAYER met3 ;
        RECT 1599.945 1869.140 1600.275 1869.145 ;
        RECT 1599.945 1869.130 1600.530 1869.140 ;
        RECT 1599.720 1868.830 1600.530 1869.130 ;
        RECT 1599.945 1868.820 1600.530 1868.830 ;
        RECT 1599.945 1868.815 1600.275 1868.820 ;
        RECT 1600.405 1865.740 1600.735 1865.745 ;
        RECT 1600.150 1865.730 1600.735 1865.740 ;
        RECT 1599.950 1865.430 1600.735 1865.730 ;
        RECT 1600.150 1865.420 1600.735 1865.430 ;
        RECT 1600.405 1865.415 1600.735 1865.420 ;
        RECT 1599.230 1863.690 1599.610 1863.700 ;
        RECT 1600.865 1863.690 1601.195 1863.705 ;
        RECT 1599.230 1863.390 1601.195 1863.690 ;
        RECT 1599.230 1863.380 1599.610 1863.390 ;
        RECT 1600.865 1863.375 1601.195 1863.390 ;
        RECT 1601.785 1863.020 1602.115 1863.025 ;
        RECT 1601.785 1863.010 1602.370 1863.020 ;
      LAYER met3 ;
        RECT 357.355 1861.440 1355.530 1862.840 ;
      LAYER met3 ;
        RECT 1601.560 1862.710 1602.370 1863.010 ;
        RECT 1601.785 1862.700 1602.370 1862.710 ;
        RECT 1601.785 1862.695 1602.115 1862.700 ;
        RECT 1355.930 1862.330 1359.930 1862.440 ;
        RECT 1372.245 1862.330 1372.575 1862.345 ;
        RECT 1355.930 1862.030 1372.575 1862.330 ;
        RECT 1355.930 1861.840 1359.930 1862.030 ;
        RECT 1372.245 1862.015 1372.575 1862.030 ;
        RECT 1603.165 1861.660 1603.495 1861.665 ;
        RECT 1602.910 1861.650 1603.495 1861.660 ;
      LAYER met3 ;
        RECT 357.355 1853.320 1355.930 1861.440 ;
      LAYER met3 ;
        RECT 1602.710 1861.350 1603.495 1861.650 ;
        RECT 1602.910 1861.340 1603.495 1861.350 ;
        RECT 1603.165 1861.335 1603.495 1861.340 ;
        RECT 1601.325 1857.580 1601.655 1857.585 ;
        RECT 1601.070 1857.570 1601.655 1857.580 ;
        RECT 1601.070 1857.270 1601.880 1857.570 ;
        RECT 1601.070 1857.260 1601.655 1857.270 ;
        RECT 1601.325 1857.255 1601.655 1857.260 ;
        RECT 1604.085 1856.220 1604.415 1856.225 ;
        RECT 1603.830 1856.210 1604.415 1856.220 ;
        RECT 1603.630 1855.910 1604.415 1856.210 ;
        RECT 1603.830 1855.900 1604.415 1855.910 ;
        RECT 1604.085 1855.895 1604.415 1855.900 ;
      LAYER met3 ;
        RECT 357.355 1851.920 1355.530 1853.320 ;
      LAYER met3 ;
        RECT 1355.930 1852.810 1359.930 1852.920 ;
        RECT 1372.245 1852.810 1372.575 1852.825 ;
        RECT 1355.930 1852.510 1372.575 1852.810 ;
        RECT 1355.930 1852.320 1359.930 1852.510 ;
        RECT 1372.245 1852.495 1372.575 1852.510 ;
      LAYER met3 ;
        RECT 357.355 1843.800 1355.930 1851.920 ;
      LAYER met3 ;
        RECT 1602.245 1848.740 1602.575 1848.745 ;
        RECT 1601.990 1848.730 1602.575 1848.740 ;
        RECT 1601.790 1848.430 1602.575 1848.730 ;
        RECT 1601.990 1848.420 1602.575 1848.430 ;
        RECT 1602.030 1848.415 1602.575 1848.420 ;
        RECT 1602.030 1847.370 1602.330 1848.415 ;
        RECT 1603.625 1847.370 1603.955 1847.385 ;
        RECT 1602.030 1847.070 1603.955 1847.370 ;
        RECT 1603.625 1847.055 1603.955 1847.070 ;
        RECT 1601.785 1846.020 1602.115 1846.025 ;
        RECT 1601.785 1846.010 1602.370 1846.020 ;
        RECT 1601.560 1845.710 1602.370 1846.010 ;
        RECT 1601.785 1845.700 1602.370 1845.710 ;
        RECT 1601.785 1845.695 1602.115 1845.700 ;
      LAYER met3 ;
        RECT 357.355 1842.400 1355.530 1843.800 ;
      LAYER met3 ;
        RECT 1355.930 1843.290 1359.930 1843.400 ;
        RECT 1368.105 1843.290 1368.435 1843.305 ;
        RECT 1355.930 1842.990 1368.435 1843.290 ;
        RECT 1355.930 1842.800 1359.930 1842.990 ;
        RECT 1368.105 1842.975 1368.435 1842.990 ;
        RECT 1599.230 1842.610 1599.610 1842.620 ;
        RECT 1600.865 1842.610 1601.195 1842.625 ;
        RECT 1604.085 1842.620 1604.415 1842.625 ;
        RECT 1603.830 1842.610 1604.415 1842.620 ;
      LAYER met3 ;
        RECT 357.355 1834.280 1355.930 1842.400 ;
      LAYER met3 ;
        RECT 1599.230 1842.310 1601.195 1842.610 ;
        RECT 1603.630 1842.310 1604.415 1842.610 ;
        RECT 1599.230 1842.300 1599.610 1842.310 ;
        RECT 1600.865 1842.295 1601.195 1842.310 ;
        RECT 1603.830 1842.300 1604.415 1842.310 ;
        RECT 1604.085 1842.295 1604.415 1842.300 ;
        RECT 1601.325 1839.900 1601.655 1839.905 ;
        RECT 1601.070 1839.890 1601.655 1839.900 ;
        RECT 1601.070 1839.590 1601.880 1839.890 ;
        RECT 1601.070 1839.580 1601.655 1839.590 ;
        RECT 1601.325 1839.575 1601.655 1839.580 ;
        RECT 1604.085 1836.500 1604.415 1836.505 ;
        RECT 1598.310 1836.490 1598.690 1836.500 ;
        RECT 1603.830 1836.490 1604.415 1836.500 ;
        RECT 1598.310 1836.190 1604.415 1836.490 ;
        RECT 1598.310 1836.180 1598.690 1836.190 ;
        RECT 1603.830 1836.180 1604.415 1836.190 ;
        RECT 1604.085 1836.175 1604.415 1836.180 ;
      LAYER met3 ;
        RECT 357.355 1832.880 1355.530 1834.280 ;
      LAYER met3 ;
        RECT 1355.930 1833.770 1359.930 1833.880 ;
        RECT 1372.705 1833.770 1373.035 1833.785 ;
        RECT 1355.930 1833.470 1373.035 1833.770 ;
        RECT 1355.930 1833.280 1359.930 1833.470 ;
        RECT 1372.705 1833.455 1373.035 1833.470 ;
      LAYER met3 ;
        RECT 357.355 1824.760 1355.930 1832.880 ;
      LAYER met3 ;
        RECT 1603.165 1831.060 1603.495 1831.065 ;
        RECT 1602.910 1831.050 1603.495 1831.060 ;
        RECT 1602.710 1830.750 1603.495 1831.050 ;
        RECT 1602.910 1830.740 1603.495 1830.750 ;
        RECT 1603.165 1830.735 1603.495 1830.740 ;
        RECT 1599.025 1828.330 1599.355 1828.345 ;
        RECT 1600.150 1828.330 1600.530 1828.340 ;
        RECT 1599.025 1828.030 1600.530 1828.330 ;
        RECT 1599.025 1828.015 1599.355 1828.030 ;
        RECT 1600.150 1828.020 1600.530 1828.030 ;
        RECT 1600.865 1824.940 1601.195 1824.945 ;
        RECT 1600.865 1824.930 1601.450 1824.940 ;
        RECT 1603.165 1824.930 1603.495 1824.945 ;
      LAYER met3 ;
        RECT 357.355 1823.360 1355.530 1824.760 ;
      LAYER met3 ;
        RECT 1600.865 1824.630 1603.495 1824.930 ;
        RECT 1600.865 1824.620 1601.450 1824.630 ;
        RECT 1600.865 1824.615 1601.195 1824.620 ;
        RECT 1603.165 1824.615 1603.495 1824.630 ;
        RECT 1355.930 1824.250 1359.930 1824.360 ;
        RECT 1369.025 1824.250 1369.355 1824.265 ;
        RECT 1355.930 1823.950 1369.355 1824.250 ;
        RECT 1355.930 1823.760 1359.930 1823.950 ;
        RECT 1369.025 1823.935 1369.355 1823.950 ;
      LAYER met3 ;
        RECT 357.355 1815.240 1355.930 1823.360 ;
      LAYER met3 ;
        RECT 1602.245 1822.220 1602.575 1822.225 ;
        RECT 1601.990 1822.210 1602.575 1822.220 ;
        RECT 1601.990 1821.910 1602.800 1822.210 ;
        RECT 1601.990 1821.900 1602.575 1821.910 ;
        RECT 1602.245 1821.895 1602.575 1821.900 ;
        RECT 1599.945 1818.820 1600.275 1818.825 ;
        RECT 1599.945 1818.810 1600.530 1818.820 ;
        RECT 1599.945 1818.510 1600.730 1818.810 ;
        RECT 1599.945 1818.500 1600.530 1818.510 ;
        RECT 1599.945 1818.495 1600.275 1818.500 ;
        RECT 1593.965 1817.450 1594.295 1817.465 ;
        RECT 1597.390 1817.450 1597.770 1817.460 ;
        RECT 1593.965 1817.150 1597.770 1817.450 ;
        RECT 1593.965 1817.135 1594.295 1817.150 ;
        RECT 1597.390 1817.140 1597.770 1817.150 ;
      LAYER met3 ;
        RECT 357.355 1813.840 1355.530 1815.240 ;
      LAYER met3 ;
        RECT 1355.930 1814.730 1359.930 1814.840 ;
        RECT 1371.785 1814.730 1372.115 1814.745 ;
        RECT 1355.930 1814.430 1372.115 1814.730 ;
        RECT 1355.930 1814.240 1359.930 1814.430 ;
        RECT 1371.785 1814.415 1372.115 1814.430 ;
      LAYER met3 ;
        RECT 357.355 1805.720 1355.930 1813.840 ;
      LAYER met3 ;
        RECT 1600.405 1813.380 1600.735 1813.385 ;
        RECT 1600.150 1813.370 1600.735 1813.380 ;
        RECT 1599.950 1813.070 1600.735 1813.370 ;
        RECT 1600.150 1813.060 1600.735 1813.070 ;
        RECT 1600.405 1813.055 1600.735 1813.060 ;
        RECT 1601.785 1810.660 1602.115 1810.665 ;
        RECT 1601.785 1810.650 1602.370 1810.660 ;
        RECT 1601.560 1810.350 1602.370 1810.650 ;
        RECT 1601.785 1810.340 1602.370 1810.350 ;
        RECT 1601.785 1810.335 1602.115 1810.340 ;
        RECT 1599.025 1807.260 1599.355 1807.265 ;
        RECT 1600.865 1807.260 1601.195 1807.265 ;
        RECT 1599.025 1807.250 1599.610 1807.260 ;
        RECT 1598.800 1806.950 1599.610 1807.250 ;
        RECT 1599.025 1806.940 1599.610 1806.950 ;
        RECT 1600.865 1807.250 1601.450 1807.260 ;
        RECT 1600.865 1806.950 1601.650 1807.250 ;
        RECT 1600.865 1806.940 1601.450 1806.950 ;
        RECT 1599.025 1806.935 1599.355 1806.940 ;
        RECT 1600.865 1806.935 1601.195 1806.940 ;
      LAYER met3 ;
        RECT 357.355 1804.320 1355.530 1805.720 ;
      LAYER met3 ;
        RECT 1355.930 1805.210 1359.930 1805.320 ;
        RECT 1367.645 1805.210 1367.975 1805.225 ;
        RECT 1601.325 1805.220 1601.655 1805.225 ;
        RECT 1355.930 1804.910 1367.975 1805.210 ;
        RECT 1355.930 1804.720 1359.930 1804.910 ;
        RECT 1367.645 1804.895 1367.975 1804.910 ;
        RECT 1601.070 1805.210 1601.655 1805.220 ;
        RECT 1601.070 1804.910 1601.880 1805.210 ;
        RECT 1601.070 1804.900 1601.655 1804.910 ;
        RECT 1601.325 1804.895 1601.655 1804.900 ;
      LAYER met3 ;
        RECT 357.355 1796.200 1355.930 1804.320 ;
      LAYER met3 ;
        RECT 1601.325 1801.820 1601.655 1801.825 ;
        RECT 1601.070 1801.810 1601.655 1801.820 ;
        RECT 1600.870 1801.510 1601.655 1801.810 ;
        RECT 1601.070 1801.500 1601.655 1801.510 ;
        RECT 1601.325 1801.495 1601.655 1801.500 ;
        RECT 1602.245 1799.100 1602.575 1799.105 ;
        RECT 1601.990 1799.090 1602.575 1799.100 ;
        RECT 1603.625 1799.090 1603.955 1799.105 ;
        RECT 1601.790 1798.790 1603.955 1799.090 ;
        RECT 1601.990 1798.780 1602.575 1798.790 ;
        RECT 1602.245 1798.775 1602.575 1798.780 ;
        RECT 1603.625 1798.775 1603.955 1798.790 ;
      LAYER met3 ;
        RECT 357.355 1794.800 1355.530 1796.200 ;
      LAYER met3 ;
        RECT 1355.930 1795.690 1359.930 1795.800 ;
        RECT 1369.025 1795.690 1369.355 1795.705 ;
        RECT 1355.930 1795.390 1369.355 1795.690 ;
        RECT 1355.930 1795.200 1359.930 1795.390 ;
        RECT 1369.025 1795.375 1369.355 1795.390 ;
      LAYER met3 ;
        RECT 357.355 1786.680 1355.930 1794.800 ;
      LAYER met3 ;
        RECT 1601.785 1792.980 1602.115 1792.985 ;
        RECT 1601.785 1792.970 1602.370 1792.980 ;
        RECT 1601.560 1792.670 1602.370 1792.970 ;
        RECT 1601.785 1792.660 1602.370 1792.670 ;
        RECT 1601.785 1792.655 1602.115 1792.660 ;
        RECT 1601.325 1789.580 1601.655 1789.585 ;
        RECT 1601.070 1789.570 1601.655 1789.580 ;
        RECT 1600.870 1789.270 1601.655 1789.570 ;
        RECT 1601.070 1789.260 1601.655 1789.270 ;
        RECT 1601.325 1789.255 1601.655 1789.260 ;
      LAYER met3 ;
        RECT 357.355 1785.280 1355.530 1786.680 ;
      LAYER met3 ;
        RECT 1355.930 1786.170 1359.930 1786.280 ;
        RECT 1369.230 1786.170 1369.610 1786.180 ;
        RECT 1355.930 1785.870 1369.610 1786.170 ;
        RECT 1355.930 1785.680 1359.930 1785.870 ;
        RECT 1369.230 1785.860 1369.610 1785.870 ;
        RECT 1602.705 1785.500 1603.035 1785.505 ;
        RECT 1602.705 1785.490 1603.290 1785.500 ;
      LAYER met3 ;
        RECT 357.355 1777.160 1355.930 1785.280 ;
      LAYER met3 ;
        RECT 1602.480 1785.190 1603.290 1785.490 ;
        RECT 1602.705 1785.180 1603.290 1785.190 ;
        RECT 1602.705 1785.175 1603.035 1785.180 ;
        RECT 1600.865 1784.140 1601.195 1784.145 ;
        RECT 1600.865 1784.130 1601.450 1784.140 ;
        RECT 1600.640 1783.830 1601.450 1784.130 ;
        RECT 1600.865 1783.820 1601.450 1783.830 ;
        RECT 1600.865 1783.815 1601.195 1783.820 ;
        RECT 1603.165 1780.060 1603.495 1780.065 ;
        RECT 1602.910 1780.050 1603.495 1780.060 ;
        RECT 1602.910 1779.750 1603.720 1780.050 ;
        RECT 1602.910 1779.740 1603.495 1779.750 ;
        RECT 1603.165 1779.735 1603.495 1779.740 ;
        RECT 1600.865 1778.020 1601.195 1778.025 ;
        RECT 1600.865 1778.010 1601.450 1778.020 ;
        RECT 1600.640 1777.710 1601.450 1778.010 ;
        RECT 1600.865 1777.700 1601.450 1777.710 ;
        RECT 1600.865 1777.695 1601.195 1777.700 ;
      LAYER met3 ;
        RECT 357.355 1775.760 1355.530 1777.160 ;
      LAYER met3 ;
        RECT 1355.930 1776.650 1359.930 1776.760 ;
        RECT 1371.785 1776.650 1372.115 1776.665 ;
        RECT 1355.930 1776.350 1372.115 1776.650 ;
        RECT 1355.930 1776.160 1359.930 1776.350 ;
        RECT 1371.785 1776.335 1372.115 1776.350 ;
      LAYER met3 ;
        RECT 357.355 1767.640 1355.930 1775.760 ;
      LAYER met3 ;
        RECT 1604.085 1773.260 1604.415 1773.265 ;
        RECT 1603.830 1773.250 1604.415 1773.260 ;
        RECT 1603.630 1772.950 1604.415 1773.250 ;
        RECT 1603.830 1772.940 1604.415 1772.950 ;
        RECT 1604.085 1772.935 1604.415 1772.940 ;
        RECT 1600.865 1772.580 1601.195 1772.585 ;
        RECT 1600.865 1772.570 1601.450 1772.580 ;
        RECT 1600.640 1772.270 1601.450 1772.570 ;
        RECT 1600.865 1772.260 1601.450 1772.270 ;
        RECT 1600.865 1772.255 1601.195 1772.260 ;
      LAYER met3 ;
        RECT 357.355 1766.240 1355.530 1767.640 ;
      LAYER met3 ;
        RECT 1355.930 1767.130 1359.930 1767.240 ;
        RECT 1369.025 1767.130 1369.355 1767.145 ;
        RECT 1355.930 1766.830 1369.355 1767.130 ;
        RECT 1355.930 1766.640 1359.930 1766.830 ;
        RECT 1369.025 1766.815 1369.355 1766.830 ;
        RECT 1599.230 1767.130 1599.610 1767.140 ;
        RECT 1601.325 1767.130 1601.655 1767.145 ;
        RECT 1599.230 1766.830 1601.655 1767.130 ;
        RECT 1599.230 1766.820 1599.610 1766.830 ;
        RECT 1601.325 1766.815 1601.655 1766.830 ;
        RECT 1601.325 1766.460 1601.655 1766.465 ;
        RECT 1604.085 1766.460 1604.415 1766.465 ;
        RECT 1601.070 1766.450 1601.655 1766.460 ;
        RECT 1603.830 1766.450 1604.415 1766.460 ;
      LAYER met3 ;
        RECT 357.355 1758.120 1355.930 1766.240 ;
      LAYER met3 ;
        RECT 1601.070 1766.150 1601.880 1766.450 ;
        RECT 1603.630 1766.150 1604.415 1766.450 ;
        RECT 1601.070 1766.140 1601.655 1766.150 ;
        RECT 1603.830 1766.140 1604.415 1766.150 ;
        RECT 1601.325 1766.135 1601.655 1766.140 ;
        RECT 1604.085 1766.135 1604.415 1766.140 ;
        RECT 1600.865 1763.060 1601.195 1763.065 ;
        RECT 1600.865 1763.050 1601.450 1763.060 ;
        RECT 1600.640 1762.750 1601.450 1763.050 ;
        RECT 1600.865 1762.740 1601.450 1762.750 ;
        RECT 1600.865 1762.735 1601.195 1762.740 ;
        RECT 1601.785 1762.380 1602.115 1762.385 ;
        RECT 1601.785 1762.370 1602.370 1762.380 ;
        RECT 1601.560 1762.070 1602.370 1762.370 ;
        RECT 1601.785 1762.060 1602.370 1762.070 ;
        RECT 1601.785 1762.055 1602.115 1762.060 ;
      LAYER met3 ;
        RECT 357.355 1756.720 1355.530 1758.120 ;
      LAYER met3 ;
        RECT 1355.930 1757.610 1359.930 1757.720 ;
        RECT 1372.705 1757.610 1373.035 1757.625 ;
        RECT 1355.930 1757.310 1373.035 1757.610 ;
        RECT 1355.930 1757.120 1359.930 1757.310 ;
        RECT 1372.705 1757.295 1373.035 1757.310 ;
      LAYER met3 ;
        RECT 357.355 1748.600 1355.930 1756.720 ;
      LAYER met3 ;
        RECT 1603.165 1756.260 1603.495 1756.265 ;
        RECT 1602.910 1756.250 1603.495 1756.260 ;
        RECT 1602.910 1755.950 1603.720 1756.250 ;
        RECT 1602.910 1755.940 1603.495 1755.950 ;
        RECT 1603.165 1755.935 1603.495 1755.940 ;
        RECT 1601.785 1754.900 1602.115 1754.905 ;
        RECT 1601.785 1754.890 1602.370 1754.900 ;
        RECT 1601.560 1754.590 1602.370 1754.890 ;
        RECT 1601.785 1754.580 1602.370 1754.590 ;
        RECT 1601.785 1754.575 1602.115 1754.580 ;
        RECT 1603.625 1750.820 1603.955 1750.825 ;
        RECT 1603.625 1750.810 1604.210 1750.820 ;
        RECT 1603.625 1750.510 1604.410 1750.810 ;
        RECT 1603.625 1750.500 1604.210 1750.510 ;
        RECT 1603.625 1750.495 1603.955 1750.500 ;
        RECT 1600.865 1748.780 1601.195 1748.785 ;
        RECT 1600.865 1748.770 1601.450 1748.780 ;
      LAYER met3 ;
        RECT 357.355 1747.200 1355.530 1748.600 ;
      LAYER met3 ;
        RECT 1600.640 1748.470 1601.450 1748.770 ;
        RECT 1600.865 1748.460 1601.450 1748.470 ;
        RECT 1600.865 1748.455 1601.195 1748.460 ;
        RECT 1355.930 1748.090 1359.930 1748.200 ;
        RECT 1367.645 1748.090 1367.975 1748.105 ;
        RECT 1355.930 1747.790 1367.975 1748.090 ;
        RECT 1355.930 1747.600 1359.930 1747.790 ;
        RECT 1367.645 1747.775 1367.975 1747.790 ;
      LAYER met3 ;
        RECT 357.355 1739.080 1355.930 1747.200 ;
      LAYER met3 ;
        RECT 1600.865 1743.340 1601.195 1743.345 ;
        RECT 1600.865 1743.330 1601.450 1743.340 ;
        RECT 1600.640 1743.030 1601.450 1743.330 ;
        RECT 1600.865 1743.020 1601.450 1743.030 ;
        RECT 1600.865 1743.015 1601.195 1743.020 ;
      LAYER met3 ;
        RECT 357.355 1737.680 1355.530 1739.080 ;
      LAYER met3 ;
        RECT 1355.930 1738.570 1359.930 1738.680 ;
        RECT 1367.645 1738.570 1367.975 1738.585 ;
        RECT 1355.930 1738.270 1367.975 1738.570 ;
        RECT 1355.930 1738.080 1359.930 1738.270 ;
        RECT 1367.645 1738.255 1367.975 1738.270 ;
      LAYER met3 ;
        RECT 357.355 1729.560 1355.930 1737.680 ;
      LAYER met3 ;
        RECT 1600.865 1731.780 1601.195 1731.785 ;
        RECT 1600.865 1731.770 1601.450 1731.780 ;
        RECT 1600.640 1731.470 1601.450 1731.770 ;
        RECT 1600.865 1731.460 1601.450 1731.470 ;
        RECT 1600.865 1731.455 1601.195 1731.460 ;
      LAYER met3 ;
        RECT 357.355 1728.160 1355.530 1729.560 ;
      LAYER met3 ;
        RECT 1355.930 1729.050 1359.930 1729.160 ;
        RECT 1367.645 1729.050 1367.975 1729.065 ;
        RECT 1355.930 1728.750 1367.975 1729.050 ;
        RECT 1355.930 1728.560 1359.930 1728.750 ;
        RECT 1367.645 1728.735 1367.975 1728.750 ;
      LAYER met3 ;
        RECT 357.355 1720.040 1355.930 1728.160 ;
        RECT 357.355 1718.640 1355.530 1720.040 ;
      LAYER met3 ;
        RECT 1355.930 1719.530 1359.930 1719.640 ;
        RECT 1368.105 1719.530 1368.435 1719.545 ;
        RECT 1355.930 1719.230 1368.435 1719.530 ;
        RECT 1355.930 1719.040 1359.930 1719.230 ;
        RECT 1368.105 1719.215 1368.435 1719.230 ;
      LAYER met3 ;
        RECT 357.355 1710.520 1355.930 1718.640 ;
        RECT 357.355 1709.120 1355.530 1710.520 ;
      LAYER met3 ;
        RECT 1355.930 1710.010 1359.930 1710.120 ;
        RECT 1367.645 1710.010 1367.975 1710.025 ;
        RECT 1355.930 1709.710 1367.975 1710.010 ;
        RECT 1355.930 1709.520 1359.930 1709.710 ;
        RECT 1367.645 1709.695 1367.975 1709.710 ;
      LAYER met3 ;
        RECT 357.355 1701.000 1355.930 1709.120 ;
        RECT 357.355 1699.600 1355.530 1701.000 ;
      LAYER met3 ;
        RECT 1355.930 1700.490 1359.930 1700.600 ;
        RECT 1367.645 1700.490 1367.975 1700.505 ;
        RECT 1355.930 1700.190 1367.975 1700.490 ;
        RECT 1355.930 1700.000 1359.930 1700.190 ;
        RECT 1367.645 1700.175 1367.975 1700.190 ;
      LAYER met3 ;
        RECT 357.355 1691.480 1355.930 1699.600 ;
        RECT 357.355 1690.080 1355.530 1691.480 ;
      LAYER met3 ;
        RECT 1355.930 1690.970 1359.930 1691.080 ;
        RECT 1369.485 1690.970 1369.815 1690.985 ;
        RECT 1355.930 1690.670 1369.815 1690.970 ;
        RECT 1355.930 1690.480 1359.930 1690.670 ;
        RECT 1369.485 1690.655 1369.815 1690.670 ;
      LAYER met3 ;
        RECT 357.355 1681.960 1355.930 1690.080 ;
        RECT 357.355 1680.560 1355.530 1681.960 ;
      LAYER met3 ;
        RECT 1355.930 1681.450 1359.930 1681.560 ;
        RECT 1366.265 1681.450 1366.595 1681.465 ;
        RECT 1355.930 1681.150 1366.595 1681.450 ;
        RECT 1355.930 1680.960 1359.930 1681.150 ;
        RECT 1366.265 1681.135 1366.595 1681.150 ;
      LAYER met3 ;
        RECT 357.355 1672.440 1355.930 1680.560 ;
        RECT 357.355 1671.040 1355.530 1672.440 ;
      LAYER met3 ;
        RECT 1355.930 1671.930 1359.930 1672.040 ;
        RECT 1369.025 1671.930 1369.355 1671.945 ;
        RECT 1355.930 1671.630 1369.355 1671.930 ;
        RECT 1355.930 1671.440 1359.930 1671.630 ;
        RECT 1369.025 1671.615 1369.355 1671.630 ;
      LAYER met3 ;
        RECT 357.355 1662.920 1355.930 1671.040 ;
        RECT 357.355 1661.520 1355.530 1662.920 ;
      LAYER met3 ;
        RECT 1355.930 1662.410 1359.930 1662.520 ;
        RECT 1371.325 1662.410 1371.655 1662.425 ;
        RECT 1355.930 1662.110 1371.655 1662.410 ;
        RECT 1355.930 1661.920 1359.930 1662.110 ;
        RECT 1371.325 1662.095 1371.655 1662.110 ;
      LAYER met3 ;
        RECT 357.355 1653.400 1355.930 1661.520 ;
        RECT 357.355 1652.000 1355.530 1653.400 ;
      LAYER met3 ;
        RECT 1355.930 1652.890 1359.930 1653.000 ;
        RECT 1366.725 1652.890 1367.055 1652.905 ;
        RECT 1355.930 1652.590 1367.055 1652.890 ;
        RECT 1355.930 1652.400 1359.930 1652.590 ;
        RECT 1366.725 1652.575 1367.055 1652.590 ;
      LAYER met3 ;
        RECT 357.355 1643.880 1355.930 1652.000 ;
        RECT 357.355 1642.480 1355.530 1643.880 ;
      LAYER met3 ;
        RECT 1355.930 1643.370 1359.930 1643.480 ;
        RECT 1369.945 1643.370 1370.275 1643.385 ;
        RECT 1355.930 1643.070 1370.275 1643.370 ;
        RECT 1355.930 1642.880 1359.930 1643.070 ;
        RECT 1369.945 1643.055 1370.275 1643.070 ;
      LAYER met3 ;
        RECT 357.355 1634.360 1355.930 1642.480 ;
        RECT 357.355 1632.960 1355.530 1634.360 ;
      LAYER met3 ;
        RECT 1355.930 1633.850 1359.930 1633.960 ;
        RECT 1367.645 1633.850 1367.975 1633.865 ;
        RECT 1355.930 1633.550 1367.975 1633.850 ;
        RECT 1355.930 1633.360 1359.930 1633.550 ;
        RECT 1367.645 1633.535 1367.975 1633.550 ;
      LAYER met3 ;
        RECT 357.355 1624.840 1355.930 1632.960 ;
        RECT 357.355 1623.440 1355.530 1624.840 ;
      LAYER met3 ;
        RECT 1355.930 1624.330 1359.930 1624.440 ;
        RECT 1367.185 1624.330 1367.515 1624.345 ;
        RECT 1355.930 1624.030 1367.515 1624.330 ;
        RECT 1355.930 1623.840 1359.930 1624.030 ;
        RECT 1367.185 1624.015 1367.515 1624.030 ;
      LAYER met3 ;
        RECT 357.355 1615.320 1355.930 1623.440 ;
        RECT 357.355 1613.920 1355.530 1615.320 ;
      LAYER met3 ;
        RECT 1355.930 1614.810 1359.930 1614.920 ;
        RECT 1367.645 1614.810 1367.975 1614.825 ;
        RECT 1355.930 1614.510 1367.975 1614.810 ;
        RECT 1355.930 1614.320 1359.930 1614.510 ;
        RECT 1367.645 1614.495 1367.975 1614.510 ;
      LAYER met3 ;
        RECT 357.355 1605.800 1355.930 1613.920 ;
        RECT 357.355 1604.935 1355.530 1605.800 ;
      LAYER met3 ;
        RECT 1355.930 1605.290 1359.930 1605.400 ;
        RECT 1367.185 1605.290 1367.515 1605.305 ;
        RECT 1355.930 1604.990 1367.515 1605.290 ;
      LAYER met3 ;
        RECT 1605.000 1605.000 2051.235 1981.480 ;
      LAYER met3 ;
        RECT 2051.235 1625.460 2052.140 1627.200 ;
        RECT 2051.235 1605.000 2052.140 1605.440 ;
        RECT 1355.930 1604.800 1359.930 1604.990 ;
        RECT 1367.185 1604.975 1367.515 1604.990 ;
        RECT 1704.490 1600.000 1704.790 1604.600 ;
        RECT 1710.130 1600.000 1710.430 1604.600 ;
        RECT 1718.630 1600.000 1718.930 1604.600 ;
        RECT 1724.270 1600.000 1724.570 1604.600 ;
        RECT 1732.770 1600.000 1733.070 1604.600 ;
        RECT 1738.410 1600.000 1738.710 1604.600 ;
        RECT 1746.910 1600.000 1747.210 1604.600 ;
        RECT 2043.600 1602.430 2044.660 1605.000 ;
        RECT 2048.265 1600.000 2048.565 1604.600 ;
        RECT 2050.400 1600.180 2052.140 1605.000 ;
      LAYER via3 ;
        RECT 784.720 3300.440 786.240 3302.050 ;
        RECT 782.500 3293.620 784.020 3294.630 ;
        RECT 1334.720 3300.440 1336.240 3302.050 ;
        RECT 1332.500 3293.620 1334.020 3294.630 ;
        RECT 517.340 2851.420 517.660 2851.740 ;
        RECT 1103.380 2850.740 1103.700 2851.060 ;
        RECT 568.940 2848.020 569.260 2848.340 ;
        RECT 592.300 2848.020 592.620 2848.340 ;
        RECT 1089.120 2848.020 1089.440 2848.340 ;
        RECT 597.380 2845.300 597.700 2845.620 ;
        RECT 604.740 2845.300 605.060 2845.620 ;
        RECT 613.020 2843.940 613.340 2844.260 ;
        RECT 573.460 2843.260 573.780 2843.580 ;
        RECT 575.300 2843.260 575.620 2843.580 ;
        RECT 432.700 2842.580 433.020 2842.900 ;
        RECT 507.220 2842.580 507.540 2842.900 ;
        RECT 523.780 2842.580 524.100 2842.900 ;
        RECT 526.540 2842.580 526.860 2842.900 ;
        RECT 529.300 2842.580 529.620 2842.900 ;
        RECT 533.900 2842.580 534.220 2842.900 ;
        RECT 543.100 2842.580 543.420 2842.900 ;
        RECT 557.820 2842.580 558.140 2842.900 ;
        RECT 642.460 2842.580 642.780 2842.900 ;
        RECT 981.020 2842.580 981.340 2842.900 ;
        RECT 988.380 2842.580 988.700 2842.900 ;
        RECT 1019.660 2842.580 1019.980 2842.900 ;
        RECT 1024.260 2842.580 1024.580 2842.900 ;
        RECT 1027.020 2842.580 1027.340 2842.900 ;
        RECT 1065.660 2842.580 1065.980 2842.900 ;
        RECT 1070.260 2842.580 1070.580 2842.900 ;
        RECT 1111.660 2842.580 1111.980 2842.900 ;
        RECT 1118.100 2842.580 1118.420 2842.900 ;
        RECT 1130.980 2842.580 1131.300 2842.900 ;
        RECT 1135.580 2842.580 1135.900 2842.900 ;
        RECT 1136.500 2842.580 1136.820 2842.900 ;
        RECT 1143.860 2842.580 1144.180 2842.900 ;
        RECT 1151.220 2842.580 1151.540 2842.900 ;
        RECT 1153.980 2842.580 1154.300 2842.900 ;
        RECT 1165.020 2842.580 1165.340 2842.900 ;
        RECT 1172.380 2842.580 1172.700 2842.900 ;
        RECT 1178.820 2842.580 1179.140 2842.900 ;
        RECT 1186.180 2842.580 1186.500 2842.900 ;
        RECT 1190.780 2842.580 1191.100 2842.900 ;
        RECT 475.940 2841.900 476.260 2842.220 ;
        RECT 549.540 2841.900 549.860 2842.220 ;
        RECT 1018.740 2841.900 1019.060 2842.220 ;
        RECT 1128.220 2841.900 1128.540 2842.220 ;
        RECT 1163.180 2841.900 1163.500 2842.220 ;
        RECT 480.540 2841.220 480.860 2841.540 ;
        RECT 504.460 2841.220 504.780 2841.540 ;
        RECT 618.540 2841.220 618.860 2841.540 ;
        RECT 621.300 2841.220 621.620 2841.540 ;
        RECT 626.820 2841.220 627.140 2841.540 ;
        RECT 647.980 2841.220 648.300 2841.540 ;
        RECT 1001.260 2840.540 1001.580 2840.860 ;
        RECT 1164.100 2840.540 1164.420 2840.860 ;
        RECT 1180.660 2840.540 1180.980 2840.860 ;
        RECT 1007.700 2839.860 1008.020 2840.180 ;
        RECT 1159.500 2839.860 1159.820 2840.180 ;
        RECT 457.540 2838.500 457.860 2838.820 ;
        RECT 488.820 2838.500 489.140 2838.820 ;
        RECT 501.700 2838.500 502.020 2838.820 ;
        RECT 551.380 2838.500 551.700 2838.820 ;
        RECT 442.820 2837.140 443.140 2837.460 ;
        RECT 437.300 2836.460 437.620 2836.780 ;
        RECT 450.180 2836.460 450.500 2836.780 ;
        RECT 621.300 2836.460 621.620 2836.780 ;
        RECT 1041.740 2836.460 1042.060 2836.780 ;
        RECT 466.740 2835.780 467.060 2836.100 ;
        RECT 471.340 2835.780 471.660 2836.100 ;
        RECT 481.460 2835.780 481.780 2836.100 ;
        RECT 494.340 2835.780 494.660 2836.100 ;
        RECT 624.060 2835.780 624.380 2836.100 ;
        RECT 633.260 2835.780 633.580 2836.100 ;
        RECT 640.620 2835.780 640.940 2836.100 ;
        RECT 1039.900 2835.780 1040.220 2836.100 ;
        RECT 1046.340 2835.780 1046.660 2836.100 ;
        RECT 1054.620 2835.780 1054.940 2836.100 ;
        RECT 1061.980 2835.780 1062.300 2836.100 ;
        RECT 1067.500 2835.780 1067.820 2836.100 ;
        RECT 1073.940 2835.780 1074.260 2836.100 ;
        RECT 1081.300 2835.780 1081.620 2836.100 ;
        RECT 1089.580 2835.780 1089.900 2836.100 ;
        RECT 1096.020 2835.780 1096.340 2836.100 ;
        RECT 1109.820 2835.780 1110.140 2836.100 ;
        RECT 1116.260 2835.780 1116.580 2836.100 ;
        RECT 1119.020 2835.780 1119.340 2836.100 ;
        RECT 586.340 2832.380 586.660 2832.700 ;
        RECT 1369.260 2582.140 1369.580 2582.460 ;
        RECT 1601.100 2560.380 1601.420 2560.700 ;
        RECT 1600.180 2545.420 1600.500 2545.740 ;
        RECT 1600.180 2539.300 1600.500 2539.620 ;
        RECT 1602.020 2537.260 1602.340 2537.580 ;
        RECT 1599.260 2531.140 1599.580 2531.460 ;
        RECT 1601.100 2531.140 1601.420 2531.460 ;
        RECT 1603.860 2523.660 1604.180 2523.980 ;
        RECT 1383.060 2518.900 1383.380 2519.220 ;
        RECT 1599.260 2518.900 1599.580 2519.220 ;
        RECT 1602.940 2518.220 1603.260 2518.540 ;
        RECT 1601.100 2515.500 1601.420 2515.820 ;
        RECT 1602.020 2512.100 1602.340 2512.420 ;
        RECT 1603.860 2506.660 1604.180 2506.980 ;
        RECT 1599.260 2504.620 1599.580 2504.940 ;
        RECT 1600.180 2503.940 1600.500 2504.260 ;
        RECT 1602.940 2500.540 1603.260 2500.860 ;
        RECT 1601.100 2497.820 1601.420 2498.140 ;
        RECT 1603.860 2494.420 1604.180 2494.740 ;
        RECT 1599.260 2489.660 1599.580 2489.980 ;
        RECT 1601.100 2488.980 1601.420 2489.300 ;
        RECT 1601.100 2486.260 1601.420 2486.580 ;
        RECT 1602.020 2482.860 1602.340 2483.180 ;
        RECT 1603.860 2477.420 1604.180 2477.740 ;
        RECT 1599.260 2476.060 1599.580 2476.380 ;
        RECT 1601.100 2474.700 1601.420 2475.020 ;
        RECT 1602.940 2472.660 1603.260 2472.980 ;
        RECT 1599.260 2468.580 1599.580 2468.900 ;
        RECT 1602.020 2467.220 1602.340 2467.540 ;
        RECT 1600.180 2463.140 1600.500 2463.460 ;
        RECT 1602.940 2461.100 1603.260 2461.420 ;
        RECT 1599.260 2455.660 1599.580 2455.980 ;
        RECT 1602.940 2454.300 1603.260 2454.620 ;
        RECT 1601.100 2451.580 1601.420 2451.900 ;
        RECT 1601.100 2448.860 1601.420 2449.180 ;
        RECT 1603.860 2442.060 1604.180 2442.380 ;
        RECT 1599.260 2439.340 1599.580 2439.660 ;
        RECT 1601.100 2439.340 1601.420 2439.660 ;
        RECT 1601.100 2436.620 1601.420 2436.940 ;
        RECT 1599.260 2433.220 1599.580 2433.540 ;
        RECT 1602.020 2430.500 1602.340 2430.820 ;
        RECT 1599.260 2427.780 1599.580 2428.100 ;
        RECT 1602.940 2424.380 1603.260 2424.700 ;
        RECT 1601.100 2422.340 1601.420 2422.660 ;
        RECT 1602.020 2420.300 1602.340 2420.620 ;
        RECT 1599.260 2414.860 1599.580 2415.180 ;
        RECT 1602.940 2412.820 1603.260 2413.140 ;
        RECT 1601.100 2410.100 1601.420 2410.420 ;
        RECT 1602.020 2407.380 1602.340 2407.700 ;
        RECT 1602.940 2401.260 1603.260 2401.580 ;
        RECT 1599.260 2398.540 1599.580 2398.860 ;
        RECT 1601.100 2398.540 1601.420 2398.860 ;
        RECT 1602.940 2395.140 1603.260 2395.460 ;
        RECT 1602.940 2389.700 1603.260 2390.020 ;
        RECT 1601.100 2383.580 1601.420 2383.900 ;
        RECT 1602.020 2383.580 1602.340 2383.900 ;
        RECT 1599.260 2378.820 1599.580 2379.140 ;
        RECT 1603.860 2378.820 1604.180 2379.140 ;
        RECT 1602.940 2378.140 1603.260 2378.460 ;
        RECT 1601.100 2372.020 1601.420 2372.340 ;
        RECT 1603.860 2372.020 1604.180 2372.340 ;
        RECT 1601.100 2365.900 1601.420 2366.220 ;
        RECT 1602.940 2365.900 1603.260 2366.220 ;
        RECT 1601.100 2361.140 1601.420 2361.460 ;
        RECT 1602.020 2360.460 1602.340 2360.780 ;
        RECT 1602.940 2355.020 1603.260 2355.340 ;
        RECT 1602.020 2354.340 1602.340 2354.660 ;
        RECT 1602.020 2350.260 1602.340 2350.580 ;
        RECT 1601.100 2348.900 1601.420 2349.220 ;
        RECT 1599.260 2345.500 1599.580 2345.820 ;
        RECT 1602.940 2344.140 1603.260 2344.460 ;
        RECT 1601.100 2342.780 1601.420 2343.100 ;
        RECT 1602.020 2338.020 1602.340 2338.340 ;
        RECT 1601.100 2325.780 1601.420 2326.100 ;
        RECT 1602.020 2325.780 1602.340 2326.100 ;
        RECT 2043.620 2202.460 2044.630 2203.980 ;
        RECT 2050.440 2200.240 2052.050 2201.760 ;
        RECT 1383.060 2023.860 1383.380 2024.180 ;
        RECT 1601.100 1959.940 1601.420 1960.260 ;
        RECT 1601.100 1949.060 1601.420 1949.380 ;
        RECT 1601.100 1944.980 1601.420 1945.300 ;
        RECT 1601.100 1937.500 1601.420 1937.820 ;
        RECT 1599.260 1932.060 1599.580 1932.380 ;
        RECT 1601.100 1931.380 1601.420 1931.700 ;
        RECT 1602.940 1923.900 1603.260 1924.220 ;
        RECT 1599.260 1918.460 1599.580 1918.780 ;
        RECT 1603.860 1917.780 1604.180 1918.100 ;
        RECT 1601.100 1915.740 1601.420 1916.060 ;
        RECT 1603.860 1912.340 1604.180 1912.660 ;
        RECT 1602.940 1906.220 1603.260 1906.540 ;
        RECT 1602.020 1904.180 1602.340 1904.500 ;
        RECT 1603.860 1900.780 1604.180 1901.100 ;
        RECT 1601.100 1898.060 1601.420 1898.380 ;
        RECT 1599.260 1897.380 1599.580 1897.700 ;
        RECT 1602.020 1894.660 1602.340 1894.980 ;
        RECT 1602.940 1891.940 1603.260 1892.260 ;
        RECT 1603.860 1888.540 1604.180 1888.860 ;
        RECT 1600.180 1883.100 1600.500 1883.420 ;
        RECT 1601.100 1880.380 1601.420 1880.700 ;
        RECT 1601.100 1876.980 1601.420 1877.300 ;
        RECT 1599.260 1875.620 1599.580 1875.940 ;
        RECT 1602.940 1871.540 1603.260 1871.860 ;
        RECT 1600.180 1868.820 1600.500 1869.140 ;
        RECT 1600.180 1865.420 1600.500 1865.740 ;
        RECT 1599.260 1863.380 1599.580 1863.700 ;
        RECT 1602.020 1862.700 1602.340 1863.020 ;
        RECT 1602.940 1861.340 1603.260 1861.660 ;
        RECT 1601.100 1857.260 1601.420 1857.580 ;
        RECT 1603.860 1855.900 1604.180 1856.220 ;
        RECT 1602.020 1848.420 1602.340 1848.740 ;
        RECT 1602.020 1845.700 1602.340 1846.020 ;
        RECT 1599.260 1842.300 1599.580 1842.620 ;
        RECT 1603.860 1842.300 1604.180 1842.620 ;
        RECT 1601.100 1839.580 1601.420 1839.900 ;
        RECT 1598.340 1836.180 1598.660 1836.500 ;
        RECT 1603.860 1836.180 1604.180 1836.500 ;
        RECT 1602.940 1830.740 1603.260 1831.060 ;
        RECT 1600.180 1828.020 1600.500 1828.340 ;
        RECT 1601.100 1824.620 1601.420 1824.940 ;
        RECT 1602.020 1821.900 1602.340 1822.220 ;
        RECT 1600.180 1818.500 1600.500 1818.820 ;
        RECT 1597.420 1817.140 1597.740 1817.460 ;
        RECT 1600.180 1813.060 1600.500 1813.380 ;
        RECT 1602.020 1810.340 1602.340 1810.660 ;
        RECT 1599.260 1806.940 1599.580 1807.260 ;
        RECT 1601.100 1806.940 1601.420 1807.260 ;
        RECT 1601.100 1804.900 1601.420 1805.220 ;
        RECT 1601.100 1801.500 1601.420 1801.820 ;
        RECT 1602.020 1798.780 1602.340 1799.100 ;
        RECT 1602.020 1792.660 1602.340 1792.980 ;
        RECT 1601.100 1789.260 1601.420 1789.580 ;
        RECT 1369.260 1785.860 1369.580 1786.180 ;
        RECT 1602.940 1785.180 1603.260 1785.500 ;
        RECT 1601.100 1783.820 1601.420 1784.140 ;
        RECT 1602.940 1779.740 1603.260 1780.060 ;
        RECT 1601.100 1777.700 1601.420 1778.020 ;
        RECT 1603.860 1772.940 1604.180 1773.260 ;
        RECT 1601.100 1772.260 1601.420 1772.580 ;
        RECT 1599.260 1766.820 1599.580 1767.140 ;
        RECT 1601.100 1766.140 1601.420 1766.460 ;
        RECT 1603.860 1766.140 1604.180 1766.460 ;
        RECT 1601.100 1762.740 1601.420 1763.060 ;
        RECT 1602.020 1762.060 1602.340 1762.380 ;
        RECT 1602.940 1755.940 1603.260 1756.260 ;
        RECT 1602.020 1754.580 1602.340 1754.900 ;
        RECT 1603.860 1750.500 1604.180 1750.820 ;
        RECT 1601.100 1748.460 1601.420 1748.780 ;
        RECT 1601.100 1743.020 1601.420 1743.340 ;
        RECT 1601.100 1731.460 1601.420 1731.780 ;
        RECT 2043.620 1602.460 2044.630 1603.980 ;
        RECT 2050.440 1600.240 2052.050 1601.760 ;
      LAYER met4 ;
        RECT 494.025 3301.635 494.325 3306.235 ;
        RECT 500.265 3301.635 500.565 3306.235 ;
        RECT 506.505 3301.635 506.805 3306.235 ;
        RECT 512.745 3301.635 513.045 3306.235 ;
        RECT 518.985 3301.635 519.285 3306.235 ;
        RECT 525.225 3301.635 525.525 3306.235 ;
        RECT 531.465 3301.635 531.765 3306.235 ;
        RECT 537.705 3301.635 538.005 3306.235 ;
        RECT 550.185 3301.635 550.485 3306.235 ;
        RECT 556.425 3301.635 556.725 3306.235 ;
        RECT 568.905 3301.635 569.205 3306.235 ;
        RECT 575.145 3301.635 575.445 3306.235 ;
        RECT 587.625 3301.635 587.925 3306.235 ;
        RECT 593.865 3301.635 594.165 3306.235 ;
        RECT 606.345 3301.635 606.645 3306.235 ;
        RECT 612.585 3301.635 612.885 3306.235 ;
        RECT 618.825 3301.635 619.125 3306.235 ;
        RECT 625.065 3301.635 625.365 3306.235 ;
        RECT 631.305 3301.635 631.605 3306.235 ;
        RECT 637.545 3301.635 637.845 3306.235 ;
        RECT 643.785 3301.635 644.085 3306.235 ;
        RECT 650.025 3301.635 650.325 3306.235 ;
        RECT 656.265 3301.635 656.565 3306.235 ;
        RECT 662.505 3301.635 662.805 3306.235 ;
        RECT 668.745 3301.635 669.045 3306.235 ;
        RECT 674.985 3301.635 675.285 3306.235 ;
        RECT 681.225 3301.635 681.525 3306.235 ;
        RECT 687.465 3301.635 687.765 3306.235 ;
        RECT 767.865 3301.635 768.165 3306.235 ;
      LAYER met4 ;
        RECT 405.000 2855.000 781.480 3301.235 ;
      LAYER met4 ;
        RECT 434.010 2851.050 434.310 2854.600 ;
        RECT 439.850 2851.050 440.150 2854.600 ;
        RECT 445.690 2851.050 445.990 2854.600 ;
        RECT 451.530 2851.050 451.830 2854.600 ;
        RECT 432.710 2850.750 434.310 2851.050 ;
        RECT 432.710 2842.905 433.010 2850.750 ;
        RECT 434.010 2850.000 434.310 2850.750 ;
        RECT 437.310 2850.750 440.150 2851.050 ;
        RECT 432.695 2842.575 433.025 2842.905 ;
        RECT 437.310 2836.785 437.610 2850.750 ;
        RECT 439.850 2850.000 440.150 2850.750 ;
        RECT 442.830 2850.750 445.990 2851.050 ;
        RECT 442.830 2837.465 443.130 2850.750 ;
        RECT 445.690 2850.000 445.990 2850.750 ;
        RECT 450.190 2850.750 451.830 2851.050 ;
        RECT 442.815 2837.135 443.145 2837.465 ;
        RECT 450.190 2836.785 450.490 2850.750 ;
        RECT 451.530 2850.000 451.830 2850.750 ;
        RECT 457.370 2851.050 457.670 2854.600 ;
        RECT 463.830 2851.050 464.130 2854.600 ;
        RECT 469.670 2851.050 469.970 2854.600 ;
        RECT 457.370 2850.000 457.850 2851.050 ;
        RECT 463.830 2850.750 467.050 2851.050 ;
        RECT 463.830 2850.000 464.130 2850.750 ;
        RECT 457.550 2838.825 457.850 2850.000 ;
        RECT 457.535 2838.495 457.865 2838.825 ;
        RECT 437.295 2836.455 437.625 2836.785 ;
        RECT 450.175 2836.455 450.505 2836.785 ;
        RECT 466.750 2836.105 467.050 2850.750 ;
        RECT 469.670 2850.750 471.650 2851.050 ;
        RECT 469.670 2850.000 469.970 2850.750 ;
        RECT 471.350 2836.105 471.650 2850.750 ;
        RECT 475.510 2847.650 475.810 2854.600 ;
        RECT 480.730 2851.050 481.030 2854.600 ;
        RECT 480.550 2850.000 481.030 2851.050 ;
        RECT 481.350 2851.050 481.650 2854.600 ;
        RECT 487.190 2851.050 487.490 2854.600 ;
        RECT 493.030 2851.050 493.330 2854.600 ;
        RECT 498.870 2851.050 499.170 2854.600 ;
        RECT 481.350 2850.000 481.770 2851.050 ;
        RECT 487.190 2850.750 489.130 2851.050 ;
        RECT 487.190 2850.000 487.490 2850.750 ;
        RECT 475.510 2847.350 476.250 2847.650 ;
        RECT 475.950 2842.225 476.250 2847.350 ;
        RECT 475.935 2841.895 476.265 2842.225 ;
        RECT 480.550 2841.545 480.850 2850.000 ;
        RECT 480.535 2841.215 480.865 2841.545 ;
        RECT 481.470 2836.105 481.770 2850.000 ;
        RECT 488.830 2838.825 489.130 2850.750 ;
        RECT 493.030 2850.750 494.650 2851.050 ;
        RECT 493.030 2850.000 493.330 2850.750 ;
        RECT 488.815 2838.495 489.145 2838.825 ;
        RECT 494.350 2836.105 494.650 2850.750 ;
        RECT 498.870 2850.750 502.010 2851.050 ;
        RECT 498.870 2850.000 499.170 2850.750 ;
        RECT 501.710 2838.825 502.010 2850.750 ;
        RECT 504.090 2847.650 504.390 2854.600 ;
        RECT 504.710 2851.050 505.010 2854.600 ;
        RECT 516.390 2852.750 516.690 2854.600 ;
        RECT 516.390 2852.450 517.650 2852.750 ;
        RECT 504.710 2850.750 507.530 2851.050 ;
        RECT 504.710 2850.000 505.010 2850.750 ;
        RECT 504.090 2847.350 504.770 2847.650 ;
        RECT 504.470 2841.545 504.770 2847.350 ;
        RECT 507.230 2842.905 507.530 2850.750 ;
        RECT 516.390 2850.000 516.690 2852.450 ;
        RECT 517.350 2851.745 517.650 2852.450 ;
        RECT 517.335 2851.415 517.665 2851.745 ;
        RECT 522.230 2851.050 522.530 2854.600 ;
        RECT 527.450 2851.050 527.750 2854.600 ;
        RECT 522.230 2850.750 524.090 2851.050 ;
        RECT 522.230 2850.000 522.530 2850.750 ;
        RECT 523.790 2842.905 524.090 2850.750 ;
        RECT 526.550 2850.750 527.750 2851.050 ;
        RECT 526.550 2842.905 526.850 2850.750 ;
        RECT 527.450 2850.000 527.750 2850.750 ;
        RECT 528.070 2851.050 528.370 2854.600 ;
        RECT 528.070 2850.750 529.610 2851.050 ;
        RECT 528.070 2850.000 528.370 2850.750 ;
        RECT 529.310 2842.905 529.610 2850.750 ;
        RECT 533.910 2842.905 534.210 2854.600 ;
        RECT 539.750 2851.050 540.050 2854.600 ;
        RECT 550.810 2852.750 551.110 2854.600 ;
        RECT 549.550 2852.450 551.110 2852.750 ;
        RECT 539.750 2850.750 543.410 2851.050 ;
        RECT 539.750 2850.000 540.050 2850.750 ;
        RECT 543.110 2842.905 543.410 2850.750 ;
        RECT 507.215 2842.575 507.545 2842.905 ;
        RECT 523.775 2842.575 524.105 2842.905 ;
        RECT 526.535 2842.575 526.865 2842.905 ;
        RECT 529.295 2842.575 529.625 2842.905 ;
        RECT 533.895 2842.575 534.225 2842.905 ;
        RECT 543.095 2842.575 543.425 2842.905 ;
        RECT 549.550 2842.225 549.850 2852.450 ;
        RECT 550.810 2850.000 551.110 2852.450 ;
        RECT 551.430 2847.650 551.730 2854.600 ;
        RECT 551.390 2847.350 551.730 2847.650 ;
        RECT 557.270 2847.650 557.570 2854.600 ;
        RECT 568.950 2848.345 569.250 2854.600 ;
        RECT 568.935 2848.015 569.265 2848.345 ;
        RECT 574.170 2847.650 574.470 2854.600 ;
        RECT 557.270 2847.350 558.130 2847.650 ;
        RECT 549.535 2841.895 549.865 2842.225 ;
        RECT 504.455 2841.215 504.785 2841.545 ;
        RECT 551.390 2838.825 551.690 2847.350 ;
        RECT 557.830 2842.905 558.130 2847.350 ;
        RECT 573.470 2847.350 574.470 2847.650 ;
        RECT 574.790 2847.650 575.090 2854.600 ;
        RECT 586.470 2847.650 586.770 2854.600 ;
        RECT 592.310 2848.345 592.610 2854.600 ;
        RECT 597.530 2851.050 597.830 2854.600 ;
        RECT 597.390 2850.000 597.830 2851.050 ;
        RECT 592.295 2848.015 592.625 2848.345 ;
        RECT 574.790 2847.350 575.610 2847.650 ;
        RECT 573.470 2843.585 573.770 2847.350 ;
        RECT 575.310 2843.585 575.610 2847.350 ;
        RECT 586.350 2847.350 586.770 2847.650 ;
        RECT 573.455 2843.255 573.785 2843.585 ;
        RECT 575.295 2843.255 575.625 2843.585 ;
        RECT 557.815 2842.575 558.145 2842.905 ;
        RECT 501.695 2838.495 502.025 2838.825 ;
        RECT 551.375 2838.495 551.705 2838.825 ;
        RECT 466.735 2835.775 467.065 2836.105 ;
        RECT 471.335 2835.775 471.665 2836.105 ;
        RECT 481.455 2835.775 481.785 2836.105 ;
        RECT 494.335 2835.775 494.665 2836.105 ;
        RECT 586.350 2832.705 586.650 2847.350 ;
        RECT 597.390 2845.625 597.690 2850.000 ;
        RECT 603.990 2849.010 604.290 2854.600 ;
        RECT 609.830 2851.050 610.130 2854.600 ;
        RECT 615.670 2851.050 615.970 2854.600 ;
        RECT 609.830 2850.750 613.330 2851.050 ;
        RECT 609.830 2850.000 610.130 2850.750 ;
        RECT 603.990 2848.710 605.050 2849.010 ;
        RECT 604.750 2845.625 605.050 2848.710 ;
        RECT 597.375 2845.295 597.705 2845.625 ;
        RECT 604.735 2845.295 605.065 2845.625 ;
        RECT 613.030 2844.265 613.330 2850.750 ;
        RECT 615.670 2850.750 618.850 2851.050 ;
        RECT 615.670 2850.000 615.970 2850.750 ;
        RECT 613.015 2843.935 613.345 2844.265 ;
        RECT 618.550 2841.545 618.850 2850.750 ;
        RECT 620.890 2847.650 621.190 2854.600 ;
        RECT 621.510 2851.050 621.810 2854.600 ;
        RECT 621.510 2850.750 624.370 2851.050 ;
        RECT 621.510 2850.000 621.810 2850.750 ;
        RECT 620.890 2847.350 621.610 2847.650 ;
        RECT 621.310 2841.545 621.610 2847.350 ;
        RECT 618.535 2841.215 618.865 2841.545 ;
        RECT 621.295 2841.215 621.625 2841.545 ;
        RECT 621.310 2836.785 621.610 2841.215 ;
        RECT 621.295 2836.455 621.625 2836.785 ;
        RECT 624.070 2836.105 624.370 2850.750 ;
        RECT 627.350 2847.650 627.650 2854.600 ;
        RECT 633.190 2851.050 633.490 2854.600 ;
        RECT 639.030 2851.050 639.330 2854.600 ;
        RECT 644.250 2851.050 644.550 2854.600 ;
        RECT 633.190 2850.000 633.570 2851.050 ;
        RECT 639.030 2850.750 640.930 2851.050 ;
        RECT 639.030 2850.000 639.330 2850.750 ;
        RECT 626.830 2847.350 627.650 2847.650 ;
        RECT 626.830 2841.545 627.130 2847.350 ;
        RECT 626.815 2841.215 627.145 2841.545 ;
        RECT 633.270 2836.105 633.570 2850.000 ;
        RECT 640.630 2836.105 640.930 2850.750 ;
        RECT 642.470 2850.750 644.550 2851.050 ;
        RECT 642.470 2842.905 642.770 2850.750 ;
        RECT 644.250 2850.000 644.550 2850.750 ;
        RECT 644.870 2851.050 645.170 2854.600 ;
        RECT 782.470 2853.670 784.070 3294.680 ;
        RECT 784.690 2854.060 786.310 3302.140 ;
        RECT 1044.025 3301.635 1044.325 3306.235 ;
        RECT 1056.505 3301.635 1056.805 3306.235 ;
        RECT 1062.745 3301.635 1063.045 3306.235 ;
        RECT 1068.985 3301.635 1069.285 3306.235 ;
        RECT 1075.225 3301.635 1075.525 3306.235 ;
        RECT 1081.465 3301.635 1081.765 3306.235 ;
        RECT 1087.705 3301.635 1088.005 3306.235 ;
        RECT 1093.945 3301.635 1094.245 3306.235 ;
        RECT 1100.185 3301.635 1100.485 3306.235 ;
        RECT 1106.425 3301.635 1106.725 3306.235 ;
        RECT 1112.665 3301.635 1112.965 3306.235 ;
        RECT 1118.905 3301.635 1119.205 3306.235 ;
        RECT 1125.145 3301.635 1125.445 3306.235 ;
        RECT 1131.385 3301.635 1131.685 3306.235 ;
        RECT 1137.625 3301.635 1137.925 3306.235 ;
        RECT 1143.865 3301.635 1144.165 3306.235 ;
        RECT 1150.105 3301.635 1150.405 3306.235 ;
        RECT 1156.345 3301.635 1156.645 3306.235 ;
        RECT 1162.585 3301.635 1162.885 3306.235 ;
        RECT 1168.825 3301.635 1169.125 3306.235 ;
        RECT 1181.305 3301.635 1181.605 3306.235 ;
        RECT 1187.545 3301.635 1187.845 3306.235 ;
        RECT 1200.025 3301.635 1200.325 3306.235 ;
        RECT 1206.265 3301.635 1206.565 3306.235 ;
        RECT 1218.745 3301.635 1219.045 3306.235 ;
        RECT 1224.985 3301.635 1225.285 3306.235 ;
        RECT 1231.225 3301.635 1231.525 3306.235 ;
        RECT 1237.465 3301.635 1237.765 3306.235 ;
        RECT 1292.890 3301.635 1293.190 3306.235 ;
      LAYER met4 ;
        RECT 955.000 2855.000 1331.480 3301.235 ;
      LAYER met4 ;
        RECT 984.010 2851.050 984.310 2854.600 ;
        RECT 989.850 2851.050 990.150 2854.600 ;
        RECT 1001.530 2851.050 1001.830 2854.600 ;
        RECT 644.870 2850.750 648.290 2851.050 ;
        RECT 644.870 2850.000 645.170 2850.750 ;
        RECT 642.455 2842.575 642.785 2842.905 ;
        RECT 647.990 2841.545 648.290 2850.750 ;
        RECT 981.030 2850.750 984.310 2851.050 ;
        RECT 981.030 2842.905 981.330 2850.750 ;
        RECT 984.010 2850.000 984.310 2850.750 ;
        RECT 988.390 2850.750 990.150 2851.050 ;
        RECT 988.390 2842.905 988.690 2850.750 ;
        RECT 989.850 2850.000 990.150 2850.750 ;
        RECT 1001.270 2850.000 1001.830 2851.050 ;
        RECT 981.015 2842.575 981.345 2842.905 ;
        RECT 988.375 2842.575 988.705 2842.905 ;
        RECT 647.975 2841.215 648.305 2841.545 ;
        RECT 1001.270 2840.865 1001.570 2850.000 ;
        RECT 1007.370 2847.650 1007.670 2854.600 ;
        RECT 1019.050 2851.050 1019.350 2854.600 ;
        RECT 1018.750 2850.000 1019.350 2851.050 ;
        RECT 1007.370 2847.350 1008.010 2847.650 ;
        RECT 1001.255 2840.535 1001.585 2840.865 ;
        RECT 1007.710 2840.185 1008.010 2847.350 ;
        RECT 1018.750 2842.225 1019.050 2850.000 ;
        RECT 1019.670 2842.905 1019.970 2854.600 ;
        RECT 1024.890 2851.050 1025.190 2854.600 ;
        RECT 1024.270 2850.750 1025.190 2851.050 ;
        RECT 1024.270 2842.905 1024.570 2850.750 ;
        RECT 1024.890 2850.000 1025.190 2850.750 ;
        RECT 1025.510 2851.050 1025.810 2854.600 ;
        RECT 1037.190 2851.050 1037.490 2854.600 ;
        RECT 1042.410 2851.050 1042.710 2854.600 ;
        RECT 1025.510 2850.750 1027.330 2851.050 ;
        RECT 1025.510 2850.000 1025.810 2850.750 ;
        RECT 1027.030 2842.905 1027.330 2850.750 ;
        RECT 1037.190 2850.750 1040.210 2851.050 ;
        RECT 1037.190 2850.000 1037.490 2850.750 ;
        RECT 1019.655 2842.575 1019.985 2842.905 ;
        RECT 1024.255 2842.575 1024.585 2842.905 ;
        RECT 1027.015 2842.575 1027.345 2842.905 ;
        RECT 1018.735 2841.895 1019.065 2842.225 ;
        RECT 1007.695 2839.855 1008.025 2840.185 ;
        RECT 1039.910 2836.105 1040.210 2850.750 ;
        RECT 1041.750 2850.750 1042.710 2851.050 ;
        RECT 1041.750 2836.785 1042.050 2850.750 ;
        RECT 1042.410 2850.000 1042.710 2850.750 ;
        RECT 1043.030 2851.050 1043.330 2854.600 ;
        RECT 1043.030 2850.750 1046.650 2851.050 ;
        RECT 1043.030 2850.000 1043.330 2850.750 ;
        RECT 1041.735 2836.455 1042.065 2836.785 ;
        RECT 1046.350 2836.105 1046.650 2850.750 ;
        RECT 1054.710 2847.650 1055.010 2854.600 ;
        RECT 1060.550 2851.050 1060.850 2854.600 ;
        RECT 1065.770 2851.050 1066.070 2854.600 ;
        RECT 1060.550 2850.750 1062.290 2851.050 ;
        RECT 1060.550 2850.000 1060.850 2850.750 ;
        RECT 1054.630 2847.350 1055.010 2847.650 ;
        RECT 1054.630 2836.105 1054.930 2847.350 ;
        RECT 1061.990 2836.105 1062.290 2850.750 ;
        RECT 1065.670 2850.000 1066.070 2851.050 ;
        RECT 1066.390 2851.050 1066.690 2854.600 ;
        RECT 1071.610 2852.750 1071.910 2854.600 ;
        RECT 1070.270 2852.450 1071.910 2852.750 ;
        RECT 1066.390 2850.750 1067.810 2851.050 ;
        RECT 1066.390 2850.000 1066.690 2850.750 ;
        RECT 1065.670 2842.905 1065.970 2850.000 ;
        RECT 1065.655 2842.575 1065.985 2842.905 ;
        RECT 1067.510 2836.105 1067.810 2850.750 ;
        RECT 1070.270 2842.905 1070.570 2852.450 ;
        RECT 1071.610 2850.000 1071.910 2852.450 ;
        RECT 1072.230 2851.050 1072.530 2854.600 ;
        RECT 1078.070 2851.050 1078.370 2854.600 ;
        RECT 1072.230 2850.750 1074.250 2851.050 ;
        RECT 1072.230 2850.000 1072.530 2850.750 ;
        RECT 1070.255 2842.575 1070.585 2842.905 ;
        RECT 1073.950 2836.105 1074.250 2850.750 ;
        RECT 1078.070 2850.750 1081.610 2851.050 ;
        RECT 1078.070 2850.000 1078.370 2850.750 ;
        RECT 1081.310 2836.105 1081.610 2850.750 ;
        RECT 1089.130 2848.345 1089.430 2854.600 ;
        RECT 1089.115 2848.015 1089.445 2848.345 ;
        RECT 1089.750 2847.650 1090.050 2854.600 ;
        RECT 1089.590 2847.350 1090.050 2847.650 ;
        RECT 1095.590 2847.650 1095.890 2854.600 ;
        RECT 1101.430 2851.050 1101.730 2854.600 ;
        RECT 1103.375 2851.050 1103.705 2851.065 ;
        RECT 1101.430 2850.750 1103.705 2851.050 ;
        RECT 1101.430 2850.000 1101.730 2850.750 ;
        RECT 1103.375 2850.735 1103.705 2850.750 ;
        RECT 1107.270 2851.050 1107.570 2854.600 ;
        RECT 1112.490 2851.050 1112.790 2854.600 ;
        RECT 1107.270 2850.750 1110.130 2851.050 ;
        RECT 1107.270 2850.000 1107.570 2850.750 ;
        RECT 1095.590 2847.350 1096.330 2847.650 ;
        RECT 1089.590 2836.105 1089.890 2847.350 ;
        RECT 1096.030 2836.105 1096.330 2847.350 ;
        RECT 1109.830 2836.105 1110.130 2850.750 ;
        RECT 1111.670 2850.750 1112.790 2851.050 ;
        RECT 1111.670 2842.905 1111.970 2850.750 ;
        RECT 1112.490 2850.000 1112.790 2850.750 ;
        RECT 1113.110 2851.050 1113.410 2854.600 ;
        RECT 1118.330 2851.050 1118.630 2854.600 ;
        RECT 1113.110 2850.750 1116.570 2851.050 ;
        RECT 1113.110 2850.000 1113.410 2850.750 ;
        RECT 1111.655 2842.575 1111.985 2842.905 ;
        RECT 1116.270 2836.105 1116.570 2850.750 ;
        RECT 1118.110 2850.000 1118.630 2851.050 ;
        RECT 1118.950 2851.050 1119.250 2854.600 ;
        RECT 1124.790 2851.050 1125.090 2854.600 ;
        RECT 1118.950 2850.000 1119.330 2851.050 ;
        RECT 1124.790 2850.750 1128.530 2851.050 ;
        RECT 1124.790 2850.000 1125.090 2850.750 ;
        RECT 1118.110 2842.905 1118.410 2850.000 ;
        RECT 1118.095 2842.575 1118.425 2842.905 ;
        RECT 1119.030 2836.105 1119.330 2850.000 ;
        RECT 1128.230 2842.225 1128.530 2850.750 ;
        RECT 1130.630 2847.650 1130.930 2854.600 ;
        RECT 1135.850 2851.050 1136.150 2854.600 ;
        RECT 1135.590 2850.000 1136.150 2851.050 ;
        RECT 1136.470 2851.050 1136.770 2854.600 ;
        RECT 1142.310 2851.050 1142.610 2854.600 ;
        RECT 1148.150 2851.050 1148.450 2854.600 ;
        RECT 1136.470 2850.000 1136.810 2851.050 ;
        RECT 1142.310 2850.750 1144.170 2851.050 ;
        RECT 1142.310 2850.000 1142.610 2850.750 ;
        RECT 1130.630 2847.350 1131.290 2847.650 ;
        RECT 1130.990 2842.905 1131.290 2847.350 ;
        RECT 1135.590 2842.905 1135.890 2850.000 ;
        RECT 1136.510 2842.905 1136.810 2850.000 ;
        RECT 1143.870 2842.905 1144.170 2850.750 ;
        RECT 1148.150 2850.750 1151.530 2851.050 ;
        RECT 1148.150 2850.000 1148.450 2850.750 ;
        RECT 1151.230 2842.905 1151.530 2850.750 ;
        RECT 1153.990 2842.905 1154.290 2854.600 ;
        RECT 1159.210 2847.650 1159.510 2854.600 ;
        RECT 1159.830 2851.050 1160.130 2854.600 ;
        RECT 1165.050 2851.050 1165.350 2854.600 ;
        RECT 1159.830 2850.750 1163.490 2851.050 ;
        RECT 1159.830 2850.000 1160.130 2850.750 ;
        RECT 1159.210 2847.350 1159.810 2847.650 ;
        RECT 1130.975 2842.575 1131.305 2842.905 ;
        RECT 1135.575 2842.575 1135.905 2842.905 ;
        RECT 1136.495 2842.575 1136.825 2842.905 ;
        RECT 1143.855 2842.575 1144.185 2842.905 ;
        RECT 1151.215 2842.575 1151.545 2842.905 ;
        RECT 1153.975 2842.575 1154.305 2842.905 ;
        RECT 1128.215 2841.895 1128.545 2842.225 ;
        RECT 1159.510 2840.185 1159.810 2847.350 ;
        RECT 1163.190 2842.225 1163.490 2850.750 ;
        RECT 1164.110 2850.750 1165.350 2851.050 ;
        RECT 1163.175 2841.895 1163.505 2842.225 ;
        RECT 1164.110 2840.865 1164.410 2850.750 ;
        RECT 1165.050 2850.000 1165.350 2850.750 ;
        RECT 1165.670 2847.650 1165.970 2854.600 ;
        RECT 1171.510 2851.050 1171.810 2854.600 ;
        RECT 1177.350 2851.050 1177.650 2854.600 ;
        RECT 1182.570 2851.050 1182.870 2854.600 ;
        RECT 1171.510 2850.750 1172.690 2851.050 ;
        RECT 1171.510 2850.000 1171.810 2850.750 ;
        RECT 1165.030 2847.350 1165.970 2847.650 ;
        RECT 1165.030 2842.905 1165.330 2847.350 ;
        RECT 1172.390 2842.905 1172.690 2850.750 ;
        RECT 1177.350 2850.750 1179.130 2851.050 ;
        RECT 1177.350 2850.000 1177.650 2850.750 ;
        RECT 1178.830 2842.905 1179.130 2850.750 ;
        RECT 1180.670 2850.750 1182.870 2851.050 ;
        RECT 1165.015 2842.575 1165.345 2842.905 ;
        RECT 1172.375 2842.575 1172.705 2842.905 ;
        RECT 1178.815 2842.575 1179.145 2842.905 ;
        RECT 1180.670 2840.865 1180.970 2850.750 ;
        RECT 1182.570 2850.000 1182.870 2850.750 ;
        RECT 1183.190 2851.050 1183.490 2854.600 ;
        RECT 1189.030 2851.050 1189.330 2854.600 ;
        RECT 1332.470 2853.670 1334.070 3294.680 ;
        RECT 1334.690 2854.060 1336.310 3302.140 ;
        RECT 1183.190 2850.750 1186.490 2851.050 ;
        RECT 1183.190 2850.000 1183.490 2850.750 ;
        RECT 1186.190 2842.905 1186.490 2850.750 ;
        RECT 1189.030 2850.750 1191.090 2851.050 ;
        RECT 1189.030 2850.000 1189.330 2850.750 ;
        RECT 1190.790 2842.905 1191.090 2850.750 ;
        RECT 1186.175 2842.575 1186.505 2842.905 ;
        RECT 1190.775 2842.575 1191.105 2842.905 ;
        RECT 1164.095 2840.535 1164.425 2840.865 ;
        RECT 1180.655 2840.535 1180.985 2840.865 ;
        RECT 1159.495 2839.855 1159.825 2840.185 ;
        RECT 624.055 2835.775 624.385 2836.105 ;
        RECT 633.255 2835.775 633.585 2836.105 ;
        RECT 640.615 2835.775 640.945 2836.105 ;
        RECT 1039.895 2835.775 1040.225 2836.105 ;
        RECT 1046.335 2835.775 1046.665 2836.105 ;
        RECT 1054.615 2835.775 1054.945 2836.105 ;
        RECT 1061.975 2835.775 1062.305 2836.105 ;
        RECT 1067.495 2835.775 1067.825 2836.105 ;
        RECT 1073.935 2835.775 1074.265 2836.105 ;
        RECT 1081.295 2835.775 1081.625 2836.105 ;
        RECT 1089.575 2835.775 1089.905 2836.105 ;
        RECT 1096.015 2835.775 1096.345 2836.105 ;
        RECT 1109.815 2835.775 1110.145 2836.105 ;
        RECT 1116.255 2835.775 1116.585 2836.105 ;
        RECT 1119.015 2835.775 1119.345 2836.105 ;
        RECT 586.335 2832.375 586.665 2832.705 ;
        RECT 370.970 1610.640 372.570 2598.480 ;
      LAYER met4 ;
        RECT 373.225 1610.640 382.020 2598.480 ;
        RECT 385.020 1610.640 400.020 2598.480 ;
        RECT 403.020 1610.640 418.020 2598.480 ;
        RECT 421.020 1610.640 447.370 2598.480 ;
      LAYER met4 ;
        RECT 447.770 1610.640 449.370 2598.480 ;
      LAYER met4 ;
        RECT 449.770 1610.640 454.020 2598.480 ;
        RECT 457.020 1610.640 472.020 2598.480 ;
        RECT 475.020 1610.640 490.020 2598.480 ;
        RECT 493.020 1610.640 508.020 2598.480 ;
        RECT 511.020 1610.640 544.020 2598.480 ;
        RECT 547.020 1610.640 562.020 2598.480 ;
        RECT 565.020 1610.640 580.020 2598.480 ;
        RECT 583.020 1610.640 598.020 2598.480 ;
        RECT 601.020 1610.640 634.020 2598.480 ;
        RECT 637.020 1610.640 652.020 2598.480 ;
        RECT 655.020 1610.640 670.020 2598.480 ;
        RECT 673.020 1610.640 688.020 2598.480 ;
        RECT 691.020 1610.640 724.020 2598.480 ;
        RECT 727.020 1610.640 742.020 2598.480 ;
        RECT 745.020 1610.640 760.020 2598.480 ;
        RECT 763.020 1610.640 778.020 2598.480 ;
        RECT 781.020 1610.640 814.020 2598.480 ;
        RECT 817.020 1610.640 832.020 2598.480 ;
        RECT 835.020 1610.640 850.020 2598.480 ;
        RECT 853.020 1610.640 868.020 2598.480 ;
        RECT 871.020 1610.640 904.020 2598.480 ;
        RECT 907.020 1610.640 922.020 2598.480 ;
        RECT 925.020 1610.640 940.020 2598.480 ;
        RECT 943.020 1610.640 958.020 2598.480 ;
        RECT 961.020 1610.640 994.020 2598.480 ;
        RECT 997.020 1610.640 1012.020 2598.480 ;
        RECT 1015.020 1610.640 1030.020 2598.480 ;
        RECT 1033.020 1610.640 1048.020 2598.480 ;
        RECT 1051.020 1610.640 1084.020 2598.480 ;
        RECT 1087.020 1610.640 1102.020 2598.480 ;
        RECT 1105.020 1610.640 1120.020 2598.480 ;
        RECT 1123.020 1610.640 1138.020 2598.480 ;
        RECT 1141.020 1610.640 1174.020 2598.480 ;
        RECT 1177.020 1610.640 1192.020 2598.480 ;
        RECT 1195.020 1610.640 1210.020 2598.480 ;
        RECT 1213.020 1610.640 1228.020 2598.480 ;
        RECT 1231.020 1610.640 1264.020 2598.480 ;
        RECT 1267.020 1610.640 1282.020 2598.480 ;
        RECT 1285.020 1610.640 1300.020 2598.480 ;
        RECT 1303.020 1610.640 1318.020 2598.480 ;
        RECT 1321.020 1610.640 1349.675 2598.480 ;
      LAYER met4 ;
        RECT 1369.255 2582.135 1369.585 2582.465 ;
        RECT 1369.270 1786.185 1369.570 2582.135 ;
        RECT 1601.095 2560.375 1601.425 2560.705 ;
        RECT 1601.110 2552.470 1601.410 2560.375 ;
        RECT 1600.000 2552.170 1604.600 2552.470 ;
        RECT 1600.000 2546.330 1604.600 2546.630 ;
        RECT 1600.190 2545.745 1600.490 2546.330 ;
        RECT 1600.175 2545.415 1600.505 2545.745 ;
        RECT 1600.000 2540.490 1604.600 2540.790 ;
        RECT 1600.190 2539.625 1600.490 2540.490 ;
        RECT 1600.175 2539.295 1600.505 2539.625 ;
        RECT 1602.015 2537.255 1602.345 2537.585 ;
        RECT 1602.030 2534.950 1602.330 2537.255 ;
        RECT 1600.000 2534.650 1604.600 2534.950 ;
        RECT 1599.255 2531.135 1599.585 2531.465 ;
        RECT 1601.095 2531.135 1601.425 2531.465 ;
        RECT 1599.270 2522.650 1599.570 2531.135 ;
        RECT 1601.110 2529.110 1601.410 2531.135 ;
        RECT 1600.000 2528.810 1604.600 2529.110 ;
        RECT 1603.855 2523.655 1604.185 2523.985 ;
        RECT 1603.870 2523.270 1604.170 2523.655 ;
        RECT 1600.000 2522.970 1604.600 2523.270 ;
        RECT 1599.270 2522.350 1604.600 2522.650 ;
        RECT 1383.055 2518.895 1383.385 2519.225 ;
        RECT 1599.255 2518.895 1599.585 2519.225 ;
        RECT 1383.070 2024.185 1383.370 2518.895 ;
        RECT 1599.270 2507.650 1599.570 2518.895 ;
        RECT 1602.935 2518.215 1603.265 2518.545 ;
        RECT 1602.950 2517.430 1603.250 2518.215 ;
        RECT 1600.000 2517.130 1604.600 2517.430 ;
        RECT 1600.000 2516.510 1604.600 2516.810 ;
        RECT 1601.110 2515.825 1601.410 2516.510 ;
        RECT 1601.095 2515.495 1601.425 2515.825 ;
        RECT 1602.015 2512.095 1602.345 2512.425 ;
        RECT 1602.030 2511.590 1602.330 2512.095 ;
        RECT 1600.000 2511.290 1604.600 2511.590 ;
        RECT 1600.000 2510.670 1604.600 2510.970 ;
        RECT 1600.190 2507.650 1600.490 2510.670 ;
        RECT 1599.270 2507.350 1600.490 2507.650 ;
        RECT 1603.855 2506.655 1604.185 2506.985 ;
        RECT 1603.870 2505.750 1604.170 2506.655 ;
        RECT 1600.000 2505.450 1604.600 2505.750 ;
        RECT 1599.255 2504.615 1599.585 2504.945 ;
        RECT 1600.000 2504.830 1604.600 2505.130 ;
        RECT 1599.270 2493.450 1599.570 2504.615 ;
        RECT 1600.190 2504.265 1600.490 2504.830 ;
        RECT 1600.175 2503.935 1600.505 2504.265 ;
        RECT 1602.935 2500.535 1603.265 2500.865 ;
        RECT 1602.950 2499.910 1603.250 2500.535 ;
        RECT 1600.000 2499.610 1604.600 2499.910 ;
        RECT 1600.000 2498.990 1604.600 2499.290 ;
        RECT 1601.110 2498.145 1601.410 2498.990 ;
        RECT 1601.095 2497.815 1601.425 2498.145 ;
        RECT 1603.855 2494.415 1604.185 2494.745 ;
        RECT 1603.870 2494.070 1604.170 2494.415 ;
        RECT 1600.000 2493.770 1604.600 2494.070 ;
        RECT 1599.270 2493.150 1604.600 2493.450 ;
        RECT 1599.255 2489.655 1599.585 2489.985 ;
        RECT 1599.270 2481.770 1599.570 2489.655 ;
        RECT 1601.095 2488.975 1601.425 2489.305 ;
        RECT 1601.110 2488.230 1601.410 2488.975 ;
        RECT 1600.000 2487.930 1604.600 2488.230 ;
        RECT 1600.000 2487.310 1604.600 2487.610 ;
        RECT 1601.110 2486.585 1601.410 2487.310 ;
        RECT 1601.095 2486.255 1601.425 2486.585 ;
        RECT 1602.015 2482.855 1602.345 2483.185 ;
        RECT 1602.030 2482.390 1602.330 2482.855 ;
        RECT 1600.000 2482.090 1604.600 2482.390 ;
        RECT 1599.270 2481.470 1604.600 2481.770 ;
        RECT 1603.855 2477.415 1604.185 2477.745 ;
        RECT 1603.870 2476.550 1604.170 2477.415 ;
        RECT 1599.255 2476.055 1599.585 2476.385 ;
        RECT 1600.000 2476.250 1604.600 2476.550 ;
        RECT 1599.270 2470.090 1599.570 2476.055 ;
        RECT 1600.000 2475.630 1604.600 2475.930 ;
        RECT 1601.110 2475.025 1601.410 2475.630 ;
        RECT 1601.095 2474.695 1601.425 2475.025 ;
        RECT 1602.935 2472.655 1603.265 2472.985 ;
        RECT 1602.950 2470.710 1603.250 2472.655 ;
        RECT 1600.000 2470.410 1604.600 2470.710 ;
        RECT 1599.270 2469.790 1604.600 2470.090 ;
        RECT 1599.255 2468.575 1599.585 2468.905 ;
        RECT 1599.270 2458.350 1599.570 2468.575 ;
        RECT 1602.015 2467.215 1602.345 2467.545 ;
        RECT 1602.030 2464.870 1602.330 2467.215 ;
        RECT 1600.000 2464.570 1604.600 2464.870 ;
        RECT 1600.000 2463.950 1604.600 2464.250 ;
        RECT 1600.190 2463.465 1600.490 2463.950 ;
        RECT 1600.175 2463.135 1600.505 2463.465 ;
        RECT 1602.935 2461.095 1603.265 2461.425 ;
        RECT 1602.950 2459.030 1603.250 2461.095 ;
        RECT 1600.000 2458.730 1604.600 2459.030 ;
        RECT 1600.000 2458.350 1604.600 2458.410 ;
        RECT 1599.270 2458.110 1604.600 2458.350 ;
        RECT 1599.270 2458.050 1600.340 2458.110 ;
        RECT 1599.255 2455.655 1599.585 2455.985 ;
        RECT 1599.270 2446.730 1599.570 2455.655 ;
        RECT 1602.935 2454.295 1603.265 2454.625 ;
        RECT 1602.950 2453.190 1603.250 2454.295 ;
        RECT 1600.000 2452.890 1604.600 2453.190 ;
        RECT 1600.000 2452.270 1604.600 2452.570 ;
        RECT 1601.110 2451.905 1601.410 2452.270 ;
        RECT 1601.095 2451.575 1601.425 2451.905 ;
        RECT 1601.095 2448.855 1601.425 2449.185 ;
        RECT 1601.110 2447.350 1601.410 2448.855 ;
        RECT 1600.000 2447.050 1604.600 2447.350 ;
        RECT 1599.270 2446.430 1604.600 2446.730 ;
        RECT 1603.855 2442.055 1604.185 2442.385 ;
        RECT 1603.870 2441.510 1604.170 2442.055 ;
        RECT 1600.000 2441.210 1604.600 2441.510 ;
        RECT 1600.000 2440.590 1604.600 2440.890 ;
        RECT 1601.110 2439.665 1601.410 2440.590 ;
        RECT 1599.255 2439.335 1599.585 2439.665 ;
        RECT 1601.095 2439.335 1601.425 2439.665 ;
        RECT 1599.270 2435.050 1599.570 2439.335 ;
        RECT 1601.095 2436.615 1601.425 2436.945 ;
        RECT 1601.110 2435.670 1601.410 2436.615 ;
        RECT 1600.000 2435.370 1604.600 2435.670 ;
        RECT 1599.270 2434.750 1604.600 2435.050 ;
        RECT 1599.255 2433.215 1599.585 2433.545 ;
        RECT 1599.270 2429.210 1599.570 2433.215 ;
        RECT 1602.015 2430.495 1602.345 2430.825 ;
        RECT 1602.030 2429.830 1602.330 2430.495 ;
        RECT 1600.000 2429.530 1604.600 2429.830 ;
        RECT 1599.270 2428.910 1604.600 2429.210 ;
        RECT 1599.255 2427.775 1599.585 2428.105 ;
        RECT 1599.270 2417.550 1599.570 2427.775 ;
        RECT 1602.935 2424.375 1603.265 2424.705 ;
        RECT 1602.950 2423.990 1603.250 2424.375 ;
        RECT 1600.000 2423.690 1604.600 2423.990 ;
        RECT 1600.000 2423.070 1604.600 2423.370 ;
        RECT 1601.110 2422.665 1601.410 2423.070 ;
        RECT 1601.095 2422.335 1601.425 2422.665 ;
        RECT 1602.015 2420.295 1602.345 2420.625 ;
        RECT 1602.030 2418.150 1602.330 2420.295 ;
        RECT 1600.000 2417.850 1604.600 2418.150 ;
        RECT 1599.270 2417.530 1600.340 2417.550 ;
        RECT 1599.270 2417.250 1604.600 2417.530 ;
        RECT 1600.000 2417.230 1604.600 2417.250 ;
        RECT 1599.255 2414.855 1599.585 2415.185 ;
        RECT 1599.270 2405.850 1599.570 2414.855 ;
        RECT 1602.935 2412.815 1603.265 2413.145 ;
        RECT 1602.950 2412.310 1603.250 2412.815 ;
        RECT 1600.000 2412.010 1604.600 2412.310 ;
        RECT 1600.000 2411.390 1604.600 2411.690 ;
        RECT 1601.110 2410.425 1601.410 2411.390 ;
        RECT 1601.095 2410.095 1601.425 2410.425 ;
        RECT 1602.015 2407.375 1602.345 2407.705 ;
        RECT 1602.030 2406.470 1602.330 2407.375 ;
        RECT 1600.000 2406.170 1604.600 2406.470 ;
        RECT 1599.270 2405.550 1604.600 2405.850 ;
        RECT 1602.935 2401.255 1603.265 2401.585 ;
        RECT 1602.950 2400.630 1603.250 2401.255 ;
        RECT 1600.000 2400.330 1604.600 2400.630 ;
        RECT 1600.000 2399.710 1604.600 2400.010 ;
        RECT 1601.110 2398.865 1601.410 2399.710 ;
        RECT 1599.255 2398.535 1599.585 2398.865 ;
        RECT 1601.095 2398.535 1601.425 2398.865 ;
        RECT 1599.270 2394.170 1599.570 2398.535 ;
        RECT 1602.935 2395.135 1603.265 2395.465 ;
        RECT 1602.950 2394.790 1603.250 2395.135 ;
        RECT 1600.000 2394.490 1604.600 2394.790 ;
        RECT 1599.270 2393.870 1604.600 2394.170 ;
        RECT 1602.935 2389.695 1603.265 2390.025 ;
        RECT 1602.950 2388.950 1603.250 2389.695 ;
        RECT 1599.270 2388.650 1604.600 2388.950 ;
        RECT 1599.270 2379.145 1599.570 2388.650 ;
        RECT 1600.000 2388.030 1604.600 2388.330 ;
        RECT 1601.110 2383.905 1601.410 2388.030 ;
        RECT 1601.095 2383.575 1601.425 2383.905 ;
        RECT 1602.015 2383.575 1602.345 2383.905 ;
        RECT 1602.030 2383.110 1602.330 2383.575 ;
        RECT 1600.000 2382.810 1604.600 2383.110 ;
        RECT 1600.000 2382.190 1604.600 2382.490 ;
        RECT 1599.255 2378.815 1599.585 2379.145 ;
        RECT 1602.950 2378.465 1603.250 2382.190 ;
        RECT 1603.855 2378.815 1604.185 2379.145 ;
        RECT 1602.935 2378.135 1603.265 2378.465 ;
        RECT 1603.870 2377.270 1604.170 2378.815 ;
        RECT 1600.000 2376.970 1604.600 2377.270 ;
        RECT 1600.000 2376.350 1604.600 2376.650 ;
        RECT 1601.110 2372.345 1601.410 2376.350 ;
        RECT 1601.095 2372.015 1601.425 2372.345 ;
        RECT 1603.855 2372.015 1604.185 2372.345 ;
        RECT 1603.870 2371.430 1604.170 2372.015 ;
        RECT 1600.000 2371.130 1604.600 2371.430 ;
        RECT 1600.000 2370.510 1604.600 2370.810 ;
        RECT 1601.110 2366.225 1601.410 2370.510 ;
        RECT 1601.095 2365.895 1601.425 2366.225 ;
        RECT 1602.935 2365.895 1603.265 2366.225 ;
        RECT 1602.950 2365.590 1603.250 2365.895 ;
        RECT 1600.000 2365.290 1604.600 2365.590 ;
        RECT 1600.000 2364.670 1604.600 2364.970 ;
        RECT 1601.095 2361.135 1601.425 2361.465 ;
        RECT 1601.110 2359.750 1601.410 2361.135 ;
        RECT 1602.030 2360.785 1602.330 2364.670 ;
        RECT 1602.015 2360.455 1602.345 2360.785 ;
        RECT 1599.270 2359.450 1604.600 2359.750 ;
        RECT 1599.270 2345.825 1599.570 2359.450 ;
        RECT 1600.000 2358.830 1604.600 2359.130 ;
        RECT 1602.030 2354.665 1602.330 2358.830 ;
        RECT 1602.935 2355.015 1603.265 2355.345 ;
        RECT 1602.015 2354.335 1602.345 2354.665 ;
        RECT 1602.950 2353.910 1603.250 2355.015 ;
        RECT 1600.000 2353.610 1604.600 2353.910 ;
        RECT 1600.000 2352.990 1604.600 2353.290 ;
        RECT 1601.110 2349.225 1601.410 2352.990 ;
        RECT 1602.015 2350.255 1602.345 2350.585 ;
        RECT 1601.095 2348.895 1601.425 2349.225 ;
        RECT 1602.030 2348.070 1602.330 2350.255 ;
        RECT 1600.000 2347.770 1604.600 2348.070 ;
        RECT 1600.000 2347.150 1604.600 2347.450 ;
        RECT 1599.255 2345.495 1599.585 2345.825 ;
        RECT 1601.110 2343.105 1601.410 2347.150 ;
        RECT 1602.935 2344.135 1603.265 2344.465 ;
        RECT 1601.095 2342.775 1601.425 2343.105 ;
        RECT 1602.950 2342.230 1603.250 2344.135 ;
        RECT 1600.000 2341.930 1604.600 2342.230 ;
        RECT 1600.000 2341.310 1604.600 2341.610 ;
        RECT 1601.110 2326.105 1601.410 2341.310 ;
        RECT 1602.015 2338.015 1602.345 2338.345 ;
        RECT 1602.030 2326.105 1602.330 2338.015 ;
        RECT 1601.095 2325.775 1601.425 2326.105 ;
        RECT 1602.015 2325.775 1602.345 2326.105 ;
      LAYER met4 ;
        RECT 1605.000 2205.000 2051.235 2581.480 ;
      LAYER met4 ;
        RECT 2051.635 2492.155 2056.235 2492.455 ;
        RECT 2051.635 2485.915 2056.235 2486.215 ;
        RECT 2051.635 2479.675 2056.235 2479.975 ;
        RECT 2051.635 2473.435 2056.235 2473.735 ;
        RECT 2051.635 2467.195 2056.235 2467.495 ;
        RECT 2051.635 2460.955 2056.235 2461.255 ;
        RECT 2051.635 2454.715 2056.235 2455.015 ;
        RECT 2051.635 2448.475 2056.235 2448.775 ;
        RECT 2051.635 2442.235 2056.235 2442.535 ;
        RECT 2051.635 2435.995 2056.235 2436.295 ;
        RECT 2051.635 2429.755 2056.235 2430.055 ;
        RECT 2051.635 2423.515 2056.235 2423.815 ;
        RECT 2051.635 2417.275 2056.235 2417.575 ;
        RECT 2051.635 2411.035 2056.235 2411.335 ;
        RECT 2051.635 2404.795 2056.235 2405.095 ;
        RECT 2051.635 2398.555 2056.235 2398.855 ;
        RECT 2051.635 2392.315 2056.235 2392.615 ;
        RECT 2051.635 2386.075 2056.235 2386.375 ;
        RECT 2051.635 2379.835 2056.235 2380.135 ;
        RECT 2051.635 2373.595 2056.235 2373.895 ;
        RECT 2051.635 2367.355 2056.235 2367.655 ;
        RECT 2051.635 2361.115 2056.235 2361.415 ;
        RECT 2051.635 2354.875 2056.235 2355.175 ;
        RECT 2051.635 2348.635 2056.235 2348.935 ;
        RECT 2051.635 2342.395 2056.235 2342.695 ;
        RECT 2051.635 2336.155 2056.235 2336.455 ;
        RECT 2051.635 2329.915 2056.235 2330.215 ;
        RECT 2051.635 2323.675 2056.235 2323.975 ;
        RECT 2051.635 2317.435 2056.235 2317.735 ;
        RECT 2051.635 2311.195 2056.235 2311.495 ;
        RECT 2051.635 2304.955 2056.235 2305.255 ;
        RECT 2051.635 2298.715 2056.235 2299.015 ;
        RECT 2051.635 2243.290 2056.235 2243.590 ;
        RECT 2051.635 2218.315 2056.235 2218.615 ;
        RECT 1603.670 2202.410 2044.680 2204.010 ;
        RECT 1604.060 2200.170 2052.140 2201.790 ;
        RECT 1383.055 2023.855 1383.385 2024.185 ;
        RECT 1601.095 1959.935 1601.425 1960.265 ;
        RECT 1601.110 1952.470 1601.410 1959.935 ;
        RECT 1600.000 1952.170 1604.600 1952.470 ;
        RECT 1601.095 1949.055 1601.425 1949.385 ;
        RECT 1601.110 1946.630 1601.410 1949.055 ;
        RECT 1600.000 1946.330 1604.600 1946.630 ;
        RECT 1601.095 1944.975 1601.425 1945.305 ;
        RECT 1601.110 1940.790 1601.410 1944.975 ;
        RECT 1600.000 1940.490 1604.600 1940.790 ;
        RECT 1601.095 1937.495 1601.425 1937.825 ;
        RECT 1601.110 1934.950 1601.410 1937.495 ;
        RECT 1600.000 1934.650 1604.600 1934.950 ;
        RECT 1599.255 1932.055 1599.585 1932.385 ;
        RECT 1599.270 1922.650 1599.570 1932.055 ;
        RECT 1601.095 1931.375 1601.425 1931.705 ;
        RECT 1601.110 1929.110 1601.410 1931.375 ;
        RECT 1600.000 1928.810 1604.600 1929.110 ;
        RECT 1602.935 1923.895 1603.265 1924.225 ;
        RECT 1602.950 1923.270 1603.250 1923.895 ;
        RECT 1600.000 1922.970 1604.600 1923.270 ;
        RECT 1599.270 1922.350 1604.600 1922.650 ;
        RECT 1599.255 1918.455 1599.585 1918.785 ;
        RECT 1599.270 1910.950 1599.570 1918.455 ;
        RECT 1603.855 1917.775 1604.185 1918.105 ;
        RECT 1603.870 1917.430 1604.170 1917.775 ;
        RECT 1600.000 1917.130 1604.600 1917.430 ;
        RECT 1600.000 1916.510 1604.600 1916.810 ;
        RECT 1601.110 1916.065 1601.410 1916.510 ;
        RECT 1601.095 1915.735 1601.425 1916.065 ;
        RECT 1603.855 1912.335 1604.185 1912.665 ;
        RECT 1603.870 1911.590 1604.170 1912.335 ;
        RECT 1600.000 1911.290 1604.600 1911.590 ;
        RECT 1600.000 1910.950 1604.600 1910.970 ;
        RECT 1599.270 1910.670 1604.600 1910.950 ;
        RECT 1599.270 1910.650 1600.340 1910.670 ;
        RECT 1602.935 1906.215 1603.265 1906.545 ;
        RECT 1602.950 1905.750 1603.250 1906.215 ;
        RECT 1600.000 1905.450 1604.600 1905.750 ;
        RECT 1600.000 1904.830 1604.600 1905.130 ;
        RECT 1602.030 1904.505 1602.330 1904.830 ;
        RECT 1602.015 1904.175 1602.345 1904.505 ;
        RECT 1603.855 1900.775 1604.185 1901.105 ;
        RECT 1603.870 1899.910 1604.170 1900.775 ;
        RECT 1600.000 1899.610 1604.600 1899.910 ;
        RECT 1600.000 1898.990 1604.600 1899.290 ;
        RECT 1601.110 1898.385 1601.410 1898.990 ;
        RECT 1601.095 1898.055 1601.425 1898.385 ;
        RECT 1599.255 1897.375 1599.585 1897.705 ;
        RECT 1599.270 1887.610 1599.570 1897.375 ;
        RECT 1602.015 1894.655 1602.345 1894.985 ;
        RECT 1602.030 1894.070 1602.330 1894.655 ;
        RECT 1600.000 1893.770 1604.600 1894.070 ;
        RECT 1600.000 1893.150 1604.600 1893.450 ;
        RECT 1602.950 1892.265 1603.250 1893.150 ;
        RECT 1602.935 1891.935 1603.265 1892.265 ;
        RECT 1603.855 1888.535 1604.185 1888.865 ;
        RECT 1603.870 1888.230 1604.170 1888.535 ;
        RECT 1600.000 1887.930 1604.600 1888.230 ;
        RECT 1599.270 1887.310 1604.600 1887.610 ;
        RECT 1600.175 1883.095 1600.505 1883.425 ;
        RECT 1600.190 1882.390 1600.490 1883.095 ;
        RECT 1598.350 1882.090 1604.600 1882.390 ;
        RECT 1598.350 1836.505 1598.650 1882.090 ;
        RECT 1600.000 1881.470 1604.600 1881.770 ;
        RECT 1601.110 1880.705 1601.410 1881.470 ;
        RECT 1601.095 1880.375 1601.425 1880.705 ;
        RECT 1601.095 1876.975 1601.425 1877.305 ;
        RECT 1601.110 1876.550 1601.410 1876.975 ;
        RECT 1600.000 1876.250 1604.600 1876.550 ;
        RECT 1599.255 1875.930 1599.585 1875.945 ;
        RECT 1599.255 1875.630 1604.600 1875.930 ;
        RECT 1599.255 1875.615 1599.585 1875.630 ;
        RECT 1602.935 1871.535 1603.265 1871.865 ;
        RECT 1602.950 1870.710 1603.250 1871.535 ;
        RECT 1600.000 1870.410 1604.600 1870.710 ;
        RECT 1600.000 1869.790 1604.600 1870.090 ;
        RECT 1600.190 1869.145 1600.490 1869.790 ;
        RECT 1600.175 1868.815 1600.505 1869.145 ;
        RECT 1600.175 1865.415 1600.505 1865.745 ;
        RECT 1600.190 1864.870 1600.490 1865.415 ;
        RECT 1600.000 1864.570 1604.600 1864.870 ;
        RECT 1600.000 1863.950 1604.600 1864.250 ;
        RECT 1599.255 1863.375 1599.585 1863.705 ;
        RECT 1599.270 1852.570 1599.570 1863.375 ;
        RECT 1602.030 1863.025 1602.330 1863.950 ;
        RECT 1602.015 1862.695 1602.345 1863.025 ;
        RECT 1602.935 1861.335 1603.265 1861.665 ;
        RECT 1602.950 1859.030 1603.250 1861.335 ;
        RECT 1600.000 1858.730 1604.600 1859.030 ;
        RECT 1600.000 1858.110 1604.600 1858.410 ;
        RECT 1601.110 1857.585 1601.410 1858.110 ;
        RECT 1601.095 1857.255 1601.425 1857.585 ;
        RECT 1603.855 1855.895 1604.185 1856.225 ;
        RECT 1603.870 1853.190 1604.170 1855.895 ;
        RECT 1600.000 1852.890 1604.600 1853.190 ;
        RECT 1599.270 1852.270 1604.600 1852.570 ;
        RECT 1602.015 1848.415 1602.345 1848.745 ;
        RECT 1602.030 1847.350 1602.330 1848.415 ;
        RECT 1600.000 1847.050 1604.600 1847.350 ;
        RECT 1600.000 1846.430 1604.600 1846.730 ;
        RECT 1602.030 1846.025 1602.330 1846.430 ;
        RECT 1602.015 1845.695 1602.345 1846.025 ;
        RECT 1599.255 1842.295 1599.585 1842.625 ;
        RECT 1603.855 1842.295 1604.185 1842.625 ;
        RECT 1598.335 1836.175 1598.665 1836.505 ;
        RECT 1599.270 1835.050 1599.570 1842.295 ;
        RECT 1603.870 1841.510 1604.170 1842.295 ;
        RECT 1600.000 1841.210 1604.600 1841.510 ;
        RECT 1600.000 1840.590 1604.600 1840.890 ;
        RECT 1601.110 1839.905 1601.410 1840.590 ;
        RECT 1601.095 1839.575 1601.425 1839.905 ;
        RECT 1603.855 1836.175 1604.185 1836.505 ;
        RECT 1603.870 1835.670 1604.170 1836.175 ;
        RECT 1600.000 1835.370 1604.600 1835.670 ;
        RECT 1599.270 1834.750 1604.600 1835.050 ;
        RECT 1602.935 1830.735 1603.265 1831.065 ;
        RECT 1602.950 1829.830 1603.250 1830.735 ;
        RECT 1600.000 1829.530 1604.600 1829.830 ;
        RECT 1600.000 1828.910 1604.600 1829.210 ;
        RECT 1600.190 1828.345 1600.490 1828.910 ;
        RECT 1600.175 1828.015 1600.505 1828.345 ;
        RECT 1601.095 1824.615 1601.425 1824.945 ;
        RECT 1601.110 1823.990 1601.410 1824.615 ;
        RECT 1600.000 1823.690 1604.600 1823.990 ;
        RECT 1600.000 1823.070 1604.600 1823.370 ;
        RECT 1602.030 1822.225 1602.330 1823.070 ;
        RECT 1602.015 1821.895 1602.345 1822.225 ;
        RECT 1600.175 1818.495 1600.505 1818.825 ;
        RECT 1600.190 1818.150 1600.490 1818.495 ;
        RECT 1600.000 1817.850 1604.600 1818.150 ;
        RECT 1597.415 1817.450 1597.745 1817.465 ;
        RECT 1600.000 1817.450 1604.600 1817.530 ;
        RECT 1597.415 1817.230 1604.600 1817.450 ;
        RECT 1597.415 1817.150 1600.340 1817.230 ;
        RECT 1597.415 1817.135 1597.745 1817.150 ;
        RECT 1600.175 1813.055 1600.505 1813.385 ;
        RECT 1600.190 1812.310 1600.490 1813.055 ;
        RECT 1600.000 1812.010 1604.600 1812.310 ;
        RECT 1600.000 1811.390 1604.600 1811.690 ;
        RECT 1602.030 1810.665 1602.330 1811.390 ;
        RECT 1602.015 1810.335 1602.345 1810.665 ;
        RECT 1599.255 1806.935 1599.585 1807.265 ;
        RECT 1601.095 1806.935 1601.425 1807.265 ;
        RECT 1599.270 1800.010 1599.570 1806.935 ;
        RECT 1601.110 1806.470 1601.410 1806.935 ;
        RECT 1600.000 1806.170 1604.600 1806.470 ;
        RECT 1600.000 1805.550 1604.600 1805.850 ;
        RECT 1601.110 1805.225 1601.410 1805.550 ;
        RECT 1601.095 1804.895 1601.425 1805.225 ;
        RECT 1601.095 1801.495 1601.425 1801.825 ;
        RECT 1601.110 1800.630 1601.410 1801.495 ;
        RECT 1600.000 1800.330 1604.600 1800.630 ;
        RECT 1599.270 1799.710 1604.600 1800.010 ;
        RECT 1602.015 1798.775 1602.345 1799.105 ;
        RECT 1602.030 1794.790 1602.330 1798.775 ;
        RECT 1600.000 1794.490 1604.600 1794.790 ;
        RECT 1600.000 1793.870 1604.600 1794.170 ;
        RECT 1602.030 1792.985 1602.330 1793.870 ;
        RECT 1602.015 1792.655 1602.345 1792.985 ;
        RECT 1601.095 1789.255 1601.425 1789.585 ;
        RECT 1601.110 1788.950 1601.410 1789.255 ;
        RECT 1600.000 1788.650 1604.600 1788.950 ;
        RECT 1600.000 1788.030 1604.600 1788.330 ;
        RECT 1369.255 1785.855 1369.585 1786.185 ;
        RECT 1601.110 1784.145 1601.410 1788.030 ;
        RECT 1602.935 1785.175 1603.265 1785.505 ;
        RECT 1601.095 1783.815 1601.425 1784.145 ;
        RECT 1602.950 1783.110 1603.250 1785.175 ;
        RECT 1600.000 1782.810 1604.600 1783.110 ;
        RECT 1600.000 1782.190 1604.600 1782.490 ;
        RECT 1601.110 1778.025 1601.410 1782.190 ;
        RECT 1602.935 1779.735 1603.265 1780.065 ;
        RECT 1601.095 1777.695 1601.425 1778.025 ;
        RECT 1602.950 1777.270 1603.250 1779.735 ;
        RECT 1600.000 1776.970 1604.600 1777.270 ;
        RECT 1600.000 1776.350 1604.600 1776.650 ;
        RECT 1601.110 1772.585 1601.410 1776.350 ;
        RECT 1603.855 1772.935 1604.185 1773.265 ;
        RECT 1601.095 1772.255 1601.425 1772.585 ;
        RECT 1603.870 1771.430 1604.170 1772.935 ;
        RECT 1600.000 1771.130 1604.600 1771.430 ;
        RECT 1600.000 1770.510 1604.600 1770.810 ;
        RECT 1599.255 1766.815 1599.585 1767.145 ;
        RECT 1599.270 1742.230 1599.570 1766.815 ;
        RECT 1601.110 1766.465 1601.410 1770.510 ;
        RECT 1601.095 1766.135 1601.425 1766.465 ;
        RECT 1603.855 1766.135 1604.185 1766.465 ;
        RECT 1603.870 1765.590 1604.170 1766.135 ;
        RECT 1600.000 1765.290 1604.600 1765.590 ;
        RECT 1600.000 1764.670 1604.600 1764.970 ;
        RECT 1601.110 1763.065 1601.410 1764.670 ;
        RECT 1601.095 1762.735 1601.425 1763.065 ;
        RECT 1602.015 1762.055 1602.345 1762.385 ;
        RECT 1602.030 1759.750 1602.330 1762.055 ;
        RECT 1600.000 1759.450 1604.600 1759.750 ;
        RECT 1600.000 1758.830 1604.600 1759.130 ;
        RECT 1602.030 1754.905 1602.330 1758.830 ;
        RECT 1602.935 1755.935 1603.265 1756.265 ;
        RECT 1602.015 1754.575 1602.345 1754.905 ;
        RECT 1602.950 1753.910 1603.250 1755.935 ;
        RECT 1600.000 1753.610 1604.600 1753.910 ;
        RECT 1600.000 1752.990 1604.600 1753.290 ;
        RECT 1601.110 1748.785 1601.410 1752.990 ;
        RECT 1603.855 1750.495 1604.185 1750.825 ;
        RECT 1601.095 1748.455 1601.425 1748.785 ;
        RECT 1603.870 1748.070 1604.170 1750.495 ;
        RECT 1600.000 1747.770 1604.600 1748.070 ;
        RECT 1600.000 1747.150 1604.600 1747.450 ;
        RECT 1601.110 1743.345 1601.410 1747.150 ;
        RECT 1601.095 1743.015 1601.425 1743.345 ;
        RECT 1599.270 1741.930 1604.600 1742.230 ;
        RECT 1600.000 1741.310 1604.600 1741.610 ;
        RECT 1601.110 1731.785 1601.410 1741.310 ;
        RECT 1601.095 1731.455 1601.425 1731.785 ;
      LAYER met4 ;
        RECT 1605.000 1605.000 2051.235 1981.480 ;
      LAYER met4 ;
        RECT 2051.635 1892.155 2056.235 1892.455 ;
        RECT 2051.635 1885.915 2056.235 1886.215 ;
        RECT 2051.635 1879.675 2056.235 1879.975 ;
        RECT 2051.635 1873.435 2056.235 1873.735 ;
        RECT 2051.635 1867.195 2056.235 1867.495 ;
        RECT 2051.635 1860.955 2056.235 1861.255 ;
        RECT 2051.635 1854.715 2056.235 1855.015 ;
        RECT 2051.635 1848.475 2056.235 1848.775 ;
        RECT 2051.635 1842.235 2056.235 1842.535 ;
        RECT 2051.635 1835.995 2056.235 1836.295 ;
        RECT 2051.635 1829.755 2056.235 1830.055 ;
        RECT 2051.635 1823.515 2056.235 1823.815 ;
        RECT 2051.635 1817.275 2056.235 1817.575 ;
        RECT 2051.635 1811.035 2056.235 1811.335 ;
        RECT 2051.635 1804.795 2056.235 1805.095 ;
        RECT 2051.635 1798.555 2056.235 1798.855 ;
        RECT 2051.635 1792.315 2056.235 1792.615 ;
        RECT 2051.635 1786.075 2056.235 1786.375 ;
        RECT 2051.635 1779.835 2056.235 1780.135 ;
        RECT 2051.635 1773.595 2056.235 1773.895 ;
        RECT 2051.635 1767.355 2056.235 1767.655 ;
        RECT 2051.635 1761.115 2056.235 1761.415 ;
        RECT 2051.635 1754.875 2056.235 1755.175 ;
        RECT 2051.635 1748.635 2056.235 1748.935 ;
        RECT 2051.635 1742.395 2056.235 1742.695 ;
        RECT 2051.635 1736.155 2056.235 1736.455 ;
        RECT 2051.635 1729.915 2056.235 1730.215 ;
        RECT 2051.635 1723.675 2056.235 1723.975 ;
        RECT 2051.635 1717.435 2056.235 1717.735 ;
        RECT 2051.635 1711.195 2056.235 1711.495 ;
        RECT 2051.635 1704.955 2056.235 1705.255 ;
        RECT 2051.635 1698.715 2056.235 1699.015 ;
        RECT 2051.635 1643.290 2056.235 1643.590 ;
        RECT 2051.635 1618.315 2056.235 1618.615 ;
        RECT 1603.670 1602.410 2044.680 1604.010 ;
        RECT 1604.060 1600.170 2052.140 1601.790 ;
      LAYER met5 ;
        RECT 405.000 3288.380 781.480 3301.235 ;
        RECT 955.000 3288.380 1331.480 3301.235 ;
        RECT 405.000 3270.380 781.480 3285.380 ;
        RECT 955.000 3270.380 1331.480 3285.380 ;
        RECT 405.000 3252.380 781.480 3267.380 ;
        RECT 955.000 3252.380 1331.480 3267.380 ;
        RECT 405.000 3216.380 781.480 3249.380 ;
        RECT 955.000 3216.380 1331.480 3249.380 ;
        RECT 405.000 3198.380 781.480 3213.380 ;
        RECT 955.000 3198.380 1331.480 3213.380 ;
        RECT 405.000 3180.380 781.480 3195.380 ;
        RECT 955.000 3180.380 1331.480 3195.380 ;
        RECT 405.000 3162.380 781.480 3177.380 ;
        RECT 955.000 3162.380 1331.480 3177.380 ;
        RECT 405.000 3126.380 781.480 3159.380 ;
        RECT 955.000 3126.380 1331.480 3159.380 ;
        RECT 405.000 3108.380 781.480 3123.380 ;
        RECT 955.000 3108.380 1331.480 3123.380 ;
        RECT 405.000 3090.380 781.480 3105.380 ;
        RECT 955.000 3090.380 1331.480 3105.380 ;
        RECT 405.000 3072.380 781.480 3087.380 ;
        RECT 955.000 3072.380 1331.480 3087.380 ;
        RECT 405.000 3036.380 781.480 3069.380 ;
        RECT 955.000 3036.380 1331.480 3069.380 ;
        RECT 405.000 3018.380 781.480 3033.380 ;
        RECT 955.000 3018.380 1331.480 3033.380 ;
        RECT 405.000 3000.380 781.480 3015.380 ;
        RECT 955.000 3000.380 1331.480 3015.380 ;
        RECT 405.000 2982.380 781.480 2997.380 ;
        RECT 955.000 2982.380 1331.480 2997.380 ;
        RECT 405.000 2946.380 781.480 2979.380 ;
        RECT 955.000 2946.380 1331.480 2979.380 ;
        RECT 405.000 2928.380 781.480 2943.380 ;
        RECT 955.000 2928.380 1331.480 2943.380 ;
        RECT 405.000 2910.380 781.480 2925.380 ;
        RECT 955.000 2910.380 1331.480 2925.380 ;
        RECT 405.000 2892.380 781.480 2907.380 ;
        RECT 955.000 2892.380 1331.480 2907.380 ;
        RECT 405.000 2856.380 781.480 2889.380 ;
        RECT 955.000 2856.380 1331.480 2889.380 ;
        RECT 1605.000 2568.380 2051.235 2581.480 ;
        RECT 1605.000 2550.380 2051.235 2565.380 ;
        RECT 1605.000 2532.380 2051.235 2547.380 ;
        RECT 1605.000 2496.380 2051.235 2529.380 ;
        RECT 1605.000 2478.380 2051.235 2493.380 ;
        RECT 1605.000 2460.380 2051.235 2475.380 ;
        RECT 1605.000 2442.380 2051.235 2457.380 ;
        RECT 1605.000 2406.380 2051.235 2439.380 ;
        RECT 1605.000 2388.380 2051.235 2403.380 ;
        RECT 1605.000 2370.380 2051.235 2385.380 ;
        RECT 1605.000 2352.380 2051.235 2367.380 ;
        RECT 1605.000 2316.380 2051.235 2349.380 ;
        RECT 1605.000 2298.380 2051.235 2313.380 ;
        RECT 1605.000 2280.380 2051.235 2295.380 ;
        RECT 1605.000 2262.380 2051.235 2277.380 ;
        RECT 1605.000 2226.380 2051.235 2259.380 ;
        RECT 1605.000 2208.380 2051.235 2223.380 ;
        RECT 1605.000 2205.000 2051.235 2205.380 ;
        RECT 1605.000 1956.380 2051.235 1981.480 ;
        RECT 1605.000 1938.380 2051.235 1953.380 ;
        RECT 1605.000 1920.380 2051.235 1935.380 ;
        RECT 1605.000 1902.380 2051.235 1917.380 ;
        RECT 1605.000 1866.380 2051.235 1899.380 ;
        RECT 1605.000 1848.380 2051.235 1863.380 ;
        RECT 1605.000 1830.380 2051.235 1845.380 ;
        RECT 1605.000 1812.380 2051.235 1827.380 ;
        RECT 1605.000 1776.380 2051.235 1809.380 ;
        RECT 1605.000 1758.380 2051.235 1773.380 ;
        RECT 1605.000 1740.380 2051.235 1755.380 ;
        RECT 1605.000 1722.380 2051.235 1737.380 ;
        RECT 1605.000 1686.380 2051.235 1719.380 ;
        RECT 1605.000 1668.380 2051.235 1683.380 ;
        RECT 1605.000 1650.380 2051.235 1665.380 ;
        RECT 1605.000 1632.380 2051.235 1647.380 ;
        RECT 1605.000 1605.000 2051.235 1629.380 ;
  END
END user_project_wrapper
END LIBRARY

