magic
tech sky130A
magscale 1 2
timestamp 1607736046
<< locali >>
rect 115397 567375 115431 568021
rect 116685 567919 116719 568497
rect 116869 567307 116903 568225
rect 116961 567443 116995 568157
rect 103161 524297 103437 524331
rect 103161 524263 103195 524297
rect 108313 524059 108347 524229
rect 105737 523515 105771 523889
rect 113189 523651 113223 524297
rect 117973 523855 118007 524025
rect 121377 523923 121411 524025
rect 122665 523855 122699 524229
rect 122757 523651 122791 524297
rect 132509 523039 132543 524297
rect 159223 524297 159373 524331
rect 132601 523107 132635 524229
rect 141985 523243 142019 524229
rect 137753 523107 137787 523209
rect 142077 523039 142111 524297
rect 156153 523583 156187 524229
rect 214021 523855 214055 524093
rect 243553 523855 243587 523957
rect 243461 523651 243495 523821
rect 243645 523719 243679 523957
rect 243737 523651 243771 523685
rect 243461 523617 243771 523651
rect 147505 523243 147539 523345
rect 147597 523039 147631 523209
rect 299489 502707 299523 502809
rect 280169 502503 280203 502605
rect 289645 502367 289679 502605
rect 289829 502367 289863 502673
rect 309057 502639 309091 502809
rect 311851 502605 311909 502639
rect 320649 490943 320683 495465
rect 320649 489923 320683 490909
rect 320833 487271 320867 489821
rect 320465 480335 320499 482817
rect 320833 478975 320867 479417
rect 320741 470475 320775 476017
rect 320373 467619 320407 467789
rect 320741 467551 320775 470441
rect 320833 467415 320867 475745
rect 320189 446811 320223 452285
rect 320281 446879 320315 457453
rect 320373 456671 320407 456909
rect 320649 452659 320683 457317
rect 320373 447015 320407 447321
rect 320649 446947 320683 449837
rect 320741 447151 320775 457453
rect 320833 456535 320867 456909
rect 320833 447083 320867 452625
rect 320649 378335 320683 379729
rect 320741 379559 320775 381361
rect 289771 376669 289829 376703
rect 298109 376635 298143 376737
rect 302893 376567 302927 376737
rect 320833 374663 320867 380273
rect 320097 372963 320131 374629
rect 320281 367863 320315 371025
rect 292589 366911 292623 366945
rect 292531 366877 292623 366911
rect 298109 366911 298143 367013
rect 307769 366843 307803 366945
rect 317429 366299 317463 366945
rect 320373 362695 320407 368577
rect 320465 363783 320499 372929
rect 320833 370515 320867 371569
rect 320281 355895 320315 360145
rect 320373 359907 320407 362661
rect 142905 318699 142939 318801
rect 152841 318699 152875 318801
rect 74365 318121 74549 318155
rect 74365 318087 74399 318121
rect 75101 318087 75135 318461
rect 75009 318019 75043 318053
rect 75285 318019 75319 318393
rect 142813 318291 142847 318665
rect 75009 317985 75319 318019
rect 84669 317611 84703 317985
rect 136925 317951 136959 318257
rect 138397 317815 138431 318121
rect 142721 317951 142755 318257
rect 84761 317611 84795 317713
rect 70409 317339 70443 317577
rect 138489 317475 138523 317781
rect 141985 317679 142019 317849
rect 142813 317747 142847 317849
rect 70869 307819 70903 309145
rect 92857 307819 92891 317373
rect 94053 307887 94087 317373
rect 139317 317339 139351 317577
rect 140789 317339 140823 317577
rect 141893 317339 141927 317645
rect 142905 317611 142939 317713
rect 145021 317679 145055 318665
rect 147505 318291 147539 318393
rect 148057 318223 148091 318665
rect 146769 317747 146803 317917
rect 145665 317339 145699 317713
rect 147321 309179 147355 317849
rect 147689 317407 147723 318189
rect 149253 317815 149287 318325
rect 150449 318223 150483 318393
rect 152749 318291 152783 318665
rect 148425 317475 148459 317781
rect 151737 317475 151771 318121
rect 153301 318087 153335 318325
rect 151829 317815 151863 317917
rect 152473 317883 152507 318053
rect 154037 317611 154071 318393
rect 157257 318155 157291 318665
rect 191021 318291 191055 318529
rect 200589 318427 200623 318801
rect 224969 318767 225003 318869
rect 162133 309179 162167 317985
rect 190009 317815 190043 318053
rect 190101 317815 190135 318257
rect 184949 317543 184983 317713
rect 195897 317679 195931 318257
rect 200681 318155 200715 318461
rect 198967 318053 199117 318087
rect 200773 317883 200807 318733
rect 201601 318563 201635 318665
rect 193873 307819 193907 309213
rect 198013 309179 198047 317849
rect 204177 317747 204211 318053
rect 204913 309179 204947 318733
rect 208593 318019 208627 318733
rect 210433 318087 210467 318325
rect 210525 318019 210559 318325
rect 212089 318155 212123 318325
rect 212549 317407 212583 317713
rect 213837 317475 213871 318733
rect 215217 318155 215251 318665
rect 220093 318495 220127 318733
rect 220001 318223 220035 318461
rect 222209 318155 222243 318665
rect 224877 318223 224911 318733
rect 224727 318189 224911 318223
rect 234353 318019 234387 318869
rect 224877 317407 224911 317713
rect 270509 317407 270543 317713
rect 236193 307819 236227 317373
rect 280077 317407 280111 317713
rect 289829 317475 289863 317713
rect 299397 317475 299431 317713
rect 309149 317611 309183 317713
rect 238953 307819 238987 317373
rect 70501 289867 70535 299421
rect 94053 298163 94087 307717
rect 105093 298163 105127 302209
rect 245577 299523 245611 309077
rect 251281 306935 251315 309553
rect 254041 299523 254075 309077
rect 70777 288439 70811 298061
rect 72157 288371 72191 296633
rect 151093 289867 151127 299421
rect 193873 288439 193907 298061
rect 227361 289867 227395 299421
rect 235733 287147 235767 296633
rect 242633 288439 242667 298061
rect 243921 288439 243955 298061
rect 246957 288439 246991 298061
rect 248245 288439 248279 298061
rect 251281 297279 251315 299421
rect 255237 298163 255271 299489
rect 255237 288439 255271 297993
rect 259285 289867 259319 297449
rect 265817 292655 265851 302141
rect 267105 299455 267139 303569
rect 324973 299523 325007 309077
rect 271521 293539 271555 299421
rect 267197 282931 267231 287725
rect 78873 278783 78907 282897
rect 324973 280211 325007 289765
rect 90005 267767 90039 273309
rect 105185 273139 105219 280109
rect 106657 273275 106691 280109
rect 151093 270555 151127 280109
rect 243829 277423 243863 278817
rect 105185 263483 105219 270453
rect 106841 260899 106875 270453
rect 234077 260899 234111 270385
rect 249625 260899 249659 270453
rect 251005 260899 251039 270453
rect 252293 260899 252327 270453
rect 259285 260899 259319 270453
rect 264621 264979 264655 274601
rect 268669 267767 268703 273241
rect 324973 260899 325007 270453
rect 70777 241519 70811 259369
rect 105185 253827 105219 260797
rect 73445 241519 73479 252569
rect 151093 251243 151127 260797
rect 70777 231863 70811 234549
rect 94053 231863 94087 244953
rect 105093 241519 105127 251141
rect 252293 241519 252327 251141
rect 324789 241587 324823 251073
rect 324881 234651 324915 241417
rect 77493 217379 77527 225641
rect 78781 219487 78815 229041
rect 105093 222207 105127 224961
rect 106473 220915 106507 230401
rect 70777 212551 70811 215237
rect 91017 212483 91051 220677
rect 266001 218059 266035 230469
rect 77493 202895 77527 205649
rect 91017 202827 91051 211089
rect 233801 208403 233835 216597
rect 105093 202895 105127 205649
rect 70777 193239 70811 195925
rect 94053 193239 94087 202793
rect 235549 200175 235583 209729
rect 252293 191879 252327 201433
rect 78781 183583 78815 186337
rect 105093 183583 105127 186337
rect 264621 185691 264655 192525
rect 70777 173927 70811 176613
rect 72341 171139 72375 174029
rect 77493 173927 77527 183481
rect 91017 180863 91051 183549
rect 91017 171139 91051 178653
rect 235641 171139 235675 180761
rect 70685 154615 70719 157437
rect 73445 144891 73479 153153
rect 81909 144823 81943 161381
rect 106657 157335 106691 164169
rect 94053 146999 94087 156621
rect 151093 154615 151127 164169
rect 193873 153255 193907 162809
rect 211905 157335 211939 164169
rect 227361 157335 227395 164169
rect 242541 162911 242575 172465
rect 266001 169779 266035 179333
rect 267289 169779 267323 179333
rect 234169 151827 234203 161381
rect 72341 124219 72375 133841
rect 73537 131563 73571 143429
rect 105093 137955 105127 143497
rect 106657 137955 106691 144857
rect 151093 135303 151127 144857
rect 193873 133943 193907 143497
rect 211905 137955 211939 144857
rect 227361 137955 227395 144857
rect 242541 143599 242575 153153
rect 243829 151827 243863 161381
rect 264621 160123 264655 169677
rect 266001 150467 266035 160021
rect 267289 150467 267323 160021
rect 78781 106335 78815 115889
rect 105093 114563 105127 124117
rect 106473 114631 106507 124049
rect 151093 115991 151127 125545
rect 193873 114563 193907 124117
rect 211905 118643 211939 125545
rect 227361 118643 227395 125545
rect 234169 124219 234203 142069
rect 242541 124219 242575 133841
rect 243829 124219 243863 133773
rect 266001 131155 266035 140709
rect 267289 131155 267323 140709
rect 234261 114631 234295 119357
rect 70777 95319 70811 104805
rect 72249 96747 72283 106233
rect 73537 95251 73571 106233
rect 90925 104907 90959 114461
rect 94053 95251 94087 104805
rect 105093 95251 105127 104805
rect 106657 93891 106691 103445
rect 151093 96679 151127 106233
rect 193873 95251 193907 104805
rect 211905 99331 211939 106233
rect 227361 99331 227395 106233
rect 234169 104907 234203 114461
rect 242541 104907 242575 114461
rect 243829 113203 243863 122757
rect 252293 114563 252327 124117
rect 255237 106335 255271 124117
rect 266001 111843 266035 121397
rect 267381 111843 267415 121397
rect 268669 113203 268703 122757
rect 234169 95251 234203 100045
rect 72157 75939 72191 85493
rect 73445 75939 73479 85493
rect 77493 75939 77527 85493
rect 78689 84303 78723 93789
rect 72157 67711 72191 72437
rect 70685 57987 70719 67541
rect 72065 56627 72099 66181
rect 78689 64923 78723 82773
rect 81725 75939 81759 85493
rect 90005 77299 90039 86853
rect 92765 77299 92799 86853
rect 106657 85595 106691 89777
rect 234169 87091 234203 91749
rect 235733 87023 235767 96577
rect 246957 95251 246991 104805
rect 252109 95251 252143 104805
rect 94053 80971 94087 85493
rect 105093 84167 105127 85493
rect 151093 77299 151127 86921
rect 193873 75939 193907 85493
rect 204729 75939 204763 85493
rect 211905 77299 211939 86921
rect 227361 77299 227395 86921
rect 242541 85595 242575 95149
rect 255237 87023 255271 104805
rect 259285 95251 259319 104805
rect 264621 102187 264655 111673
rect 266001 92531 266035 102085
rect 267289 92531 267323 102085
rect 268577 93891 268611 103445
rect 234169 75939 234203 85493
rect 90005 58055 90039 67541
rect 92765 58055 92799 67541
rect 94145 64923 94179 74477
rect 105001 66283 105035 74545
rect 106473 66351 106507 75837
rect 211905 70363 211939 75837
rect 235733 67643 235767 77197
rect 246957 75939 246991 85493
rect 252293 75939 252327 85493
rect 255237 75939 255271 85493
rect 259285 75939 259319 85493
rect 264621 82875 264655 92361
rect 90925 55267 90959 56661
rect 72065 37315 72099 46869
rect 73445 37315 73479 46869
rect 81725 38675 81759 51765
rect 94145 50643 94179 59993
rect 151093 57987 151127 67541
rect 242541 66283 242575 75837
rect 266001 73219 266035 82773
rect 267289 73219 267323 82773
rect 324973 67643 325007 77197
rect 193873 56627 193907 66181
rect 204913 56627 204947 66181
rect 96997 47039 97031 56525
rect 211905 50711 211939 57885
rect 227361 51051 227395 57885
rect 234077 57851 234111 66181
rect 235733 48331 235767 57885
rect 246957 56627 246991 66181
rect 252293 56627 252327 66181
rect 255237 56627 255271 66181
rect 259285 56627 259319 66181
rect 78781 37315 78815 38641
rect 96997 37315 97031 46869
rect 151093 38675 151127 48229
rect 242541 46971 242575 56525
rect 267289 53839 267323 63461
rect 73445 29019 73479 36261
rect 106841 31603 106875 38573
rect 193873 29019 193907 46869
rect 204913 37315 204947 46869
rect 234077 38675 234111 46869
rect 211905 29019 211939 38573
rect 235733 29019 235767 38573
rect 246957 37315 246991 46869
rect 251005 37315 251039 46869
rect 252293 37315 252327 46869
rect 255237 37315 255271 46869
rect 259285 37315 259319 46869
rect 264621 44319 264655 53737
rect 77493 18003 77527 27557
rect 78873 18003 78907 27557
rect 90005 19363 90039 28917
rect 91109 18003 91143 27557
rect 96997 21947 97031 28917
rect 151093 19363 151127 28917
rect 242541 27659 242575 37213
rect 267289 35819 267323 44081
rect 324881 38539 324915 46869
rect 261953 29699 261987 33133
rect 73353 8347 73387 17901
rect 193781 12427 193815 19261
rect 204913 18003 204947 27557
rect 227361 11883 227395 19261
rect 235733 15895 235767 19261
rect 248245 18003 248279 27557
rect 249625 18003 249659 27557
rect 255237 18003 255271 27557
rect 259193 13175 259227 22729
rect 260389 13107 260423 26197
rect 255145 11067 255179 13073
rect 81633 3927 81667 4097
rect 70317 3689 70443 3723
rect 70317 3655 70351 3689
rect 70409 3655 70443 3689
rect 70501 3451 70535 3757
rect 70685 3723 70719 3893
rect 45385 3043 45419 3349
rect 45477 3111 45511 3281
rect 55229 2839 55263 3349
rect 55321 3043 55355 3281
rect 61117 2703 61151 3009
rect 62313 2771 62347 3077
rect 64613 2703 64647 3281
rect 64705 2771 64739 3213
rect 64797 2839 64831 3349
rect 71513 3247 71547 3417
rect 71513 3213 71881 3247
rect 73721 1003 73755 3689
rect 75101 3485 75319 3519
rect 75101 3247 75135 3485
rect 75285 3451 75319 3485
rect 76205 3451 76239 3757
rect 79977 3723 80011 3893
rect 79885 3451 79919 3689
rect 79885 3417 79977 3451
rect 75193 3247 75227 3417
rect 82461 3383 82495 3825
rect 89177 3247 89211 4029
rect 89269 3179 89303 3961
rect 91569 3383 91603 4029
rect 91661 3791 91695 4029
rect 91477 3247 91511 3349
rect 94237 2907 94271 9605
rect 161305 8823 161339 8925
rect 167009 8619 167043 8789
rect 176577 8619 176611 8789
rect 186329 8415 186363 8789
rect 195805 8789 195897 8823
rect 193229 8279 193263 8585
rect 195805 8483 195839 8789
rect 238861 8687 238895 9605
rect 239321 9435 239355 9537
rect 239229 8891 239263 9401
rect 239413 9367 239447 9605
rect 239505 8551 239539 9469
rect 244841 8755 244875 9469
rect 246681 9299 246715 9469
rect 248981 9401 249291 9435
rect 248981 9231 249015 9401
rect 249257 9367 249291 9401
rect 248981 8483 249015 8857
rect 196081 8279 196115 8449
rect 197185 8211 197219 8381
rect 205591 8381 205649 8415
rect 202889 8211 202923 8381
rect 205499 8313 205741 8347
rect 215125 8007 215159 8449
rect 249073 8483 249107 8789
rect 249165 8551 249199 9333
rect 249257 8687 249291 9061
rect 249349 8755 249383 9265
rect 249441 8687 249475 9401
rect 254961 8891 254995 9265
rect 255053 8891 255087 9129
rect 258733 8891 258767 9333
rect 259009 9163 259043 9401
rect 259101 9095 259135 9129
rect 258825 9061 259135 9095
rect 258641 8823 258675 8857
rect 258825 8823 258859 9061
rect 258641 8789 258859 8823
rect 215217 8075 215251 8381
rect 215309 8075 215343 8381
rect 215401 8007 215435 8449
rect 157349 4811 157383 5525
rect 127483 3961 127817 3995
rect 127725 3655 127759 3893
rect 123251 3553 123585 3587
rect 122021 3179 122055 3349
rect 127541 3179 127575 3485
rect 127633 3315 127667 3485
rect 127817 3247 127851 3621
rect 127909 3383 127943 4165
rect 132509 4063 132543 4233
rect 136189 3519 136223 4165
rect 153703 4097 153945 4131
rect 127909 3179 127943 3213
rect 127541 3145 127943 3179
rect 132969 2771 133003 3485
rect 133061 2975 133095 3417
rect 138673 3043 138707 3485
rect 148885 3043 148919 3485
rect 149069 3247 149103 3349
rect 148977 3043 149011 3213
rect 153025 3179 153059 4029
rect 155233 3383 155267 3893
rect 157257 3179 157291 4097
rect 157349 4063 157383 4165
rect 161213 3179 161247 7429
rect 162133 3315 162167 6613
rect 171793 4199 171827 4777
rect 181453 4199 181487 4777
rect 162041 3179 162075 3281
rect 162409 3247 162443 3553
rect 164801 3383 164835 4029
rect 195897 3995 195931 4777
rect 195989 3995 196023 4777
rect 201601 4335 201635 7021
rect 205189 4403 205223 7021
rect 215435 4777 215527 4811
rect 211721 4505 212365 4539
rect 211721 4471 211755 4505
rect 215217 4471 215251 4777
rect 215493 4743 215527 4777
rect 215343 4709 215435 4743
rect 219081 4709 219357 4743
rect 215401 4539 215435 4709
rect 219081 4539 219115 4709
rect 219173 4539 219207 4641
rect 223037 4607 223071 4709
rect 229569 4471 229603 4777
rect 229753 4607 229787 4777
rect 239137 4539 239171 4709
rect 204821 4267 204855 4301
rect 225889 4267 225923 4437
rect 204821 4233 205373 4267
rect 229661 4199 229695 4505
rect 234445 4505 234629 4539
rect 234445 4471 234479 4505
rect 239229 4471 239263 4641
rect 232639 4369 232697 4403
rect 231961 4267 231995 4369
rect 231903 4233 231995 4267
rect 239413 4199 239447 4505
rect 241437 4199 241471 6885
rect 247877 4743 247911 5117
rect 244139 4369 244381 4403
rect 248889 4267 248923 5049
rect 249349 4335 249383 4981
rect 249441 4403 249475 5457
rect 249625 4539 249659 6885
rect 254869 4811 254903 5049
rect 255053 4743 255087 4981
rect 257445 4811 257479 4981
rect 257537 4811 257571 4913
rect 258089 4913 258273 4947
rect 258089 4879 258123 4913
rect 258733 4607 258767 5321
rect 258825 5151 258859 5321
rect 268059 4981 268301 5015
rect 268485 4879 268519 5117
rect 340153 3995 340187 4097
rect 369041 3927 369075 4097
rect 369041 3893 369225 3927
rect 378609 3893 378827 3927
rect 169033 3247 169067 3553
rect 162501 3179 162535 3213
rect 162041 3145 162535 3179
rect 169953 3281 170137 3315
rect 137385 2839 137419 3009
rect 151829 2907 151863 3077
rect 158637 2975 158671 3145
rect 153979 2805 154071 2839
rect 154037 2771 154071 2805
rect 158821 2771 158855 2941
rect 163421 2839 163455 3213
rect 169953 3179 169987 3281
rect 180257 2907 180291 3689
rect 357817 3383 357851 3893
rect 189733 2839 189767 3009
rect 314761 2975 314795 3349
rect 347697 3043 347731 3281
rect 349169 2975 349203 3281
rect 359381 3111 359415 3281
rect 163421 2805 163697 2839
rect 348341 2771 348375 2941
rect 350365 2771 350399 3077
rect 353861 2907 353895 3077
rect 359565 3043 359599 3349
rect 378609 3179 378643 3893
rect 378793 3859 378827 3893
rect 378793 3825 378885 3859
rect 378701 3179 378735 3825
rect 353861 2873 354045 2907
<< viali >>
rect 116685 568497 116719 568531
rect 115397 568021 115431 568055
rect 116685 567885 116719 567919
rect 116869 568225 116903 568259
rect 115397 567341 115431 567375
rect 116961 568157 116995 568191
rect 116961 567409 116995 567443
rect 116869 567273 116903 567307
rect 103437 524297 103471 524331
rect 113189 524297 113223 524331
rect 103161 524229 103195 524263
rect 108313 524229 108347 524263
rect 108313 524025 108347 524059
rect 105737 523889 105771 523923
rect 122757 524297 122791 524331
rect 122665 524229 122699 524263
rect 117973 524025 118007 524059
rect 121377 524025 121411 524059
rect 121377 523889 121411 523923
rect 117973 523821 118007 523855
rect 122665 523821 122699 523855
rect 113189 523617 113223 523651
rect 122757 523617 122791 523651
rect 132509 524297 132543 524331
rect 105737 523481 105771 523515
rect 142077 524297 142111 524331
rect 159189 524297 159223 524331
rect 159373 524297 159407 524331
rect 132601 524229 132635 524263
rect 141985 524229 142019 524263
rect 132601 523073 132635 523107
rect 137753 523209 137787 523243
rect 141985 523209 142019 523243
rect 137753 523073 137787 523107
rect 132509 523005 132543 523039
rect 156153 524229 156187 524263
rect 214021 524093 214055 524127
rect 243553 523957 243587 523991
rect 214021 523821 214055 523855
rect 243461 523821 243495 523855
rect 243553 523821 243587 523855
rect 243645 523957 243679 523991
rect 243645 523685 243679 523719
rect 243737 523685 243771 523719
rect 156153 523549 156187 523583
rect 147505 523345 147539 523379
rect 147505 523209 147539 523243
rect 147597 523209 147631 523243
rect 142077 523005 142111 523039
rect 147597 523005 147631 523039
rect 299489 502809 299523 502843
rect 289829 502673 289863 502707
rect 299489 502673 299523 502707
rect 309057 502809 309091 502843
rect 280169 502605 280203 502639
rect 280169 502469 280203 502503
rect 289645 502605 289679 502639
rect 289645 502333 289679 502367
rect 309057 502605 309091 502639
rect 311817 502605 311851 502639
rect 311909 502605 311943 502639
rect 289829 502333 289863 502367
rect 320649 495465 320683 495499
rect 320649 490909 320683 490943
rect 320649 489889 320683 489923
rect 320833 489821 320867 489855
rect 320833 487237 320867 487271
rect 320465 482817 320499 482851
rect 320465 480301 320499 480335
rect 320833 479417 320867 479451
rect 320833 478941 320867 478975
rect 320741 476017 320775 476051
rect 320741 470441 320775 470475
rect 320373 467789 320407 467823
rect 320373 467585 320407 467619
rect 320741 467517 320775 467551
rect 320833 475745 320867 475779
rect 320833 467381 320867 467415
rect 320281 457453 320315 457487
rect 320189 452285 320223 452319
rect 320741 457453 320775 457487
rect 320649 457317 320683 457351
rect 320373 456909 320407 456943
rect 320373 456637 320407 456671
rect 320649 452625 320683 452659
rect 320649 449837 320683 449871
rect 320373 447321 320407 447355
rect 320373 446981 320407 447015
rect 320833 456909 320867 456943
rect 320833 456501 320867 456535
rect 320741 447117 320775 447151
rect 320833 452625 320867 452659
rect 320833 447049 320867 447083
rect 320649 446913 320683 446947
rect 320281 446845 320315 446879
rect 320189 446777 320223 446811
rect 320741 381361 320775 381395
rect 320649 379729 320683 379763
rect 320741 379525 320775 379559
rect 320833 380273 320867 380307
rect 320649 378301 320683 378335
rect 298109 376737 298143 376771
rect 289737 376669 289771 376703
rect 289829 376669 289863 376703
rect 298109 376601 298143 376635
rect 302893 376737 302927 376771
rect 302893 376533 302927 376567
rect 320097 374629 320131 374663
rect 320833 374629 320867 374663
rect 320097 372929 320131 372963
rect 320465 372929 320499 372963
rect 320281 371025 320315 371059
rect 320281 367829 320315 367863
rect 320373 368577 320407 368611
rect 298109 367013 298143 367047
rect 292589 366945 292623 366979
rect 292497 366877 292531 366911
rect 298109 366877 298143 366911
rect 307769 366945 307803 366979
rect 307769 366809 307803 366843
rect 317429 366945 317463 366979
rect 317429 366265 317463 366299
rect 320833 371569 320867 371603
rect 320833 370481 320867 370515
rect 320465 363749 320499 363783
rect 320373 362661 320407 362695
rect 320281 360145 320315 360179
rect 320373 359873 320407 359907
rect 320281 355861 320315 355895
rect 224969 318869 225003 318903
rect 142905 318801 142939 318835
rect 152841 318801 152875 318835
rect 200589 318801 200623 318835
rect 142813 318665 142847 318699
rect 142905 318665 142939 318699
rect 145021 318665 145055 318699
rect 75101 318461 75135 318495
rect 74549 318121 74583 318155
rect 74365 318053 74399 318087
rect 75009 318053 75043 318087
rect 75101 318053 75135 318087
rect 75285 318393 75319 318427
rect 136925 318257 136959 318291
rect 84669 317985 84703 318019
rect 142721 318257 142755 318291
rect 142813 318257 142847 318291
rect 136925 317917 136959 317951
rect 138397 318121 138431 318155
rect 142721 317917 142755 317951
rect 141985 317849 142019 317883
rect 138397 317781 138431 317815
rect 138489 317781 138523 317815
rect 70409 317577 70443 317611
rect 84669 317577 84703 317611
rect 84761 317713 84795 317747
rect 84761 317577 84795 317611
rect 142813 317849 142847 317883
rect 142813 317713 142847 317747
rect 142905 317713 142939 317747
rect 141893 317645 141927 317679
rect 141985 317645 142019 317679
rect 138489 317441 138523 317475
rect 139317 317577 139351 317611
rect 70409 317305 70443 317339
rect 92857 317373 92891 317407
rect 70869 309145 70903 309179
rect 70869 307785 70903 307819
rect 94053 317373 94087 317407
rect 139317 317305 139351 317339
rect 140789 317577 140823 317611
rect 140789 317305 140823 317339
rect 148057 318665 148091 318699
rect 147505 318393 147539 318427
rect 147505 318257 147539 318291
rect 152749 318665 152783 318699
rect 152841 318665 152875 318699
rect 157257 318665 157291 318699
rect 150449 318393 150483 318427
rect 147689 318189 147723 318223
rect 148057 318189 148091 318223
rect 149253 318325 149287 318359
rect 146769 317917 146803 317951
rect 145021 317645 145055 317679
rect 145665 317713 145699 317747
rect 146769 317713 146803 317747
rect 147321 317849 147355 317883
rect 142905 317577 142939 317611
rect 141893 317305 141927 317339
rect 145665 317305 145699 317339
rect 154037 318393 154071 318427
rect 152749 318257 152783 318291
rect 153301 318325 153335 318359
rect 150449 318189 150483 318223
rect 148425 317781 148459 317815
rect 149253 317781 149287 317815
rect 151737 318121 151771 318155
rect 148425 317441 148459 317475
rect 152473 318053 152507 318087
rect 153301 318053 153335 318087
rect 151829 317917 151863 317951
rect 152473 317849 152507 317883
rect 151829 317781 151863 317815
rect 191021 318529 191055 318563
rect 200773 318733 200807 318767
rect 200589 318393 200623 318427
rect 200681 318461 200715 318495
rect 157257 318121 157291 318155
rect 190101 318257 190135 318291
rect 191021 318257 191055 318291
rect 195897 318257 195931 318291
rect 190009 318053 190043 318087
rect 154037 317577 154071 317611
rect 162133 317985 162167 318019
rect 151737 317441 151771 317475
rect 147689 317373 147723 317407
rect 147321 309145 147355 309179
rect 190009 317781 190043 317815
rect 190101 317781 190135 317815
rect 184949 317713 184983 317747
rect 200681 318121 200715 318155
rect 198933 318053 198967 318087
rect 199117 318053 199151 318087
rect 204913 318733 204947 318767
rect 201601 318665 201635 318699
rect 201601 318529 201635 318563
rect 195897 317645 195931 317679
rect 198013 317849 198047 317883
rect 200773 317849 200807 317883
rect 204177 318053 204211 318087
rect 184949 317509 184983 317543
rect 162133 309145 162167 309179
rect 193873 309213 193907 309247
rect 94053 307853 94087 307887
rect 92857 307785 92891 307819
rect 204177 317713 204211 317747
rect 198013 309145 198047 309179
rect 208593 318733 208627 318767
rect 213837 318733 213871 318767
rect 210433 318325 210467 318359
rect 210433 318053 210467 318087
rect 210525 318325 210559 318359
rect 208593 317985 208627 318019
rect 212089 318325 212123 318359
rect 212089 318121 212123 318155
rect 210525 317985 210559 318019
rect 212549 317713 212583 317747
rect 220093 318733 220127 318767
rect 215217 318665 215251 318699
rect 224877 318733 224911 318767
rect 224969 318733 225003 318767
rect 234353 318869 234387 318903
rect 220001 318461 220035 318495
rect 220093 318461 220127 318495
rect 222209 318665 222243 318699
rect 220001 318189 220035 318223
rect 215217 318121 215251 318155
rect 224693 318189 224727 318223
rect 222209 318121 222243 318155
rect 234353 317985 234387 318019
rect 213837 317441 213871 317475
rect 224877 317713 224911 317747
rect 212549 317373 212583 317407
rect 270509 317713 270543 317747
rect 224877 317373 224911 317407
rect 236193 317373 236227 317407
rect 204913 309145 204947 309179
rect 193873 307785 193907 307819
rect 236193 307785 236227 307819
rect 238953 317373 238987 317407
rect 270509 317373 270543 317407
rect 280077 317713 280111 317747
rect 289829 317713 289863 317747
rect 289829 317441 289863 317475
rect 299397 317713 299431 317747
rect 309149 317713 309183 317747
rect 309149 317577 309183 317611
rect 299397 317441 299431 317475
rect 280077 317373 280111 317407
rect 251281 309553 251315 309587
rect 238953 307785 238987 307819
rect 245577 309077 245611 309111
rect 94053 307717 94087 307751
rect 70501 299421 70535 299455
rect 94053 298129 94087 298163
rect 105093 302209 105127 302243
rect 251281 306901 251315 306935
rect 254041 309077 254075 309111
rect 245577 299489 245611 299523
rect 324973 309077 325007 309111
rect 267105 303569 267139 303603
rect 265817 302141 265851 302175
rect 254041 299489 254075 299523
rect 255237 299489 255271 299523
rect 105093 298129 105127 298163
rect 151093 299421 151127 299455
rect 70501 289833 70535 289867
rect 70777 298061 70811 298095
rect 70777 288405 70811 288439
rect 72157 296633 72191 296667
rect 227361 299421 227395 299455
rect 151093 289833 151127 289867
rect 193873 298061 193907 298095
rect 251281 299421 251315 299455
rect 242633 298061 242667 298095
rect 227361 289833 227395 289867
rect 235733 296633 235767 296667
rect 193873 288405 193907 288439
rect 72157 288337 72191 288371
rect 242633 288405 242667 288439
rect 243921 298061 243955 298095
rect 243921 288405 243955 288439
rect 246957 298061 246991 298095
rect 246957 288405 246991 288439
rect 248245 298061 248279 298095
rect 255237 298129 255271 298163
rect 251281 297245 251315 297279
rect 255237 297993 255271 298027
rect 248245 288405 248279 288439
rect 259285 297449 259319 297483
rect 324973 299489 325007 299523
rect 267105 299421 267139 299455
rect 271521 299421 271555 299455
rect 271521 293505 271555 293539
rect 265817 292621 265851 292655
rect 259285 289833 259319 289867
rect 255237 288405 255271 288439
rect 324973 289765 325007 289799
rect 235733 287113 235767 287147
rect 267197 287725 267231 287759
rect 78873 282897 78907 282931
rect 267197 282897 267231 282931
rect 324973 280177 325007 280211
rect 78873 278749 78907 278783
rect 105185 280109 105219 280143
rect 90005 273309 90039 273343
rect 106657 280109 106691 280143
rect 106657 273241 106691 273275
rect 151093 280109 151127 280143
rect 105185 273105 105219 273139
rect 243829 278817 243863 278851
rect 243829 277389 243863 277423
rect 151093 270521 151127 270555
rect 264621 274601 264655 274635
rect 90005 267733 90039 267767
rect 105185 270453 105219 270487
rect 105185 263449 105219 263483
rect 106841 270453 106875 270487
rect 249625 270453 249659 270487
rect 106841 260865 106875 260899
rect 234077 270385 234111 270419
rect 234077 260865 234111 260899
rect 249625 260865 249659 260899
rect 251005 270453 251039 270487
rect 251005 260865 251039 260899
rect 252293 270453 252327 270487
rect 252293 260865 252327 260899
rect 259285 270453 259319 270487
rect 268669 273241 268703 273275
rect 268669 267733 268703 267767
rect 324973 270453 325007 270487
rect 264621 264945 264655 264979
rect 259285 260865 259319 260899
rect 324973 260865 325007 260899
rect 105185 260797 105219 260831
rect 70777 259369 70811 259403
rect 105185 253793 105219 253827
rect 151093 260797 151127 260831
rect 70777 241485 70811 241519
rect 73445 252569 73479 252603
rect 151093 251209 151127 251243
rect 105093 251141 105127 251175
rect 73445 241485 73479 241519
rect 94053 244953 94087 244987
rect 70777 234549 70811 234583
rect 70777 231829 70811 231863
rect 105093 241485 105127 241519
rect 252293 251141 252327 251175
rect 324789 251073 324823 251107
rect 324789 241553 324823 241587
rect 252293 241485 252327 241519
rect 324881 241417 324915 241451
rect 324881 234617 324915 234651
rect 94053 231829 94087 231863
rect 266001 230469 266035 230503
rect 106473 230401 106507 230435
rect 78781 229041 78815 229075
rect 77493 225641 77527 225675
rect 105093 224961 105127 224995
rect 105093 222173 105127 222207
rect 106473 220881 106507 220915
rect 78781 219453 78815 219487
rect 91017 220677 91051 220711
rect 77493 217345 77527 217379
rect 70777 215237 70811 215271
rect 70777 212517 70811 212551
rect 266001 218025 266035 218059
rect 91017 212449 91051 212483
rect 233801 216597 233835 216631
rect 91017 211089 91051 211123
rect 77493 205649 77527 205683
rect 77493 202861 77527 202895
rect 233801 208369 233835 208403
rect 235549 209729 235583 209763
rect 105093 205649 105127 205683
rect 105093 202861 105127 202895
rect 91017 202793 91051 202827
rect 94053 202793 94087 202827
rect 70777 195925 70811 195959
rect 70777 193205 70811 193239
rect 235549 200141 235583 200175
rect 252293 201433 252327 201467
rect 94053 193205 94087 193239
rect 252293 191845 252327 191879
rect 264621 192525 264655 192559
rect 78781 186337 78815 186371
rect 105093 186337 105127 186371
rect 264621 185657 264655 185691
rect 78781 183549 78815 183583
rect 91017 183549 91051 183583
rect 105093 183549 105127 183583
rect 77493 183481 77527 183515
rect 70777 176613 70811 176647
rect 70777 173893 70811 173927
rect 72341 174029 72375 174063
rect 91017 180829 91051 180863
rect 235641 180761 235675 180795
rect 77493 173893 77527 173927
rect 91017 178653 91051 178687
rect 72341 171105 72375 171139
rect 91017 171105 91051 171139
rect 266001 179333 266035 179367
rect 235641 171105 235675 171139
rect 242541 172465 242575 172499
rect 106657 164169 106691 164203
rect 81909 161381 81943 161415
rect 70685 157437 70719 157471
rect 70685 154581 70719 154615
rect 73445 153153 73479 153187
rect 73445 144857 73479 144891
rect 106657 157301 106691 157335
rect 151093 164169 151127 164203
rect 94053 156621 94087 156655
rect 211905 164169 211939 164203
rect 151093 154581 151127 154615
rect 193873 162809 193907 162843
rect 211905 157301 211939 157335
rect 227361 164169 227395 164203
rect 266001 169745 266035 169779
rect 267289 179333 267323 179367
rect 267289 169745 267323 169779
rect 242541 162877 242575 162911
rect 264621 169677 264655 169711
rect 227361 157301 227395 157335
rect 234169 161381 234203 161415
rect 193873 153221 193907 153255
rect 243829 161381 243863 161415
rect 234169 151793 234203 151827
rect 242541 153153 242575 153187
rect 94053 146965 94087 146999
rect 81909 144789 81943 144823
rect 106657 144857 106691 144891
rect 105093 143497 105127 143531
rect 73537 143429 73571 143463
rect 72341 133841 72375 133875
rect 105093 137921 105127 137955
rect 106657 137921 106691 137955
rect 151093 144857 151127 144891
rect 211905 144857 211939 144891
rect 151093 135269 151127 135303
rect 193873 143497 193907 143531
rect 211905 137921 211939 137955
rect 227361 144857 227395 144891
rect 264621 160089 264655 160123
rect 243829 151793 243863 151827
rect 266001 160021 266035 160055
rect 266001 150433 266035 150467
rect 267289 160021 267323 160055
rect 267289 150433 267323 150467
rect 242541 143565 242575 143599
rect 227361 137921 227395 137955
rect 234169 142069 234203 142103
rect 193873 133909 193907 133943
rect 73537 131529 73571 131563
rect 72341 124185 72375 124219
rect 151093 125545 151127 125579
rect 105093 124117 105127 124151
rect 78781 115889 78815 115923
rect 106473 124049 106507 124083
rect 211905 125545 211939 125579
rect 151093 115957 151127 115991
rect 193873 124117 193907 124151
rect 106473 114597 106507 114631
rect 105093 114529 105127 114563
rect 211905 118609 211939 118643
rect 227361 125545 227395 125579
rect 266001 140709 266035 140743
rect 234169 124185 234203 124219
rect 242541 133841 242575 133875
rect 242541 124185 242575 124219
rect 243829 133773 243863 133807
rect 266001 131121 266035 131155
rect 267289 140709 267323 140743
rect 267289 131121 267323 131155
rect 243829 124185 243863 124219
rect 252293 124117 252327 124151
rect 243829 122757 243863 122791
rect 227361 118609 227395 118643
rect 234261 119357 234295 119391
rect 234261 114597 234295 114631
rect 193873 114529 193907 114563
rect 78781 106301 78815 106335
rect 90925 114461 90959 114495
rect 72249 106233 72283 106267
rect 70777 104805 70811 104839
rect 72249 96713 72283 96747
rect 73537 106233 73571 106267
rect 70777 95285 70811 95319
rect 234169 114461 234203 114495
rect 90925 104873 90959 104907
rect 151093 106233 151127 106267
rect 73537 95217 73571 95251
rect 94053 104805 94087 104839
rect 94053 95217 94087 95251
rect 105093 104805 105127 104839
rect 105093 95217 105127 95251
rect 106657 103445 106691 103479
rect 211905 106233 211939 106267
rect 151093 96645 151127 96679
rect 193873 104805 193907 104839
rect 211905 99297 211939 99331
rect 227361 106233 227395 106267
rect 234169 104873 234203 104907
rect 242541 114461 242575 114495
rect 252293 114529 252327 114563
rect 255237 124117 255271 124151
rect 243829 113169 243863 113203
rect 268669 122757 268703 122791
rect 266001 121397 266035 121431
rect 266001 111809 266035 111843
rect 267381 121397 267415 121431
rect 268669 113169 268703 113203
rect 267381 111809 267415 111843
rect 255237 106301 255271 106335
rect 264621 111673 264655 111707
rect 242541 104873 242575 104907
rect 246957 104805 246991 104839
rect 227361 99297 227395 99331
rect 234169 100045 234203 100079
rect 193873 95217 193907 95251
rect 234169 95217 234203 95251
rect 235733 96577 235767 96611
rect 106657 93857 106691 93891
rect 78689 93789 78723 93823
rect 72157 85493 72191 85527
rect 72157 75905 72191 75939
rect 73445 85493 73479 85527
rect 73445 75905 73479 75939
rect 77493 85493 77527 85527
rect 234169 91749 234203 91783
rect 106657 89777 106691 89811
rect 90005 86853 90039 86887
rect 78689 84269 78723 84303
rect 81725 85493 81759 85527
rect 77493 75905 77527 75939
rect 78689 82773 78723 82807
rect 72157 72437 72191 72471
rect 72157 67677 72191 67711
rect 70685 67541 70719 67575
rect 70685 57953 70719 57987
rect 72065 66181 72099 66215
rect 90005 77265 90039 77299
rect 92765 86853 92799 86887
rect 234169 87057 234203 87091
rect 246957 95217 246991 95251
rect 252109 104805 252143 104839
rect 252109 95217 252143 95251
rect 255237 104805 255271 104839
rect 235733 86989 235767 87023
rect 242541 95149 242575 95183
rect 106657 85561 106691 85595
rect 151093 86921 151127 86955
rect 94053 85493 94087 85527
rect 105093 85493 105127 85527
rect 105093 84133 105127 84167
rect 94053 80937 94087 80971
rect 92765 77265 92799 77299
rect 211905 86921 211939 86955
rect 151093 77265 151127 77299
rect 193873 85493 193907 85527
rect 81725 75905 81759 75939
rect 193873 75905 193907 75939
rect 204729 85493 204763 85527
rect 211905 77265 211939 77299
rect 227361 86921 227395 86955
rect 259285 104805 259319 104839
rect 264621 102153 264655 102187
rect 268577 103445 268611 103479
rect 259285 95217 259319 95251
rect 266001 102085 266035 102119
rect 266001 92497 266035 92531
rect 267289 102085 267323 102119
rect 268577 93857 268611 93891
rect 267289 92497 267323 92531
rect 255237 86989 255271 87023
rect 264621 92361 264655 92395
rect 242541 85561 242575 85595
rect 227361 77265 227395 77299
rect 234169 85493 234203 85527
rect 204729 75905 204763 75939
rect 246957 85493 246991 85527
rect 234169 75905 234203 75939
rect 235733 77197 235767 77231
rect 106473 75837 106507 75871
rect 105001 74545 105035 74579
rect 94145 74477 94179 74511
rect 78689 64889 78723 64923
rect 90005 67541 90039 67575
rect 90005 58021 90039 58055
rect 92765 67541 92799 67575
rect 211905 75837 211939 75871
rect 211905 70329 211939 70363
rect 246957 75905 246991 75939
rect 252293 85493 252327 85527
rect 252293 75905 252327 75939
rect 255237 85493 255271 85527
rect 255237 75905 255271 75939
rect 259285 85493 259319 85527
rect 264621 82841 264655 82875
rect 259285 75905 259319 75939
rect 266001 82773 266035 82807
rect 235733 67609 235767 67643
rect 242541 75837 242575 75871
rect 106473 66317 106507 66351
rect 151093 67541 151127 67575
rect 105001 66249 105035 66283
rect 94145 64889 94179 64923
rect 92765 58021 92799 58055
rect 94145 59993 94179 60027
rect 72065 56593 72099 56627
rect 90925 56661 90959 56695
rect 90925 55233 90959 55267
rect 81725 51765 81759 51799
rect 72065 46869 72099 46903
rect 72065 37281 72099 37315
rect 73445 46869 73479 46903
rect 266001 73185 266035 73219
rect 267289 82773 267323 82807
rect 267289 73185 267323 73219
rect 324973 77197 325007 77231
rect 324973 67609 325007 67643
rect 242541 66249 242575 66283
rect 151093 57953 151127 57987
rect 193873 66181 193907 66215
rect 193873 56593 193907 56627
rect 204913 66181 204947 66215
rect 234077 66181 234111 66215
rect 204913 56593 204947 56627
rect 211905 57885 211939 57919
rect 94145 50609 94179 50643
rect 96997 56525 97031 56559
rect 227361 57885 227395 57919
rect 246957 66181 246991 66215
rect 234077 57817 234111 57851
rect 235733 57885 235767 57919
rect 227361 51017 227395 51051
rect 211905 50677 211939 50711
rect 246957 56593 246991 56627
rect 252293 66181 252327 66215
rect 252293 56593 252327 56627
rect 255237 66181 255271 66215
rect 255237 56593 255271 56627
rect 259285 66181 259319 66215
rect 259285 56593 259319 56627
rect 267289 63461 267323 63495
rect 235733 48297 235767 48331
rect 242541 56525 242575 56559
rect 96997 47005 97031 47039
rect 151093 48229 151127 48263
rect 73445 37281 73479 37315
rect 78781 38641 78815 38675
rect 81725 38641 81759 38675
rect 96997 46869 97031 46903
rect 78781 37281 78815 37315
rect 267289 53805 267323 53839
rect 242541 46937 242575 46971
rect 264621 53737 264655 53771
rect 151093 38641 151127 38675
rect 193873 46869 193907 46903
rect 96997 37281 97031 37315
rect 106841 38573 106875 38607
rect 73445 36261 73479 36295
rect 106841 31569 106875 31603
rect 73445 28985 73479 29019
rect 204913 46869 204947 46903
rect 234077 46869 234111 46903
rect 234077 38641 234111 38675
rect 246957 46869 246991 46903
rect 204913 37281 204947 37315
rect 211905 38573 211939 38607
rect 193873 28985 193907 29019
rect 211905 28985 211939 29019
rect 235733 38573 235767 38607
rect 246957 37281 246991 37315
rect 251005 46869 251039 46903
rect 251005 37281 251039 37315
rect 252293 46869 252327 46903
rect 252293 37281 252327 37315
rect 255237 46869 255271 46903
rect 255237 37281 255271 37315
rect 259285 46869 259319 46903
rect 264621 44285 264655 44319
rect 324881 46869 324915 46903
rect 259285 37281 259319 37315
rect 267289 44081 267323 44115
rect 235733 28985 235767 29019
rect 242541 37213 242575 37247
rect 90005 28917 90039 28951
rect 77493 27557 77527 27591
rect 77493 17969 77527 18003
rect 78873 27557 78907 27591
rect 96997 28917 97031 28951
rect 90005 19329 90039 19363
rect 91109 27557 91143 27591
rect 78873 17969 78907 18003
rect 96997 21913 97031 21947
rect 151093 28917 151127 28951
rect 324881 38505 324915 38539
rect 267289 35785 267323 35819
rect 261953 33133 261987 33167
rect 261953 29665 261987 29699
rect 242541 27625 242575 27659
rect 151093 19329 151127 19363
rect 204913 27557 204947 27591
rect 91109 17969 91143 18003
rect 193781 19261 193815 19295
rect 73353 17901 73387 17935
rect 248245 27557 248279 27591
rect 204913 17969 204947 18003
rect 227361 19261 227395 19295
rect 193781 12393 193815 12427
rect 235733 19261 235767 19295
rect 248245 17969 248279 18003
rect 249625 27557 249659 27591
rect 249625 17969 249659 18003
rect 255237 27557 255271 27591
rect 260389 26197 260423 26231
rect 255237 17969 255271 18003
rect 259193 22729 259227 22763
rect 235733 15861 235767 15895
rect 259193 13141 259227 13175
rect 227361 11849 227395 11883
rect 255145 13073 255179 13107
rect 260389 13073 260423 13107
rect 255145 11033 255179 11067
rect 73353 8313 73387 8347
rect 94237 9605 94271 9639
rect 81633 4097 81667 4131
rect 70685 3893 70719 3927
rect 70501 3757 70535 3791
rect 70317 3621 70351 3655
rect 70409 3621 70443 3655
rect 79977 3893 80011 3927
rect 81633 3893 81667 3927
rect 89177 4029 89211 4063
rect 76205 3757 76239 3791
rect 70685 3689 70719 3723
rect 73721 3689 73755 3723
rect 70501 3417 70535 3451
rect 71513 3417 71547 3451
rect 45385 3349 45419 3383
rect 55229 3349 55263 3383
rect 45477 3281 45511 3315
rect 45477 3077 45511 3111
rect 45385 3009 45419 3043
rect 64797 3349 64831 3383
rect 55321 3281 55355 3315
rect 64613 3281 64647 3315
rect 62313 3077 62347 3111
rect 55321 3009 55355 3043
rect 61117 3009 61151 3043
rect 55229 2805 55263 2839
rect 62313 2737 62347 2771
rect 61117 2669 61151 2703
rect 64705 3213 64739 3247
rect 71881 3213 71915 3247
rect 64797 2805 64831 2839
rect 64705 2737 64739 2771
rect 64613 2669 64647 2703
rect 75101 3213 75135 3247
rect 75193 3417 75227 3451
rect 75285 3417 75319 3451
rect 76205 3417 76239 3451
rect 79885 3689 79919 3723
rect 79977 3689 80011 3723
rect 82461 3825 82495 3859
rect 79977 3417 80011 3451
rect 82461 3349 82495 3383
rect 75193 3213 75227 3247
rect 91569 4029 91603 4063
rect 89177 3213 89211 3247
rect 89269 3961 89303 3995
rect 91661 4029 91695 4063
rect 91661 3757 91695 3791
rect 91477 3349 91511 3383
rect 91569 3349 91603 3383
rect 91477 3213 91511 3247
rect 89269 3145 89303 3179
rect 238861 9605 238895 9639
rect 161305 8925 161339 8959
rect 161305 8789 161339 8823
rect 167009 8789 167043 8823
rect 167009 8585 167043 8619
rect 176577 8789 176611 8823
rect 176577 8585 176611 8619
rect 186329 8789 186363 8823
rect 195897 8789 195931 8823
rect 186329 8381 186363 8415
rect 193229 8585 193263 8619
rect 239413 9605 239447 9639
rect 239321 9537 239355 9571
rect 239229 9401 239263 9435
rect 239321 9401 239355 9435
rect 239413 9333 239447 9367
rect 239505 9469 239539 9503
rect 239229 8857 239263 8891
rect 238861 8653 238895 8687
rect 244841 9469 244875 9503
rect 246681 9469 246715 9503
rect 246681 9265 246715 9299
rect 248981 9197 249015 9231
rect 249165 9333 249199 9367
rect 249257 9333 249291 9367
rect 249441 9401 249475 9435
rect 244841 8721 244875 8755
rect 248981 8857 249015 8891
rect 239505 8517 239539 8551
rect 195805 8449 195839 8483
rect 196081 8449 196115 8483
rect 193229 8245 193263 8279
rect 215125 8449 215159 8483
rect 196081 8245 196115 8279
rect 197185 8381 197219 8415
rect 197185 8177 197219 8211
rect 202889 8381 202923 8415
rect 205557 8381 205591 8415
rect 205649 8381 205683 8415
rect 205465 8313 205499 8347
rect 205741 8313 205775 8347
rect 202889 8177 202923 8211
rect 215401 8449 215435 8483
rect 248981 8449 249015 8483
rect 249073 8789 249107 8823
rect 249349 9265 249383 9299
rect 249257 9061 249291 9095
rect 249349 8721 249383 8755
rect 249257 8653 249291 8687
rect 259009 9401 259043 9435
rect 258733 9333 258767 9367
rect 254961 9265 254995 9299
rect 254961 8857 254995 8891
rect 255053 9129 255087 9163
rect 259009 9129 259043 9163
rect 259101 9129 259135 9163
rect 255053 8857 255087 8891
rect 258641 8857 258675 8891
rect 258733 8857 258767 8891
rect 249441 8653 249475 8687
rect 249165 8517 249199 8551
rect 249073 8449 249107 8483
rect 215217 8381 215251 8415
rect 215217 8041 215251 8075
rect 215309 8381 215343 8415
rect 215309 8041 215343 8075
rect 215125 7973 215159 8007
rect 215401 7973 215435 8007
rect 161213 7429 161247 7463
rect 157349 5525 157383 5559
rect 157349 4777 157383 4811
rect 132509 4233 132543 4267
rect 127909 4165 127943 4199
rect 127449 3961 127483 3995
rect 127817 3961 127851 3995
rect 127725 3893 127759 3927
rect 127725 3621 127759 3655
rect 127817 3621 127851 3655
rect 123217 3553 123251 3587
rect 123585 3553 123619 3587
rect 127541 3485 127575 3519
rect 122021 3349 122055 3383
rect 122021 3145 122055 3179
rect 127633 3485 127667 3519
rect 127633 3281 127667 3315
rect 132509 4029 132543 4063
rect 136189 4165 136223 4199
rect 157349 4165 157383 4199
rect 153669 4097 153703 4131
rect 153945 4097 153979 4131
rect 157257 4097 157291 4131
rect 153025 4029 153059 4063
rect 127909 3349 127943 3383
rect 132969 3485 133003 3519
rect 136189 3485 136223 3519
rect 138673 3485 138707 3519
rect 127817 3213 127851 3247
rect 127909 3213 127943 3247
rect 94237 2873 94271 2907
rect 133061 3417 133095 3451
rect 133061 2941 133095 2975
rect 137385 3009 137419 3043
rect 138673 3009 138707 3043
rect 148885 3485 148919 3519
rect 149069 3349 149103 3383
rect 148885 3009 148919 3043
rect 148977 3213 149011 3247
rect 149069 3213 149103 3247
rect 155233 3893 155267 3927
rect 155233 3349 155267 3383
rect 153025 3145 153059 3179
rect 157349 4029 157383 4063
rect 201601 7021 201635 7055
rect 162133 6613 162167 6647
rect 171793 4777 171827 4811
rect 171793 4165 171827 4199
rect 181453 4777 181487 4811
rect 181453 4165 181487 4199
rect 195897 4777 195931 4811
rect 164801 4029 164835 4063
rect 157257 3145 157291 3179
rect 158637 3145 158671 3179
rect 161213 3145 161247 3179
rect 162041 3281 162075 3315
rect 162133 3281 162167 3315
rect 162409 3553 162443 3587
rect 195897 3961 195931 3995
rect 195989 4777 196023 4811
rect 205189 7021 205223 7055
rect 241437 6885 241471 6919
rect 215217 4777 215251 4811
rect 215401 4777 215435 4811
rect 212365 4505 212399 4539
rect 211721 4437 211755 4471
rect 229569 4777 229603 4811
rect 215309 4709 215343 4743
rect 215493 4709 215527 4743
rect 219357 4709 219391 4743
rect 223037 4709 223071 4743
rect 215401 4505 215435 4539
rect 219081 4505 219115 4539
rect 219173 4641 219207 4675
rect 223037 4573 223071 4607
rect 219173 4505 219207 4539
rect 229753 4777 229787 4811
rect 229753 4573 229787 4607
rect 239137 4709 239171 4743
rect 215217 4437 215251 4471
rect 225889 4437 225923 4471
rect 229569 4437 229603 4471
rect 229661 4505 229695 4539
rect 205189 4369 205223 4403
rect 201601 4301 201635 4335
rect 204821 4301 204855 4335
rect 205373 4233 205407 4267
rect 225889 4233 225923 4267
rect 234629 4505 234663 4539
rect 239137 4505 239171 4539
rect 239229 4641 239263 4675
rect 234445 4437 234479 4471
rect 239229 4437 239263 4471
rect 239413 4505 239447 4539
rect 231961 4369 231995 4403
rect 232605 4369 232639 4403
rect 232697 4369 232731 4403
rect 231869 4233 231903 4267
rect 229661 4165 229695 4199
rect 239413 4165 239447 4199
rect 249625 6885 249659 6919
rect 249441 5457 249475 5491
rect 247877 5117 247911 5151
rect 247877 4709 247911 4743
rect 248889 5049 248923 5083
rect 244105 4369 244139 4403
rect 244381 4369 244415 4403
rect 249349 4981 249383 5015
rect 258733 5321 258767 5355
rect 254869 5049 254903 5083
rect 254869 4777 254903 4811
rect 255053 4981 255087 5015
rect 257445 4981 257479 5015
rect 257445 4777 257479 4811
rect 257537 4913 257571 4947
rect 258273 4913 258307 4947
rect 258089 4845 258123 4879
rect 257537 4777 257571 4811
rect 255053 4709 255087 4743
rect 258825 5321 258859 5355
rect 258825 5117 258859 5151
rect 268485 5117 268519 5151
rect 268025 4981 268059 5015
rect 268301 4981 268335 5015
rect 268485 4845 268519 4879
rect 258733 4573 258767 4607
rect 249625 4505 249659 4539
rect 249441 4369 249475 4403
rect 249349 4301 249383 4335
rect 248889 4233 248923 4267
rect 241437 4165 241471 4199
rect 195989 3961 196023 3995
rect 340153 4097 340187 4131
rect 340153 3961 340187 3995
rect 369041 4097 369075 4131
rect 357817 3893 357851 3927
rect 369225 3893 369259 3927
rect 180257 3689 180291 3723
rect 164801 3349 164835 3383
rect 169033 3553 169067 3587
rect 162409 3213 162443 3247
rect 162501 3213 162535 3247
rect 163421 3213 163455 3247
rect 169033 3213 169067 3247
rect 170137 3281 170171 3315
rect 148977 3009 149011 3043
rect 151829 3077 151863 3111
rect 158637 2941 158671 2975
rect 158821 2941 158855 2975
rect 151829 2873 151863 2907
rect 137385 2805 137419 2839
rect 153945 2805 153979 2839
rect 132969 2737 133003 2771
rect 154037 2737 154071 2771
rect 169953 3145 169987 3179
rect 314761 3349 314795 3383
rect 357817 3349 357851 3383
rect 359565 3349 359599 3383
rect 180257 2873 180291 2907
rect 189733 3009 189767 3043
rect 347697 3281 347731 3315
rect 347697 3009 347731 3043
rect 349169 3281 349203 3315
rect 359381 3281 359415 3315
rect 314761 2941 314795 2975
rect 348341 2941 348375 2975
rect 349169 2941 349203 2975
rect 350365 3077 350399 3111
rect 163697 2805 163731 2839
rect 189733 2805 189767 2839
rect 158821 2737 158855 2771
rect 348341 2737 348375 2771
rect 353861 3077 353895 3111
rect 359381 3077 359415 3111
rect 378609 3145 378643 3179
rect 378701 3825 378735 3859
rect 378885 3825 378919 3859
rect 378701 3145 378735 3179
rect 359565 3009 359599 3043
rect 354045 2873 354079 2907
rect 350365 2737 350399 2771
rect 73721 969 73755 1003
<< metal1 >>
rect 156598 655528 156604 655580
rect 156656 655568 156662 655580
rect 187694 655568 187700 655580
rect 156656 655540 187700 655568
rect 156656 655528 156662 655540
rect 187694 655528 187700 655540
rect 187752 655528 187758 655580
rect 95142 568488 95148 568540
rect 95200 568528 95206 568540
rect 103146 568528 103152 568540
rect 95200 568500 103152 568528
rect 95200 568488 95206 568500
rect 103146 568488 103152 568500
rect 103204 568488 103210 568540
rect 116673 568531 116731 568537
rect 116673 568497 116685 568531
rect 116719 568528 116731 568531
rect 119430 568528 119436 568540
rect 116719 568500 119436 568528
rect 116719 568497 116731 568500
rect 116673 568491 116731 568497
rect 119430 568488 119436 568500
rect 119488 568528 119494 568540
rect 128446 568528 128452 568540
rect 119488 568500 128452 568528
rect 119488 568488 119494 568500
rect 128446 568488 128452 568500
rect 128504 568488 128510 568540
rect 132402 568488 132408 568540
rect 132460 568528 132466 568540
rect 209590 568528 209596 568540
rect 132460 568500 209596 568528
rect 132460 568488 132466 568500
rect 209590 568488 209596 568500
rect 209648 568488 209654 568540
rect 110322 568420 110328 568472
rect 110380 568460 110386 568472
rect 135898 568460 135904 568472
rect 110380 568432 135904 568460
rect 110380 568420 110386 568432
rect 135898 568420 135904 568432
rect 135956 568420 135962 568472
rect 117958 568352 117964 568404
rect 118016 568392 118022 568404
rect 137278 568392 137284 568404
rect 118016 568364 137284 568392
rect 118016 568352 118022 568364
rect 137278 568352 137284 568364
rect 137336 568352 137342 568404
rect 98362 568284 98368 568336
rect 98420 568324 98426 568336
rect 107746 568324 107752 568336
rect 98420 568296 107752 568324
rect 98420 568284 98426 568296
rect 107746 568284 107752 568296
rect 107804 568324 107810 568336
rect 117130 568324 117136 568336
rect 107804 568296 117136 568324
rect 107804 568284 107810 568296
rect 117130 568284 117136 568296
rect 117188 568284 117194 568336
rect 120994 568284 121000 568336
rect 121052 568324 121058 568336
rect 140038 568324 140044 568336
rect 121052 568296 140044 568324
rect 121052 568284 121058 568296
rect 140038 568284 140044 568296
rect 140096 568284 140102 568336
rect 217134 568284 217140 568336
rect 217192 568324 217198 568336
rect 225874 568324 225880 568336
rect 217192 568296 225880 568324
rect 217192 568284 217198 568296
rect 225874 568284 225880 568296
rect 225932 568324 225938 568336
rect 234614 568324 234620 568336
rect 225932 568296 234620 568324
rect 225932 568284 225938 568296
rect 234614 568284 234620 568296
rect 234672 568284 234678 568336
rect 100662 568216 100668 568268
rect 100720 568256 100726 568268
rect 109034 568256 109040 568268
rect 100720 568228 109040 568256
rect 100720 568216 100726 568228
rect 109034 568216 109040 568228
rect 109092 568256 109098 568268
rect 116857 568259 116915 568265
rect 116857 568256 116869 568259
rect 109092 568228 116869 568256
rect 109092 568216 109098 568228
rect 116857 568225 116869 568228
rect 116903 568225 116915 568259
rect 124306 568256 124312 568268
rect 116857 568219 116915 568225
rect 117056 568228 124312 568256
rect 97902 568148 97908 568200
rect 97960 568188 97966 568200
rect 106642 568188 106648 568200
rect 97960 568160 106648 568188
rect 97960 568148 97966 568160
rect 106642 568148 106648 568160
rect 106700 568188 106706 568200
rect 115842 568188 115848 568200
rect 106700 568160 115848 568188
rect 106700 568148 106706 568160
rect 115842 568148 115848 568160
rect 115900 568188 115906 568200
rect 116949 568191 117007 568197
rect 116949 568188 116961 568191
rect 115900 568160 116961 568188
rect 115900 568148 115906 568160
rect 116949 568157 116961 568160
rect 116995 568157 117007 568191
rect 116949 568151 117007 568157
rect 93762 568080 93768 568132
rect 93820 568120 93826 568132
rect 101766 568120 101772 568132
rect 93820 568092 101772 568120
rect 93820 568080 93826 568092
rect 101766 568080 101772 568092
rect 101824 568120 101830 568132
rect 110690 568120 110696 568132
rect 101824 568092 110696 568120
rect 101824 568080 101830 568092
rect 110690 568080 110696 568092
rect 110748 568080 110754 568132
rect 103146 568012 103152 568064
rect 103204 568052 103210 568064
rect 112254 568052 112260 568064
rect 103204 568024 112260 568052
rect 103204 568012 103210 568024
rect 112254 568012 112260 568024
rect 112312 568052 112318 568064
rect 115385 568055 115443 568061
rect 115385 568052 115397 568055
rect 112312 568024 115397 568052
rect 112312 568012 112318 568024
rect 115385 568021 115397 568024
rect 115431 568021 115443 568055
rect 115385 568015 115443 568021
rect 96522 567944 96528 567996
rect 96580 567984 96586 567996
rect 105262 567984 105268 567996
rect 96580 567956 105268 567984
rect 96580 567944 96586 567956
rect 105262 567944 105268 567956
rect 105320 567984 105326 567996
rect 114738 567984 114744 567996
rect 105320 567956 114744 567984
rect 105320 567944 105326 567956
rect 114738 567944 114744 567956
rect 114796 567984 114802 567996
rect 117056 567984 117084 568228
rect 124306 568216 124312 568228
rect 124364 568216 124370 568268
rect 126606 568256 126612 568268
rect 124508 568228 126612 568256
rect 117130 568148 117136 568200
rect 117188 568188 117194 568200
rect 124508 568188 124536 568228
rect 126606 568216 126612 568228
rect 126664 568256 126670 568268
rect 144914 568256 144920 568268
rect 126664 568228 144920 568256
rect 126664 568216 126670 568228
rect 144914 568216 144920 568228
rect 144972 568216 144978 568268
rect 215570 568216 215576 568268
rect 215628 568256 215634 568268
rect 224770 568256 224776 568268
rect 215628 568228 224776 568256
rect 215628 568216 215634 568228
rect 224770 568216 224776 568228
rect 224828 568256 224834 568268
rect 233234 568256 233240 568268
rect 224828 568228 233240 568256
rect 224828 568216 224834 568228
rect 233234 568216 233240 568228
rect 233292 568216 233298 568268
rect 117188 568160 124536 568188
rect 117188 568148 117194 568160
rect 128446 568148 128452 568200
rect 128504 568188 128510 568200
rect 149054 568188 149060 568200
rect 128504 568160 149060 568188
rect 128504 568148 128510 568160
rect 149054 568148 149060 568160
rect 149112 568148 149118 568200
rect 209590 568148 209596 568200
rect 209648 568188 209654 568200
rect 218974 568188 218980 568200
rect 209648 568160 218980 568188
rect 209648 568148 209654 568160
rect 218974 568148 218980 568160
rect 219032 568188 219038 568200
rect 228358 568188 228364 568200
rect 219032 568160 228364 568188
rect 219032 568148 219038 568160
rect 228358 568148 228364 568160
rect 228416 568188 228422 568200
rect 237374 568188 237380 568200
rect 228416 568160 237380 568188
rect 228416 568148 228422 568160
rect 237374 568148 237380 568160
rect 237432 568148 237438 568200
rect 123478 568120 123484 568132
rect 114796 567956 117084 567984
rect 117976 568092 123484 568120
rect 114796 567944 114802 567956
rect 102042 567876 102048 567928
rect 102100 567916 102106 567928
rect 109862 567916 109868 567928
rect 102100 567888 109868 567916
rect 102100 567876 102106 567888
rect 109862 567876 109868 567888
rect 109920 567916 109926 567928
rect 116673 567919 116731 567925
rect 116673 567916 116685 567919
rect 109920 567888 116685 567916
rect 109920 567876 109926 567888
rect 116673 567885 116685 567888
rect 116719 567885 116731 567919
rect 116673 567879 116731 567885
rect 94866 567808 94872 567860
rect 94924 567848 94930 567860
rect 104066 567848 104072 567860
rect 94924 567820 104072 567848
rect 94924 567808 94930 567820
rect 104066 567808 104072 567820
rect 104124 567848 104130 567860
rect 113634 567848 113640 567860
rect 104124 567820 113640 567848
rect 104124 567808 104130 567820
rect 113634 567808 113640 567820
rect 113692 567848 113698 567860
rect 117976 567848 118004 568092
rect 123478 568080 123484 568092
rect 123536 568080 123542 568132
rect 124122 568080 124128 568132
rect 124180 568120 124186 568132
rect 146938 568120 146944 568132
rect 124180 568092 146944 568120
rect 124180 568080 124186 568092
rect 146938 568080 146944 568092
rect 146996 568080 147002 568132
rect 217870 568080 217876 568132
rect 217928 568120 217934 568132
rect 227162 568120 227168 568132
rect 217928 568092 227168 568120
rect 217928 568080 217934 568092
rect 227162 568080 227168 568092
rect 227220 568120 227226 568132
rect 235994 568120 236000 568132
rect 227220 568092 236000 568120
rect 227220 568080 227226 568092
rect 235994 568080 236000 568092
rect 236052 568080 236058 568132
rect 120074 568012 120080 568064
rect 120132 568052 120138 568064
rect 144178 568052 144184 568064
rect 120132 568024 144184 568052
rect 120132 568012 120138 568024
rect 144178 568012 144184 568024
rect 144236 568012 144242 568064
rect 202230 568012 202236 568064
rect 202288 568052 202294 568064
rect 211890 568052 211896 568064
rect 202288 568024 211896 568052
rect 202288 568012 202294 568024
rect 211890 568012 211896 568024
rect 211948 568052 211954 568064
rect 221458 568052 221464 568064
rect 211948 568024 221464 568052
rect 211948 568012 211954 568024
rect 221458 568012 221464 568024
rect 221516 568052 221522 568064
rect 230474 568052 230480 568064
rect 221516 568024 230480 568052
rect 221516 568012 221522 568024
rect 230474 568012 230480 568024
rect 230532 568012 230538 568064
rect 119246 567944 119252 567996
rect 119304 567984 119310 567996
rect 142890 567984 142896 567996
rect 119304 567956 142896 567984
rect 119304 567944 119310 567956
rect 142890 567944 142896 567956
rect 142948 567944 142954 567996
rect 203702 567944 203708 567996
rect 203760 567984 203766 567996
rect 213086 567984 213092 567996
rect 203760 567956 213092 567984
rect 203760 567944 203766 567956
rect 213086 567944 213092 567956
rect 213144 567984 213150 567996
rect 222378 567984 222384 567996
rect 213144 567956 222384 567984
rect 213144 567944 213150 567956
rect 222378 567944 222384 567956
rect 222436 567984 222442 567996
rect 231854 567984 231860 567996
rect 222436 567956 231860 567984
rect 222436 567944 222442 567956
rect 231854 567944 231860 567956
rect 231912 567944 231918 567996
rect 125502 567876 125508 567928
rect 125560 567916 125566 567928
rect 152458 567916 152464 567928
rect 125560 567888 152464 567916
rect 125560 567876 125566 567888
rect 152458 567876 152464 567888
rect 152516 567876 152522 567928
rect 204806 567876 204812 567928
rect 204864 567916 204870 567928
rect 214098 567916 214104 567928
rect 204864 567888 214104 567916
rect 204864 567876 204870 567888
rect 214098 567876 214104 567888
rect 214156 567916 214162 567928
rect 223666 567916 223672 567928
rect 214156 567888 223672 567916
rect 214156 567876 214162 567888
rect 223666 567876 223672 567888
rect 223724 567916 223730 567928
rect 231946 567916 231952 567928
rect 223724 567888 231952 567916
rect 223724 567876 223730 567888
rect 231946 567876 231952 567888
rect 232004 567876 232010 567928
rect 113692 567820 118004 567848
rect 113692 567808 113698 567820
rect 118050 567808 118056 567860
rect 118108 567848 118114 567860
rect 142798 567848 142804 567860
rect 118108 567820 142804 567848
rect 118108 567808 118114 567820
rect 142798 567808 142804 567820
rect 142856 567808 142862 567860
rect 208302 567808 208308 567860
rect 208360 567848 208366 567860
rect 217134 567848 217140 567860
rect 208360 567820 217140 567848
rect 208360 567808 208366 567820
rect 217134 567808 217140 567820
rect 217192 567808 217198 567860
rect 220078 567808 220084 567860
rect 220136 567848 220142 567860
rect 229370 567848 229376 567860
rect 220136 567820 229376 567848
rect 220136 567808 220142 567820
rect 229370 567808 229376 567820
rect 229428 567848 229434 567860
rect 238754 567848 238760 567860
rect 229428 567820 238760 567848
rect 229428 567808 229434 567820
rect 238754 567808 238760 567820
rect 238812 567808 238818 567860
rect 102962 567740 102968 567792
rect 103020 567780 103026 567792
rect 156690 567780 156696 567792
rect 103020 567752 156696 567780
rect 103020 567740 103026 567752
rect 156690 567740 156696 567752
rect 156748 567740 156754 567792
rect 85482 567672 85488 567724
rect 85540 567712 85546 567724
rect 91094 567712 91100 567724
rect 85540 567684 91100 567712
rect 85540 567672 85546 567684
rect 91094 567672 91100 567684
rect 91152 567672 91158 567724
rect 100662 567672 100668 567724
rect 100720 567712 100726 567724
rect 156782 567712 156788 567724
rect 100720 567684 156788 567712
rect 100720 567672 100726 567684
rect 156782 567672 156788 567684
rect 156840 567672 156846 567724
rect 97902 567604 97908 567656
rect 97960 567644 97966 567656
rect 155218 567644 155224 567656
rect 97960 567616 155224 567644
rect 97960 567604 97966 567616
rect 155218 567604 155224 567616
rect 155276 567604 155282 567656
rect 95142 567536 95148 567588
rect 95200 567576 95206 567588
rect 153838 567576 153844 567588
rect 95200 567548 153844 567576
rect 95200 567536 95206 567548
rect 153838 567536 153844 567548
rect 153896 567536 153902 567588
rect 194410 567536 194416 567588
rect 194468 567576 194474 567588
rect 252186 567576 252192 567588
rect 194468 567548 252192 567576
rect 194468 567536 194474 567548
rect 252186 567536 252192 567548
rect 252244 567536 252250 567588
rect 110322 567468 110328 567520
rect 110380 567508 110386 567520
rect 138658 567508 138664 567520
rect 110380 567480 138664 567508
rect 110380 567468 110386 567480
rect 138658 567468 138664 567480
rect 138716 567468 138722 567520
rect 116949 567443 117007 567449
rect 116949 567409 116961 567443
rect 116995 567440 117007 567443
rect 124858 567440 124864 567452
rect 116995 567412 124864 567440
rect 116995 567409 117007 567412
rect 116949 567403 117007 567409
rect 124858 567400 124864 567412
rect 124916 567400 124922 567452
rect 127618 567440 127624 567452
rect 124968 567412 127624 567440
rect 81342 567332 81348 567384
rect 81400 567372 81406 567384
rect 88334 567372 88340 567384
rect 81400 567344 88340 567372
rect 81400 567332 81406 567344
rect 88334 567332 88340 567344
rect 88392 567332 88398 567384
rect 115385 567375 115443 567381
rect 115385 567341 115397 567375
rect 115431 567372 115443 567375
rect 120626 567372 120632 567384
rect 115431 567344 120632 567372
rect 115431 567341 115443 567344
rect 115385 567335 115443 567341
rect 120626 567332 120632 567344
rect 120684 567332 120690 567384
rect 124968 567372 124996 567412
rect 127618 567400 127624 567412
rect 127676 567400 127682 567452
rect 128262 567400 128268 567452
rect 128320 567440 128326 567452
rect 207014 567440 207020 567452
rect 128320 567412 207020 567440
rect 128320 567400 128326 567412
rect 207014 567400 207020 567412
rect 207072 567440 207078 567452
rect 208302 567440 208308 567452
rect 207072 567412 208308 567440
rect 207072 567400 207078 567412
rect 208302 567400 208308 567412
rect 208360 567400 208366 567452
rect 120736 567344 124996 567372
rect 82722 567264 82728 567316
rect 82780 567304 82786 567316
rect 89990 567304 89996 567316
rect 82780 567276 89996 567304
rect 82780 567264 82786 567276
rect 89990 567264 89996 567276
rect 90048 567264 90054 567316
rect 116857 567307 116915 567313
rect 116857 567273 116869 567307
rect 116903 567304 116915 567307
rect 118326 567304 118332 567316
rect 116903 567276 118332 567304
rect 116903 567273 116915 567276
rect 116857 567267 116915 567273
rect 118326 567264 118332 567276
rect 118384 567304 118390 567316
rect 120736 567304 120764 567344
rect 125410 567332 125416 567384
rect 125468 567372 125474 567384
rect 204806 567372 204812 567384
rect 125468 567344 204812 567372
rect 125468 567332 125474 567344
rect 204806 567332 204812 567344
rect 204864 567332 204870 567384
rect 209038 567332 209044 567384
rect 209096 567372 209102 567384
rect 217870 567372 217876 567384
rect 209096 567344 217876 567372
rect 209096 567332 209102 567344
rect 217870 567332 217876 567344
rect 217928 567332 217934 567384
rect 118384 567276 120764 567304
rect 118384 567264 118390 567276
rect 121270 567264 121276 567316
rect 121328 567304 121334 567316
rect 202230 567304 202236 567316
rect 121328 567276 202236 567304
rect 121328 567264 121334 567276
rect 202230 567264 202236 567276
rect 202288 567264 202294 567316
rect 210418 567264 210424 567316
rect 210476 567304 210482 567316
rect 220078 567304 220084 567316
rect 210476 567276 220084 567304
rect 210476 567264 210482 567276
rect 220078 567264 220084 567276
rect 220136 567264 220142 567316
rect 78122 567196 78128 567248
rect 78180 567236 78186 567248
rect 86954 567236 86960 567248
rect 78180 567208 86960 567236
rect 78180 567196 78186 567208
rect 86954 567196 86960 567208
rect 87012 567196 87018 567248
rect 110690 567196 110696 567248
rect 110748 567236 110754 567248
rect 120718 567236 120724 567248
rect 110748 567208 120724 567236
rect 110748 567196 110754 567208
rect 120718 567196 120724 567208
rect 120776 567196 120782 567248
rect 122650 567196 122656 567248
rect 122708 567236 122714 567248
rect 203702 567236 203708 567248
rect 122708 567208 203708 567236
rect 122708 567196 122714 567208
rect 203702 567196 203708 567208
rect 203760 567196 203766 567248
rect 206278 567196 206284 567248
rect 206336 567236 206342 567248
rect 215570 567236 215576 567248
rect 206336 567208 215576 567236
rect 206336 567196 206342 567208
rect 215570 567196 215576 567208
rect 215628 567196 215634 567248
rect 252554 557540 252560 557592
rect 252612 557580 252618 557592
rect 252612 557552 253980 557580
rect 252612 557540 252618 557552
rect 253952 557512 253980 557552
rect 257982 557512 257988 557524
rect 253952 557484 257988 557512
rect 257982 557472 257988 557484
rect 258040 557472 258046 557524
rect 258074 551624 258080 551676
rect 258132 551664 258138 551676
rect 259730 551664 259736 551676
rect 258132 551636 259736 551664
rect 258132 551624 258138 551636
rect 259730 551624 259736 551636
rect 259788 551624 259794 551676
rect 259730 549176 259736 549228
rect 259788 549216 259794 549228
rect 261478 549216 261484 549228
rect 259788 549188 261484 549216
rect 259788 549176 259794 549188
rect 261478 549176 261484 549188
rect 261536 549176 261542 549228
rect 261478 540948 261484 541000
rect 261536 540988 261542 541000
rect 261536 540960 262260 540988
rect 261536 540948 261542 540960
rect 262232 540920 262260 540960
rect 263594 540920 263600 540932
rect 262232 540892 263600 540920
rect 263594 540880 263600 540892
rect 263652 540880 263658 540932
rect 263594 538840 263600 538892
rect 263652 538880 263658 538892
rect 272058 538880 272064 538892
rect 263652 538852 272064 538880
rect 263652 538840 263658 538852
rect 272058 538840 272064 538852
rect 272116 538840 272122 538892
rect 272058 534556 272064 534608
rect 272116 534596 272122 534608
rect 273898 534596 273904 534608
rect 272116 534568 273904 534596
rect 272116 534556 272122 534568
rect 273898 534556 273904 534568
rect 273956 534556 273962 534608
rect 111702 525716 111708 525768
rect 111760 525756 111766 525768
rect 181438 525756 181444 525768
rect 111760 525728 181444 525756
rect 111760 525716 111766 525728
rect 181438 525716 181444 525728
rect 181496 525716 181502 525768
rect 119982 525648 119988 525700
rect 120040 525688 120046 525700
rect 194778 525688 194784 525700
rect 120040 525660 194784 525688
rect 120040 525648 120046 525660
rect 194778 525648 194784 525660
rect 194836 525648 194842 525700
rect 128170 525580 128176 525632
rect 128228 525620 128234 525632
rect 208118 525620 208124 525632
rect 128228 525592 208124 525620
rect 128228 525580 128234 525592
rect 208118 525580 208124 525592
rect 208176 525580 208182 525632
rect 101398 525512 101404 525564
rect 101456 525552 101462 525564
rect 188338 525552 188344 525564
rect 101456 525524 188344 525552
rect 101456 525512 101462 525524
rect 188338 525512 188344 525524
rect 188396 525512 188402 525564
rect 99466 525444 99472 525496
rect 99524 525484 99530 525496
rect 188430 525484 188436 525496
rect 99524 525456 188436 525484
rect 99524 525444 99530 525456
rect 188430 525444 188436 525456
rect 188488 525444 188494 525496
rect 97626 525376 97632 525428
rect 97684 525416 97690 525428
rect 188522 525416 188528 525428
rect 97684 525388 188528 525416
rect 97684 525376 97690 525388
rect 188522 525376 188528 525388
rect 188580 525376 188586 525428
rect 95694 525308 95700 525360
rect 95752 525348 95758 525360
rect 188614 525348 188620 525360
rect 95752 525320 188620 525348
rect 95752 525308 95758 525320
rect 188614 525308 188620 525320
rect 188672 525308 188678 525360
rect 93762 525240 93768 525292
rect 93820 525280 93826 525292
rect 188706 525280 188712 525292
rect 93820 525252 188712 525280
rect 93820 525240 93826 525252
rect 188706 525240 188712 525252
rect 188764 525240 188770 525292
rect 91830 525172 91836 525224
rect 91888 525212 91894 525224
rect 188798 525212 188804 525224
rect 91888 525184 188804 525212
rect 91888 525172 91894 525184
rect 188798 525172 188804 525184
rect 188856 525172 188862 525224
rect 86126 525104 86132 525156
rect 86184 525144 86190 525156
rect 188890 525144 188896 525156
rect 86184 525116 188896 525144
rect 86184 525104 86190 525116
rect 188890 525104 188896 525116
rect 188948 525104 188954 525156
rect 89990 525036 89996 525088
rect 90048 525076 90054 525088
rect 195974 525076 195980 525088
rect 90048 525048 195980 525076
rect 90048 525036 90054 525048
rect 195974 525036 195980 525048
rect 196032 525036 196038 525088
rect 108942 524968 108948 525020
rect 109000 525008 109006 525020
rect 175734 525008 175740 525020
rect 109000 524980 175740 525008
rect 109000 524968 109006 524980
rect 175734 524968 175740 524980
rect 175792 524968 175798 525020
rect 107562 524900 107568 524952
rect 107620 524940 107626 524952
rect 173802 524940 173808 524952
rect 107620 524912 173808 524940
rect 107620 524900 107626 524912
rect 173802 524900 173808 524912
rect 173860 524900 173866 524952
rect 104802 524832 104808 524884
rect 104860 524872 104866 524884
rect 170030 524872 170036 524884
rect 104860 524844 170036 524872
rect 104860 524832 104866 524844
rect 170030 524832 170036 524844
rect 170088 524832 170094 524884
rect 106182 524764 106188 524816
rect 106240 524804 106246 524816
rect 171962 524804 171968 524816
rect 106240 524776 171968 524804
rect 106240 524764 106246 524776
rect 171962 524764 171968 524776
rect 172020 524764 172026 524816
rect 93670 524696 93676 524748
rect 93728 524736 93734 524748
rect 150986 524736 150992 524748
rect 93728 524708 150992 524736
rect 93728 524696 93734 524708
rect 150986 524696 150992 524708
rect 151044 524696 151050 524748
rect 74718 524356 74724 524408
rect 74776 524396 74782 524408
rect 75822 524396 75828 524408
rect 74776 524368 75828 524396
rect 74776 524356 74782 524368
rect 75822 524356 75828 524368
rect 75880 524356 75886 524408
rect 80422 524356 80428 524408
rect 80480 524396 80486 524408
rect 81342 524396 81348 524408
rect 80480 524368 81348 524396
rect 80480 524356 80486 524368
rect 81342 524356 81348 524368
rect 81400 524356 81406 524408
rect 84286 524356 84292 524408
rect 84344 524396 84350 524408
rect 85482 524396 85488 524408
rect 84344 524368 85488 524396
rect 84344 524356 84350 524368
rect 85482 524356 85488 524368
rect 85540 524356 85546 524408
rect 95050 524356 95056 524408
rect 95108 524396 95114 524408
rect 152826 524396 152832 524408
rect 95108 524368 152832 524396
rect 95108 524356 95114 524368
rect 152826 524356 152832 524368
rect 152884 524356 152890 524408
rect 153838 524356 153844 524408
rect 153896 524396 153902 524408
rect 154758 524396 154764 524408
rect 153896 524368 154764 524396
rect 153896 524356 153902 524368
rect 154758 524356 154764 524368
rect 154816 524356 154822 524408
rect 155218 524356 155224 524408
rect 155276 524396 155282 524408
rect 158530 524396 158536 524408
rect 155276 524368 158536 524396
rect 155276 524356 155282 524368
rect 158530 524356 158536 524368
rect 158588 524356 158594 524408
rect 162394 524396 162400 524408
rect 159284 524368 162400 524396
rect 99190 524288 99196 524340
rect 99248 524328 99254 524340
rect 103425 524331 103483 524337
rect 99248 524300 103284 524328
rect 99248 524288 99254 524300
rect 96430 524220 96436 524272
rect 96488 524260 96494 524272
rect 103149 524263 103207 524269
rect 103149 524260 103161 524263
rect 96488 524232 103161 524260
rect 96488 524220 96494 524232
rect 103149 524229 103161 524232
rect 103195 524229 103207 524263
rect 103256 524260 103284 524300
rect 103425 524297 103437 524331
rect 103471 524328 103483 524331
rect 113177 524331 113235 524337
rect 113177 524328 113189 524331
rect 103471 524300 113189 524328
rect 103471 524297 103483 524300
rect 103425 524291 103483 524297
rect 113177 524297 113189 524300
rect 113223 524297 113235 524331
rect 113177 524291 113235 524297
rect 122745 524331 122803 524337
rect 122745 524297 122757 524331
rect 122791 524328 122803 524331
rect 132497 524331 132555 524337
rect 132497 524328 132509 524331
rect 122791 524300 132509 524328
rect 122791 524297 122803 524300
rect 122745 524291 122803 524297
rect 132497 524297 132509 524300
rect 132543 524297 132555 524331
rect 132497 524291 132555 524297
rect 142065 524331 142123 524337
rect 142065 524297 142077 524331
rect 142111 524328 142123 524331
rect 156414 524328 156420 524340
rect 142111 524300 156420 524328
rect 142111 524297 142123 524300
rect 142065 524291 142123 524297
rect 156414 524288 156420 524300
rect 156472 524288 156478 524340
rect 156690 524288 156696 524340
rect 156748 524328 156754 524340
rect 159177 524331 159235 524337
rect 159177 524328 159189 524331
rect 156748 524300 159189 524328
rect 156748 524288 156754 524300
rect 159177 524297 159189 524300
rect 159223 524297 159235 524331
rect 159177 524291 159235 524297
rect 108301 524263 108359 524269
rect 108301 524260 108313 524263
rect 103256 524232 108313 524260
rect 103149 524223 103207 524229
rect 108301 524229 108313 524232
rect 108347 524229 108359 524263
rect 108301 524223 108359 524229
rect 122653 524263 122711 524269
rect 122653 524229 122665 524263
rect 122699 524260 122711 524263
rect 132589 524263 132647 524269
rect 132589 524260 132601 524263
rect 122699 524232 132601 524260
rect 122699 524229 122711 524232
rect 122653 524223 122711 524229
rect 132589 524229 132601 524232
rect 132635 524229 132647 524263
rect 132589 524223 132647 524229
rect 141973 524263 142031 524269
rect 141973 524229 141985 524263
rect 142019 524260 142031 524263
rect 156141 524263 156199 524269
rect 156141 524260 156153 524263
rect 142019 524232 156153 524260
rect 142019 524229 142031 524232
rect 141973 524223 142031 524229
rect 156141 524229 156153 524232
rect 156187 524229 156199 524263
rect 156141 524223 156199 524229
rect 156782 524220 156788 524272
rect 156840 524260 156846 524272
rect 159284 524260 159312 524368
rect 162394 524356 162400 524368
rect 162452 524356 162458 524408
rect 208302 524356 208308 524408
rect 208360 524396 208366 524408
rect 219526 524396 219532 524408
rect 208360 524368 219532 524396
rect 208360 524356 208366 524368
rect 219526 524356 219532 524368
rect 219584 524356 219590 524408
rect 229002 524356 229008 524408
rect 229060 524396 229066 524408
rect 253842 524396 253848 524408
rect 229060 524368 253848 524396
rect 229060 524356 229066 524368
rect 253842 524356 253848 524368
rect 253900 524356 253906 524408
rect 159361 524331 159419 524337
rect 159361 524297 159373 524331
rect 159407 524328 159419 524331
rect 166166 524328 166172 524340
rect 159407 524300 166172 524328
rect 159407 524297 159419 524300
rect 159361 524291 159419 524297
rect 166166 524288 166172 524300
rect 166224 524288 166230 524340
rect 211062 524288 211068 524340
rect 211120 524328 211126 524340
rect 223390 524328 223396 524340
rect 211120 524300 223396 524328
rect 211120 524288 211126 524300
rect 223390 524288 223396 524300
rect 223448 524288 223454 524340
rect 227622 524288 227628 524340
rect 227680 524328 227686 524340
rect 252002 524328 252008 524340
rect 227680 524300 252008 524328
rect 227680 524288 227686 524300
rect 252002 524288 252008 524300
rect 252060 524288 252066 524340
rect 156840 524232 159312 524260
rect 156840 524220 156846 524232
rect 209682 524220 209688 524272
rect 209740 524260 209746 524272
rect 221458 524260 221464 524272
rect 209740 524232 221464 524260
rect 209740 524220 209746 524232
rect 221458 524220 221464 524232
rect 221516 524220 221522 524272
rect 231762 524220 231768 524272
rect 231820 524260 231826 524272
rect 257706 524260 257712 524272
rect 231820 524232 257712 524260
rect 231820 524220 231826 524232
rect 257706 524220 257712 524232
rect 257764 524220 257770 524272
rect 101950 524152 101956 524204
rect 102008 524192 102014 524204
rect 164326 524192 164332 524204
rect 102008 524164 164332 524192
rect 102008 524152 102014 524164
rect 164326 524152 164332 524164
rect 164384 524152 164390 524204
rect 212442 524152 212448 524204
rect 212500 524192 212506 524204
rect 227162 524192 227168 524204
rect 212500 524164 227168 524192
rect 212500 524152 212506 524164
rect 227162 524152 227168 524164
rect 227220 524152 227226 524204
rect 230382 524152 230388 524204
rect 230440 524192 230446 524204
rect 255774 524192 255780 524204
rect 230440 524164 255780 524192
rect 230440 524152 230446 524164
rect 255774 524152 255780 524164
rect 255832 524152 255838 524204
rect 78858 524084 78864 524136
rect 78916 524124 78922 524136
rect 88058 524124 88064 524136
rect 78916 524096 88064 524124
rect 78916 524084 78922 524096
rect 88058 524084 88064 524096
rect 88116 524084 88122 524136
rect 103330 524084 103336 524136
rect 103388 524124 103394 524136
rect 168098 524124 168104 524136
rect 103388 524096 168104 524124
rect 103388 524084 103394 524096
rect 168098 524084 168104 524096
rect 168156 524084 168162 524136
rect 214009 524127 214067 524133
rect 214009 524093 214021 524127
rect 214055 524124 214067 524127
rect 225322 524124 225328 524136
rect 214055 524096 225328 524124
rect 214055 524093 214067 524096
rect 214009 524087 214067 524093
rect 225322 524084 225328 524096
rect 225380 524084 225386 524136
rect 233142 524084 233148 524136
rect 233200 524124 233206 524136
rect 259546 524124 259552 524136
rect 233200 524096 259552 524124
rect 233200 524084 233206 524096
rect 259546 524084 259552 524096
rect 259604 524084 259610 524136
rect 78766 524016 78772 524068
rect 78824 524056 78830 524068
rect 108301 524059 108359 524065
rect 78824 524028 106320 524056
rect 78824 524016 78830 524028
rect 78674 523948 78680 524000
rect 78732 523988 78738 524000
rect 106292 523988 106320 524028
rect 108301 524025 108313 524059
rect 108347 524056 108359 524059
rect 117961 524059 118019 524065
rect 117961 524056 117973 524059
rect 108347 524028 117973 524056
rect 108347 524025 108359 524028
rect 108301 524019 108359 524025
rect 117961 524025 117973 524028
rect 118007 524025 118019 524059
rect 117961 524019 118019 524025
rect 120442 524016 120448 524068
rect 120500 524056 120506 524068
rect 121270 524056 121276 524068
rect 120500 524028 121276 524056
rect 120500 524016 120506 524028
rect 121270 524016 121276 524028
rect 121328 524016 121334 524068
rect 121365 524059 121423 524065
rect 121365 524025 121377 524059
rect 121411 524056 121423 524059
rect 185302 524056 185308 524068
rect 121411 524028 185308 524056
rect 121411 524025 121423 524028
rect 121365 524019 121423 524025
rect 185302 524016 185308 524028
rect 185360 524016 185366 524068
rect 204162 524016 204168 524068
rect 204220 524056 204226 524068
rect 213822 524056 213828 524068
rect 204220 524028 213828 524056
rect 204220 524016 204226 524028
rect 213822 524016 213828 524028
rect 213880 524016 213886 524068
rect 213914 524016 213920 524068
rect 213972 524056 213978 524068
rect 229094 524056 229100 524068
rect 213972 524028 229100 524056
rect 213972 524016 213978 524028
rect 229094 524016 229100 524028
rect 229152 524016 229158 524068
rect 234522 524016 234528 524068
rect 234580 524056 234586 524068
rect 263410 524056 263416 524068
rect 234580 524028 263416 524056
rect 234580 524016 234586 524028
rect 263410 524016 263416 524028
rect 263468 524016 263474 524068
rect 109034 523988 109040 524000
rect 78732 523960 105860 523988
rect 106292 523960 109040 523988
rect 78732 523948 78738 523960
rect 78306 523880 78312 523932
rect 78364 523920 78370 523932
rect 105725 523923 105783 523929
rect 105725 523920 105737 523923
rect 78364 523892 105737 523920
rect 78364 523880 78370 523892
rect 105725 523889 105737 523892
rect 105771 523889 105783 523923
rect 105832 523920 105860 523960
rect 109034 523948 109040 523960
rect 109092 523948 109098 524000
rect 118510 523948 118516 524000
rect 118568 523988 118574 524000
rect 191006 523988 191012 524000
rect 118568 523960 191012 523988
rect 118568 523948 118574 523960
rect 191006 523948 191012 523960
rect 191064 523948 191070 524000
rect 205542 523948 205548 524000
rect 205600 523988 205606 524000
rect 215754 523988 215760 524000
rect 205600 523960 215760 523988
rect 205600 523948 205606 523960
rect 215754 523948 215760 523960
rect 215812 523948 215818 524000
rect 216582 523948 216588 524000
rect 216640 523988 216646 524000
rect 232866 523988 232872 524000
rect 216640 523960 232872 523988
rect 216640 523948 216646 523960
rect 232866 523948 232872 523960
rect 232924 523948 232930 524000
rect 235902 523948 235908 524000
rect 235960 523988 235966 524000
rect 243541 523991 243599 523997
rect 243541 523988 243553 523991
rect 235960 523960 243553 523988
rect 235960 523948 235966 523960
rect 243541 523957 243553 523960
rect 243587 523957 243599 523991
rect 243541 523951 243599 523957
rect 243633 523991 243691 523997
rect 243633 523957 243645 523991
rect 243679 523988 243691 523991
rect 261478 523988 261484 524000
rect 243679 523960 261484 523988
rect 243679 523957 243691 523960
rect 243633 523951 243691 523957
rect 261478 523948 261484 523960
rect 261536 523948 261542 524000
rect 110966 523920 110972 523932
rect 105832 523892 110972 523920
rect 105725 523883 105783 523889
rect 110966 523880 110972 523892
rect 111024 523880 111030 523932
rect 114462 523880 114468 523932
rect 114520 523920 114526 523932
rect 121365 523923 121423 523929
rect 121365 523920 121377 523923
rect 114520 523892 121377 523920
rect 114520 523880 114526 523892
rect 121365 523889 121377 523892
rect 121411 523889 121423 523923
rect 121365 523883 121423 523889
rect 122742 523880 122748 523932
rect 122800 523920 122806 523932
rect 198642 523920 198648 523932
rect 122800 523892 198648 523920
rect 122800 523880 122806 523892
rect 198642 523880 198648 523892
rect 198700 523880 198706 523932
rect 202782 523880 202788 523932
rect 202840 523920 202846 523932
rect 211982 523920 211988 523932
rect 202840 523892 211988 523920
rect 202840 523880 202846 523892
rect 211982 523880 211988 523892
rect 212040 523880 212046 523932
rect 215202 523880 215208 523932
rect 215260 523920 215266 523932
rect 231026 523920 231032 523932
rect 215260 523892 231032 523920
rect 215260 523880 215266 523892
rect 231026 523880 231032 523892
rect 231084 523880 231090 523932
rect 233050 523880 233056 523932
rect 233108 523920 233114 523932
rect 233108 523892 235028 523920
rect 233108 523880 233114 523892
rect 78398 523812 78404 523864
rect 78456 523852 78462 523864
rect 114738 523852 114744 523864
rect 78456 523824 114744 523852
rect 78456 523812 78462 523824
rect 114738 523812 114744 523824
rect 114796 523812 114802 523864
rect 117961 523855 118019 523861
rect 117961 523821 117973 523855
rect 118007 523852 118019 523855
rect 122653 523855 122711 523861
rect 122653 523852 122665 523855
rect 118007 523824 122665 523852
rect 118007 523821 118019 523824
rect 117961 523815 118019 523821
rect 122653 523821 122665 523824
rect 122699 523821 122711 523855
rect 122653 523815 122711 523821
rect 124306 523812 124312 523864
rect 124364 523852 124370 523864
rect 125410 523852 125416 523864
rect 124364 523824 125416 523852
rect 124364 523812 124370 523824
rect 125410 523812 125416 523824
rect 125468 523812 125474 523864
rect 133782 523812 133788 523864
rect 133840 523852 133846 523864
rect 210418 523852 210424 523864
rect 133840 523824 210424 523852
rect 133840 523812 133846 523824
rect 210418 523812 210424 523824
rect 210476 523812 210482 523864
rect 210970 523812 210976 523864
rect 211028 523852 211034 523864
rect 214009 523855 214067 523861
rect 214009 523852 214021 523855
rect 211028 523824 214021 523852
rect 211028 523812 211034 523824
rect 214009 523821 214021 523824
rect 214055 523821 214067 523855
rect 214009 523815 214067 523821
rect 217962 523812 217968 523864
rect 218020 523852 218026 523864
rect 234798 523852 234804 523864
rect 218020 523824 234804 523852
rect 218020 523812 218026 523824
rect 234798 523812 234804 523824
rect 234856 523812 234862 523864
rect 235000 523852 235028 523892
rect 237282 523880 237288 523932
rect 237340 523920 237346 523932
rect 267182 523920 267188 523932
rect 237340 523892 267188 523920
rect 237340 523880 237346 523892
rect 267182 523880 267188 523892
rect 267240 523880 267246 523932
rect 235000 523824 238432 523852
rect 78490 523744 78496 523796
rect 78548 523784 78554 523796
rect 116670 523784 116676 523796
rect 78548 523756 116676 523784
rect 78548 523744 78554 523756
rect 116670 523744 116676 523756
rect 116728 523744 116734 523796
rect 130010 523744 130016 523796
rect 130068 523784 130074 523796
rect 209038 523784 209044 523796
rect 130068 523756 209044 523784
rect 130068 523744 130074 523756
rect 209038 523744 209044 523756
rect 209096 523744 209102 523796
rect 219342 523744 219348 523796
rect 219400 523784 219406 523796
rect 238294 523784 238300 523796
rect 219400 523756 238300 523784
rect 219400 523744 219406 523756
rect 238294 523744 238300 523756
rect 238352 523744 238358 523796
rect 78582 523676 78588 523728
rect 78640 523716 78646 523728
rect 118510 523716 118516 523728
rect 78640 523688 118516 523716
rect 78640 523676 78646 523688
rect 118510 523676 118516 523688
rect 118568 523676 118574 523728
rect 126146 523676 126152 523728
rect 126204 523716 126210 523728
rect 206278 523716 206284 523728
rect 126204 523688 206284 523716
rect 126204 523676 126210 523688
rect 206278 523676 206284 523688
rect 206336 523676 206342 523728
rect 206922 523676 206928 523728
rect 206980 523716 206986 523728
rect 217686 523716 217692 523728
rect 206980 523688 217692 523716
rect 206980 523676 206986 523688
rect 217686 523676 217692 523688
rect 217744 523676 217750 523728
rect 217870 523676 217876 523728
rect 217928 523716 217934 523728
rect 236730 523716 236736 523728
rect 217928 523688 236736 523716
rect 217928 523676 217934 523688
rect 236730 523676 236736 523688
rect 236788 523676 236794 523728
rect 238404 523716 238432 523824
rect 238662 523812 238668 523864
rect 238720 523852 238726 523864
rect 238720 523824 239996 523852
rect 238720 523812 238726 523824
rect 239968 523784 239996 523824
rect 240042 523812 240048 523864
rect 240100 523852 240106 523864
rect 243449 523855 243507 523861
rect 243449 523852 243461 523855
rect 240100 523824 243461 523852
rect 240100 523812 240106 523824
rect 243449 523821 243461 523824
rect 243495 523821 243507 523855
rect 243449 523815 243507 523821
rect 243541 523855 243599 523861
rect 243541 523821 243553 523855
rect 243587 523852 243599 523855
rect 265342 523852 265348 523864
rect 243587 523824 265348 523852
rect 243587 523821 243599 523824
rect 243541 523815 243599 523821
rect 265342 523812 265348 523824
rect 265400 523812 265406 523864
rect 269114 523784 269120 523796
rect 239968 523756 269120 523784
rect 269114 523744 269120 523756
rect 269172 523744 269178 523796
rect 273898 523744 273904 523796
rect 273956 523784 273962 523796
rect 275370 523784 275376 523796
rect 273956 523756 275376 523784
rect 273956 523744 273962 523756
rect 275370 523744 275376 523756
rect 275428 523744 275434 523796
rect 243633 523719 243691 523725
rect 243633 523716 243645 523719
rect 238404 523688 243645 523716
rect 243633 523685 243645 523688
rect 243679 523685 243691 523719
rect 243633 523679 243691 523685
rect 243725 523719 243783 523725
rect 243725 523685 243737 523719
rect 243771 523716 243783 523719
rect 271046 523716 271052 523728
rect 243771 523688 271052 523716
rect 243771 523685 243783 523688
rect 243725 523679 243783 523685
rect 271046 523676 271052 523688
rect 271104 523676 271110 523728
rect 78214 523608 78220 523660
rect 78272 523648 78278 523660
rect 107102 523648 107108 523660
rect 78272 523620 107108 523648
rect 78272 523608 78278 523620
rect 107102 523608 107108 523620
rect 107160 523608 107166 523660
rect 113177 523651 113235 523657
rect 113177 523617 113189 523651
rect 113223 523648 113235 523651
rect 122745 523651 122803 523657
rect 122745 523648 122757 523651
rect 113223 523620 122757 523648
rect 113223 523617 113235 523620
rect 113177 523611 113235 523617
rect 122745 523617 122757 523620
rect 122791 523617 122803 523651
rect 122745 523611 122803 523617
rect 123478 523608 123484 523660
rect 123536 523648 123542 523660
rect 139486 523648 139492 523660
rect 123536 523620 139492 523648
rect 123536 523608 123542 523620
rect 139486 523608 139492 523620
rect 139544 523608 139550 523660
rect 140038 523608 140044 523660
rect 140096 523648 140102 523660
rect 196710 523648 196716 523660
rect 140096 523620 196716 523648
rect 140096 523608 140102 523620
rect 196710 523608 196716 523620
rect 196768 523608 196774 523660
rect 226242 523608 226248 523660
rect 226300 523648 226306 523660
rect 250070 523648 250076 523660
rect 226300 523620 250076 523648
rect 226300 523608 226306 523620
rect 250070 523608 250076 523620
rect 250128 523608 250134 523660
rect 103330 523540 103336 523592
rect 103388 523580 103394 523592
rect 155954 523580 155960 523592
rect 103388 523552 155960 523580
rect 103388 523540 103394 523552
rect 155954 523540 155960 523552
rect 156012 523540 156018 523592
rect 156141 523583 156199 523589
rect 156141 523549 156153 523583
rect 156187 523580 156199 523583
rect 160462 523580 160468 523592
rect 156187 523552 160468 523580
rect 156187 523549 156199 523552
rect 156141 523543 156199 523549
rect 160462 523540 160468 523552
rect 160520 523540 160526 523592
rect 226150 523540 226156 523592
rect 226208 523580 226214 523592
rect 248138 523580 248144 523592
rect 226208 523552 248144 523580
rect 226208 523540 226214 523552
rect 248138 523540 248144 523552
rect 248196 523540 248202 523592
rect 86770 523472 86776 523524
rect 86828 523512 86834 523524
rect 105170 523512 105176 523524
rect 86828 523484 105176 523512
rect 86828 523472 86834 523484
rect 105170 523472 105176 523484
rect 105228 523472 105234 523524
rect 105725 523515 105783 523521
rect 105725 523481 105737 523515
rect 105771 523512 105783 523515
rect 112806 523512 112812 523524
rect 105771 523484 112812 523512
rect 105771 523481 105783 523484
rect 105725 523475 105783 523481
rect 112806 523472 112812 523484
rect 112864 523472 112870 523524
rect 127618 523472 127624 523524
rect 127676 523512 127682 523524
rect 147122 523512 147128 523524
rect 127676 523484 147128 523512
rect 127676 523472 127682 523484
rect 147122 523472 147128 523484
rect 147180 523472 147186 523524
rect 200482 523512 200488 523524
rect 147324 523484 200488 523512
rect 124858 523404 124864 523456
rect 124916 523444 124922 523456
rect 143350 523444 143356 523456
rect 124916 523416 143356 523444
rect 124916 523404 124922 523416
rect 143350 523404 143356 523416
rect 143408 523404 143414 523456
rect 146938 523404 146944 523456
rect 146996 523444 147002 523456
rect 147324 523444 147352 523484
rect 200482 523472 200488 523484
rect 200540 523472 200546 523524
rect 223482 523472 223488 523524
rect 223540 523512 223546 523524
rect 244366 523512 244372 523524
rect 223540 523484 244372 523512
rect 223540 523472 223546 523484
rect 244366 523472 244372 523484
rect 244424 523472 244430 523524
rect 192846 523444 192852 523456
rect 146996 523416 147352 523444
rect 147416 523416 192852 523444
rect 146996 523404 147002 523416
rect 125042 523336 125048 523388
rect 125100 523376 125106 523388
rect 141418 523376 141424 523388
rect 125100 523348 141424 523376
rect 125100 523336 125106 523348
rect 141418 523336 141424 523348
rect 141476 523336 141482 523388
rect 144178 523336 144184 523388
rect 144236 523376 144242 523388
rect 147416 523376 147444 523416
rect 192846 523404 192852 523416
rect 192904 523404 192910 523456
rect 224862 523404 224868 523456
rect 224920 523444 224926 523456
rect 246206 523444 246212 523456
rect 224920 523416 246212 523444
rect 224920 523404 224926 523416
rect 246206 523404 246212 523416
rect 246264 523404 246270 523456
rect 144236 523348 147444 523376
rect 147493 523379 147551 523385
rect 144236 523336 144242 523348
rect 147493 523345 147505 523379
rect 147539 523376 147551 523379
rect 189074 523376 189080 523388
rect 147539 523348 189080 523376
rect 147539 523345 147551 523348
rect 147493 523339 147551 523345
rect 189074 523336 189080 523348
rect 189132 523336 189138 523388
rect 222102 523336 222108 523388
rect 222160 523376 222166 523388
rect 242434 523376 242440 523388
rect 222160 523348 242440 523376
rect 222160 523336 222166 523348
rect 242434 523336 242440 523348
rect 242492 523336 242498 523388
rect 120718 523268 120724 523320
rect 120776 523308 120782 523320
rect 135714 523308 135720 523320
rect 120776 523280 135720 523308
rect 120776 523268 120782 523280
rect 135714 523268 135720 523280
rect 135772 523268 135778 523320
rect 137278 523268 137284 523320
rect 137336 523308 137342 523320
rect 183370 523308 183376 523320
rect 137336 523280 183376 523308
rect 137336 523268 137342 523280
rect 183370 523268 183376 523280
rect 183428 523268 183434 523320
rect 220722 523268 220728 523320
rect 220780 523308 220786 523320
rect 240502 523308 240508 523320
rect 220780 523280 240508 523308
rect 220780 523268 220786 523280
rect 240502 523268 240508 523280
rect 240560 523268 240566 523320
rect 122098 523200 122104 523252
rect 122156 523240 122162 523252
rect 137646 523240 137652 523252
rect 122156 523212 137652 523240
rect 122156 523200 122162 523212
rect 137646 523200 137652 523212
rect 137704 523200 137710 523252
rect 137741 523243 137799 523249
rect 137741 523209 137753 523243
rect 137787 523240 137799 523243
rect 141973 523243 142031 523249
rect 141973 523240 141985 523243
rect 137787 523212 141985 523240
rect 137787 523209 137799 523212
rect 137741 523203 137799 523209
rect 141973 523209 141985 523212
rect 142019 523209 142031 523243
rect 141973 523203 142031 523209
rect 142890 523200 142896 523252
rect 142948 523240 142954 523252
rect 147493 523243 147551 523249
rect 147493 523240 147505 523243
rect 142948 523212 147505 523240
rect 142948 523200 142954 523212
rect 147493 523209 147505 523212
rect 147539 523209 147551 523243
rect 147493 523203 147551 523209
rect 147585 523243 147643 523249
rect 147585 523209 147597 523243
rect 147631 523240 147643 523243
rect 187142 523240 187148 523252
rect 147631 523212 187148 523240
rect 147631 523209 147643 523212
rect 147585 523203 147643 523209
rect 187142 523200 187148 523212
rect 187200 523200 187206 523252
rect 135898 523132 135904 523184
rect 135956 523172 135962 523184
rect 177666 523172 177672 523184
rect 135956 523144 177672 523172
rect 135956 523132 135962 523144
rect 177666 523132 177672 523144
rect 177724 523132 177730 523184
rect 132589 523107 132647 523113
rect 132589 523073 132601 523107
rect 132635 523104 132647 523107
rect 137741 523107 137799 523113
rect 137741 523104 137753 523107
rect 132635 523076 137753 523104
rect 132635 523073 132647 523076
rect 132589 523067 132647 523073
rect 137741 523073 137753 523076
rect 137787 523073 137799 523107
rect 137741 523067 137799 523073
rect 138658 523064 138664 523116
rect 138716 523104 138722 523116
rect 179506 523104 179512 523116
rect 138716 523076 179512 523104
rect 138716 523064 138722 523076
rect 179506 523064 179512 523076
rect 179564 523064 179570 523116
rect 132497 523039 132555 523045
rect 132497 523005 132509 523039
rect 132543 523036 132555 523039
rect 142065 523039 142123 523045
rect 142065 523036 142077 523039
rect 132543 523008 142077 523036
rect 132543 523005 132555 523008
rect 132497 522999 132555 523005
rect 142065 523005 142077 523008
rect 142111 523005 142123 523039
rect 142065 522999 142123 523005
rect 142798 522996 142804 523048
rect 142856 523036 142862 523048
rect 147585 523039 147643 523045
rect 147585 523036 147597 523039
rect 142856 523008 147597 523036
rect 142856 522996 142862 523008
rect 147585 523005 147597 523008
rect 147631 523005 147643 523039
rect 147585 522999 147643 523005
rect 275370 518984 275376 519036
rect 275428 519024 275434 519036
rect 278774 519024 278780 519036
rect 275428 518996 278780 519024
rect 275428 518984 275434 518996
rect 278774 518984 278780 518996
rect 278832 518984 278838 519036
rect 274266 518916 274272 518968
rect 274324 518956 274330 518968
rect 301498 518956 301504 518968
rect 274324 518928 301504 518956
rect 274324 518916 274330 518928
rect 301498 518916 301504 518928
rect 301556 518916 301562 518968
rect 278774 517012 278780 517064
rect 278832 517052 278838 517064
rect 280062 517052 280068 517064
rect 278832 517024 280068 517052
rect 278832 517012 278838 517024
rect 280062 517012 280068 517024
rect 280120 517012 280126 517064
rect 280062 516808 280068 516860
rect 280120 516848 280126 516860
rect 320174 516848 320180 516860
rect 280120 516820 320180 516848
rect 280120 516808 280126 516820
rect 320174 516808 320180 516820
rect 320232 516808 320238 516860
rect 273898 516740 273904 516792
rect 273956 516780 273962 516792
rect 337746 516780 337752 516792
rect 273956 516752 337752 516780
rect 273956 516740 273962 516752
rect 337746 516740 337752 516752
rect 337804 516740 337810 516792
rect 338390 516740 338396 516792
rect 338448 516780 338454 516792
rect 340874 516780 340880 516792
rect 338448 516752 340880 516780
rect 338448 516740 338454 516752
rect 340874 516740 340880 516752
rect 340932 516740 340938 516792
rect 275370 516672 275376 516724
rect 275428 516712 275434 516724
rect 398834 516712 398840 516724
rect 275428 516684 398840 516712
rect 275428 516672 275434 516684
rect 398834 516672 398840 516684
rect 398892 516672 398898 516724
rect 275462 516604 275468 516656
rect 275520 516644 275526 516656
rect 400214 516644 400220 516656
rect 275520 516616 400220 516644
rect 275520 516604 275526 516616
rect 400214 516604 400220 516616
rect 400272 516604 400278 516656
rect 274358 516536 274364 516588
rect 274416 516576 274422 516588
rect 401594 516576 401600 516588
rect 274416 516548 401600 516576
rect 274416 516536 274422 516548
rect 401594 516536 401600 516548
rect 401652 516536 401658 516588
rect 274450 516468 274456 516520
rect 274508 516508 274514 516520
rect 403342 516508 403348 516520
rect 274508 516480 403348 516508
rect 274508 516468 274514 516480
rect 403342 516468 403348 516480
rect 403400 516468 403406 516520
rect 274542 516400 274548 516452
rect 274600 516440 274606 516452
rect 404354 516440 404360 516452
rect 274600 516412 404360 516440
rect 274600 516400 274606 516412
rect 404354 516400 404360 516412
rect 404412 516400 404418 516452
rect 406010 516400 406016 516452
rect 406068 516400 406074 516452
rect 273806 516332 273812 516384
rect 273864 516372 273870 516384
rect 406028 516372 406056 516400
rect 273864 516344 406056 516372
rect 273864 516332 273870 516344
rect 273622 514768 273628 514820
rect 273680 514808 273686 514820
rect 298738 514808 298744 514820
rect 273680 514780 298744 514808
rect 273680 514768 273686 514780
rect 298738 514768 298744 514780
rect 298796 514768 298802 514820
rect 275278 511980 275284 512032
rect 275336 512020 275342 512032
rect 320174 512020 320180 512032
rect 275336 511992 320180 512020
rect 275336 511980 275342 511992
rect 320174 511980 320180 511992
rect 320232 511980 320238 512032
rect 273530 510620 273536 510672
rect 273588 510660 273594 510672
rect 297358 510660 297364 510672
rect 273588 510632 297364 510660
rect 273588 510620 273594 510632
rect 297358 510620 297364 510632
rect 297416 510620 297422 510672
rect 279418 509260 279424 509312
rect 279476 509300 279482 509312
rect 320358 509300 320364 509312
rect 279476 509272 320364 509300
rect 279476 509260 279482 509272
rect 320358 509260 320364 509272
rect 320416 509260 320422 509312
rect 302878 507832 302884 507884
rect 302936 507872 302942 507884
rect 320174 507872 320180 507884
rect 302936 507844 320180 507872
rect 302936 507832 302942 507844
rect 320174 507832 320180 507844
rect 320232 507832 320238 507884
rect 273714 506540 273720 506592
rect 273772 506580 273778 506592
rect 294598 506580 294604 506592
rect 273772 506552 294604 506580
rect 273772 506540 273778 506552
rect 294598 506540 294604 506552
rect 294656 506540 294662 506592
rect 275554 506472 275560 506524
rect 275612 506512 275618 506524
rect 319806 506512 319812 506524
rect 275612 506484 319812 506512
rect 275612 506472 275618 506484
rect 319806 506472 319812 506484
rect 319864 506472 319870 506524
rect 273530 505180 273536 505232
rect 273588 505220 273594 505232
rect 291838 505220 291844 505232
rect 273588 505192 291844 505220
rect 273588 505180 273594 505192
rect 291838 505180 291844 505192
rect 291896 505180 291902 505232
rect 275646 505112 275652 505164
rect 275704 505152 275710 505164
rect 320174 505152 320180 505164
rect 275704 505124 320180 505152
rect 275704 505112 275710 505124
rect 320174 505112 320180 505124
rect 320232 505112 320238 505164
rect 276658 503684 276664 503736
rect 276716 503724 276722 503736
rect 319990 503724 319996 503736
rect 276716 503696 319996 503724
rect 276716 503684 276722 503696
rect 319990 503684 319996 503696
rect 320048 503684 320054 503736
rect 299477 502843 299535 502849
rect 299477 502809 299489 502843
rect 299523 502840 299535 502843
rect 309045 502843 309103 502849
rect 309045 502840 309057 502843
rect 299523 502812 309057 502840
rect 299523 502809 299535 502812
rect 299477 502803 299535 502809
rect 309045 502809 309057 502812
rect 309091 502809 309103 502843
rect 309045 502803 309103 502809
rect 289817 502707 289875 502713
rect 289817 502673 289829 502707
rect 289863 502704 289875 502707
rect 299477 502707 299535 502713
rect 299477 502704 299489 502707
rect 289863 502676 299489 502704
rect 289863 502673 289875 502676
rect 289817 502667 289875 502673
rect 299477 502673 299489 502676
rect 299523 502673 299535 502707
rect 299477 502667 299535 502673
rect 280157 502639 280215 502645
rect 280157 502605 280169 502639
rect 280203 502636 280215 502639
rect 289633 502639 289691 502645
rect 289633 502636 289645 502639
rect 280203 502608 289645 502636
rect 280203 502605 280215 502608
rect 280157 502599 280215 502605
rect 289633 502605 289645 502608
rect 289679 502605 289691 502639
rect 289633 502599 289691 502605
rect 309045 502639 309103 502645
rect 309045 502605 309057 502639
rect 309091 502636 309103 502639
rect 311805 502639 311863 502645
rect 311805 502636 311817 502639
rect 309091 502608 311817 502636
rect 309091 502605 309103 502608
rect 309045 502599 309103 502605
rect 311805 502605 311817 502608
rect 311851 502605 311863 502639
rect 311805 502599 311863 502605
rect 311897 502639 311955 502645
rect 311897 502605 311909 502639
rect 311943 502636 311955 502639
rect 311943 502608 312124 502636
rect 311943 502605 311955 502608
rect 311897 502599 311955 502605
rect 312096 502568 312124 502608
rect 320266 502568 320272 502580
rect 312096 502540 320272 502568
rect 320266 502528 320272 502540
rect 320324 502528 320330 502580
rect 276750 502460 276756 502512
rect 276808 502500 276814 502512
rect 280157 502503 280215 502509
rect 280157 502500 280169 502503
rect 276808 502472 280169 502500
rect 276808 502460 276814 502472
rect 280157 502469 280169 502472
rect 280203 502469 280215 502503
rect 280157 502463 280215 502469
rect 289633 502367 289691 502373
rect 289633 502333 289645 502367
rect 289679 502364 289691 502367
rect 289817 502367 289875 502373
rect 289817 502364 289829 502367
rect 289679 502336 289829 502364
rect 289679 502333 289691 502336
rect 289633 502327 289691 502333
rect 289817 502333 289829 502336
rect 289863 502333 289875 502367
rect 289817 502327 289875 502333
rect 273622 501032 273628 501084
rect 273680 501072 273686 501084
rect 290458 501072 290464 501084
rect 273680 501044 290464 501072
rect 273680 501032 273686 501044
rect 290458 501032 290464 501044
rect 290516 501032 290522 501084
rect 276842 500964 276848 501016
rect 276900 501004 276906 501016
rect 319806 501004 319812 501016
rect 276900 500976 319812 501004
rect 276900 500964 276906 500976
rect 319806 500964 319812 500976
rect 319864 500964 319870 501016
rect 273714 499604 273720 499656
rect 273772 499644 273778 499656
rect 287698 499644 287704 499656
rect 273772 499616 287704 499644
rect 273772 499604 273778 499616
rect 287698 499604 287704 499616
rect 287756 499604 287762 499656
rect 276934 499536 276940 499588
rect 276992 499576 276998 499588
rect 320174 499576 320180 499588
rect 276992 499548 320180 499576
rect 276992 499536 276998 499548
rect 320174 499536 320180 499548
rect 320232 499536 320238 499588
rect 277026 498176 277032 498228
rect 277084 498216 277090 498228
rect 319806 498216 319812 498228
rect 277084 498188 319812 498216
rect 277084 498176 277090 498188
rect 319806 498176 319812 498188
rect 319864 498176 319870 498228
rect 273714 496884 273720 496936
rect 273772 496924 273778 496936
rect 286318 496924 286324 496936
rect 273772 496896 286324 496924
rect 273772 496884 273778 496896
rect 286318 496884 286324 496896
rect 286376 496884 286382 496936
rect 278590 496816 278596 496868
rect 278648 496856 278654 496868
rect 320174 496856 320180 496868
rect 278648 496828 320180 496856
rect 278648 496816 278654 496828
rect 320174 496816 320180 496828
rect 320232 496816 320238 496868
rect 273714 495592 273720 495644
rect 273772 495632 273778 495644
rect 284938 495632 284944 495644
rect 273772 495604 284944 495632
rect 273772 495592 273778 495604
rect 284938 495592 284944 495604
rect 284996 495592 285002 495644
rect 279510 495524 279516 495576
rect 279568 495564 279574 495576
rect 319806 495564 319812 495576
rect 279568 495536 319812 495564
rect 279568 495524 279574 495536
rect 319806 495524 319812 495536
rect 319864 495524 319870 495576
rect 275738 495456 275744 495508
rect 275796 495496 275802 495508
rect 319990 495496 319996 495508
rect 275796 495468 319996 495496
rect 275796 495456 275802 495468
rect 319990 495456 319996 495468
rect 320048 495456 320054 495508
rect 320634 495496 320640 495508
rect 320595 495468 320640 495496
rect 320634 495456 320640 495468
rect 320692 495456 320698 495508
rect 273622 494096 273628 494148
rect 273680 494136 273686 494148
rect 278038 494136 278044 494148
rect 273680 494108 278044 494136
rect 273680 494096 273686 494108
rect 278038 494096 278044 494108
rect 278096 494096 278102 494148
rect 275830 494028 275836 494080
rect 275888 494068 275894 494080
rect 319806 494068 319812 494080
rect 275888 494040 319812 494068
rect 275888 494028 275894 494040
rect 319806 494028 319812 494040
rect 319864 494028 319870 494080
rect 275922 492668 275928 492720
rect 275980 492708 275986 492720
rect 320174 492708 320180 492720
rect 275980 492680 320180 492708
rect 275980 492668 275986 492680
rect 320174 492668 320180 492680
rect 320232 492668 320238 492720
rect 320726 492328 320732 492380
rect 320784 492328 320790 492380
rect 320818 492328 320824 492380
rect 320876 492328 320882 492380
rect 320744 492176 320772 492328
rect 320836 492176 320864 492328
rect 320726 492124 320732 492176
rect 320784 492124 320790 492176
rect 320818 492124 320824 492176
rect 320876 492124 320882 492176
rect 273622 491376 273628 491428
rect 273680 491416 273686 491428
rect 283558 491416 283564 491428
rect 273680 491388 283564 491416
rect 273680 491376 273686 491388
rect 283558 491376 283564 491388
rect 283616 491376 283622 491428
rect 275186 491308 275192 491360
rect 275244 491348 275250 491360
rect 319806 491348 319812 491360
rect 275244 491320 319812 491348
rect 275244 491308 275250 491320
rect 319806 491308 319812 491320
rect 319864 491308 319870 491360
rect 320634 490940 320640 490952
rect 320595 490912 320640 490940
rect 320634 490900 320640 490912
rect 320692 490900 320698 490952
rect 273438 489948 273444 490000
rect 273496 489988 273502 490000
rect 280798 489988 280804 490000
rect 273496 489960 280804 489988
rect 273496 489948 273502 489960
rect 280798 489948 280804 489960
rect 280856 489948 280862 490000
rect 275094 489880 275100 489932
rect 275152 489920 275158 489932
rect 320174 489920 320180 489932
rect 275152 489892 320180 489920
rect 275152 489880 275158 489892
rect 320174 489880 320180 489892
rect 320232 489880 320238 489932
rect 320634 489920 320640 489932
rect 320595 489892 320640 489920
rect 320634 489880 320640 489892
rect 320692 489880 320698 489932
rect 320082 489812 320088 489864
rect 320140 489852 320146 489864
rect 320726 489852 320732 489864
rect 320140 489824 320732 489852
rect 320140 489812 320146 489824
rect 320726 489812 320732 489824
rect 320784 489812 320790 489864
rect 320818 489812 320824 489864
rect 320876 489852 320882 489864
rect 320876 489824 320921 489852
rect 320876 489812 320882 489824
rect 320744 489716 320772 489812
rect 320744 489688 320864 489716
rect 320836 489456 320864 489688
rect 320818 489404 320824 489456
rect 320876 489404 320882 489456
rect 273622 488656 273628 488708
rect 273680 488696 273686 488708
rect 278130 488696 278136 488708
rect 273680 488668 278136 488696
rect 273680 488656 273686 488668
rect 278130 488656 278136 488668
rect 278188 488656 278194 488708
rect 275002 488588 275008 488640
rect 275060 488628 275066 488640
rect 319806 488628 319812 488640
rect 275060 488600 319812 488628
rect 275060 488588 275066 488600
rect 319806 488588 319812 488600
rect 319864 488588 319870 488640
rect 274910 488520 274916 488572
rect 274968 488560 274974 488572
rect 319714 488560 319720 488572
rect 274968 488532 319720 488560
rect 274968 488520 274974 488532
rect 319714 488520 319720 488532
rect 319772 488520 319778 488572
rect 320450 487228 320456 487280
rect 320508 487268 320514 487280
rect 320821 487271 320879 487277
rect 320821 487268 320833 487271
rect 320508 487240 320833 487268
rect 320508 487228 320514 487240
rect 320821 487237 320833 487240
rect 320867 487237 320879 487271
rect 320821 487231 320879 487237
rect 274818 487160 274824 487212
rect 274876 487200 274882 487212
rect 320174 487200 320180 487212
rect 274876 487172 320180 487200
rect 274876 487160 274882 487172
rect 320174 487160 320180 487172
rect 320232 487160 320238 487212
rect 320542 486208 320548 486260
rect 320600 486208 320606 486260
rect 320634 486208 320640 486260
rect 320692 486208 320698 486260
rect 320560 486056 320588 486208
rect 320652 486056 320680 486208
rect 320542 486004 320548 486056
rect 320600 486004 320606 486056
rect 320634 486004 320640 486056
rect 320692 486004 320698 486056
rect 273530 485868 273536 485920
rect 273588 485908 273594 485920
rect 278222 485908 278228 485920
rect 273588 485880 278228 485908
rect 273588 485868 273594 485880
rect 278222 485868 278228 485880
rect 278280 485868 278286 485920
rect 274726 485800 274732 485852
rect 274784 485840 274790 485852
rect 319806 485840 319812 485852
rect 274784 485812 319812 485840
rect 274784 485800 274790 485812
rect 319806 485800 319812 485812
rect 319864 485800 319870 485852
rect 273622 484440 273628 484492
rect 273680 484480 273686 484492
rect 278314 484480 278320 484492
rect 273680 484452 278320 484480
rect 273680 484440 273686 484452
rect 278314 484440 278320 484452
rect 278372 484440 278378 484492
rect 274634 484372 274640 484424
rect 274692 484412 274698 484424
rect 320174 484412 320180 484424
rect 274692 484384 320180 484412
rect 274692 484372 274698 484384
rect 320174 484372 320180 484384
rect 320232 484372 320238 484424
rect 277210 483012 277216 483064
rect 277268 483052 277274 483064
rect 319806 483052 319812 483064
rect 277268 483024 319812 483052
rect 277268 483012 277274 483024
rect 319806 483012 319812 483024
rect 319864 483012 319870 483064
rect 320450 482848 320456 482860
rect 320411 482820 320456 482848
rect 320450 482808 320456 482820
rect 320508 482808 320514 482860
rect 320450 482672 320456 482724
rect 320508 482712 320514 482724
rect 320634 482712 320640 482724
rect 320508 482684 320640 482712
rect 320508 482672 320514 482684
rect 320634 482672 320640 482684
rect 320692 482672 320698 482724
rect 320818 482672 320824 482724
rect 320876 482672 320882 482724
rect 320542 482332 320548 482384
rect 320600 482372 320606 482384
rect 320836 482372 320864 482672
rect 320600 482344 320864 482372
rect 320600 482332 320606 482344
rect 273622 481720 273628 481772
rect 273680 481760 273686 481772
rect 278406 481760 278412 481772
rect 273680 481732 278412 481760
rect 273680 481720 273686 481732
rect 278406 481720 278412 481732
rect 278464 481720 278470 481772
rect 277302 481652 277308 481704
rect 277360 481692 277366 481704
rect 320174 481692 320180 481704
rect 277360 481664 320180 481692
rect 277360 481652 277366 481664
rect 320174 481652 320180 481664
rect 320232 481652 320238 481704
rect 320266 480428 320272 480480
rect 320324 480468 320330 480480
rect 320818 480468 320824 480480
rect 320324 480440 320824 480468
rect 320324 480428 320330 480440
rect 320818 480428 320824 480440
rect 320876 480428 320882 480480
rect 273622 480292 273628 480344
rect 273680 480332 273686 480344
rect 278498 480332 278504 480344
rect 273680 480304 278504 480332
rect 273680 480292 273686 480304
rect 278498 480292 278504 480304
rect 278556 480292 278562 480344
rect 320266 480292 320272 480344
rect 320324 480332 320330 480344
rect 320453 480335 320511 480341
rect 320453 480332 320465 480335
rect 320324 480304 320465 480332
rect 320324 480292 320330 480304
rect 320453 480301 320465 480304
rect 320499 480301 320511 480335
rect 320453 480295 320511 480301
rect 276566 480224 276572 480276
rect 276624 480264 276630 480276
rect 319806 480264 319812 480276
rect 276624 480236 319812 480264
rect 276624 480224 276630 480236
rect 319806 480224 319812 480236
rect 319864 480224 319870 480276
rect 320818 479448 320824 479460
rect 320779 479420 320824 479448
rect 320818 479408 320824 479420
rect 320876 479408 320882 479460
rect 320174 479272 320180 479324
rect 320232 479312 320238 479324
rect 320818 479312 320824 479324
rect 320232 479284 320824 479312
rect 320232 479272 320238 479284
rect 320818 479272 320824 479284
rect 320876 479272 320882 479324
rect 320634 478932 320640 478984
rect 320692 478972 320698 478984
rect 320821 478975 320879 478981
rect 320821 478972 320833 478975
rect 320692 478944 320833 478972
rect 320692 478932 320698 478944
rect 320821 478941 320833 478944
rect 320867 478941 320879 478975
rect 320821 478935 320879 478941
rect 273622 478864 273628 478916
rect 273680 478904 273686 478916
rect 315298 478904 315304 478916
rect 273680 478876 315304 478904
rect 273680 478864 273686 478876
rect 315298 478864 315304 478876
rect 315356 478864 315362 478916
rect 320450 476960 320456 477012
rect 320508 477000 320514 477012
rect 320634 477000 320640 477012
rect 320508 476972 320640 477000
rect 320508 476960 320514 476972
rect 320634 476960 320640 476972
rect 320692 476960 320698 477012
rect 320174 476824 320180 476876
rect 320232 476824 320238 476876
rect 320192 476660 320220 476824
rect 320266 476660 320272 476672
rect 320192 476632 320272 476660
rect 320266 476620 320272 476632
rect 320324 476620 320330 476672
rect 273622 476076 273628 476128
rect 273680 476116 273686 476128
rect 312538 476116 312544 476128
rect 273680 476088 312544 476116
rect 273680 476076 273686 476088
rect 312538 476076 312544 476088
rect 312596 476076 312602 476128
rect 320726 476048 320732 476060
rect 320687 476020 320732 476048
rect 320726 476008 320732 476020
rect 320784 476008 320790 476060
rect 320634 475872 320640 475924
rect 320692 475872 320698 475924
rect 320450 475804 320456 475856
rect 320508 475844 320514 475856
rect 320652 475844 320680 475872
rect 320508 475816 320680 475844
rect 320508 475804 320514 475816
rect 320818 475776 320824 475788
rect 320779 475748 320824 475776
rect 320818 475736 320824 475748
rect 320876 475736 320882 475788
rect 273622 474784 273628 474836
rect 273680 474824 273686 474836
rect 309778 474824 309784 474836
rect 273680 474796 309784 474824
rect 273680 474784 273686 474796
rect 309778 474784 309784 474796
rect 309836 474784 309842 474836
rect 276474 474716 276480 474768
rect 276532 474756 276538 474768
rect 320174 474756 320180 474768
rect 276532 474728 320180 474756
rect 276532 474716 276538 474728
rect 320174 474716 320180 474728
rect 320232 474716 320238 474768
rect 273530 473968 273536 474020
rect 273588 474008 273594 474020
rect 320358 474008 320364 474020
rect 273588 473980 320364 474008
rect 273588 473968 273594 473980
rect 320358 473968 320364 473980
rect 320416 473968 320422 474020
rect 273622 473356 273628 473408
rect 273680 473396 273686 473408
rect 308398 473396 308404 473408
rect 273680 473368 308404 473396
rect 273680 473356 273686 473368
rect 308398 473356 308404 473368
rect 308456 473356 308462 473408
rect 273438 471996 273444 472048
rect 273496 472036 273502 472048
rect 320174 472036 320180 472048
rect 273496 472008 320180 472036
rect 273496 471996 273502 472008
rect 320174 471996 320180 472008
rect 320232 471996 320238 472048
rect 273530 470636 273536 470688
rect 273588 470676 273594 470688
rect 305638 470676 305644 470688
rect 273588 470648 305644 470676
rect 273588 470636 273594 470648
rect 305638 470636 305644 470648
rect 305696 470636 305702 470688
rect 273346 470568 273352 470620
rect 273404 470608 273410 470620
rect 320266 470608 320272 470620
rect 273404 470580 320272 470608
rect 273404 470568 273410 470580
rect 320266 470568 320272 470580
rect 320324 470568 320330 470620
rect 320266 470432 320272 470484
rect 320324 470472 320330 470484
rect 320729 470475 320787 470481
rect 320729 470472 320741 470475
rect 320324 470444 320741 470472
rect 320324 470432 320330 470444
rect 320729 470441 320741 470444
rect 320775 470441 320787 470475
rect 320729 470435 320787 470441
rect 273530 469276 273536 469328
rect 273588 469316 273594 469328
rect 304258 469316 304264 469328
rect 273588 469288 304264 469316
rect 273588 469276 273594 469288
rect 304258 469276 304264 469288
rect 304316 469276 304322 469328
rect 276382 469208 276388 469260
rect 276440 469248 276446 469260
rect 320358 469248 320364 469260
rect 276440 469220 320364 469248
rect 276440 469208 276446 469220
rect 320358 469208 320364 469220
rect 320416 469208 320422 469260
rect 276290 467916 276296 467968
rect 276348 467956 276354 467968
rect 320450 467956 320456 467968
rect 276348 467928 320456 467956
rect 276348 467916 276354 467928
rect 320450 467916 320456 467928
rect 320508 467916 320514 467968
rect 276198 467848 276204 467900
rect 276256 467888 276262 467900
rect 320266 467888 320272 467900
rect 276256 467860 320272 467888
rect 276256 467848 276262 467860
rect 320266 467848 320272 467860
rect 320324 467848 320330 467900
rect 320361 467823 320419 467829
rect 320361 467789 320373 467823
rect 320407 467820 320419 467823
rect 320542 467820 320548 467832
rect 320407 467792 320548 467820
rect 320407 467789 320419 467792
rect 320361 467783 320419 467789
rect 320542 467780 320548 467792
rect 320600 467780 320606 467832
rect 320266 467712 320272 467764
rect 320324 467752 320330 467764
rect 320726 467752 320732 467764
rect 320324 467724 320732 467752
rect 320324 467712 320330 467724
rect 320726 467712 320732 467724
rect 320784 467712 320790 467764
rect 320082 467644 320088 467696
rect 320140 467684 320146 467696
rect 320542 467684 320548 467696
rect 320140 467656 320548 467684
rect 320140 467644 320146 467656
rect 320542 467644 320548 467656
rect 320600 467644 320606 467696
rect 320358 467616 320364 467628
rect 320319 467588 320364 467616
rect 320358 467576 320364 467588
rect 320416 467576 320422 467628
rect 320634 467508 320640 467560
rect 320692 467548 320698 467560
rect 320729 467551 320787 467557
rect 320729 467548 320741 467551
rect 320692 467520 320741 467548
rect 320692 467508 320698 467520
rect 320729 467517 320741 467520
rect 320775 467517 320787 467551
rect 320729 467511 320787 467517
rect 320726 467372 320732 467424
rect 320784 467412 320790 467424
rect 320821 467415 320879 467421
rect 320821 467412 320833 467415
rect 320784 467384 320833 467412
rect 320784 467372 320790 467384
rect 320821 467381 320833 467384
rect 320867 467381 320879 467415
rect 320821 467375 320879 467381
rect 273530 466488 273536 466540
rect 273588 466528 273594 466540
rect 302970 466528 302976 466540
rect 273588 466500 302976 466528
rect 273588 466488 273594 466500
rect 302970 466488 302976 466500
rect 303028 466488 303034 466540
rect 276106 466420 276112 466472
rect 276164 466460 276170 466472
rect 320174 466460 320180 466472
rect 276164 466432 320180 466460
rect 276164 466420 276170 466432
rect 320174 466420 320180 466432
rect 320232 466420 320238 466472
rect 276014 465060 276020 465112
rect 276072 465100 276078 465112
rect 320174 465100 320180 465112
rect 276072 465072 320180 465100
rect 276072 465060 276078 465072
rect 320174 465060 320180 465072
rect 320232 465060 320238 465112
rect 273254 463700 273260 463752
rect 273312 463740 273318 463752
rect 277118 463740 277124 463752
rect 273312 463712 277124 463740
rect 273312 463700 273318 463712
rect 277118 463700 277124 463712
rect 277176 463700 277182 463752
rect 273254 460912 273260 460964
rect 273312 460952 273318 460964
rect 278682 460952 278688 460964
rect 273312 460924 278688 460952
rect 273312 460912 273318 460924
rect 278682 460912 278688 460924
rect 278740 460912 278746 460964
rect 273254 460028 273260 460080
rect 273312 460068 273318 460080
rect 276014 460068 276020 460080
rect 273312 460040 276020 460068
rect 273312 460028 273318 460040
rect 276014 460028 276020 460040
rect 276072 460028 276078 460080
rect 273254 458124 273260 458176
rect 273312 458164 273318 458176
rect 276106 458164 276112 458176
rect 273312 458136 276112 458164
rect 273312 458124 273318 458136
rect 276106 458124 276112 458136
rect 276164 458124 276170 458176
rect 320269 457487 320327 457493
rect 320269 457453 320281 457487
rect 320315 457484 320327 457487
rect 320450 457484 320456 457496
rect 320315 457456 320456 457484
rect 320315 457453 320327 457456
rect 320269 457447 320327 457453
rect 320450 457444 320456 457456
rect 320508 457444 320514 457496
rect 320634 457444 320640 457496
rect 320692 457484 320698 457496
rect 320729 457487 320787 457493
rect 320729 457484 320741 457487
rect 320692 457456 320741 457484
rect 320692 457444 320698 457456
rect 320729 457453 320741 457456
rect 320775 457453 320787 457487
rect 320729 457447 320787 457453
rect 320637 457351 320695 457357
rect 320637 457317 320649 457351
rect 320683 457348 320695 457351
rect 320818 457348 320824 457360
rect 320683 457320 320824 457348
rect 320683 457317 320695 457320
rect 320637 457311 320695 457317
rect 320818 457308 320824 457320
rect 320876 457308 320882 457360
rect 320174 457104 320180 457156
rect 320232 457104 320238 457156
rect 320192 456872 320220 457104
rect 320358 456940 320364 456952
rect 320319 456912 320364 456940
rect 320358 456900 320364 456912
rect 320416 456900 320422 456952
rect 320726 456900 320732 456952
rect 320784 456940 320790 456952
rect 320821 456943 320879 456949
rect 320821 456940 320833 456943
rect 320784 456912 320833 456940
rect 320784 456900 320790 456912
rect 320821 456909 320833 456912
rect 320867 456909 320879 456943
rect 320821 456903 320879 456909
rect 320192 456844 320772 456872
rect 320358 456668 320364 456680
rect 320319 456640 320364 456668
rect 320358 456628 320364 456640
rect 320416 456628 320422 456680
rect 320450 456628 320456 456680
rect 320508 456668 320514 456680
rect 320744 456668 320772 456844
rect 320508 456640 320772 456668
rect 320508 456628 320514 456640
rect 320634 456492 320640 456544
rect 320692 456532 320698 456544
rect 320821 456535 320879 456541
rect 320821 456532 320833 456535
rect 320692 456504 320833 456532
rect 320692 456492 320698 456504
rect 320821 456501 320833 456504
rect 320867 456501 320879 456535
rect 320821 456495 320879 456501
rect 273254 456220 273260 456272
rect 273312 456260 273318 456272
rect 276198 456260 276204 456272
rect 273312 456232 276204 456260
rect 273312 456220 273318 456232
rect 276198 456220 276204 456232
rect 276256 456220 276262 456272
rect 273254 454316 273260 454368
rect 273312 454356 273318 454368
rect 276290 454356 276296 454368
rect 273312 454328 276296 454356
rect 273312 454316 273318 454328
rect 276290 454316 276296 454328
rect 276348 454316 276354 454368
rect 320637 452659 320695 452665
rect 320637 452625 320649 452659
rect 320683 452656 320695 452659
rect 320821 452659 320879 452665
rect 320821 452656 320833 452659
rect 320683 452628 320833 452656
rect 320683 452625 320695 452628
rect 320637 452619 320695 452625
rect 320821 452625 320833 452628
rect 320867 452625 320879 452659
rect 320821 452619 320879 452625
rect 273254 452412 273260 452464
rect 273312 452452 273318 452464
rect 276382 452452 276388 452464
rect 273312 452424 276388 452452
rect 273312 452412 273318 452424
rect 276382 452412 276388 452424
rect 276440 452412 276446 452464
rect 320174 452316 320180 452328
rect 320135 452288 320180 452316
rect 320174 452276 320180 452288
rect 320232 452276 320238 452328
rect 320634 449868 320640 449880
rect 320595 449840 320640 449868
rect 320634 449828 320640 449840
rect 320692 449828 320698 449880
rect 320358 447352 320364 447364
rect 320319 447324 320364 447352
rect 320358 447312 320364 447324
rect 320416 447312 320422 447364
rect 320450 447312 320456 447364
rect 320508 447312 320514 447364
rect 320542 447312 320548 447364
rect 320600 447312 320606 447364
rect 320468 447228 320496 447312
rect 320560 447228 320588 447312
rect 320450 447176 320456 447228
rect 320508 447176 320514 447228
rect 320542 447176 320548 447228
rect 320600 447176 320606 447228
rect 320634 447108 320640 447160
rect 320692 447148 320698 447160
rect 320729 447151 320787 447157
rect 320729 447148 320741 447151
rect 320692 447120 320741 447148
rect 320692 447108 320698 447120
rect 320729 447117 320741 447120
rect 320775 447117 320787 447151
rect 320729 447111 320787 447117
rect 273438 447040 273444 447092
rect 273496 447080 273502 447092
rect 320821 447083 320879 447089
rect 320821 447080 320833 447083
rect 273496 447052 320833 447080
rect 273496 447040 273502 447052
rect 320821 447049 320833 447052
rect 320867 447049 320879 447083
rect 320821 447043 320879 447049
rect 320358 447012 320364 447024
rect 320319 446984 320364 447012
rect 320358 446972 320364 446984
rect 320416 446972 320422 447024
rect 320637 446947 320695 446953
rect 320637 446913 320649 446947
rect 320683 446944 320695 446947
rect 320818 446944 320824 446956
rect 320683 446916 320824 446944
rect 320683 446913 320695 446916
rect 320637 446907 320695 446913
rect 320818 446904 320824 446916
rect 320876 446904 320882 446956
rect 320269 446879 320327 446885
rect 320269 446845 320281 446879
rect 320315 446876 320327 446879
rect 320726 446876 320732 446888
rect 320315 446848 320732 446876
rect 320315 446845 320327 446848
rect 320269 446839 320327 446845
rect 320726 446836 320732 446848
rect 320784 446836 320790 446888
rect 320177 446811 320235 446817
rect 320177 446777 320189 446811
rect 320223 446808 320235 446811
rect 320818 446808 320824 446820
rect 320223 446780 320824 446808
rect 320223 446777 320235 446780
rect 320177 446771 320235 446777
rect 320818 446768 320824 446780
rect 320876 446768 320882 446820
rect 273438 444796 273444 444848
rect 273496 444836 273502 444848
rect 276474 444836 276480 444848
rect 273496 444808 276480 444836
rect 273496 444796 273502 444808
rect 276474 444796 276480 444808
rect 276532 444796 276538 444848
rect 273438 442892 273444 442944
rect 273496 442932 273502 442944
rect 276566 442932 276572 442944
rect 273496 442904 276572 442932
rect 273496 442892 273502 442904
rect 276566 442892 276572 442904
rect 276624 442892 276630 442944
rect 320542 442416 320548 442468
rect 320600 442416 320606 442468
rect 320726 442416 320732 442468
rect 320784 442416 320790 442468
rect 320560 442196 320588 442416
rect 320542 442144 320548 442196
rect 320600 442144 320606 442196
rect 320450 442008 320456 442060
rect 320508 442048 320514 442060
rect 320744 442048 320772 442416
rect 320508 442020 320772 442048
rect 320508 442008 320514 442020
rect 273438 441260 273444 441312
rect 273496 441300 273502 441312
rect 277302 441300 277308 441312
rect 273496 441272 277308 441300
rect 273496 441260 273502 441272
rect 277302 441260 277308 441272
rect 277360 441260 277366 441312
rect 273438 439696 273444 439748
rect 273496 439736 273502 439748
rect 277210 439736 277216 439748
rect 273496 439708 277216 439736
rect 273496 439696 273502 439708
rect 277210 439696 277216 439708
rect 277268 439696 277274 439748
rect 273254 433372 273260 433424
rect 273312 433412 273318 433424
rect 274818 433412 274824 433424
rect 273312 433384 274824 433412
rect 273312 433372 273318 433384
rect 274818 433372 274824 433384
rect 274876 433372 274882 433424
rect 320266 431944 320272 431996
rect 320324 431984 320330 431996
rect 320818 431984 320824 431996
rect 320324 431956 320824 431984
rect 320324 431944 320330 431956
rect 320818 431944 320824 431956
rect 320876 431944 320882 431996
rect 273254 431468 273260 431520
rect 273312 431508 273318 431520
rect 274910 431508 274916 431520
rect 273312 431480 274916 431508
rect 273312 431468 273318 431480
rect 274910 431468 274916 431480
rect 274968 431468 274974 431520
rect 273254 429564 273260 429616
rect 273312 429604 273318 429616
rect 275002 429604 275008 429616
rect 273312 429576 275008 429604
rect 273312 429564 273318 429576
rect 275002 429564 275008 429576
rect 275060 429564 275066 429616
rect 320266 427728 320272 427780
rect 320324 427768 320330 427780
rect 320818 427768 320824 427780
rect 320324 427740 320824 427768
rect 320324 427728 320330 427740
rect 320818 427728 320824 427740
rect 320876 427728 320882 427780
rect 273254 427660 273260 427712
rect 273312 427700 273318 427712
rect 275094 427700 275100 427712
rect 273312 427672 275100 427700
rect 273312 427660 273318 427672
rect 275094 427660 275100 427672
rect 275152 427660 275158 427712
rect 273254 425756 273260 425808
rect 273312 425796 273318 425808
rect 275186 425796 275192 425808
rect 273312 425768 275192 425796
rect 273312 425756 273318 425768
rect 275186 425756 275192 425768
rect 275244 425756 275250 425808
rect 273438 423988 273444 424040
rect 273496 424028 273502 424040
rect 275922 424028 275928 424040
rect 273496 424000 275928 424028
rect 273496 423988 273502 424000
rect 275922 423988 275928 424000
rect 275980 423988 275986 424040
rect 273438 422016 273444 422068
rect 273496 422056 273502 422068
rect 275830 422056 275836 422068
rect 273496 422028 275836 422056
rect 273496 422016 273502 422028
rect 275830 422016 275836 422028
rect 275888 422016 275894 422068
rect 273438 420044 273444 420096
rect 273496 420084 273502 420096
rect 275738 420084 275744 420096
rect 273496 420056 275744 420084
rect 273496 420044 273502 420056
rect 275738 420044 275744 420056
rect 275796 420044 275802 420096
rect 273438 418072 273444 418124
rect 273496 418112 273502 418124
rect 279510 418112 279516 418124
rect 273496 418084 279516 418112
rect 273496 418072 273502 418084
rect 279510 418072 279516 418084
rect 279568 418072 279574 418124
rect 273438 416236 273444 416288
rect 273496 416276 273502 416288
rect 278590 416276 278596 416288
rect 273496 416248 278596 416276
rect 273496 416236 273502 416248
rect 278590 416236 278596 416248
rect 278648 416236 278654 416288
rect 273438 414332 273444 414384
rect 273496 414372 273502 414384
rect 277026 414372 277032 414384
rect 273496 414344 277032 414372
rect 273496 414332 273502 414344
rect 277026 414332 277032 414344
rect 277084 414332 277090 414384
rect 273438 412428 273444 412480
rect 273496 412468 273502 412480
rect 276934 412468 276940 412480
rect 273496 412440 276940 412468
rect 273496 412428 273502 412440
rect 276934 412428 276940 412440
rect 276992 412428 276998 412480
rect 273438 410524 273444 410576
rect 273496 410564 273502 410576
rect 276842 410564 276848 410576
rect 273496 410536 276848 410564
rect 273496 410524 273502 410536
rect 276842 410524 276848 410536
rect 276900 410524 276906 410576
rect 273438 408620 273444 408672
rect 273496 408660 273502 408672
rect 276750 408660 276756 408672
rect 273496 408632 276756 408660
rect 273496 408620 273502 408632
rect 276750 408620 276756 408632
rect 276808 408620 276814 408672
rect 273438 406716 273444 406768
rect 273496 406756 273502 406768
rect 276658 406756 276664 406768
rect 273496 406728 276664 406756
rect 273496 406716 273502 406728
rect 276658 406716 276664 406728
rect 276716 406716 276722 406768
rect 273438 402908 273444 402960
rect 273496 402948 273502 402960
rect 275646 402948 275652 402960
rect 273496 402920 275652 402948
rect 273496 402908 273502 402920
rect 275646 402908 275652 402920
rect 275704 402908 275710 402960
rect 273438 401004 273444 401056
rect 273496 401044 273502 401056
rect 275554 401044 275560 401056
rect 273496 401016 275560 401044
rect 273496 401004 273502 401016
rect 275554 401004 275560 401016
rect 275612 401004 275618 401056
rect 273438 400120 273444 400172
rect 273496 400160 273502 400172
rect 320726 400160 320732 400172
rect 273496 400132 320732 400160
rect 273496 400120 273502 400132
rect 320726 400120 320732 400132
rect 320784 400120 320790 400172
rect 320174 398828 320180 398880
rect 320232 398868 320238 398880
rect 320818 398868 320824 398880
rect 320232 398840 320824 398868
rect 320232 398828 320238 398840
rect 320818 398828 320824 398840
rect 320876 398828 320882 398880
rect 273438 397400 273444 397452
rect 273496 397440 273502 397452
rect 320634 397440 320640 397452
rect 273496 397412 320640 397440
rect 273496 397400 273502 397412
rect 320634 397400 320640 397412
rect 320692 397400 320698 397452
rect 273254 396788 273260 396840
rect 273312 396828 273318 396840
rect 338666 396828 338672 396840
rect 273312 396800 338672 396828
rect 273312 396788 273318 396800
rect 338666 396788 338672 396800
rect 338724 396788 338730 396840
rect 275738 396720 275744 396772
rect 275796 396760 275802 396772
rect 397454 396760 397460 396772
rect 275796 396732 397460 396760
rect 275796 396720 275802 396732
rect 397454 396720 397460 396732
rect 397512 396720 397518 396772
rect 275922 396652 275928 396704
rect 275980 396692 275986 396704
rect 398834 396692 398840 396704
rect 275980 396664 398840 396692
rect 275980 396652 275986 396664
rect 398834 396652 398840 396664
rect 398892 396652 398898 396704
rect 275186 396584 275192 396636
rect 275244 396624 275250 396636
rect 400214 396624 400220 396636
rect 275244 396596 400220 396624
rect 275244 396584 275250 396596
rect 400214 396584 400220 396596
rect 400272 396584 400278 396636
rect 275094 396516 275100 396568
rect 275152 396556 275158 396568
rect 401594 396556 401600 396568
rect 275152 396528 401600 396556
rect 275152 396516 275158 396528
rect 401594 396516 401600 396528
rect 401652 396516 401658 396568
rect 275002 396448 275008 396500
rect 275060 396488 275066 396500
rect 403342 396488 403348 396500
rect 275060 396460 403348 396488
rect 275060 396448 275066 396460
rect 403342 396448 403348 396460
rect 403400 396448 403406 396500
rect 274910 396380 274916 396432
rect 274968 396420 274974 396432
rect 404354 396420 404360 396432
rect 274968 396392 404360 396420
rect 274968 396380 274974 396392
rect 404354 396380 404360 396392
rect 404412 396380 404418 396432
rect 406010 396380 406016 396432
rect 406068 396380 406074 396432
rect 274818 396312 274824 396364
rect 274876 396352 274882 396364
rect 406028 396352 406056 396380
rect 274876 396324 406056 396352
rect 274876 396312 274882 396324
rect 273438 395972 273444 396024
rect 273496 396012 273502 396024
rect 320542 396012 320548 396024
rect 273496 395984 320548 396012
rect 273496 395972 273502 395984
rect 320542 395972 320548 395984
rect 320600 395972 320606 396024
rect 273438 394612 273444 394664
rect 273496 394652 273502 394664
rect 320450 394652 320456 394664
rect 273496 394624 320456 394652
rect 273496 394612 273502 394624
rect 320450 394612 320456 394624
rect 320508 394612 320514 394664
rect 275830 392028 275836 392080
rect 275888 392068 275894 392080
rect 320174 392068 320180 392080
rect 275888 392040 320180 392068
rect 275888 392028 275894 392040
rect 320174 392028 320180 392040
rect 320232 392028 320238 392080
rect 275554 391960 275560 392012
rect 275612 392000 275618 392012
rect 320266 392000 320272 392012
rect 275612 391972 320272 392000
rect 275612 391960 275618 391972
rect 320266 391960 320272 391972
rect 320324 391960 320330 392012
rect 273438 391892 273444 391944
rect 273496 391932 273502 391944
rect 320358 391932 320364 391944
rect 273496 391904 320364 391932
rect 273496 391892 273502 391904
rect 320358 391892 320364 391904
rect 320416 391892 320422 391944
rect 275646 390532 275652 390584
rect 275704 390572 275710 390584
rect 320082 390572 320088 390584
rect 275704 390544 320088 390572
rect 275704 390532 275710 390544
rect 320082 390532 320088 390544
rect 320140 390532 320146 390584
rect 273530 390464 273536 390516
rect 273588 390504 273594 390516
rect 320174 390504 320180 390516
rect 273588 390476 320180 390504
rect 273588 390464 273594 390476
rect 320174 390464 320180 390476
rect 320232 390464 320238 390516
rect 273438 389172 273444 389224
rect 273496 389212 273502 389224
rect 320266 389212 320272 389224
rect 273496 389184 320272 389212
rect 273496 389172 273502 389184
rect 320266 389172 320272 389184
rect 320324 389172 320330 389224
rect 273346 388016 273352 388068
rect 273404 388056 273410 388068
rect 273530 388056 273536 388068
rect 273404 388028 273536 388056
rect 273404 388016 273410 388028
rect 273530 388016 273536 388028
rect 273588 388016 273594 388068
rect 320174 387852 320180 387864
rect 273548 387824 320180 387852
rect 273548 387580 273576 387824
rect 320174 387812 320180 387824
rect 320232 387812 320238 387864
rect 273622 387744 273628 387796
rect 273680 387784 273686 387796
rect 320818 387784 320824 387796
rect 273680 387756 320824 387784
rect 273680 387744 273686 387756
rect 320818 387744 320824 387756
rect 320876 387744 320882 387796
rect 278682 387676 278688 387728
rect 278740 387716 278746 387728
rect 320358 387716 320364 387728
rect 278740 387688 320364 387716
rect 278740 387676 278746 387688
rect 320358 387676 320364 387688
rect 320416 387676 320422 387728
rect 273622 387580 273628 387592
rect 273548 387552 273628 387580
rect 273622 387540 273628 387552
rect 273680 387540 273686 387592
rect 277118 386316 277124 386368
rect 277176 386356 277182 386368
rect 320266 386356 320272 386368
rect 277176 386328 320272 386356
rect 277176 386316 277182 386328
rect 320266 386316 320272 386328
rect 320324 386316 320330 386368
rect 273346 384956 273352 385008
rect 273404 384996 273410 385008
rect 320174 384996 320180 385008
rect 273404 384968 320180 384996
rect 273404 384956 273410 384968
rect 320174 384956 320180 384968
rect 320232 384956 320238 385008
rect 302970 384888 302976 384940
rect 303028 384928 303034 384940
rect 320358 384928 320364 384940
rect 303028 384900 320364 384928
rect 303028 384888 303034 384900
rect 320358 384888 320364 384900
rect 320416 384888 320422 384940
rect 304258 383596 304264 383648
rect 304316 383636 304322 383648
rect 320174 383636 320180 383648
rect 304316 383608 320180 383636
rect 304316 383596 304322 383608
rect 320174 383596 320180 383608
rect 320232 383596 320238 383648
rect 273346 383528 273352 383580
rect 273404 383528 273410 383580
rect 273364 383364 273392 383528
rect 273438 383364 273444 383376
rect 273364 383336 273444 383364
rect 273438 383324 273444 383336
rect 273496 383324 273502 383376
rect 305638 382168 305644 382220
rect 305696 382208 305702 382220
rect 320542 382208 320548 382220
rect 305696 382180 320548 382208
rect 305696 382168 305702 382180
rect 320542 382168 320548 382180
rect 320600 382168 320606 382220
rect 320634 381352 320640 381404
rect 320692 381392 320698 381404
rect 320729 381395 320787 381401
rect 320729 381392 320741 381395
rect 320692 381364 320741 381392
rect 320692 381352 320698 381364
rect 320729 381361 320741 381364
rect 320775 381361 320787 381395
rect 320729 381355 320787 381361
rect 308398 380808 308404 380860
rect 308456 380848 308462 380860
rect 320174 380848 320180 380860
rect 308456 380820 320180 380848
rect 308456 380808 308462 380820
rect 320174 380808 320180 380820
rect 320232 380808 320238 380860
rect 320818 380304 320824 380316
rect 320779 380276 320824 380304
rect 320818 380264 320824 380276
rect 320876 380264 320882 380316
rect 273530 380196 273536 380248
rect 273588 380236 273594 380248
rect 320082 380236 320088 380248
rect 273588 380208 320088 380236
rect 273588 380196 273594 380208
rect 320082 380196 320088 380208
rect 320140 380196 320146 380248
rect 273622 380128 273628 380180
rect 273680 380168 273686 380180
rect 320450 380168 320456 380180
rect 273680 380140 320456 380168
rect 273680 380128 273686 380140
rect 320450 380128 320456 380140
rect 320508 380128 320514 380180
rect 320634 379760 320640 379772
rect 320595 379732 320640 379760
rect 320634 379720 320640 379732
rect 320692 379720 320698 379772
rect 320726 379556 320732 379568
rect 320687 379528 320732 379556
rect 320726 379516 320732 379528
rect 320784 379516 320790 379568
rect 309778 379448 309784 379500
rect 309836 379488 309842 379500
rect 320266 379488 320272 379500
rect 309836 379460 320272 379488
rect 309836 379448 309842 379460
rect 320266 379448 320272 379460
rect 320324 379448 320330 379500
rect 273530 378904 273536 378956
rect 273588 378944 273594 378956
rect 274450 378944 274456 378956
rect 273588 378916 274456 378944
rect 273588 378904 273594 378916
rect 274450 378904 274456 378916
rect 274508 378904 274514 378956
rect 274634 378836 274640 378888
rect 274692 378876 274698 378888
rect 320358 378876 320364 378888
rect 274692 378848 320364 378876
rect 274692 378836 274698 378848
rect 320358 378836 320364 378848
rect 320416 378836 320422 378888
rect 274450 378768 274456 378820
rect 274508 378808 274514 378820
rect 320818 378808 320824 378820
rect 274508 378780 320824 378808
rect 274508 378768 274514 378780
rect 320818 378768 320824 378780
rect 320876 378768 320882 378820
rect 320542 378292 320548 378344
rect 320600 378332 320606 378344
rect 320637 378335 320695 378341
rect 320637 378332 320649 378335
rect 320600 378304 320649 378332
rect 320600 378292 320606 378304
rect 320637 378301 320649 378304
rect 320683 378301 320695 378335
rect 320637 378295 320695 378301
rect 315298 376796 315304 376848
rect 315356 376836 315362 376848
rect 319990 376836 319996 376848
rect 315356 376808 319996 376836
rect 315356 376796 315362 376808
rect 319990 376796 319996 376808
rect 320048 376796 320054 376848
rect 298097 376771 298155 376777
rect 298097 376737 298109 376771
rect 298143 376768 298155 376771
rect 302881 376771 302939 376777
rect 302881 376768 302893 376771
rect 298143 376740 302893 376768
rect 298143 376737 298155 376740
rect 298097 376731 298155 376737
rect 302881 376737 302893 376740
rect 302927 376737 302939 376771
rect 302881 376731 302939 376737
rect 312538 376728 312544 376780
rect 312596 376768 312602 376780
rect 319806 376768 319812 376780
rect 312596 376740 319812 376768
rect 312596 376728 312602 376740
rect 319806 376728 319812 376740
rect 319864 376728 319870 376780
rect 278590 376660 278596 376712
rect 278648 376700 278654 376712
rect 289725 376703 289783 376709
rect 289725 376700 289737 376703
rect 278648 376672 289737 376700
rect 278648 376660 278654 376672
rect 289725 376669 289737 376672
rect 289771 376669 289783 376703
rect 289725 376663 289783 376669
rect 289817 376703 289875 376709
rect 289817 376669 289829 376703
rect 289863 376700 289875 376703
rect 289863 376672 293264 376700
rect 289863 376669 289875 376672
rect 289817 376663 289875 376669
rect 293236 376632 293264 376672
rect 298097 376635 298155 376641
rect 298097 376632 298109 376635
rect 293236 376604 298109 376632
rect 298097 376601 298109 376604
rect 298143 376601 298155 376635
rect 298097 376595 298155 376601
rect 302881 376567 302939 376573
rect 302881 376533 302893 376567
rect 302927 376564 302939 376567
rect 320358 376564 320364 376576
rect 302927 376536 320364 376564
rect 302927 376533 302939 376536
rect 302881 376527 302939 376533
rect 320358 376524 320364 376536
rect 320416 376524 320422 376576
rect 274450 375980 274456 376032
rect 274508 376020 274514 376032
rect 320542 376020 320548 376032
rect 274508 375992 320548 376020
rect 274508 375980 274514 375992
rect 320542 375980 320548 375992
rect 320600 375980 320606 376032
rect 278406 375300 278412 375352
rect 278464 375340 278470 375352
rect 320266 375340 320272 375352
rect 278464 375312 320272 375340
rect 278464 375300 278470 375312
rect 320266 375300 320272 375312
rect 320324 375300 320330 375352
rect 273622 374620 273628 374672
rect 273680 374660 273686 374672
rect 273806 374660 273812 374672
rect 273680 374632 273812 374660
rect 273680 374620 273686 374632
rect 273806 374620 273812 374632
rect 273864 374620 273870 374672
rect 274450 374620 274456 374672
rect 274508 374660 274514 374672
rect 320085 374663 320143 374669
rect 320085 374660 320097 374663
rect 274508 374632 320097 374660
rect 274508 374620 274514 374632
rect 320085 374629 320097 374632
rect 320131 374660 320143 374663
rect 320821 374663 320879 374669
rect 320821 374660 320833 374663
rect 320131 374632 320833 374660
rect 320131 374629 320143 374632
rect 320085 374623 320143 374629
rect 320821 374629 320833 374632
rect 320867 374629 320879 374663
rect 320821 374623 320879 374629
rect 273530 374484 273536 374536
rect 273588 374524 273594 374536
rect 273806 374524 273812 374536
rect 273588 374496 273812 374524
rect 273588 374484 273594 374496
rect 273806 374484 273812 374496
rect 273864 374484 273870 374536
rect 320542 374416 320548 374468
rect 320600 374416 320606 374468
rect 320560 374252 320588 374416
rect 320634 374252 320640 374264
rect 320560 374224 320640 374252
rect 320634 374212 320640 374224
rect 320692 374212 320698 374264
rect 278314 373940 278320 373992
rect 278372 373980 278378 373992
rect 320174 373980 320180 373992
rect 278372 373952 320180 373980
rect 278372 373940 278378 373952
rect 320174 373940 320180 373952
rect 320232 373940 320238 373992
rect 320082 372960 320088 372972
rect 319995 372932 320088 372960
rect 320082 372920 320088 372932
rect 320140 372960 320146 372972
rect 320453 372963 320511 372969
rect 320453 372960 320465 372963
rect 320140 372932 320465 372960
rect 320140 372920 320146 372932
rect 320453 372929 320465 372932
rect 320499 372929 320511 372963
rect 320453 372923 320511 372929
rect 278222 372512 278228 372564
rect 278280 372552 278286 372564
rect 278280 372524 320404 372552
rect 278280 372512 278286 372524
rect 320376 372496 320404 372524
rect 320358 372444 320364 372496
rect 320416 372444 320422 372496
rect 274450 371832 274456 371884
rect 274508 371872 274514 371884
rect 319898 371872 319904 371884
rect 274508 371844 319904 371872
rect 274508 371832 274514 371844
rect 319898 371832 319904 371844
rect 319956 371872 319962 371884
rect 320542 371872 320548 371884
rect 319956 371844 320548 371872
rect 319956 371832 319962 371844
rect 320542 371832 320548 371844
rect 320600 371832 320606 371884
rect 320818 371600 320824 371612
rect 320779 371572 320824 371600
rect 320818 371560 320824 371572
rect 320876 371560 320882 371612
rect 278130 371152 278136 371204
rect 278188 371192 278194 371204
rect 320266 371192 320272 371204
rect 278188 371164 320272 371192
rect 278188 371152 278194 371164
rect 320266 371152 320272 371164
rect 320324 371152 320330 371204
rect 320269 371059 320327 371065
rect 320269 371025 320281 371059
rect 320315 371056 320327 371059
rect 320818 371056 320824 371068
rect 320315 371028 320824 371056
rect 320315 371025 320327 371028
rect 320269 371019 320327 371025
rect 320818 371016 320824 371028
rect 320876 371016 320882 371068
rect 274450 370472 274456 370524
rect 274508 370512 274514 370524
rect 319990 370512 319996 370524
rect 274508 370484 319996 370512
rect 274508 370472 274514 370484
rect 319990 370472 319996 370484
rect 320048 370472 320054 370524
rect 320634 370472 320640 370524
rect 320692 370472 320698 370524
rect 320818 370512 320824 370524
rect 320779 370484 320824 370512
rect 320818 370472 320824 370484
rect 320876 370472 320882 370524
rect 320652 370320 320680 370472
rect 320634 370268 320640 370320
rect 320692 370268 320698 370320
rect 280798 369792 280804 369844
rect 280856 369832 280862 369844
rect 320174 369832 320180 369844
rect 280856 369804 320180 369832
rect 280856 369792 280862 369804
rect 320174 369792 320180 369804
rect 320232 369792 320238 369844
rect 283558 369724 283564 369776
rect 283616 369764 283622 369776
rect 319806 369764 319812 369776
rect 283616 369736 319812 369764
rect 283616 369724 283622 369736
rect 319806 369724 319812 369736
rect 319864 369724 319870 369776
rect 319990 369452 319996 369504
rect 320048 369492 320054 369504
rect 320634 369492 320640 369504
rect 320048 369464 320640 369492
rect 320048 369452 320054 369464
rect 320634 369452 320640 369464
rect 320692 369452 320698 369504
rect 319898 369044 319904 369096
rect 319956 369084 319962 369096
rect 320358 369084 320364 369096
rect 319956 369056 320364 369084
rect 319956 369044 319962 369056
rect 320358 369044 320364 369056
rect 320416 369044 320422 369096
rect 320361 368611 320419 368617
rect 320361 368577 320373 368611
rect 320407 368608 320419 368611
rect 320450 368608 320456 368620
rect 320407 368580 320456 368608
rect 320407 368577 320419 368580
rect 320361 368571 320419 368577
rect 320450 368568 320456 368580
rect 320508 368568 320514 368620
rect 278038 368432 278044 368484
rect 278096 368472 278102 368484
rect 320450 368472 320456 368484
rect 278096 368444 320456 368472
rect 278096 368432 278102 368444
rect 320450 368432 320456 368444
rect 320508 368432 320514 368484
rect 320266 367860 320272 367872
rect 320227 367832 320272 367860
rect 320266 367820 320272 367832
rect 320324 367820 320330 367872
rect 298097 367047 298155 367053
rect 298097 367044 298109 367047
rect 292776 367016 298109 367044
rect 292577 366979 292635 366985
rect 292577 366945 292589 366979
rect 292623 366976 292635 366979
rect 292776 366976 292804 367016
rect 298097 367013 298109 367016
rect 298143 367013 298155 367047
rect 298097 367007 298155 367013
rect 292623 366948 292804 366976
rect 307757 366979 307815 366985
rect 292623 366945 292635 366948
rect 292577 366939 292635 366945
rect 307757 366945 307769 366979
rect 307803 366976 307815 366979
rect 317417 366979 317475 366985
rect 317417 366976 317429 366979
rect 307803 366948 317429 366976
rect 307803 366945 307815 366948
rect 307757 366939 307815 366945
rect 317417 366945 317429 366948
rect 317463 366945 317475 366979
rect 317417 366939 317475 366945
rect 284938 366868 284944 366920
rect 284996 366908 285002 366920
rect 292485 366911 292543 366917
rect 292485 366908 292497 366911
rect 284996 366880 292497 366908
rect 284996 366868 285002 366880
rect 292485 366877 292497 366880
rect 292531 366877 292543 366911
rect 292485 366871 292543 366877
rect 298097 366911 298155 366917
rect 298097 366877 298109 366911
rect 298143 366908 298155 366911
rect 298143 366880 307708 366908
rect 298143 366877 298155 366880
rect 298097 366871 298155 366877
rect 307680 366840 307708 366880
rect 307757 366843 307815 366849
rect 307757 366840 307769 366843
rect 307680 366812 307769 366840
rect 307757 366809 307769 366812
rect 307803 366809 307815 366843
rect 307757 366803 307815 366809
rect 317417 366299 317475 366305
rect 317417 366265 317429 366299
rect 317463 366296 317475 366299
rect 318794 366296 318800 366308
rect 317463 366268 318800 366296
rect 317463 366265 317475 366268
rect 317417 366259 317475 366265
rect 318794 366256 318800 366268
rect 318852 366256 318858 366308
rect 320358 365820 320364 365832
rect 320192 365792 320364 365820
rect 320192 365764 320220 365792
rect 320358 365780 320364 365792
rect 320416 365780 320422 365832
rect 320174 365712 320180 365764
rect 320232 365712 320238 365764
rect 286318 365644 286324 365696
rect 286376 365684 286382 365696
rect 320358 365684 320364 365696
rect 286376 365656 320364 365684
rect 286376 365644 286382 365656
rect 320358 365644 320364 365656
rect 320416 365644 320422 365696
rect 287698 364284 287704 364336
rect 287756 364324 287762 364336
rect 320266 364324 320272 364336
rect 287756 364296 320272 364324
rect 287756 364284 287762 364296
rect 320266 364284 320272 364296
rect 320324 364284 320330 364336
rect 319990 363740 319996 363792
rect 320048 363780 320054 363792
rect 320453 363783 320511 363789
rect 320453 363780 320465 363783
rect 320048 363752 320465 363780
rect 320048 363740 320054 363752
rect 320453 363749 320465 363752
rect 320499 363749 320511 363783
rect 320453 363743 320511 363749
rect 273714 362856 273720 362908
rect 273772 362896 273778 362908
rect 320450 362896 320456 362908
rect 273772 362868 320456 362896
rect 273772 362856 273778 362868
rect 320450 362856 320456 362868
rect 320508 362856 320514 362908
rect 290458 362788 290464 362840
rect 290516 362828 290522 362840
rect 319806 362828 319812 362840
rect 290516 362800 319812 362828
rect 290516 362788 290522 362800
rect 319806 362788 319812 362800
rect 319864 362788 319870 362840
rect 320082 362652 320088 362704
rect 320140 362692 320146 362704
rect 320361 362695 320419 362701
rect 320361 362692 320373 362695
rect 320140 362664 320373 362692
rect 320140 362652 320146 362664
rect 320361 362661 320373 362664
rect 320407 362661 320419 362695
rect 320361 362655 320419 362661
rect 273530 361020 273536 361072
rect 273588 361060 273594 361072
rect 275462 361060 275468 361072
rect 273588 361032 275468 361060
rect 273588 361020 273594 361032
rect 275462 361020 275468 361032
rect 275520 361020 275526 361072
rect 320266 360884 320272 360936
rect 320324 360924 320330 360936
rect 320726 360924 320732 360936
rect 320324 360896 320732 360924
rect 320324 360884 320330 360896
rect 320726 360884 320732 360896
rect 320784 360884 320790 360936
rect 320818 360312 320824 360324
rect 320468 360284 320824 360312
rect 320468 360256 320496 360284
rect 320818 360272 320824 360284
rect 320876 360272 320882 360324
rect 320450 360204 320456 360256
rect 320508 360204 320514 360256
rect 320266 360136 320272 360188
rect 320324 360176 320330 360188
rect 320324 360148 320369 360176
rect 320324 360136 320330 360148
rect 320266 360000 320272 360052
rect 320324 360040 320330 360052
rect 320726 360040 320732 360052
rect 320324 360012 320732 360040
rect 320324 360000 320330 360012
rect 320726 360000 320732 360012
rect 320784 360000 320790 360052
rect 320361 359907 320419 359913
rect 320361 359873 320373 359907
rect 320407 359904 320419 359907
rect 320726 359904 320732 359916
rect 320407 359876 320732 359904
rect 320407 359873 320419 359876
rect 320361 359867 320419 359873
rect 320726 359864 320732 359876
rect 320784 359864 320790 359916
rect 319990 359796 319996 359848
rect 320048 359836 320054 359848
rect 320818 359836 320824 359848
rect 320048 359808 320824 359836
rect 320048 359796 320054 359808
rect 320818 359796 320824 359808
rect 320876 359796 320882 359848
rect 273806 359660 273812 359712
rect 273864 359700 273870 359712
rect 275370 359700 275376 359712
rect 273864 359672 275376 359700
rect 273864 359660 273870 359672
rect 275370 359660 275376 359672
rect 275428 359660 275434 359712
rect 320174 356872 320180 356924
rect 320232 356912 320238 356924
rect 320358 356912 320364 356924
rect 320232 356884 320364 356912
rect 320232 356872 320238 356884
rect 320358 356872 320364 356884
rect 320416 356872 320422 356924
rect 291838 355988 291844 356040
rect 291896 356028 291902 356040
rect 320174 356028 320180 356040
rect 291896 356000 320180 356028
rect 291896 355988 291902 356000
rect 320174 355988 320180 356000
rect 320232 355988 320238 356040
rect 274358 355920 274364 355972
rect 274416 355960 274422 355972
rect 275278 355960 275284 355972
rect 274416 355932 275284 355960
rect 274416 355920 274422 355932
rect 275278 355920 275284 355932
rect 275336 355920 275342 355972
rect 320269 355895 320327 355901
rect 320269 355861 320281 355895
rect 320315 355892 320327 355895
rect 320634 355892 320640 355904
rect 320315 355864 320640 355892
rect 320315 355861 320327 355864
rect 320269 355855 320327 355861
rect 320634 355852 320640 355864
rect 320692 355852 320698 355904
rect 294598 354628 294604 354680
rect 294656 354668 294662 354680
rect 320174 354668 320180 354680
rect 294656 354640 320180 354668
rect 294656 354628 294662 354640
rect 320174 354628 320180 354640
rect 320232 354628 320238 354680
rect 273806 353404 273812 353456
rect 273864 353444 273870 353456
rect 274818 353444 274824 353456
rect 273864 353416 274824 353444
rect 273864 353404 273870 353416
rect 274818 353404 274824 353416
rect 274876 353404 274882 353456
rect 274266 353200 274272 353252
rect 274324 353240 274330 353252
rect 320174 353240 320180 353252
rect 274324 353212 320180 353240
rect 274324 353200 274330 353212
rect 320174 353200 320180 353212
rect 320232 353200 320238 353252
rect 297358 351840 297364 351892
rect 297416 351880 297422 351892
rect 320266 351880 320272 351892
rect 297416 351852 320272 351880
rect 297416 351840 297422 351852
rect 320266 351840 320272 351852
rect 320324 351840 320330 351892
rect 274174 350412 274180 350464
rect 274232 350452 274238 350464
rect 320266 350452 320272 350464
rect 274232 350424 320272 350452
rect 274232 350412 274238 350424
rect 320266 350412 320272 350424
rect 320324 350412 320330 350464
rect 273530 349596 273536 349648
rect 273588 349636 273594 349648
rect 275002 349636 275008 349648
rect 273588 349608 275008 349636
rect 273588 349596 273594 349608
rect 275002 349596 275008 349608
rect 275060 349596 275066 349648
rect 274082 349052 274088 349104
rect 274140 349092 274146 349104
rect 320174 349092 320180 349104
rect 274140 349064 320180 349092
rect 274140 349052 274146 349064
rect 320174 349052 320180 349064
rect 320232 349052 320238 349104
rect 298738 348984 298744 349036
rect 298796 349024 298802 349036
rect 320358 349024 320364 349036
rect 298796 348996 320364 349024
rect 298796 348984 298802 348996
rect 320358 348984 320364 348996
rect 320416 348984 320422 349036
rect 273530 347692 273536 347744
rect 273588 347732 273594 347744
rect 275094 347732 275100 347744
rect 273588 347704 275100 347732
rect 273588 347692 273594 347704
rect 275094 347692 275100 347704
rect 275152 347692 275158 347744
rect 301498 347692 301504 347744
rect 301556 347732 301562 347744
rect 320174 347732 320180 347744
rect 301556 347704 320180 347732
rect 301556 347692 301562 347704
rect 320174 347692 320180 347704
rect 320232 347692 320238 347744
rect 273990 346332 273996 346384
rect 274048 346372 274054 346384
rect 320174 346372 320180 346384
rect 274048 346344 320180 346372
rect 274048 346332 274054 346344
rect 320174 346332 320180 346344
rect 320232 346332 320238 346384
rect 273530 345856 273536 345908
rect 273588 345896 273594 345908
rect 275186 345896 275192 345908
rect 273588 345868 275192 345896
rect 273588 345856 273594 345868
rect 275186 345856 275192 345868
rect 275244 345856 275250 345908
rect 273622 343952 273628 344004
rect 273680 343992 273686 344004
rect 275922 343992 275928 344004
rect 273680 343964 275928 343992
rect 273680 343952 273686 343964
rect 275922 343952 275928 343964
rect 275980 343952 275986 344004
rect 273530 342116 273536 342168
rect 273588 342156 273594 342168
rect 275738 342156 275744 342168
rect 273588 342128 275744 342156
rect 273588 342116 273594 342128
rect 275738 342116 275744 342128
rect 275796 342116 275802 342168
rect 273530 340076 273536 340128
rect 273588 340116 273594 340128
rect 275830 340116 275836 340128
rect 273588 340088 275836 340116
rect 273588 340076 273594 340088
rect 275830 340076 275836 340088
rect 275888 340076 275894 340128
rect 273806 335248 273812 335300
rect 273864 335288 273870 335300
rect 302878 335288 302884 335300
rect 273864 335260 302884 335288
rect 273864 335248 273870 335260
rect 302878 335248 302884 335260
rect 302936 335248 302942 335300
rect 274266 332460 274272 332512
rect 274324 332500 274330 332512
rect 279418 332500 279424 332512
rect 274324 332472 279424 332500
rect 274324 332460 274330 332472
rect 279418 332460 279424 332472
rect 279476 332460 279482 332512
rect 273346 331304 273352 331356
rect 273404 331344 273410 331356
rect 273530 331344 273536 331356
rect 273404 331316 273536 331344
rect 273404 331304 273410 331316
rect 273530 331304 273536 331316
rect 273588 331304 273594 331356
rect 273346 331168 273352 331220
rect 273404 331208 273410 331220
rect 319438 331208 319444 331220
rect 273404 331180 319444 331208
rect 273404 331168 273410 331180
rect 319438 331168 319444 331180
rect 319496 331168 319502 331220
rect 273990 329740 273996 329792
rect 274048 329780 274054 329792
rect 316678 329780 316684 329792
rect 274048 329752 316684 329780
rect 274048 329740 274054 329752
rect 316678 329740 316684 329752
rect 316736 329740 316742 329792
rect 273530 323280 273536 323332
rect 273588 323320 273594 323332
rect 275646 323320 275652 323332
rect 273588 323292 275652 323320
rect 273588 323280 273594 323292
rect 275646 323280 275652 323292
rect 275704 323280 275710 323332
rect 273438 321240 273444 321292
rect 273496 321280 273502 321292
rect 275554 321280 275560 321292
rect 273496 321252 275560 321280
rect 273496 321240 273502 321252
rect 275554 321240 275560 321252
rect 275612 321240 275618 321292
rect 230658 320152 230664 320204
rect 230716 320192 230722 320204
rect 231486 320192 231492 320204
rect 230716 320164 231492 320192
rect 230716 320152 230722 320164
rect 231486 320152 231492 320164
rect 231544 320152 231550 320204
rect 235626 320192 235632 320204
rect 235460 320164 235632 320192
rect 235460 319932 235488 320164
rect 235626 320152 235632 320164
rect 235684 320152 235690 320204
rect 240686 320152 240692 320204
rect 240744 320192 240750 320204
rect 241330 320192 241336 320204
rect 240744 320164 241336 320192
rect 240744 320152 240750 320164
rect 241330 320152 241336 320164
rect 241388 320152 241394 320204
rect 241882 320152 241888 320204
rect 241940 320192 241946 320204
rect 242710 320192 242716 320204
rect 241940 320164 242716 320192
rect 241940 320152 241946 320164
rect 242710 320152 242716 320164
rect 242768 320152 242774 320204
rect 244274 320152 244280 320204
rect 244332 320192 244338 320204
rect 245102 320192 245108 320204
rect 244332 320164 245108 320192
rect 244332 320152 244338 320164
rect 245102 320152 245108 320164
rect 245160 320152 245166 320204
rect 245654 320152 245660 320204
rect 245712 320192 245718 320204
rect 246390 320192 246396 320204
rect 245712 320164 246396 320192
rect 245712 320152 245718 320164
rect 246390 320152 246396 320164
rect 246448 320152 246454 320204
rect 247126 320152 247132 320204
rect 247184 320192 247190 320204
rect 248046 320192 248052 320204
rect 247184 320164 248052 320192
rect 247184 320152 247190 320164
rect 248046 320152 248052 320164
rect 248104 320152 248110 320204
rect 253014 320152 253020 320204
rect 253072 320192 253078 320204
rect 253750 320192 253756 320204
rect 253072 320164 253756 320192
rect 253072 320152 253078 320164
rect 253750 320152 253756 320164
rect 253808 320152 253814 320204
rect 255958 320152 255964 320204
rect 256016 320192 256022 320204
rect 256326 320192 256332 320204
rect 256016 320164 256332 320192
rect 256016 320152 256022 320164
rect 256326 320152 256332 320164
rect 256384 320152 256390 320204
rect 260834 320152 260840 320204
rect 260892 320192 260898 320204
rect 261570 320192 261576 320204
rect 260892 320164 261576 320192
rect 260892 320152 260898 320164
rect 261570 320152 261576 320164
rect 261628 320152 261634 320204
rect 263594 320152 263600 320204
rect 263652 320192 263658 320204
rect 264054 320192 264060 320204
rect 263652 320164 264060 320192
rect 263652 320152 263658 320164
rect 264054 320152 264060 320164
rect 264112 320152 264118 320204
rect 266630 320152 266636 320204
rect 266688 320192 266694 320204
rect 267458 320192 267464 320204
rect 266688 320164 267464 320192
rect 266688 320152 266694 320164
rect 267458 320152 267464 320164
rect 267516 320152 267522 320204
rect 269114 320152 269120 320204
rect 269172 320192 269178 320204
rect 269850 320192 269856 320204
rect 269172 320164 269856 320192
rect 269172 320152 269178 320164
rect 269850 320152 269856 320164
rect 269908 320152 269914 320204
rect 235442 319880 235448 319932
rect 235500 319880 235506 319932
rect 251450 319404 251456 319456
rect 251508 319444 251514 319456
rect 251634 319444 251640 319456
rect 251508 319416 251640 319444
rect 251508 319404 251514 319416
rect 251634 319404 251640 319416
rect 251692 319404 251698 319456
rect 267366 319404 267372 319456
rect 267424 319444 267430 319456
rect 267550 319444 267556 319456
rect 267424 319416 267556 319444
rect 267424 319404 267430 319416
rect 267550 319404 267556 319416
rect 267608 319404 267614 319456
rect 271690 319404 271696 319456
rect 271748 319444 271754 319456
rect 271874 319444 271880 319456
rect 271748 319416 271880 319444
rect 271748 319404 271754 319416
rect 271874 319404 271880 319416
rect 271932 319404 271938 319456
rect 224957 318903 225015 318909
rect 224957 318869 224969 318903
rect 225003 318900 225015 318903
rect 234341 318903 234399 318909
rect 234341 318900 234353 318903
rect 225003 318872 234353 318900
rect 225003 318869 225015 318872
rect 224957 318863 225015 318869
rect 234341 318869 234353 318872
rect 234387 318869 234399 318903
rect 234341 318863 234399 318869
rect 142062 318792 142068 318844
rect 142120 318832 142126 318844
rect 142893 318835 142951 318841
rect 142893 318832 142905 318835
rect 142120 318804 142905 318832
rect 142120 318792 142126 318804
rect 142893 318801 142905 318804
rect 142939 318801 142951 318835
rect 142893 318795 142951 318801
rect 150802 318792 150808 318844
rect 150860 318832 150866 318844
rect 152829 318835 152887 318841
rect 152829 318832 152841 318835
rect 150860 318804 152841 318832
rect 150860 318792 150866 318804
rect 152829 318801 152841 318804
rect 152875 318801 152887 318835
rect 152829 318795 152887 318801
rect 200577 318835 200635 318841
rect 200577 318801 200589 318835
rect 200623 318832 200635 318835
rect 200623 318804 200896 318832
rect 200623 318801 200635 318804
rect 200577 318795 200635 318801
rect 49602 318724 49608 318776
rect 49660 318764 49666 318776
rect 87046 318764 87052 318776
rect 49660 318736 87052 318764
rect 49660 318724 49666 318736
rect 87046 318724 87052 318736
rect 87104 318724 87110 318776
rect 118418 318724 118424 318776
rect 118476 318764 118482 318776
rect 133138 318764 133144 318776
rect 118476 318736 133144 318764
rect 118476 318724 118482 318736
rect 133138 318724 133144 318736
rect 133196 318724 133202 318776
rect 135714 318724 135720 318776
rect 135772 318764 135778 318776
rect 159450 318764 159456 318776
rect 135772 318736 159456 318764
rect 135772 318724 135778 318736
rect 159450 318724 159456 318736
rect 159508 318724 159514 318776
rect 164234 318724 164240 318776
rect 164292 318724 164298 318776
rect 166994 318724 167000 318776
rect 167052 318764 167058 318776
rect 167052 318736 191236 318764
rect 167052 318724 167058 318736
rect 46842 318656 46848 318708
rect 46900 318696 46906 318708
rect 85850 318696 85856 318708
rect 46900 318668 85856 318696
rect 46900 318656 46906 318668
rect 85850 318656 85856 318668
rect 85908 318656 85914 318708
rect 126606 318656 126612 318708
rect 126664 318696 126670 318708
rect 142801 318699 142859 318705
rect 142801 318696 142813 318699
rect 126664 318668 142813 318696
rect 126664 318656 126670 318668
rect 142801 318665 142813 318668
rect 142847 318665 142859 318699
rect 142801 318659 142859 318665
rect 142893 318699 142951 318705
rect 142893 318665 142905 318699
rect 142939 318696 142951 318699
rect 145009 318699 145067 318705
rect 145009 318696 145021 318699
rect 142939 318668 145021 318696
rect 142939 318665 142951 318668
rect 142893 318659 142951 318665
rect 145009 318665 145021 318668
rect 145055 318665 145067 318699
rect 145009 318659 145067 318665
rect 145650 318656 145656 318708
rect 145708 318696 145714 318708
rect 148045 318699 148103 318705
rect 148045 318696 148057 318699
rect 145708 318668 148057 318696
rect 145708 318656 145714 318668
rect 148045 318665 148057 318668
rect 148091 318665 148103 318699
rect 148045 318659 148103 318665
rect 148134 318656 148140 318708
rect 148192 318696 148198 318708
rect 152737 318699 152795 318705
rect 152737 318696 152749 318699
rect 148192 318668 152749 318696
rect 148192 318656 148198 318668
rect 152737 318665 152749 318668
rect 152783 318665 152795 318699
rect 152737 318659 152795 318665
rect 152829 318699 152887 318705
rect 152829 318665 152841 318699
rect 152875 318696 152887 318699
rect 157245 318699 157303 318705
rect 157245 318696 157257 318699
rect 152875 318668 157257 318696
rect 152875 318665 152887 318668
rect 152829 318659 152887 318665
rect 157245 318665 157257 318668
rect 157291 318665 157303 318699
rect 157245 318659 157303 318665
rect 164142 318656 164148 318708
rect 164200 318696 164206 318708
rect 164252 318696 164280 318724
rect 164200 318668 164280 318696
rect 164200 318656 164206 318668
rect 39942 318588 39948 318640
rect 40000 318628 40006 318640
rect 83734 318628 83740 318640
rect 40000 318600 83740 318628
rect 40000 318588 40006 318600
rect 83734 318588 83740 318600
rect 83792 318588 83798 318640
rect 91002 318588 91008 318640
rect 91060 318628 91066 318640
rect 101490 318628 101496 318640
rect 91060 318600 101496 318628
rect 91060 318588 91066 318600
rect 101490 318588 101496 318600
rect 101548 318588 101554 318640
rect 117130 318588 117136 318640
rect 117188 318628 117194 318640
rect 133230 318628 133236 318640
rect 117188 318600 133236 318628
rect 117188 318588 117194 318600
rect 133230 318588 133236 318600
rect 133288 318588 133294 318640
rect 134518 318588 134524 318640
rect 134576 318628 134582 318640
rect 159358 318628 159364 318640
rect 134576 318600 159364 318628
rect 134576 318588 134582 318600
rect 159358 318588 159364 318600
rect 159416 318588 159422 318640
rect 162946 318588 162952 318640
rect 163004 318628 163010 318640
rect 164050 318628 164056 318640
rect 163004 318600 164056 318628
rect 163004 318588 163010 318600
rect 164050 318588 164056 318600
rect 164108 318588 164114 318640
rect 41322 318520 41328 318572
rect 41380 318560 41386 318572
rect 84194 318560 84200 318572
rect 41380 318532 84200 318560
rect 41380 318520 41386 318532
rect 84194 318520 84200 318532
rect 84252 318520 84258 318572
rect 93118 318520 93124 318572
rect 93176 318560 93182 318572
rect 99466 318560 99472 318572
rect 93176 318532 99472 318560
rect 93176 318520 93182 318532
rect 99466 318520 99472 318532
rect 99524 318520 99530 318572
rect 127894 318520 127900 318572
rect 127952 318560 127958 318572
rect 164878 318560 164884 318572
rect 127952 318532 164884 318560
rect 127952 318520 127958 318532
rect 164878 318520 164884 318532
rect 164936 318520 164942 318572
rect 185210 318520 185216 318572
rect 185268 318560 185274 318572
rect 191009 318563 191067 318569
rect 191009 318560 191021 318563
rect 185268 318532 191021 318560
rect 185268 318520 185274 318532
rect 191009 318529 191021 318532
rect 191055 318529 191067 318563
rect 191208 318560 191236 318736
rect 192662 318724 192668 318776
rect 192720 318764 192726 318776
rect 200761 318767 200819 318773
rect 200761 318764 200773 318767
rect 192720 318736 200773 318764
rect 192720 318724 192726 318736
rect 200761 318733 200773 318736
rect 200807 318733 200819 318767
rect 200868 318764 200896 318804
rect 224788 318804 225092 318832
rect 204901 318767 204959 318773
rect 204901 318764 204913 318767
rect 200868 318736 204913 318764
rect 200761 318727 200819 318733
rect 204901 318733 204913 318736
rect 204947 318733 204959 318767
rect 204901 318727 204959 318733
rect 204990 318724 204996 318776
rect 205048 318764 205054 318776
rect 208581 318767 208639 318773
rect 208581 318764 208593 318767
rect 205048 318736 208593 318764
rect 205048 318724 205054 318736
rect 208581 318733 208593 318736
rect 208627 318733 208639 318767
rect 208581 318727 208639 318733
rect 208670 318724 208676 318776
rect 208728 318764 208734 318776
rect 213825 318767 213883 318773
rect 213825 318764 213837 318767
rect 208728 318736 213837 318764
rect 208728 318724 208734 318736
rect 213825 318733 213837 318736
rect 213871 318733 213883 318767
rect 213825 318727 213883 318733
rect 214926 318724 214932 318776
rect 214984 318764 214990 318776
rect 220081 318767 220139 318773
rect 220081 318764 220093 318767
rect 214984 318736 220093 318764
rect 214984 318724 214990 318736
rect 220081 318733 220093 318736
rect 220127 318733 220139 318767
rect 220081 318727 220139 318733
rect 220170 318724 220176 318776
rect 220228 318764 220234 318776
rect 224788 318764 224816 318804
rect 220228 318736 224816 318764
rect 224865 318767 224923 318773
rect 220228 318724 220234 318736
rect 224865 318733 224877 318767
rect 224911 318764 224923 318767
rect 224957 318767 225015 318773
rect 224957 318764 224969 318767
rect 224911 318736 224969 318764
rect 224911 318733 224923 318736
rect 224865 318727 224923 318733
rect 224957 318733 224969 318736
rect 225003 318733 225015 318767
rect 225064 318764 225092 318804
rect 237650 318792 237656 318844
rect 237708 318832 237714 318844
rect 238018 318832 238024 318844
rect 237708 318804 238024 318832
rect 237708 318792 237714 318804
rect 238018 318792 238024 318804
rect 238076 318792 238082 318844
rect 240502 318792 240508 318844
rect 240560 318832 240566 318844
rect 240870 318832 240876 318844
rect 240560 318804 240876 318832
rect 240560 318792 240566 318804
rect 240870 318792 240876 318804
rect 240928 318792 240934 318844
rect 241606 318792 241612 318844
rect 241664 318832 241670 318844
rect 242066 318832 242072 318844
rect 241664 318804 242072 318832
rect 241664 318792 241670 318804
rect 242066 318792 242072 318804
rect 242124 318792 242130 318844
rect 245010 318792 245016 318844
rect 245068 318832 245074 318844
rect 245562 318832 245568 318844
rect 245068 318804 245568 318832
rect 245068 318792 245074 318804
rect 245562 318792 245568 318804
rect 245620 318792 245626 318844
rect 245746 318792 245752 318844
rect 245804 318832 245810 318844
rect 245838 318832 245844 318844
rect 245804 318804 245844 318832
rect 245804 318792 245810 318804
rect 245838 318792 245844 318804
rect 245896 318792 245902 318844
rect 256418 318792 256424 318844
rect 256476 318832 256482 318844
rect 256602 318832 256608 318844
rect 256476 318804 256608 318832
rect 256476 318792 256482 318804
rect 256602 318792 256608 318804
rect 256660 318792 256666 318844
rect 261570 318792 261576 318844
rect 261628 318832 261634 318844
rect 261662 318832 261668 318844
rect 261628 318804 261668 318832
rect 261628 318792 261634 318804
rect 261662 318792 261668 318804
rect 261720 318792 261726 318844
rect 269206 318792 269212 318844
rect 269264 318832 269270 318844
rect 269390 318832 269396 318844
rect 269264 318804 269396 318832
rect 269264 318792 269270 318804
rect 269390 318792 269396 318804
rect 269448 318792 269454 318844
rect 353938 318764 353944 318776
rect 225064 318736 353944 318764
rect 224957 318727 225015 318733
rect 353938 318724 353944 318736
rect 353996 318724 354002 318776
rect 197538 318656 197544 318708
rect 197596 318696 197602 318708
rect 201589 318699 201647 318705
rect 201589 318696 201601 318699
rect 197596 318668 201601 318696
rect 197596 318656 197602 318668
rect 201589 318665 201601 318668
rect 201635 318665 201647 318699
rect 201589 318659 201647 318665
rect 202138 318656 202144 318708
rect 202196 318696 202202 318708
rect 202690 318696 202696 318708
rect 202196 318668 202696 318696
rect 202196 318656 202202 318668
rect 202690 318656 202696 318668
rect 202748 318656 202754 318708
rect 214466 318656 214472 318708
rect 214524 318696 214530 318708
rect 215110 318696 215116 318708
rect 214524 318668 215116 318696
rect 214524 318656 214530 318668
rect 215110 318656 215116 318668
rect 215168 318656 215174 318708
rect 215205 318699 215263 318705
rect 215205 318665 215217 318699
rect 215251 318696 215263 318699
rect 222197 318699 222255 318705
rect 222197 318696 222209 318699
rect 215251 318668 222209 318696
rect 215251 318665 215263 318668
rect 215205 318659 215263 318665
rect 222197 318665 222209 318668
rect 222243 318665 222255 318699
rect 222197 318659 222255 318665
rect 222286 318656 222292 318708
rect 222344 318696 222350 318708
rect 356698 318696 356704 318708
rect 222344 318668 356704 318696
rect 222344 318656 222350 318668
rect 356698 318656 356704 318668
rect 356756 318656 356762 318708
rect 195054 318588 195060 318640
rect 195112 318628 195118 318640
rect 329098 318628 329104 318640
rect 195112 318600 329104 318628
rect 195112 318588 195118 318600
rect 329098 318588 329104 318600
rect 329156 318588 329162 318640
rect 201589 318563 201647 318569
rect 191208 318532 200804 318560
rect 191009 318523 191067 318529
rect 38562 318452 38568 318504
rect 38620 318492 38626 318504
rect 75089 318495 75147 318501
rect 75089 318492 75101 318495
rect 38620 318464 75101 318492
rect 38620 318452 38626 318464
rect 75089 318461 75101 318464
rect 75135 318461 75147 318495
rect 81710 318492 81716 318504
rect 75089 318455 75147 318461
rect 75196 318464 81716 318492
rect 34422 318384 34428 318436
rect 34480 318424 34486 318436
rect 75196 318424 75224 318464
rect 81710 318452 81716 318464
rect 81768 318452 81774 318504
rect 93762 318452 93768 318504
rect 93820 318492 93826 318504
rect 102318 318492 102324 318504
rect 93820 318464 102324 318492
rect 93820 318452 93826 318464
rect 102318 318452 102324 318464
rect 102376 318452 102382 318504
rect 132126 318452 132132 318504
rect 132184 318492 132190 318504
rect 132402 318492 132408 318504
rect 132184 318464 132408 318492
rect 132184 318452 132190 318464
rect 132402 318452 132408 318464
rect 132460 318452 132466 318504
rect 133506 318452 133512 318504
rect 133564 318492 133570 318504
rect 157978 318492 157984 318504
rect 133564 318464 157984 318492
rect 133564 318452 133570 318464
rect 157978 318452 157984 318464
rect 158036 318452 158042 318504
rect 161658 318452 161664 318504
rect 161716 318492 161722 318504
rect 200669 318495 200727 318501
rect 200669 318492 200681 318495
rect 161716 318464 200681 318492
rect 161716 318452 161722 318464
rect 200669 318461 200681 318464
rect 200715 318461 200727 318495
rect 200776 318492 200804 318532
rect 201589 318529 201601 318563
rect 201635 318560 201647 318563
rect 331858 318560 331864 318572
rect 201635 318532 331864 318560
rect 201635 318529 201647 318532
rect 201589 318523 201647 318529
rect 331858 318520 331864 318532
rect 331916 318520 331922 318572
rect 215938 318492 215944 318504
rect 200776 318464 215944 318492
rect 200669 318455 200727 318461
rect 215938 318452 215944 318464
rect 215996 318452 216002 318504
rect 217318 318452 217324 318504
rect 217376 318492 217382 318504
rect 219989 318495 220047 318501
rect 219989 318492 220001 318495
rect 217376 318464 220001 318492
rect 217376 318452 217382 318464
rect 219989 318461 220001 318464
rect 220035 318461 220047 318495
rect 219989 318455 220047 318461
rect 220081 318495 220139 318501
rect 220081 318461 220093 318495
rect 220127 318492 220139 318495
rect 348418 318492 348424 318504
rect 220127 318464 348424 318492
rect 220127 318461 220139 318464
rect 220081 318455 220139 318461
rect 348418 318452 348424 318464
rect 348476 318452 348482 318504
rect 34480 318396 75224 318424
rect 75273 318427 75331 318433
rect 34480 318384 34486 318396
rect 75273 318393 75285 318427
rect 75319 318424 75331 318427
rect 78858 318424 78864 318436
rect 75319 318396 78864 318424
rect 75319 318393 75331 318396
rect 75273 318387 75331 318393
rect 78858 318384 78864 318396
rect 78916 318384 78922 318436
rect 81342 318424 81348 318436
rect 78968 318396 81348 318424
rect 33042 318316 33048 318368
rect 33100 318356 33106 318368
rect 78968 318356 78996 318396
rect 81342 318384 81348 318396
rect 81400 318384 81406 318436
rect 88978 318384 88984 318436
rect 89036 318424 89042 318436
rect 98178 318424 98184 318436
rect 89036 318396 98184 318424
rect 89036 318384 89042 318396
rect 98178 318384 98184 318396
rect 98236 318384 98242 318436
rect 123754 318384 123760 318436
rect 123812 318424 123818 318436
rect 147398 318424 147404 318436
rect 123812 318396 147404 318424
rect 123812 318384 123818 318396
rect 147398 318384 147404 318396
rect 147456 318384 147462 318436
rect 147493 318427 147551 318433
rect 147493 318393 147505 318427
rect 147539 318424 147551 318427
rect 149698 318424 149704 318436
rect 147539 318396 149704 318424
rect 147539 318393 147551 318396
rect 147493 318387 147551 318393
rect 149698 318384 149704 318396
rect 149756 318384 149762 318436
rect 149790 318384 149796 318436
rect 149848 318424 149854 318436
rect 150250 318424 150256 318436
rect 149848 318396 150256 318424
rect 149848 318384 149854 318396
rect 150250 318384 150256 318396
rect 150308 318384 150314 318436
rect 150437 318427 150495 318433
rect 150437 318393 150449 318427
rect 150483 318424 150495 318427
rect 154025 318427 154083 318433
rect 154025 318424 154037 318427
rect 150483 318396 154037 318424
rect 150483 318393 150495 318396
rect 150437 318387 150495 318393
rect 154025 318393 154037 318396
rect 154071 318393 154083 318427
rect 154025 318387 154083 318393
rect 159266 318384 159272 318436
rect 159324 318424 159330 318436
rect 200577 318427 200635 318433
rect 200577 318424 200589 318427
rect 159324 318396 200589 318424
rect 159324 318384 159330 318396
rect 200577 318393 200589 318396
rect 200623 318393 200635 318427
rect 209038 318424 209044 318436
rect 200577 318387 200635 318393
rect 200776 318396 209044 318424
rect 33100 318328 78996 318356
rect 33100 318316 33106 318328
rect 91738 318316 91744 318368
rect 91796 318356 91802 318368
rect 101122 318356 101128 318368
rect 91796 318328 101128 318356
rect 91796 318316 91802 318328
rect 101122 318316 101128 318328
rect 101180 318316 101186 318368
rect 124214 318316 124220 318368
rect 124272 318356 124278 318368
rect 149241 318359 149299 318365
rect 149241 318356 149253 318359
rect 124272 318328 149253 318356
rect 124272 318316 124278 318328
rect 149241 318325 149253 318328
rect 149287 318325 149299 318359
rect 149241 318319 149299 318325
rect 149330 318316 149336 318368
rect 149388 318356 149394 318368
rect 153289 318359 153347 318365
rect 153289 318356 153301 318359
rect 149388 318328 153301 318356
rect 149388 318316 149394 318328
rect 153289 318325 153301 318328
rect 153335 318325 153347 318359
rect 153289 318319 153347 318325
rect 153838 318316 153844 318368
rect 153896 318356 153902 318368
rect 154298 318356 154304 318368
rect 153896 318328 154304 318356
rect 153896 318316 153902 318328
rect 154298 318316 154304 318328
rect 154356 318316 154362 318368
rect 160462 318316 160468 318368
rect 160520 318356 160526 318368
rect 200776 318356 200804 318396
rect 209038 318384 209044 318396
rect 209096 318384 209102 318436
rect 209958 318384 209964 318436
rect 210016 318424 210022 318436
rect 210016 318396 212396 318424
rect 210016 318384 210022 318396
rect 160520 318328 200804 318356
rect 160520 318316 160526 318328
rect 202506 318316 202512 318368
rect 202564 318356 202570 318368
rect 210421 318359 210479 318365
rect 210421 318356 210433 318359
rect 202564 318328 210433 318356
rect 202564 318316 202570 318328
rect 210421 318325 210433 318328
rect 210467 318325 210479 318359
rect 210421 318319 210479 318325
rect 210513 318359 210571 318365
rect 210513 318325 210525 318359
rect 210559 318356 210571 318359
rect 212077 318359 212135 318365
rect 212077 318356 212089 318359
rect 210559 318328 212089 318356
rect 210559 318325 210571 318328
rect 210513 318319 210571 318325
rect 212077 318325 212089 318328
rect 212123 318325 212135 318359
rect 212368 318356 212396 318396
rect 212442 318384 212448 318436
rect 212500 318424 212506 318436
rect 347038 318424 347044 318436
rect 212500 318396 347044 318424
rect 212500 318384 212506 318396
rect 347038 318384 347044 318396
rect 347096 318384 347102 318436
rect 345658 318356 345664 318368
rect 212368 318328 345664 318356
rect 212077 318319 212135 318325
rect 345658 318316 345664 318328
rect 345716 318316 345722 318368
rect 27522 318248 27528 318300
rect 27580 318288 27586 318300
rect 79226 318288 79232 318300
rect 27580 318260 79232 318288
rect 27580 318248 27586 318260
rect 79226 318248 79232 318260
rect 79284 318248 79290 318300
rect 89070 318248 89076 318300
rect 89128 318288 89134 318300
rect 99834 318288 99840 318300
rect 89128 318260 99840 318288
rect 89128 318248 89134 318260
rect 99834 318248 99840 318260
rect 99892 318248 99898 318300
rect 108942 318248 108948 318300
rect 109000 318288 109006 318300
rect 111058 318288 111064 318300
rect 109000 318260 111064 318288
rect 109000 318248 109006 318260
rect 111058 318248 111064 318260
rect 111116 318248 111122 318300
rect 120074 318248 120080 318300
rect 120132 318288 120138 318300
rect 136913 318291 136971 318297
rect 136913 318288 136925 318291
rect 120132 318260 136925 318288
rect 120132 318248 120138 318260
rect 136913 318257 136925 318260
rect 136959 318257 136971 318291
rect 136913 318251 136971 318257
rect 140682 318248 140688 318300
rect 140740 318288 140746 318300
rect 142709 318291 142767 318297
rect 142709 318288 142721 318291
rect 140740 318260 142721 318288
rect 140740 318248 140746 318260
rect 142709 318257 142721 318260
rect 142755 318257 142767 318291
rect 142709 318251 142767 318257
rect 142801 318291 142859 318297
rect 142801 318257 142813 318291
rect 142847 318288 142859 318291
rect 147493 318291 147551 318297
rect 147493 318288 147505 318291
rect 142847 318260 147505 318288
rect 142847 318257 142859 318260
rect 142801 318251 142859 318257
rect 147493 318257 147505 318260
rect 147539 318257 147551 318291
rect 152458 318288 152464 318300
rect 147493 318251 147551 318257
rect 147784 318260 152464 318288
rect 31662 318180 31668 318232
rect 31720 318220 31726 318232
rect 100294 318220 100300 318232
rect 31720 318192 78536 318220
rect 31720 318180 31726 318192
rect 26142 318112 26148 318164
rect 26200 318152 26206 318164
rect 74537 318155 74595 318161
rect 26200 318124 74488 318152
rect 26200 318112 26206 318124
rect 24762 318044 24768 318096
rect 24820 318084 24826 318096
rect 74353 318087 74411 318093
rect 74353 318084 74365 318087
rect 24820 318056 74365 318084
rect 24820 318044 24826 318056
rect 74353 318053 74365 318056
rect 74399 318053 74411 318087
rect 74460 318084 74488 318124
rect 74537 318121 74549 318155
rect 74583 318152 74595 318155
rect 78398 318152 78404 318164
rect 74583 318124 78404 318152
rect 74583 318121 74595 318124
rect 74537 318115 74595 318121
rect 78398 318112 78404 318124
rect 78456 318112 78462 318164
rect 78508 318152 78536 318192
rect 94516 318192 100300 318220
rect 80882 318152 80888 318164
rect 78508 318124 80888 318152
rect 80882 318112 80888 318124
rect 80940 318112 80946 318164
rect 88242 318112 88248 318164
rect 88300 318152 88306 318164
rect 94516 318152 94544 318192
rect 100294 318180 100300 318192
rect 100352 318180 100358 318232
rect 113082 318180 113088 318232
rect 113140 318220 113146 318232
rect 123478 318220 123484 318232
rect 113140 318192 123484 318220
rect 113140 318180 113146 318192
rect 123478 318180 123484 318192
rect 123536 318180 123542 318232
rect 128262 318180 128268 318232
rect 128320 318220 128326 318232
rect 147677 318223 147735 318229
rect 147677 318220 147689 318223
rect 128320 318192 147689 318220
rect 128320 318180 128326 318192
rect 147677 318189 147689 318192
rect 147723 318189 147735 318223
rect 147677 318183 147735 318189
rect 88300 318124 94544 318152
rect 88300 318112 88306 318124
rect 97258 318112 97264 318164
rect 97316 318152 97322 318164
rect 100662 318152 100668 318164
rect 97316 318124 100668 318152
rect 97316 318112 97322 318124
rect 100662 318112 100668 318124
rect 100720 318112 100726 318164
rect 110138 318112 110144 318164
rect 110196 318152 110202 318164
rect 111150 318152 111156 318164
rect 110196 318124 111156 318152
rect 110196 318112 110202 318124
rect 111150 318112 111156 318124
rect 111208 318112 111214 318164
rect 112254 318112 112260 318164
rect 112312 318152 112318 318164
rect 116578 318152 116584 318164
rect 112312 318124 116584 318152
rect 112312 318112 112318 318124
rect 116578 318112 116584 318124
rect 116636 318112 116642 318164
rect 121270 318112 121276 318164
rect 121328 318152 121334 318164
rect 138385 318155 138443 318161
rect 121328 318124 138336 318152
rect 121328 318112 121334 318124
rect 74997 318087 75055 318093
rect 74997 318084 75009 318087
rect 74460 318056 75009 318084
rect 74353 318047 74411 318053
rect 74997 318053 75009 318056
rect 75043 318053 75055 318087
rect 74997 318047 75055 318053
rect 75089 318087 75147 318093
rect 75089 318053 75101 318087
rect 75135 318084 75147 318087
rect 83366 318084 83372 318096
rect 75135 318056 83372 318084
rect 75135 318053 75147 318056
rect 75089 318047 75147 318053
rect 83366 318044 83372 318056
rect 83424 318044 83430 318096
rect 86218 318084 86224 318096
rect 83476 318056 86224 318084
rect 48130 317976 48136 318028
rect 48188 318016 48194 318028
rect 83476 318016 83504 318056
rect 86218 318044 86224 318056
rect 86276 318044 86282 318096
rect 111794 318044 111800 318096
rect 111852 318084 111858 318096
rect 111852 318056 113404 318084
rect 111852 318044 111858 318056
rect 48188 317988 83504 318016
rect 84657 318019 84715 318025
rect 48188 317976 48194 317988
rect 84657 317985 84669 318019
rect 84703 318016 84715 318019
rect 92842 318016 92848 318028
rect 84703 317988 92848 318016
rect 84703 317985 84715 317988
rect 84657 317979 84715 317985
rect 92842 317976 92848 317988
rect 92900 317976 92906 318028
rect 110966 317976 110972 318028
rect 111024 318016 111030 318028
rect 111702 318016 111708 318028
rect 111024 317988 111708 318016
rect 111024 317976 111030 317988
rect 111702 317976 111708 317988
rect 111760 317976 111766 318028
rect 112622 317976 112628 318028
rect 112680 318016 112686 318028
rect 113082 318016 113088 318028
rect 112680 317988 113088 318016
rect 112680 317976 112686 317988
rect 113082 317976 113088 317988
rect 113140 317976 113146 318028
rect 50982 317908 50988 317960
rect 51040 317948 51046 317960
rect 87506 317948 87512 317960
rect 51040 317920 87512 317948
rect 51040 317908 51046 317920
rect 87506 317908 87512 317920
rect 87564 317908 87570 317960
rect 109310 317908 109316 317960
rect 109368 317948 109374 317960
rect 110230 317948 110236 317960
rect 109368 317920 110236 317948
rect 109368 317908 109374 317920
rect 110230 317908 110236 317920
rect 110288 317908 110294 317960
rect 113376 317948 113404 318056
rect 113910 318044 113916 318096
rect 113968 318084 113974 318096
rect 114370 318084 114376 318096
rect 113968 318056 114376 318084
rect 113968 318044 113974 318056
rect 114370 318044 114376 318056
rect 114428 318044 114434 318096
rect 114738 318044 114744 318096
rect 114796 318084 114802 318096
rect 115658 318084 115664 318096
rect 114796 318056 115664 318084
rect 114796 318044 114802 318056
rect 115658 318044 115664 318056
rect 115716 318044 115722 318096
rect 116302 318044 116308 318096
rect 116360 318084 116366 318096
rect 117222 318084 117228 318096
rect 116360 318056 117228 318084
rect 116360 318044 116366 318056
rect 117222 318044 117228 318056
rect 117280 318044 117286 318096
rect 119246 318044 119252 318096
rect 119304 318084 119310 318096
rect 119890 318084 119896 318096
rect 119304 318056 119896 318084
rect 119304 318044 119310 318056
rect 119890 318044 119896 318056
rect 119948 318044 119954 318096
rect 121730 318044 121736 318096
rect 121788 318084 121794 318096
rect 122558 318084 122564 318096
rect 121788 318056 122564 318084
rect 121788 318044 121794 318056
rect 122558 318044 122564 318056
rect 122616 318044 122622 318096
rect 138308 318084 138336 318124
rect 138385 318121 138397 318155
rect 138431 318152 138443 318155
rect 147784 318152 147812 318260
rect 152458 318248 152464 318260
rect 152516 318248 152522 318300
rect 152737 318291 152795 318297
rect 152737 318257 152749 318291
rect 152783 318288 152795 318291
rect 190089 318291 190147 318297
rect 190089 318288 190101 318291
rect 152783 318260 190101 318288
rect 152783 318257 152795 318260
rect 152737 318251 152795 318257
rect 190089 318257 190101 318260
rect 190135 318257 190147 318291
rect 190089 318251 190147 318257
rect 191009 318291 191067 318297
rect 191009 318257 191021 318291
rect 191055 318288 191067 318291
rect 195885 318291 195943 318297
rect 195885 318288 195897 318291
rect 191055 318260 195897 318288
rect 191055 318257 191067 318260
rect 191009 318251 191067 318257
rect 195885 318257 195897 318260
rect 195931 318257 195943 318291
rect 195885 318251 195943 318257
rect 200022 318248 200028 318300
rect 200080 318288 200086 318300
rect 335998 318288 336004 318300
rect 200080 318260 336004 318288
rect 200080 318248 200086 318260
rect 335998 318248 336004 318260
rect 336056 318248 336062 318300
rect 148045 318223 148103 318229
rect 148045 318189 148057 318223
rect 148091 318220 148103 318223
rect 150437 318223 150495 318229
rect 150437 318220 150449 318223
rect 148091 318192 150449 318220
rect 148091 318189 148103 318192
rect 148045 318183 148103 318189
rect 150437 318189 150449 318192
rect 150483 318189 150495 318223
rect 150437 318183 150495 318189
rect 163958 318180 163964 318232
rect 164016 318220 164022 318232
rect 218698 318220 218704 318232
rect 164016 318192 218704 318220
rect 164016 318180 164022 318192
rect 218698 318180 218704 318192
rect 218756 318180 218762 318232
rect 219989 318223 220047 318229
rect 219989 318189 220001 318223
rect 220035 318220 220047 318223
rect 224681 318223 224739 318229
rect 224681 318220 224693 318223
rect 220035 318192 224693 318220
rect 220035 318189 220047 318192
rect 219989 318183 220047 318189
rect 224681 318189 224693 318192
rect 224727 318189 224739 318223
rect 224681 318183 224739 318189
rect 224770 318180 224776 318232
rect 224828 318220 224834 318232
rect 360838 318220 360844 318232
rect 224828 318192 360844 318220
rect 224828 318180 224834 318192
rect 360838 318180 360844 318192
rect 360896 318180 360902 318232
rect 138431 318124 147812 318152
rect 138431 318121 138443 318124
rect 138385 318115 138443 318121
rect 147858 318112 147864 318164
rect 147916 318152 147922 318164
rect 150894 318152 150900 318164
rect 147916 318124 150900 318152
rect 147916 318112 147922 318124
rect 150894 318112 150900 318124
rect 150952 318112 150958 318164
rect 151725 318155 151783 318161
rect 151725 318121 151737 318155
rect 151771 318152 151783 318155
rect 156598 318152 156604 318164
rect 151771 318124 156604 318152
rect 151771 318121 151783 318124
rect 151725 318115 151783 318121
rect 156598 318112 156604 318124
rect 156656 318112 156662 318164
rect 157245 318155 157303 318161
rect 157245 318121 157257 318155
rect 157291 318152 157303 318155
rect 200669 318155 200727 318161
rect 157291 318124 199056 318152
rect 157291 318121 157303 318124
rect 157245 318115 157303 318121
rect 145650 318084 145656 318096
rect 122668 318056 138244 318084
rect 138308 318056 145656 318084
rect 113450 317976 113456 318028
rect 113508 318016 113514 318028
rect 114462 318016 114468 318028
rect 113508 317988 114468 318016
rect 113508 317976 113514 317988
rect 114462 317976 114468 317988
rect 114520 317976 114526 318028
rect 115934 317976 115940 318028
rect 115992 318016 115998 318028
rect 117130 318016 117136 318028
rect 115992 317988 117136 318016
rect 115992 317976 115998 317988
rect 117130 317976 117136 317988
rect 117188 317976 117194 318028
rect 118786 317976 118792 318028
rect 118844 318016 118850 318028
rect 119982 318016 119988 318028
rect 118844 317988 119988 318016
rect 118844 317976 118850 317988
rect 119982 317976 119988 317988
rect 120040 317976 120046 318028
rect 120902 317976 120908 318028
rect 120960 318016 120966 318028
rect 122668 318016 122696 318056
rect 120960 317988 122696 318016
rect 122760 317988 132816 318016
rect 120960 317976 120966 317988
rect 120258 317948 120264 317960
rect 113376 317920 120264 317948
rect 120258 317908 120264 317920
rect 120316 317908 120322 317960
rect 122760 317948 122788 317988
rect 122668 317920 122788 317948
rect 56410 317840 56416 317892
rect 56468 317880 56474 317892
rect 89530 317880 89536 317892
rect 56468 317852 89536 317880
rect 56468 317840 56474 317852
rect 89530 317840 89536 317852
rect 89588 317840 89594 317892
rect 96522 317840 96528 317892
rect 96580 317880 96586 317892
rect 103146 317880 103152 317892
rect 96580 317852 103152 317880
rect 96580 317840 96586 317852
rect 103146 317840 103152 317852
rect 103204 317840 103210 317892
rect 115106 317840 115112 317892
rect 115164 317880 115170 317892
rect 115842 317880 115848 317892
rect 115164 317852 115848 317880
rect 115164 317840 115170 317852
rect 115842 317840 115848 317852
rect 115900 317840 115906 317892
rect 119614 317840 119620 317892
rect 119672 317880 119678 317892
rect 122668 317880 122696 317920
rect 122926 317908 122932 317960
rect 122984 317948 122990 317960
rect 124122 317948 124128 317960
rect 122984 317920 124128 317948
rect 122984 317908 122990 317920
rect 124122 317908 124128 317920
rect 124180 317908 124186 317960
rect 124582 317908 124588 317960
rect 124640 317948 124646 317960
rect 125502 317948 125508 317960
rect 124640 317920 125508 317948
rect 124640 317908 124646 317920
rect 125502 317908 125508 317920
rect 125560 317908 125566 317960
rect 126238 317908 126244 317960
rect 126296 317948 126302 317960
rect 126882 317948 126888 317960
rect 126296 317920 126888 317948
rect 126296 317908 126302 317920
rect 126882 317908 126888 317920
rect 126940 317908 126946 317960
rect 127434 317908 127440 317960
rect 127492 317948 127498 317960
rect 128262 317948 128268 317960
rect 127492 317920 128268 317948
rect 127492 317908 127498 317920
rect 128262 317908 128268 317920
rect 128320 317908 128326 317960
rect 128722 317908 128728 317960
rect 128780 317948 128786 317960
rect 129642 317948 129648 317960
rect 128780 317920 129648 317948
rect 128780 317908 128786 317920
rect 129642 317908 129648 317920
rect 129700 317908 129706 317960
rect 129918 317908 129924 317960
rect 129976 317948 129982 317960
rect 131022 317948 131028 317960
rect 129976 317920 131028 317948
rect 129976 317908 129982 317920
rect 131022 317908 131028 317920
rect 131080 317908 131086 317960
rect 132788 317948 132816 317988
rect 132862 317976 132868 318028
rect 132920 318016 132926 318028
rect 133782 318016 133788 318028
rect 132920 317988 133788 318016
rect 132920 317976 132926 317988
rect 133782 317976 133788 317988
rect 133840 317976 133846 318028
rect 135346 317976 135352 318028
rect 135404 318016 135410 318028
rect 136542 318016 136548 318028
rect 135404 317988 136548 318016
rect 135404 317976 135410 317988
rect 136542 317976 136548 317988
rect 136600 317976 136606 318028
rect 137002 317976 137008 318028
rect 137060 318016 137066 318028
rect 137922 318016 137928 318028
rect 137060 317988 137928 318016
rect 137060 317976 137066 317988
rect 137922 317976 137928 317988
rect 137980 317976 137986 318028
rect 138216 318016 138244 318056
rect 145650 318044 145656 318056
rect 145708 318044 145714 318096
rect 146846 318044 146852 318096
rect 146904 318084 146910 318096
rect 152461 318087 152519 318093
rect 152461 318084 152473 318087
rect 146904 318056 152473 318084
rect 146904 318044 146910 318056
rect 152461 318053 152473 318056
rect 152507 318053 152519 318087
rect 152461 318047 152519 318053
rect 153289 318087 153347 318093
rect 153289 318053 153301 318087
rect 153335 318084 153347 318087
rect 189997 318087 190055 318093
rect 153335 318056 187648 318084
rect 153335 318053 153347 318056
rect 153289 318047 153347 318053
rect 146570 318016 146576 318028
rect 138216 317988 146576 318016
rect 146570 317976 146576 317988
rect 146628 317976 146634 318028
rect 162121 318019 162179 318025
rect 162121 318016 162133 318019
rect 146680 317988 162133 318016
rect 134518 317948 134524 317960
rect 131132 317920 132724 317948
rect 132788 317920 134524 317948
rect 119672 317852 122696 317880
rect 119672 317840 119678 317852
rect 125870 317840 125876 317892
rect 125928 317880 125934 317892
rect 131132 317880 131160 317920
rect 125928 317852 131160 317880
rect 125928 317840 125934 317852
rect 131206 317840 131212 317892
rect 131264 317880 131270 317892
rect 132402 317880 132408 317892
rect 131264 317852 132408 317880
rect 131264 317840 131270 317852
rect 132402 317840 132408 317852
rect 132460 317840 132466 317892
rect 57882 317772 57888 317824
rect 57940 317812 57946 317824
rect 57940 317784 84884 317812
rect 57940 317772 57946 317784
rect 64782 317704 64788 317756
rect 64840 317744 64846 317756
rect 84749 317747 84807 317753
rect 84749 317744 84761 317747
rect 64840 317716 84761 317744
rect 64840 317704 64846 317716
rect 84749 317713 84761 317716
rect 84795 317713 84807 317747
rect 84856 317744 84884 317784
rect 84930 317772 84936 317824
rect 84988 317812 84994 317824
rect 84988 317784 92152 317812
rect 84988 317772 84994 317784
rect 89990 317744 89996 317756
rect 84856 317716 89996 317744
rect 84749 317707 84807 317713
rect 89990 317704 89996 317716
rect 90048 317704 90054 317756
rect 92124 317744 92152 317784
rect 96338 317772 96344 317824
rect 96396 317812 96402 317824
rect 102778 317812 102784 317824
rect 96396 317784 102784 317812
rect 96396 317772 96402 317784
rect 102778 317772 102784 317784
rect 102836 317772 102842 317824
rect 122098 317772 122104 317824
rect 122156 317812 122162 317824
rect 122742 317812 122748 317824
rect 122156 317784 122748 317812
rect 122156 317772 122162 317784
rect 122742 317772 122748 317784
rect 122800 317772 122806 317824
rect 129090 317772 129096 317824
rect 129148 317812 129154 317824
rect 129458 317812 129464 317824
rect 129148 317784 129464 317812
rect 129148 317772 129154 317784
rect 129458 317772 129464 317784
rect 129516 317772 129522 317824
rect 130378 317772 130384 317824
rect 130436 317812 130442 317824
rect 130838 317812 130844 317824
rect 130436 317784 130844 317812
rect 130436 317772 130442 317784
rect 130838 317772 130844 317784
rect 130896 317772 130902 317824
rect 131574 317772 131580 317824
rect 131632 317812 131638 317824
rect 132218 317812 132224 317824
rect 131632 317784 132224 317812
rect 131632 317772 131638 317784
rect 132218 317772 132224 317784
rect 132276 317772 132282 317824
rect 98638 317744 98644 317756
rect 92124 317716 98644 317744
rect 98638 317704 98644 317716
rect 98696 317704 98702 317756
rect 123386 317704 123392 317756
rect 123444 317744 123450 317756
rect 124030 317744 124036 317756
rect 123444 317716 124036 317744
rect 123444 317704 123450 317716
rect 124030 317704 124036 317716
rect 124088 317704 124094 317756
rect 127066 317704 127072 317756
rect 127124 317744 127130 317756
rect 128170 317744 128176 317756
rect 127124 317716 128176 317744
rect 127124 317704 127130 317716
rect 128170 317704 128176 317716
rect 128228 317704 128234 317756
rect 63402 317636 63408 317688
rect 63460 317676 63466 317688
rect 91646 317676 91652 317688
rect 63460 317648 91652 317676
rect 63460 317636 63466 317648
rect 91646 317636 91652 317648
rect 91704 317636 91710 317688
rect 97902 317636 97908 317688
rect 97960 317676 97966 317688
rect 103606 317676 103612 317688
rect 97960 317648 103612 317676
rect 97960 317636 97966 317648
rect 103606 317636 103612 317648
rect 103664 317636 103670 317688
rect 132126 317636 132132 317688
rect 132184 317676 132190 317688
rect 132696 317676 132724 317920
rect 134518 317908 134524 317920
rect 134576 317908 134582 317960
rect 136913 317951 136971 317957
rect 136913 317917 136925 317951
rect 136959 317948 136971 317951
rect 141418 317948 141424 317960
rect 136959 317920 141424 317948
rect 136959 317917 136971 317920
rect 136913 317911 136971 317917
rect 141418 317908 141424 317920
rect 141476 317908 141482 317960
rect 142709 317951 142767 317957
rect 142709 317917 142721 317951
rect 142755 317948 142767 317951
rect 146680 317948 146708 317988
rect 162121 317985 162133 317988
rect 162167 317985 162179 318019
rect 162121 317979 162179 317985
rect 142755 317920 146708 317948
rect 146757 317951 146815 317957
rect 142755 317917 142767 317920
rect 142709 317911 142767 317917
rect 146757 317917 146769 317951
rect 146803 317948 146815 317951
rect 151817 317951 151875 317957
rect 151817 317948 151829 317951
rect 146803 317920 151829 317948
rect 146803 317917 146815 317920
rect 146757 317911 146815 317917
rect 151817 317917 151829 317920
rect 151863 317917 151875 317951
rect 153838 317948 153844 317960
rect 151817 317911 151875 317917
rect 151924 317920 153844 317948
rect 136174 317840 136180 317892
rect 136232 317880 136238 317892
rect 141973 317883 142031 317889
rect 141973 317880 141985 317883
rect 136232 317852 141985 317880
rect 136232 317840 136238 317852
rect 141973 317849 141985 317852
rect 142019 317849 142031 317883
rect 141973 317843 142031 317849
rect 142801 317883 142859 317889
rect 142801 317849 142813 317883
rect 142847 317880 142859 317883
rect 147309 317883 147367 317889
rect 147309 317880 147321 317883
rect 142847 317852 147321 317880
rect 142847 317849 142859 317852
rect 142801 317843 142859 317849
rect 147309 317849 147321 317852
rect 147355 317849 147367 317883
rect 151924 317880 151952 317920
rect 153838 317908 153844 317920
rect 153896 317908 153902 317960
rect 147309 317843 147367 317849
rect 151096 317852 151952 317880
rect 152461 317883 152519 317889
rect 134058 317772 134064 317824
rect 134116 317812 134122 317824
rect 135162 317812 135168 317824
rect 134116 317784 135168 317812
rect 134116 317772 134122 317784
rect 135162 317772 135168 317784
rect 135220 317772 135226 317824
rect 137370 317772 137376 317824
rect 137428 317812 137434 317824
rect 138385 317815 138443 317821
rect 138385 317812 138397 317815
rect 137428 317784 138397 317812
rect 137428 317772 137434 317784
rect 138385 317781 138397 317784
rect 138431 317781 138443 317815
rect 138385 317775 138443 317781
rect 138477 317815 138535 317821
rect 138477 317781 138489 317815
rect 138523 317812 138535 317815
rect 148318 317812 148324 317824
rect 138523 317784 148324 317812
rect 138523 317781 138535 317784
rect 138477 317775 138535 317781
rect 148318 317772 148324 317784
rect 148376 317772 148382 317824
rect 148413 317815 148471 317821
rect 148413 317781 148425 317815
rect 148459 317812 148471 317815
rect 149241 317815 149299 317821
rect 148459 317784 148916 317812
rect 148459 317781 148471 317784
rect 148413 317775 148471 317781
rect 134886 317704 134892 317756
rect 134944 317744 134950 317756
rect 142801 317747 142859 317753
rect 142801 317744 142813 317747
rect 134944 317716 142813 317744
rect 134944 317704 134950 317716
rect 142801 317713 142813 317716
rect 142847 317713 142859 317747
rect 142801 317707 142859 317713
rect 142893 317747 142951 317753
rect 142893 317713 142905 317747
rect 142939 317744 142951 317747
rect 145558 317744 145564 317756
rect 142939 317716 145564 317744
rect 142939 317713 142951 317716
rect 142893 317707 142951 317713
rect 145558 317704 145564 317716
rect 145616 317704 145622 317756
rect 145653 317747 145711 317753
rect 145653 317713 145665 317747
rect 145699 317744 145711 317747
rect 146757 317747 146815 317753
rect 146757 317744 146769 317747
rect 145699 317716 146769 317744
rect 145699 317713 145711 317716
rect 145653 317707 145711 317713
rect 146757 317713 146769 317716
rect 146803 317713 146815 317747
rect 146757 317707 146815 317713
rect 147674 317704 147680 317756
rect 147732 317744 147738 317756
rect 148778 317744 148784 317756
rect 147732 317716 148784 317744
rect 147732 317704 147738 317716
rect 148778 317704 148784 317716
rect 148836 317704 148842 317756
rect 148888 317744 148916 317784
rect 149241 317781 149253 317815
rect 149287 317812 149299 317815
rect 151096 317812 151124 317852
rect 152461 317849 152473 317883
rect 152507 317880 152519 317883
rect 167638 317880 167644 317892
rect 152507 317852 167644 317880
rect 152507 317849 152519 317852
rect 152461 317843 152519 317849
rect 167638 317840 167644 317852
rect 167696 317840 167702 317892
rect 187620 317880 187648 318056
rect 189997 318053 190009 318087
rect 190043 318084 190055 318087
rect 198921 318087 198979 318093
rect 198921 318084 198933 318087
rect 190043 318056 198933 318084
rect 190043 318053 190055 318056
rect 189997 318047 190055 318053
rect 198921 318053 198933 318056
rect 198967 318053 198979 318087
rect 198921 318047 198979 318053
rect 199028 318016 199056 318124
rect 200669 318121 200681 318155
rect 200715 318152 200727 318155
rect 211982 318152 211988 318164
rect 200715 318124 211988 318152
rect 200715 318121 200727 318124
rect 200669 318115 200727 318121
rect 211982 318112 211988 318124
rect 212040 318112 212046 318164
rect 212077 318155 212135 318161
rect 212077 318121 212089 318155
rect 212123 318152 212135 318155
rect 215205 318155 215263 318161
rect 215205 318152 215217 318155
rect 212123 318124 215217 318152
rect 212123 318121 212135 318124
rect 212077 318115 212135 318121
rect 215205 318121 215217 318124
rect 215251 318121 215263 318155
rect 215205 318115 215263 318121
rect 215294 318112 215300 318164
rect 215352 318152 215358 318164
rect 216490 318152 216496 318164
rect 215352 318124 216496 318152
rect 215352 318112 215358 318124
rect 216490 318112 216496 318124
rect 216548 318112 216554 318164
rect 218606 318112 218612 318164
rect 218664 318152 218670 318164
rect 219342 318152 219348 318164
rect 218664 318124 219348 318152
rect 218664 318112 218670 318124
rect 219342 318112 219348 318124
rect 219400 318112 219406 318164
rect 220262 318112 220268 318164
rect 220320 318152 220326 318164
rect 220722 318152 220728 318164
rect 220320 318124 220728 318152
rect 220320 318112 220326 318124
rect 220722 318112 220728 318124
rect 220780 318112 220786 318164
rect 221090 318112 221096 318164
rect 221148 318152 221154 318164
rect 222102 318152 222108 318164
rect 221148 318124 222108 318152
rect 221148 318112 221154 318124
rect 222102 318112 222108 318124
rect 222160 318112 222166 318164
rect 222197 318155 222255 318161
rect 222197 318121 222209 318155
rect 222243 318152 222255 318155
rect 342898 318152 342904 318164
rect 222243 318124 342904 318152
rect 222243 318121 222255 318124
rect 222197 318115 222255 318121
rect 342898 318112 342904 318124
rect 342956 318112 342962 318164
rect 199105 318087 199163 318093
rect 199105 318053 199117 318087
rect 199151 318084 199163 318087
rect 204165 318087 204223 318093
rect 204165 318084 204177 318087
rect 199151 318056 204177 318084
rect 199151 318053 199163 318056
rect 199105 318047 199163 318053
rect 204165 318053 204177 318056
rect 204211 318053 204223 318087
rect 204165 318047 204223 318053
rect 207842 318044 207848 318096
rect 207900 318084 207906 318096
rect 208302 318084 208308 318096
rect 207900 318056 208308 318084
rect 207900 318044 207906 318056
rect 208302 318044 208308 318056
rect 208360 318044 208366 318096
rect 210421 318087 210479 318093
rect 210421 318053 210433 318087
rect 210467 318084 210479 318087
rect 340138 318084 340144 318096
rect 210467 318056 340144 318084
rect 210467 318053 210479 318056
rect 210421 318047 210479 318053
rect 340138 318044 340144 318056
rect 340196 318044 340202 318096
rect 202138 318016 202144 318028
rect 199028 317988 202144 318016
rect 202138 317976 202144 317988
rect 202196 317976 202202 318028
rect 203334 317976 203340 318028
rect 203392 318016 203398 318028
rect 203886 318016 203892 318028
rect 203392 317988 203892 318016
rect 203392 317976 203398 317988
rect 203886 317976 203892 317988
rect 203944 317976 203950 318028
rect 206186 317976 206192 318028
rect 206244 318016 206250 318028
rect 206646 318016 206652 318028
rect 206244 317988 206652 318016
rect 206244 317976 206250 317988
rect 206646 317976 206652 317988
rect 206704 317976 206710 318028
rect 207474 317976 207480 318028
rect 207532 318016 207538 318028
rect 208210 318016 208216 318028
rect 207532 317988 208216 318016
rect 207532 317976 207538 317988
rect 208210 317976 208216 317988
rect 208268 317976 208274 318028
rect 208581 318019 208639 318025
rect 208581 317985 208593 318019
rect 208627 318016 208639 318019
rect 210513 318019 210571 318025
rect 210513 318016 210525 318019
rect 208627 317988 210525 318016
rect 208627 317985 208639 317988
rect 208581 317979 208639 317985
rect 210513 317985 210525 317988
rect 210559 317985 210571 318019
rect 210513 317979 210571 317985
rect 211614 317976 211620 318028
rect 211672 318016 211678 318028
rect 212442 318016 212448 318028
rect 211672 317988 212448 318016
rect 211672 317976 211678 317988
rect 212442 317976 212448 317988
rect 212500 317976 212506 318028
rect 213270 317976 213276 318028
rect 213328 318016 213334 318028
rect 213638 318016 213644 318028
rect 213328 317988 213644 318016
rect 213328 317976 213334 317988
rect 213638 317976 213644 317988
rect 213696 317976 213702 318028
rect 214098 317976 214104 318028
rect 214156 318016 214162 318028
rect 215202 318016 215208 318028
rect 214156 317988 215208 318016
rect 214156 317976 214162 317988
rect 215202 317976 215208 317988
rect 215260 317976 215266 318028
rect 215754 317976 215760 318028
rect 215812 318016 215818 318028
rect 216398 318016 216404 318028
rect 215812 317988 216404 318016
rect 215812 317976 215818 317988
rect 216398 317976 216404 317988
rect 216456 317976 216462 318028
rect 216950 317976 216956 318028
rect 217008 318016 217014 318028
rect 217870 318016 217876 318028
rect 217008 317988 217876 318016
rect 217008 317976 217014 317988
rect 217870 317976 217876 317988
rect 217928 317976 217934 318028
rect 218146 317976 218152 318028
rect 218204 318016 218210 318028
rect 219158 318016 219164 318028
rect 218204 317988 219164 318016
rect 218204 317976 218210 317988
rect 219158 317976 219164 317988
rect 219216 317976 219222 318028
rect 219434 317976 219440 318028
rect 219492 318016 219498 318028
rect 220538 318016 220544 318028
rect 219492 317988 220544 318016
rect 219492 317976 219498 317988
rect 220538 317976 220544 317988
rect 220596 317976 220602 318028
rect 221458 317976 221464 318028
rect 221516 318016 221522 318028
rect 222010 318016 222016 318028
rect 221516 317988 222016 318016
rect 221516 317976 221522 317988
rect 222010 317976 222016 317988
rect 222068 317976 222074 318028
rect 222746 317976 222752 318028
rect 222804 318016 222810 318028
rect 223482 318016 223488 318028
rect 222804 317988 223488 318016
rect 222804 317976 222810 317988
rect 223482 317976 223488 317988
rect 223540 317976 223546 318028
rect 223942 317976 223948 318028
rect 224000 318016 224006 318028
rect 224770 318016 224776 318028
rect 224000 317988 224776 318016
rect 224000 317976 224006 317988
rect 224770 317976 224776 317988
rect 224828 317976 224834 318028
rect 226426 317976 226432 318028
rect 226484 318016 226490 318028
rect 227622 318016 227628 318028
rect 226484 317988 227628 318016
rect 226484 317976 226490 317988
rect 227622 317976 227628 317988
rect 227680 317976 227686 318028
rect 228082 317976 228088 318028
rect 228140 318016 228146 318028
rect 228818 318016 228824 318028
rect 228140 317988 228824 318016
rect 228140 317976 228146 317988
rect 228818 317976 228824 317988
rect 228876 317976 228882 318028
rect 229278 317976 229284 318028
rect 229336 318016 229342 318028
rect 230290 318016 230296 318028
rect 229336 317988 230296 318016
rect 229336 317976 229342 317988
rect 230290 317976 230296 317988
rect 230348 317976 230354 318028
rect 231854 317976 231860 318028
rect 231912 318016 231918 318028
rect 233050 318016 233056 318028
rect 231912 317988 233056 318016
rect 231912 317976 231918 317988
rect 233050 317976 233056 317988
rect 233108 317976 233114 318028
rect 233326 317976 233332 318028
rect 233384 318016 233390 318028
rect 234246 318016 234252 318028
rect 233384 317988 234252 318016
rect 233384 317976 233390 317988
rect 234246 317976 234252 317988
rect 234304 317976 234310 318028
rect 234341 318019 234399 318025
rect 234341 317985 234353 318019
rect 234387 318016 234399 318019
rect 349798 318016 349804 318028
rect 234387 317988 349804 318016
rect 234387 317985 234399 317988
rect 234341 317979 234399 317985
rect 349798 317976 349804 317988
rect 349856 317976 349862 318028
rect 190178 317908 190184 317960
rect 190236 317948 190242 317960
rect 322198 317948 322204 317960
rect 190236 317920 322204 317948
rect 190236 317908 190242 317920
rect 322198 317908 322204 317920
rect 322256 317908 322262 317960
rect 198001 317883 198059 317889
rect 198001 317880 198013 317883
rect 187620 317852 198013 317880
rect 198001 317849 198013 317852
rect 198047 317849 198059 317883
rect 198001 317843 198059 317849
rect 200761 317883 200819 317889
rect 200761 317849 200773 317883
rect 200807 317880 200819 317883
rect 325050 317880 325056 317892
rect 200807 317852 325056 317880
rect 200807 317849 200819 317852
rect 200761 317843 200819 317849
rect 325050 317840 325056 317852
rect 325108 317840 325114 317892
rect 149287 317784 151124 317812
rect 151817 317815 151875 317821
rect 149287 317781 149299 317784
rect 149241 317775 149299 317781
rect 151817 317781 151829 317815
rect 151863 317812 151875 317815
rect 160738 317812 160744 317824
rect 151863 317784 160744 317812
rect 151863 317781 151875 317784
rect 151817 317775 151875 317781
rect 160738 317772 160744 317784
rect 160796 317772 160802 317824
rect 182726 317772 182732 317824
rect 182784 317812 182790 317824
rect 189997 317815 190055 317821
rect 189997 317812 190009 317815
rect 182784 317784 190009 317812
rect 182784 317772 182790 317784
rect 189997 317781 190009 317784
rect 190043 317781 190055 317815
rect 189997 317775 190055 317781
rect 190089 317815 190147 317821
rect 190089 317781 190101 317815
rect 190135 317812 190147 317815
rect 193766 317812 193772 317824
rect 190135 317784 193772 317812
rect 190135 317781 190147 317784
rect 190089 317775 190147 317781
rect 193766 317772 193772 317784
rect 193824 317772 193830 317824
rect 318058 317812 318064 317824
rect 193876 317784 318064 317812
rect 155218 317744 155224 317756
rect 148888 317716 155224 317744
rect 155218 317704 155224 317716
rect 155276 317704 155282 317756
rect 177758 317704 177764 317756
rect 177816 317744 177822 317756
rect 184937 317747 184995 317753
rect 184937 317744 184949 317747
rect 177816 317716 184949 317744
rect 177816 317704 177822 317716
rect 184937 317713 184949 317716
rect 184983 317713 184995 317747
rect 184937 317707 184995 317713
rect 187694 317704 187700 317756
rect 187752 317744 187758 317756
rect 193876 317744 193904 317784
rect 318058 317772 318064 317784
rect 318116 317772 318122 317824
rect 187752 317716 193904 317744
rect 187752 317704 187758 317716
rect 196342 317704 196348 317756
rect 196400 317744 196406 317756
rect 197170 317744 197176 317756
rect 196400 317716 197176 317744
rect 196400 317704 196406 317716
rect 197170 317704 197176 317716
rect 197228 317704 197234 317756
rect 198826 317704 198832 317756
rect 198884 317744 198890 317756
rect 200022 317744 200028 317756
rect 198884 317716 200028 317744
rect 198884 317704 198890 317716
rect 200022 317704 200028 317716
rect 200080 317704 200086 317756
rect 202966 317704 202972 317756
rect 203024 317744 203030 317756
rect 204070 317744 204076 317756
rect 203024 317716 204076 317744
rect 203024 317704 203030 317716
rect 204070 317704 204076 317716
rect 204128 317704 204134 317756
rect 204165 317747 204223 317753
rect 204165 317713 204177 317747
rect 204211 317744 204223 317747
rect 212537 317747 212595 317753
rect 212537 317744 212549 317747
rect 204211 317716 212549 317744
rect 204211 317713 204223 317716
rect 204165 317707 204223 317713
rect 212537 317713 212549 317716
rect 212583 317713 212595 317747
rect 212537 317707 212595 317713
rect 224865 317747 224923 317753
rect 224865 317713 224877 317747
rect 224911 317744 224923 317747
rect 270497 317747 270555 317753
rect 270497 317744 270509 317747
rect 224911 317716 270509 317744
rect 224911 317713 224923 317716
rect 224865 317707 224923 317713
rect 270497 317713 270509 317716
rect 270543 317713 270555 317747
rect 270497 317707 270555 317713
rect 280065 317747 280123 317753
rect 280065 317713 280077 317747
rect 280111 317744 280123 317747
rect 289817 317747 289875 317753
rect 289817 317744 289829 317747
rect 280111 317716 289829 317744
rect 280111 317713 280123 317716
rect 280065 317707 280123 317713
rect 289817 317713 289829 317716
rect 289863 317713 289875 317747
rect 289817 317707 289875 317713
rect 299385 317747 299443 317753
rect 299385 317713 299397 317747
rect 299431 317744 299443 317747
rect 309137 317747 309195 317753
rect 309137 317744 309149 317747
rect 299431 317716 309149 317744
rect 299431 317713 299443 317716
rect 299385 317707 299443 317713
rect 309137 317713 309149 317716
rect 309183 317713 309195 317747
rect 309137 317707 309195 317713
rect 135898 317676 135904 317688
rect 132184 317648 132540 317676
rect 132696 317648 135904 317676
rect 132184 317636 132190 317648
rect 70397 317611 70455 317617
rect 70397 317577 70409 317611
rect 70443 317608 70455 317611
rect 84657 317611 84715 317617
rect 84657 317608 84669 317611
rect 70443 317580 84669 317608
rect 70443 317577 70455 317580
rect 70397 317571 70455 317577
rect 84657 317577 84669 317580
rect 84703 317577 84715 317611
rect 84657 317571 84715 317577
rect 84749 317611 84807 317617
rect 84749 317577 84761 317611
rect 84795 317608 84807 317611
rect 92474 317608 92480 317620
rect 84795 317580 92480 317608
rect 84795 317577 84807 317580
rect 84749 317571 84807 317577
rect 92474 317568 92480 317580
rect 92532 317568 92538 317620
rect 100018 317568 100024 317620
rect 100076 317608 100082 317620
rect 104342 317608 104348 317620
rect 100076 317580 104348 317608
rect 100076 317568 100082 317580
rect 104342 317568 104348 317580
rect 104400 317568 104406 317620
rect 117590 317568 117596 317620
rect 117648 317608 117654 317620
rect 118510 317608 118516 317620
rect 117648 317580 118516 317608
rect 117648 317568 117654 317580
rect 118510 317568 118516 317580
rect 118568 317568 118574 317620
rect 120442 317568 120448 317620
rect 120500 317608 120506 317620
rect 121362 317608 121368 317620
rect 120500 317580 121368 317608
rect 120500 317568 120506 317580
rect 121362 317568 121368 317580
rect 121420 317568 121426 317620
rect 132512 317608 132540 317648
rect 135898 317636 135904 317648
rect 135956 317636 135962 317688
rect 138198 317636 138204 317688
rect 138256 317676 138262 317688
rect 141881 317679 141939 317685
rect 141881 317676 141893 317679
rect 138256 317648 141893 317676
rect 138256 317636 138262 317648
rect 141881 317645 141893 317648
rect 141927 317645 141939 317679
rect 141881 317639 141939 317645
rect 141973 317679 142031 317685
rect 141973 317645 141985 317679
rect 142019 317676 142031 317679
rect 145009 317679 145067 317685
rect 142019 317648 144960 317676
rect 142019 317645 142031 317648
rect 141973 317639 142031 317645
rect 139305 317611 139363 317617
rect 139305 317608 139317 317611
rect 132512 317580 139317 317608
rect 139305 317577 139317 317580
rect 139351 317577 139363 317611
rect 139305 317571 139363 317577
rect 139394 317568 139400 317620
rect 139452 317608 139458 317620
rect 140682 317608 140688 317620
rect 139452 317580 140688 317608
rect 139452 317568 139458 317580
rect 140682 317568 140688 317580
rect 140740 317568 140746 317620
rect 140777 317611 140835 317617
rect 140777 317577 140789 317611
rect 140823 317608 140835 317611
rect 142893 317611 142951 317617
rect 142893 317608 142905 317611
rect 140823 317580 142905 317608
rect 140823 317577 140835 317580
rect 140777 317571 140835 317577
rect 142893 317577 142905 317580
rect 142939 317577 142951 317611
rect 142893 317571 142951 317577
rect 144362 317568 144368 317620
rect 144420 317608 144426 317620
rect 144822 317608 144828 317620
rect 144420 317580 144828 317608
rect 144420 317568 144426 317580
rect 144822 317568 144828 317580
rect 144880 317568 144886 317620
rect 144932 317608 144960 317648
rect 145009 317645 145021 317679
rect 145055 317676 145067 317679
rect 158070 317676 158076 317688
rect 145055 317648 158076 317676
rect 145055 317645 145067 317648
rect 145009 317639 145067 317645
rect 158070 317636 158076 317648
rect 158128 317636 158134 317688
rect 180242 317636 180248 317688
rect 180300 317676 180306 317688
rect 180300 317648 184980 317676
rect 180300 317636 180306 317648
rect 151078 317608 151084 317620
rect 144932 317580 151084 317608
rect 151078 317568 151084 317580
rect 151136 317568 151142 317620
rect 153930 317608 153936 317620
rect 151188 317580 153936 317608
rect 64690 317500 64696 317552
rect 64748 317540 64754 317552
rect 92014 317540 92020 317552
rect 64748 317512 92020 317540
rect 64748 317500 64754 317512
rect 92014 317500 92020 317512
rect 92072 317500 92078 317552
rect 103422 317500 103428 317552
rect 103480 317540 103486 317552
rect 105630 317540 105636 317552
rect 103480 317512 105636 317540
rect 103480 317500 103486 317512
rect 105630 317500 105636 317512
rect 105688 317500 105694 317552
rect 137738 317500 137744 317552
rect 137796 317540 137802 317552
rect 151188 317540 151216 317580
rect 153930 317568 153936 317580
rect 153988 317568 153994 317620
rect 154025 317611 154083 317617
rect 154025 317577 154037 317611
rect 154071 317608 154083 317611
rect 166166 317608 166172 317620
rect 154071 317580 166172 317608
rect 154071 317577 154083 317580
rect 154025 317571 154083 317577
rect 166166 317568 166172 317580
rect 166224 317568 166230 317620
rect 171594 317568 171600 317620
rect 171652 317608 171658 317620
rect 172146 317608 172152 317620
rect 171652 317580 172152 317608
rect 171652 317568 171658 317580
rect 172146 317568 172152 317580
rect 172204 317568 172210 317620
rect 183922 317568 183928 317620
rect 183980 317608 183986 317620
rect 184842 317608 184848 317620
rect 183980 317580 184848 317608
rect 183980 317568 183986 317580
rect 184842 317568 184848 317580
rect 184900 317568 184906 317620
rect 184952 317608 184980 317648
rect 186406 317636 186412 317688
rect 186464 317676 186470 317688
rect 187602 317676 187608 317688
rect 186464 317648 187608 317676
rect 186464 317636 186470 317648
rect 187602 317636 187608 317648
rect 187660 317636 187666 317688
rect 189718 317636 189724 317688
rect 189776 317676 189782 317688
rect 190270 317676 190276 317688
rect 189776 317648 190276 317676
rect 189776 317636 189782 317648
rect 190270 317636 190276 317648
rect 190328 317636 190334 317688
rect 191006 317636 191012 317688
rect 191064 317676 191070 317688
rect 191558 317676 191564 317688
rect 191064 317648 191564 317676
rect 191064 317636 191070 317648
rect 191558 317636 191564 317648
rect 191616 317636 191622 317688
rect 191834 317636 191840 317688
rect 191892 317676 191898 317688
rect 193030 317676 193036 317688
rect 191892 317648 193036 317676
rect 191892 317636 191898 317648
rect 193030 317636 193036 317648
rect 193088 317636 193094 317688
rect 193858 317636 193864 317688
rect 193916 317676 193922 317688
rect 194502 317676 194508 317688
rect 193916 317648 194508 317676
rect 193916 317636 193922 317648
rect 194502 317636 194508 317648
rect 194560 317636 194566 317688
rect 194686 317636 194692 317688
rect 194744 317676 194750 317688
rect 195790 317676 195796 317688
rect 194744 317648 195796 317676
rect 194744 317636 194750 317648
rect 195790 317636 195796 317648
rect 195848 317636 195854 317688
rect 195885 317679 195943 317685
rect 195885 317645 195897 317679
rect 195931 317676 195943 317679
rect 313918 317676 313924 317688
rect 195931 317648 313924 317676
rect 195931 317645 195943 317648
rect 195885 317639 195943 317645
rect 313918 317636 313924 317648
rect 313976 317636 313982 317688
rect 307018 317608 307024 317620
rect 184952 317580 307024 317608
rect 307018 317568 307024 317580
rect 307076 317568 307082 317620
rect 309137 317611 309195 317617
rect 309137 317577 309149 317611
rect 309183 317608 309195 317611
rect 311158 317608 311164 317620
rect 309183 317580 311164 317608
rect 309183 317577 309195 317580
rect 309137 317571 309195 317577
rect 311158 317568 311164 317580
rect 311216 317568 311222 317620
rect 137796 317512 151216 317540
rect 137796 317500 137802 317512
rect 152182 317500 152188 317552
rect 152240 317540 152246 317552
rect 153102 317540 153108 317552
rect 152240 317512 153108 317540
rect 152240 317500 152246 317512
rect 153102 317500 153108 317512
rect 153160 317500 153166 317552
rect 154666 317500 154672 317552
rect 154724 317540 154730 317552
rect 155862 317540 155868 317552
rect 154724 317512 155868 317540
rect 154724 317500 154730 317512
rect 155862 317500 155868 317512
rect 155920 317500 155926 317552
rect 155954 317500 155960 317552
rect 156012 317540 156018 317552
rect 157242 317540 157248 317552
rect 156012 317512 157248 317540
rect 156012 317500 156018 317512
rect 157242 317500 157248 317512
rect 157300 317500 157306 317552
rect 158806 317500 158812 317552
rect 158864 317540 158870 317552
rect 159910 317540 159916 317552
rect 158864 317512 159916 317540
rect 158864 317500 158870 317512
rect 159910 317500 159916 317512
rect 159968 317500 159974 317552
rect 163774 317500 163780 317552
rect 163832 317540 163838 317552
rect 164050 317540 164056 317552
rect 163832 317512 164056 317540
rect 163832 317500 163838 317512
rect 164050 317500 164056 317512
rect 164108 317500 164114 317552
rect 164970 317500 164976 317552
rect 165028 317540 165034 317552
rect 165522 317540 165528 317552
rect 165028 317512 165528 317540
rect 165028 317500 165034 317512
rect 165522 317500 165528 317512
rect 165580 317500 165586 317552
rect 165798 317500 165804 317552
rect 165856 317540 165862 317552
rect 166902 317540 166908 317552
rect 165856 317512 166908 317540
rect 165856 317500 165862 317512
rect 166902 317500 166908 317512
rect 166960 317500 166966 317552
rect 167454 317500 167460 317552
rect 167512 317540 167518 317552
rect 168282 317540 168288 317552
rect 167512 317512 168288 317540
rect 167512 317500 167518 317512
rect 168282 317500 168288 317512
rect 168340 317500 168346 317552
rect 171962 317500 171968 317552
rect 172020 317540 172026 317552
rect 172422 317540 172428 317552
rect 172020 317512 172428 317540
rect 172020 317500 172026 317512
rect 172422 317500 172428 317512
rect 172480 317500 172486 317552
rect 173250 317500 173256 317552
rect 173308 317540 173314 317552
rect 173802 317540 173808 317552
rect 173308 317512 173808 317540
rect 173308 317500 173314 317512
rect 173802 317500 173808 317512
rect 173860 317500 173866 317552
rect 174078 317500 174084 317552
rect 174136 317540 174142 317552
rect 175182 317540 175188 317552
rect 174136 317512 175188 317540
rect 174136 317500 174142 317512
rect 175182 317500 175188 317512
rect 175240 317500 175246 317552
rect 175734 317500 175740 317552
rect 175792 317540 175798 317552
rect 176562 317540 176568 317552
rect 175792 317512 176568 317540
rect 175792 317500 175798 317512
rect 176562 317500 176568 317512
rect 176620 317500 176626 317552
rect 177390 317500 177396 317552
rect 177448 317540 177454 317552
rect 177850 317540 177856 317552
rect 177448 317512 177856 317540
rect 177448 317500 177454 317512
rect 177850 317500 177856 317512
rect 177908 317500 177914 317552
rect 178586 317500 178592 317552
rect 178644 317540 178650 317552
rect 179046 317540 179052 317552
rect 178644 317512 179052 317540
rect 178644 317500 178650 317512
rect 179046 317500 179052 317512
rect 179104 317500 179110 317552
rect 179414 317500 179420 317552
rect 179472 317540 179478 317552
rect 180702 317540 180708 317552
rect 179472 317512 180708 317540
rect 179472 317500 179478 317512
rect 180702 317500 180708 317512
rect 180760 317500 180766 317552
rect 183554 317500 183560 317552
rect 183612 317540 183618 317552
rect 184658 317540 184664 317552
rect 183612 317512 184664 317540
rect 183612 317500 183618 317512
rect 184658 317500 184664 317512
rect 184716 317500 184722 317552
rect 184937 317543 184995 317549
rect 184937 317509 184949 317543
rect 184983 317540 184995 317543
rect 300118 317540 300124 317552
rect 184983 317512 300124 317540
rect 184983 317509 184995 317512
rect 184937 317503 184995 317509
rect 300118 317500 300124 317512
rect 300176 317500 300182 317552
rect 68278 317432 68284 317484
rect 68336 317472 68342 317484
rect 68336 317444 69612 317472
rect 68336 317432 68342 317444
rect 69584 317336 69612 317444
rect 69658 317432 69664 317484
rect 69716 317472 69722 317484
rect 88334 317472 88340 317484
rect 69716 317444 88340 317472
rect 69716 317432 69722 317444
rect 88334 317432 88340 317444
rect 88392 317432 88398 317484
rect 100110 317432 100116 317484
rect 100168 317472 100174 317484
rect 101950 317472 101956 317484
rect 100168 317444 101956 317472
rect 100168 317432 100174 317444
rect 101950 317432 101956 317444
rect 102008 317432 102014 317484
rect 102778 317432 102784 317484
rect 102836 317472 102842 317484
rect 103974 317472 103980 317484
rect 102836 317444 103980 317472
rect 102836 317432 102842 317444
rect 103974 317432 103980 317444
rect 104032 317432 104038 317484
rect 104802 317432 104808 317484
rect 104860 317472 104866 317484
rect 105998 317472 106004 317484
rect 104860 317444 106004 317472
rect 104860 317432 104866 317444
rect 105998 317432 106004 317444
rect 106056 317432 106062 317484
rect 108114 317432 108120 317484
rect 108172 317472 108178 317484
rect 108850 317472 108856 317484
rect 108172 317444 108856 317472
rect 108172 317432 108178 317444
rect 108850 317432 108856 317444
rect 108908 317432 108914 317484
rect 110598 317432 110604 317484
rect 110656 317472 110662 317484
rect 113818 317472 113824 317484
rect 110656 317444 113824 317472
rect 110656 317432 110662 317444
rect 113818 317432 113824 317444
rect 113876 317432 113882 317484
rect 133690 317432 133696 317484
rect 133748 317472 133754 317484
rect 138477 317475 138535 317481
rect 138477 317472 138489 317475
rect 133748 317444 138489 317472
rect 133748 317432 133754 317444
rect 138477 317441 138489 317444
rect 138523 317441 138535 317475
rect 138477 317435 138535 317441
rect 138566 317432 138572 317484
rect 138624 317472 138630 317484
rect 139302 317472 139308 317484
rect 138624 317444 139308 317472
rect 138624 317432 138630 317444
rect 139302 317432 139308 317444
rect 139360 317432 139366 317484
rect 139854 317432 139860 317484
rect 139912 317472 139918 317484
rect 140590 317472 140596 317484
rect 139912 317444 140596 317472
rect 139912 317432 139918 317444
rect 140590 317432 140596 317444
rect 140648 317432 140654 317484
rect 141050 317432 141056 317484
rect 141108 317472 141114 317484
rect 142062 317472 142068 317484
rect 141108 317444 142068 317472
rect 141108 317432 141114 317444
rect 142062 317432 142068 317444
rect 142120 317432 142126 317484
rect 142338 317432 142344 317484
rect 142396 317472 142402 317484
rect 143442 317472 143448 317484
rect 142396 317444 143448 317472
rect 142396 317432 142402 317444
rect 143442 317432 143448 317444
rect 143500 317432 143506 317484
rect 143534 317432 143540 317484
rect 143592 317472 143598 317484
rect 144638 317472 144644 317484
rect 143592 317444 144644 317472
rect 143592 317432 143598 317444
rect 144638 317432 144644 317444
rect 144696 317432 144702 317484
rect 145190 317432 145196 317484
rect 145248 317472 145254 317484
rect 146110 317472 146116 317484
rect 145248 317444 146116 317472
rect 145248 317432 145254 317444
rect 146110 317432 146116 317444
rect 146168 317432 146174 317484
rect 146478 317432 146484 317484
rect 146536 317472 146542 317484
rect 147398 317472 147404 317484
rect 146536 317444 147404 317472
rect 146536 317432 146542 317444
rect 147398 317432 147404 317444
rect 147456 317432 147462 317484
rect 148413 317475 148471 317481
rect 148413 317472 148425 317475
rect 147508 317444 148425 317472
rect 92845 317407 92903 317413
rect 92845 317373 92857 317407
rect 92891 317404 92903 317407
rect 93026 317404 93032 317416
rect 92891 317376 93032 317404
rect 92891 317373 92903 317376
rect 92845 317367 92903 317373
rect 93026 317364 93032 317376
rect 93084 317364 93090 317416
rect 94038 317404 94044 317416
rect 93999 317376 94044 317404
rect 94038 317364 94044 317376
rect 94096 317364 94102 317416
rect 139210 317364 139216 317416
rect 139268 317404 139274 317416
rect 147508 317404 147536 317444
rect 148413 317441 148425 317444
rect 148459 317441 148471 317475
rect 148413 317435 148471 317441
rect 148502 317432 148508 317484
rect 148560 317472 148566 317484
rect 148962 317472 148968 317484
rect 148560 317444 148968 317472
rect 148560 317432 148566 317444
rect 148962 317432 148968 317444
rect 149020 317432 149026 317484
rect 151725 317475 151783 317481
rect 151725 317472 151737 317475
rect 149072 317444 151737 317472
rect 139268 317376 147536 317404
rect 147677 317407 147735 317413
rect 139268 317364 139274 317376
rect 147677 317373 147689 317407
rect 147723 317404 147735 317407
rect 149072 317404 149100 317444
rect 151725 317441 151737 317444
rect 151771 317441 151783 317475
rect 151725 317435 151783 317441
rect 151814 317432 151820 317484
rect 151872 317472 151878 317484
rect 152642 317472 152648 317484
rect 151872 317444 152648 317472
rect 151872 317432 151878 317444
rect 152642 317432 152648 317444
rect 152700 317432 152706 317484
rect 153470 317432 153476 317484
rect 153528 317472 153534 317484
rect 154482 317472 154488 317484
rect 153528 317444 154488 317472
rect 153528 317432 153534 317444
rect 154482 317432 154488 317444
rect 154540 317432 154546 317484
rect 155126 317432 155132 317484
rect 155184 317472 155190 317484
rect 155770 317472 155776 317484
rect 155184 317444 155776 317472
rect 155184 317432 155190 317444
rect 155770 317432 155776 317444
rect 155828 317432 155834 317484
rect 156322 317432 156328 317484
rect 156380 317472 156386 317484
rect 157058 317472 157064 317484
rect 156380 317444 157064 317472
rect 156380 317432 156386 317444
rect 157058 317432 157064 317444
rect 157116 317432 157122 317484
rect 159634 317432 159640 317484
rect 159692 317472 159698 317484
rect 160002 317472 160008 317484
rect 159692 317444 160008 317472
rect 159692 317432 159698 317444
rect 160002 317432 160008 317444
rect 160060 317432 160066 317484
rect 160830 317432 160836 317484
rect 160888 317472 160894 317484
rect 161382 317472 161388 317484
rect 160888 317444 161388 317472
rect 160888 317432 160894 317444
rect 161382 317432 161388 317444
rect 161440 317432 161446 317484
rect 162118 317432 162124 317484
rect 162176 317472 162182 317484
rect 162762 317472 162768 317484
rect 162176 317444 162768 317472
rect 162176 317432 162182 317444
rect 162762 317432 162768 317444
rect 162820 317432 162826 317484
rect 163314 317432 163320 317484
rect 163372 317472 163378 317484
rect 164142 317472 164148 317484
rect 163372 317444 164148 317472
rect 163372 317432 163378 317444
rect 164142 317432 164148 317444
rect 164200 317432 164206 317484
rect 164602 317432 164608 317484
rect 164660 317472 164666 317484
rect 165338 317472 165344 317484
rect 164660 317444 165344 317472
rect 164660 317432 164666 317444
rect 165338 317432 165344 317444
rect 165396 317432 165402 317484
rect 166258 317432 166264 317484
rect 166316 317472 166322 317484
rect 166810 317472 166816 317484
rect 166316 317444 166816 317472
rect 166316 317432 166322 317444
rect 166810 317432 166816 317444
rect 166868 317432 166874 317484
rect 167086 317432 167092 317484
rect 167144 317472 167150 317484
rect 168098 317472 168104 317484
rect 167144 317444 168104 317472
rect 167144 317432 167150 317444
rect 168098 317432 168104 317444
rect 168156 317432 168162 317484
rect 168742 317432 168748 317484
rect 168800 317472 168806 317484
rect 169570 317472 169576 317484
rect 168800 317444 169576 317472
rect 168800 317432 168806 317444
rect 169570 317432 169576 317444
rect 169628 317432 169634 317484
rect 169938 317432 169944 317484
rect 169996 317472 170002 317484
rect 170950 317472 170956 317484
rect 169996 317444 170956 317472
rect 169996 317432 170002 317444
rect 170950 317432 170956 317444
rect 171008 317432 171014 317484
rect 171226 317432 171232 317484
rect 171284 317472 171290 317484
rect 172238 317472 172244 317484
rect 171284 317444 172244 317472
rect 171284 317432 171290 317444
rect 172238 317432 172244 317444
rect 172296 317432 172302 317484
rect 172790 317432 172796 317484
rect 172848 317472 172854 317484
rect 173618 317472 173624 317484
rect 172848 317444 173624 317472
rect 172848 317432 172854 317444
rect 173618 317432 173624 317444
rect 173676 317432 173682 317484
rect 174446 317432 174452 317484
rect 174504 317472 174510 317484
rect 175090 317472 175096 317484
rect 174504 317444 175096 317472
rect 174504 317432 174510 317444
rect 175090 317432 175096 317444
rect 175148 317432 175154 317484
rect 175274 317432 175280 317484
rect 175332 317472 175338 317484
rect 176286 317472 176292 317484
rect 175332 317444 176292 317472
rect 175332 317432 175338 317444
rect 176286 317432 176292 317444
rect 176344 317432 176350 317484
rect 176930 317432 176936 317484
rect 176988 317472 176994 317484
rect 177942 317472 177948 317484
rect 176988 317444 177948 317472
rect 176988 317432 176994 317444
rect 177942 317432 177948 317444
rect 178000 317432 178006 317484
rect 178218 317432 178224 317484
rect 178276 317472 178282 317484
rect 179138 317472 179144 317484
rect 178276 317444 179144 317472
rect 178276 317432 178282 317444
rect 179138 317432 179144 317444
rect 179196 317432 179202 317484
rect 179874 317432 179880 317484
rect 179932 317472 179938 317484
rect 180518 317472 180524 317484
rect 179932 317444 180524 317472
rect 179932 317432 179938 317444
rect 180518 317432 180524 317444
rect 180576 317432 180582 317484
rect 181070 317432 181076 317484
rect 181128 317472 181134 317484
rect 181622 317472 181628 317484
rect 181128 317444 181628 317472
rect 181128 317432 181134 317444
rect 181622 317432 181628 317444
rect 181680 317432 181686 317484
rect 182358 317432 182364 317484
rect 182416 317472 182422 317484
rect 183186 317472 183192 317484
rect 182416 317444 183192 317472
rect 182416 317432 182422 317444
rect 183186 317432 183192 317444
rect 183244 317432 183250 317484
rect 184382 317432 184388 317484
rect 184440 317472 184446 317484
rect 184750 317472 184756 317484
rect 184440 317444 184756 317472
rect 184440 317432 184446 317444
rect 184750 317432 184756 317444
rect 184808 317432 184814 317484
rect 185578 317432 185584 317484
rect 185636 317472 185642 317484
rect 186222 317472 186228 317484
rect 185636 317444 186228 317472
rect 185636 317432 185642 317444
rect 186222 317432 186228 317444
rect 186280 317432 186286 317484
rect 186866 317432 186872 317484
rect 186924 317472 186930 317484
rect 187510 317472 187516 317484
rect 186924 317444 187516 317472
rect 186924 317432 186930 317444
rect 187510 317432 187516 317444
rect 187568 317432 187574 317484
rect 188062 317432 188068 317484
rect 188120 317472 188126 317484
rect 188890 317472 188896 317484
rect 188120 317444 188896 317472
rect 188120 317432 188126 317444
rect 188890 317432 188896 317444
rect 188948 317432 188954 317484
rect 189350 317432 189356 317484
rect 189408 317472 189414 317484
rect 190362 317472 190368 317484
rect 189408 317444 190368 317472
rect 189408 317432 189414 317444
rect 190362 317432 190368 317444
rect 190420 317432 190426 317484
rect 190546 317432 190552 317484
rect 190604 317472 190610 317484
rect 191742 317472 191748 317484
rect 190604 317444 191748 317472
rect 190604 317432 190610 317444
rect 191742 317432 191748 317444
rect 191800 317432 191806 317484
rect 192202 317432 192208 317484
rect 192260 317472 192266 317484
rect 192938 317472 192944 317484
rect 192260 317444 192944 317472
rect 192260 317432 192266 317444
rect 192938 317432 192944 317444
rect 192996 317432 193002 317484
rect 193490 317432 193496 317484
rect 193548 317472 193554 317484
rect 194318 317472 194324 317484
rect 193548 317444 194324 317472
rect 193548 317432 193554 317444
rect 194318 317432 194324 317444
rect 194376 317432 194382 317484
rect 195514 317432 195520 317484
rect 195572 317472 195578 317484
rect 195882 317472 195888 317484
rect 195572 317444 195888 317472
rect 195572 317432 195578 317444
rect 195882 317432 195888 317444
rect 195940 317432 195946 317484
rect 196710 317432 196716 317484
rect 196768 317472 196774 317484
rect 197262 317472 197268 317484
rect 196768 317444 197268 317472
rect 196768 317432 196774 317444
rect 197262 317432 197268 317444
rect 197320 317432 197326 317484
rect 197998 317432 198004 317484
rect 198056 317472 198062 317484
rect 198642 317472 198648 317484
rect 198056 317444 198648 317472
rect 198056 317432 198062 317444
rect 198642 317432 198648 317444
rect 198700 317432 198706 317484
rect 199194 317432 199200 317484
rect 199252 317472 199258 317484
rect 199930 317472 199936 317484
rect 199252 317444 199936 317472
rect 199252 317432 199258 317444
rect 199930 317432 199936 317444
rect 199988 317432 199994 317484
rect 200482 317432 200488 317484
rect 200540 317472 200546 317484
rect 201218 317472 201224 317484
rect 200540 317444 201224 317472
rect 200540 317432 200546 317444
rect 201218 317432 201224 317444
rect 201276 317432 201282 317484
rect 201678 317432 201684 317484
rect 201736 317472 201742 317484
rect 202782 317472 202788 317484
rect 201736 317444 202788 317472
rect 201736 317432 201742 317444
rect 202782 317432 202788 317444
rect 202840 317432 202846 317484
rect 203794 317432 203800 317484
rect 203852 317472 203858 317484
rect 204162 317472 204168 317484
rect 203852 317444 204168 317472
rect 203852 317432 203858 317444
rect 204162 317432 204168 317444
rect 204220 317432 204226 317484
rect 204622 317432 204628 317484
rect 204680 317472 204686 317484
rect 205450 317472 205456 317484
rect 204680 317444 205456 317472
rect 204680 317432 204686 317444
rect 205450 317432 205456 317444
rect 205508 317432 205514 317484
rect 205818 317432 205824 317484
rect 205876 317472 205882 317484
rect 206738 317472 206744 317484
rect 205876 317444 206744 317472
rect 205876 317432 205882 317444
rect 206738 317432 206744 317444
rect 206796 317432 206802 317484
rect 207014 317432 207020 317484
rect 207072 317472 207078 317484
rect 208026 317472 208032 317484
rect 207072 317444 208032 317472
rect 207072 317432 207078 317444
rect 208026 317432 208032 317444
rect 208084 317432 208090 317484
rect 209130 317432 209136 317484
rect 209188 317472 209194 317484
rect 209682 317472 209688 317484
rect 209188 317444 209688 317472
rect 209188 317432 209194 317444
rect 209682 317432 209688 317444
rect 209740 317432 209746 317484
rect 210326 317432 210332 317484
rect 210384 317472 210390 317484
rect 211062 317472 211068 317484
rect 210384 317444 211068 317472
rect 210384 317432 210390 317444
rect 211062 317432 211068 317444
rect 211120 317432 211126 317484
rect 211154 317432 211160 317484
rect 211212 317472 211218 317484
rect 212074 317472 212080 317484
rect 211212 317444 212080 317472
rect 211212 317432 211218 317444
rect 212074 317432 212080 317444
rect 212132 317432 212138 317484
rect 212810 317432 212816 317484
rect 212868 317472 212874 317484
rect 213730 317472 213736 317484
rect 212868 317444 213736 317472
rect 212868 317432 212874 317444
rect 213730 317432 213736 317444
rect 213788 317432 213794 317484
rect 213825 317475 213883 317481
rect 213825 317441 213837 317475
rect 213871 317472 213883 317475
rect 276658 317472 276664 317484
rect 213871 317444 276664 317472
rect 213871 317441 213883 317444
rect 213825 317435 213883 317441
rect 276658 317432 276664 317444
rect 276716 317432 276722 317484
rect 289817 317475 289875 317481
rect 289817 317441 289829 317475
rect 289863 317472 289875 317475
rect 299385 317475 299443 317481
rect 299385 317472 299397 317475
rect 289863 317444 299397 317472
rect 289863 317441 289875 317444
rect 289817 317435 289875 317441
rect 299385 317441 299397 317444
rect 299431 317441 299443 317475
rect 299385 317435 299443 317441
rect 147723 317376 149100 317404
rect 212537 317407 212595 317413
rect 147723 317373 147735 317376
rect 147677 317367 147735 317373
rect 212537 317373 212549 317407
rect 212583 317404 212595 317407
rect 224865 317407 224923 317413
rect 224865 317404 224877 317407
rect 212583 317376 224877 317404
rect 212583 317373 212595 317376
rect 212537 317367 212595 317373
rect 224865 317373 224877 317376
rect 224911 317373 224923 317407
rect 236178 317404 236184 317416
rect 236139 317376 236184 317404
rect 224865 317367 224923 317373
rect 236178 317364 236184 317376
rect 236236 317364 236242 317416
rect 237650 317364 237656 317416
rect 237708 317404 237714 317416
rect 238570 317404 238576 317416
rect 237708 317376 238576 317404
rect 237708 317364 237714 317376
rect 238570 317364 238576 317376
rect 238628 317364 238634 317416
rect 238938 317404 238944 317416
rect 238899 317376 238944 317404
rect 238938 317364 238944 317376
rect 238996 317364 239002 317416
rect 240502 317364 240508 317416
rect 240560 317404 240566 317416
rect 241238 317404 241244 317416
rect 240560 317376 241244 317404
rect 240560 317364 240566 317376
rect 241238 317364 241244 317376
rect 241296 317364 241302 317416
rect 248138 317364 248144 317416
rect 248196 317404 248202 317416
rect 248322 317404 248328 317416
rect 248196 317376 248328 317404
rect 248196 317364 248202 317376
rect 248322 317364 248328 317376
rect 248380 317364 248386 317416
rect 266906 317364 266912 317416
rect 266964 317404 266970 317416
rect 267642 317404 267648 317416
rect 266964 317376 267648 317404
rect 266964 317364 266970 317376
rect 267642 317364 267648 317376
rect 267700 317364 267706 317416
rect 267734 317364 267740 317416
rect 267792 317404 267798 317416
rect 268930 317404 268936 317416
rect 267792 317376 268936 317404
rect 267792 317364 267798 317376
rect 268930 317364 268936 317376
rect 268988 317364 268994 317416
rect 270497 317407 270555 317413
rect 270497 317373 270509 317407
rect 270543 317404 270555 317407
rect 280065 317407 280123 317413
rect 280065 317404 280077 317407
rect 270543 317376 280077 317404
rect 270543 317373 270555 317376
rect 270497 317367 270555 317373
rect 280065 317373 280077 317376
rect 280111 317373 280123 317407
rect 280065 317367 280123 317373
rect 70397 317339 70455 317345
rect 70397 317336 70409 317339
rect 69584 317308 70409 317336
rect 70397 317305 70409 317308
rect 70443 317305 70455 317339
rect 70397 317299 70455 317305
rect 139305 317339 139363 317345
rect 139305 317305 139317 317339
rect 139351 317336 139363 317339
rect 140777 317339 140835 317345
rect 140777 317336 140789 317339
rect 139351 317308 140789 317336
rect 139351 317305 139363 317308
rect 139305 317299 139363 317305
rect 140777 317305 140789 317308
rect 140823 317305 140835 317339
rect 140777 317299 140835 317305
rect 141881 317339 141939 317345
rect 141881 317305 141893 317339
rect 141927 317336 141939 317339
rect 145653 317339 145711 317345
rect 145653 317336 145665 317339
rect 141927 317308 145665 317336
rect 141927 317305 141939 317308
rect 141881 317299 141939 317305
rect 145653 317305 145665 317308
rect 145699 317305 145711 317339
rect 145653 317299 145711 317305
rect 238846 316140 238852 316192
rect 238904 316180 238910 316192
rect 239950 316180 239956 316192
rect 238904 316152 239956 316180
rect 238904 316140 238910 316152
rect 239950 316140 239956 316152
rect 240008 316140 240014 316192
rect 251358 316140 251364 316192
rect 251416 316180 251422 316192
rect 252462 316180 252468 316192
rect 251416 316152 252468 316180
rect 251416 316140 251422 316152
rect 252462 316140 252468 316152
rect 252520 316140 252526 316192
rect 95234 316072 95240 316124
rect 95292 316112 95298 316124
rect 95878 316112 95884 316124
rect 95292 316084 95884 316112
rect 95292 316072 95298 316084
rect 95878 316072 95884 316084
rect 95936 316072 95942 316124
rect 244090 316072 244096 316124
rect 244148 316072 244154 316124
rect 256970 316072 256976 316124
rect 257028 316112 257034 316124
rect 257798 316112 257804 316124
rect 257028 316084 257804 316112
rect 257028 316072 257034 316084
rect 257798 316072 257804 316084
rect 257856 316072 257862 316124
rect 75914 316004 75920 316056
rect 75972 316044 75978 316056
rect 76466 316044 76472 316056
rect 75972 316016 76472 316044
rect 75972 316004 75978 316016
rect 76466 316004 76472 316016
rect 76524 316004 76530 316056
rect 93946 316004 93952 316056
rect 94004 316044 94010 316056
rect 94590 316044 94596 316056
rect 94004 316016 94596 316044
rect 94004 316004 94010 316016
rect 94590 316004 94596 316016
rect 94648 316004 94654 316056
rect 234890 316004 234896 316056
rect 234948 316044 234954 316056
rect 235626 316044 235632 316056
rect 234948 316016 235632 316044
rect 234948 316004 234954 316016
rect 235626 316004 235632 316016
rect 235684 316004 235690 316056
rect 238846 316004 238852 316056
rect 238904 316044 238910 316056
rect 239766 316044 239772 316056
rect 238904 316016 239772 316044
rect 238904 316004 238910 316016
rect 239766 316004 239772 316016
rect 239824 316004 239830 316056
rect 70394 315936 70400 315988
rect 70452 315976 70458 315988
rect 71038 315976 71044 315988
rect 70452 315948 71044 315976
rect 70452 315936 70458 315948
rect 71038 315936 71044 315948
rect 71096 315936 71102 315988
rect 71866 315936 71872 315988
rect 71924 315976 71930 315988
rect 72694 315976 72700 315988
rect 71924 315948 72700 315976
rect 71924 315936 71930 315948
rect 72694 315936 72700 315948
rect 72752 315936 72758 315988
rect 73154 315936 73160 315988
rect 73212 315976 73218 315988
rect 73982 315976 73988 315988
rect 73212 315948 73988 315976
rect 73212 315936 73218 315948
rect 73982 315936 73988 315948
rect 74040 315936 74046 315988
rect 76006 315936 76012 315988
rect 76064 315976 76070 315988
rect 76926 315976 76932 315988
rect 76064 315948 76932 315976
rect 76064 315936 76070 315948
rect 76926 315936 76932 315948
rect 76984 315936 76990 315988
rect 81526 315936 81532 315988
rect 81584 315976 81590 315988
rect 82262 315976 82268 315988
rect 81584 315948 82268 315976
rect 81584 315936 81590 315948
rect 82262 315936 82268 315948
rect 82320 315936 82326 315988
rect 88426 315936 88432 315988
rect 88484 315976 88490 315988
rect 88886 315976 88892 315988
rect 88484 315948 88892 315976
rect 88484 315936 88490 315948
rect 88886 315936 88892 315948
rect 88944 315936 88950 315988
rect 92566 315936 92572 315988
rect 92624 315976 92630 315988
rect 93302 315976 93308 315988
rect 92624 315948 93308 315976
rect 92624 315936 92630 315948
rect 93302 315936 93308 315948
rect 93360 315936 93366 315988
rect 93854 315936 93860 315988
rect 93912 315976 93918 315988
rect 94222 315976 94228 315988
rect 93912 315948 94228 315976
rect 93912 315936 93918 315948
rect 94222 315936 94228 315948
rect 94280 315936 94286 315988
rect 96614 315936 96620 315988
rect 96672 315976 96678 315988
rect 97534 315976 97540 315988
rect 96672 315948 97540 315976
rect 96672 315936 96678 315948
rect 97534 315936 97540 315948
rect 97592 315936 97598 315988
rect 228726 315936 228732 315988
rect 228784 315976 228790 315988
rect 229002 315976 229008 315988
rect 228784 315948 229008 315976
rect 228784 315936 228790 315948
rect 229002 315936 229008 315948
rect 229060 315936 229066 315988
rect 234614 315936 234620 315988
rect 234672 315976 234678 315988
rect 235442 315976 235448 315988
rect 234672 315948 235448 315976
rect 234672 315936 234678 315948
rect 235442 315936 235448 315948
rect 235500 315936 235506 315988
rect 235994 315936 236000 315988
rect 236052 315976 236058 315988
rect 236454 315976 236460 315988
rect 236052 315948 236460 315976
rect 236052 315936 236058 315948
rect 236454 315936 236460 315948
rect 236512 315936 236518 315988
rect 237466 315936 237472 315988
rect 237524 315976 237530 315988
rect 238110 315976 238116 315988
rect 237524 315948 238116 315976
rect 237524 315936 237530 315948
rect 238110 315936 238116 315948
rect 238168 315936 238174 315988
rect 238754 315936 238760 315988
rect 238812 315976 238818 315988
rect 239306 315976 239312 315988
rect 238812 315948 239312 315976
rect 238812 315936 238818 315948
rect 239306 315936 239312 315948
rect 239364 315936 239370 315988
rect 240134 315936 240140 315988
rect 240192 315976 240198 315988
rect 240962 315976 240968 315988
rect 240192 315948 240968 315976
rect 240192 315936 240198 315948
rect 240962 315936 240968 315948
rect 241020 315936 241026 315988
rect 241514 315936 241520 315988
rect 241572 315976 241578 315988
rect 242158 315976 242164 315988
rect 241572 315948 242164 315976
rect 241572 315936 241578 315948
rect 242158 315936 242164 315948
rect 242216 315936 242222 315988
rect 242894 315936 242900 315988
rect 242952 315976 242958 315988
rect 243078 315976 243084 315988
rect 242952 315948 243084 315976
rect 242952 315936 242958 315948
rect 243078 315936 243084 315948
rect 243136 315936 243142 315988
rect 244108 315920 244136 316072
rect 270494 316004 270500 316056
rect 270552 316044 270558 316056
rect 271690 316044 271696 316056
rect 270552 316016 271696 316044
rect 270552 316004 270558 316016
rect 271690 316004 271696 316016
rect 271748 316004 271754 316056
rect 252554 315936 252560 315988
rect 252612 315976 252618 315988
rect 253382 315976 253388 315988
rect 252612 315948 253388 315976
rect 252612 315936 252618 315948
rect 253382 315936 253388 315948
rect 253440 315936 253446 315988
rect 258810 315936 258816 315988
rect 258868 315976 258874 315988
rect 259362 315976 259368 315988
rect 258868 315948 259368 315976
rect 258868 315936 258874 315948
rect 259362 315936 259368 315948
rect 259420 315936 259426 315988
rect 259454 315936 259460 315988
rect 259512 315976 259518 315988
rect 260006 315976 260012 315988
rect 259512 315948 260012 315976
rect 259512 315936 259518 315948
rect 260006 315936 260012 315948
rect 260064 315936 260070 315988
rect 261294 315936 261300 315988
rect 261352 315976 261358 315988
rect 262122 315976 262128 315988
rect 261352 315948 262128 315976
rect 261352 315936 261358 315948
rect 262122 315936 262128 315948
rect 262180 315936 262186 315988
rect 262306 315936 262312 315988
rect 262364 315976 262370 315988
rect 262364 315948 262444 315976
rect 262364 315936 262370 315948
rect 157794 315868 157800 315920
rect 157852 315908 157858 315920
rect 158438 315908 158444 315920
rect 157852 315880 158444 315908
rect 157852 315868 157858 315880
rect 158438 315868 158444 315880
rect 158496 315868 158502 315920
rect 244090 315868 244096 315920
rect 244148 315868 244154 315920
rect 262416 315784 262444 315948
rect 265250 315936 265256 315988
rect 265308 315976 265314 315988
rect 266078 315976 266084 315988
rect 265308 315948 266084 315976
rect 265308 315936 265314 315948
rect 266078 315936 266084 315948
rect 266136 315936 266142 315988
rect 271230 315936 271236 315988
rect 271288 315976 271294 315988
rect 271782 315976 271788 315988
rect 271288 315948 271788 315976
rect 271288 315936 271294 315948
rect 271782 315936 271788 315948
rect 271840 315936 271846 315988
rect 266446 315868 266452 315920
rect 266504 315908 266510 315920
rect 267550 315908 267556 315920
rect 266504 315880 267556 315908
rect 266504 315868 266510 315880
rect 267550 315868 267556 315880
rect 267608 315868 267614 315920
rect 262398 315732 262404 315784
rect 262456 315732 262462 315784
rect 230566 315324 230572 315376
rect 230624 315364 230630 315376
rect 231486 315364 231492 315376
rect 230624 315336 231492 315364
rect 230624 315324 230630 315336
rect 231486 315324 231492 315336
rect 231544 315324 231550 315376
rect 73246 315256 73252 315308
rect 73304 315296 73310 315308
rect 73614 315296 73620 315308
rect 73304 315268 73620 315296
rect 73304 315256 73310 315268
rect 73614 315256 73620 315268
rect 73672 315256 73678 315308
rect 246482 315188 246488 315240
rect 246540 315228 246546 315240
rect 246942 315228 246948 315240
rect 246540 315200 246948 315228
rect 246540 315188 246546 315200
rect 246942 315188 246948 315200
rect 247000 315188 247006 315240
rect 255314 314984 255320 315036
rect 255372 315024 255378 315036
rect 256418 315024 256424 315036
rect 255372 314996 256424 315024
rect 255372 314984 255378 314996
rect 256418 314984 256424 314996
rect 256476 314984 256482 315036
rect 257430 314984 257436 315036
rect 257488 315024 257494 315036
rect 257890 315024 257896 315036
rect 257488 314996 257896 315024
rect 257488 314984 257494 314996
rect 257890 314984 257896 314996
rect 257948 314984 257954 315036
rect 267826 314644 267832 314696
rect 267884 314684 267890 314696
rect 268102 314684 268108 314696
rect 267884 314656 268108 314684
rect 267884 314644 267890 314656
rect 268102 314644 268108 314656
rect 268160 314644 268166 314696
rect 241606 314100 241612 314152
rect 241664 314140 241670 314152
rect 242618 314140 242624 314152
rect 241664 314112 242624 314140
rect 241664 314100 241670 314112
rect 242618 314100 242624 314112
rect 242676 314100 242682 314152
rect 250530 313896 250536 313948
rect 250588 313936 250594 313948
rect 250990 313936 250996 313948
rect 250588 313908 250996 313936
rect 250588 313896 250594 313908
rect 250990 313896 250996 313908
rect 251048 313896 251054 313948
rect 264146 313896 264152 313948
rect 264204 313936 264210 313948
rect 264698 313936 264704 313948
rect 264204 313908 264704 313936
rect 264204 313896 264210 313908
rect 264698 313896 264704 313908
rect 264756 313896 264762 313948
rect 262306 312740 262312 312792
rect 262364 312780 262370 312792
rect 262766 312780 262772 312792
rect 262364 312752 262772 312780
rect 262364 312740 262370 312752
rect 262766 312740 262772 312752
rect 262824 312740 262830 312792
rect 262214 312672 262220 312724
rect 262272 312712 262278 312724
rect 262490 312712 262496 312724
rect 262272 312684 262496 312712
rect 262272 312672 262278 312684
rect 262490 312672 262496 312684
rect 262548 312672 262554 312724
rect 150894 312604 150900 312656
rect 150952 312644 150958 312656
rect 151170 312644 151176 312656
rect 150952 312616 151176 312644
rect 150952 312604 150958 312616
rect 151170 312604 151176 312616
rect 151228 312604 151234 312656
rect 105078 311924 105084 311976
rect 105136 311924 105142 311976
rect 105096 311760 105124 311924
rect 233326 311788 233332 311840
rect 233384 311828 233390 311840
rect 234338 311828 234344 311840
rect 233384 311800 234344 311828
rect 233384 311788 233390 311800
rect 234338 311788 234344 311800
rect 234396 311788 234402 311840
rect 105170 311760 105176 311772
rect 105096 311732 105176 311760
rect 105170 311720 105176 311732
rect 105228 311720 105234 311772
rect 248506 311584 248512 311636
rect 248564 311624 248570 311636
rect 249426 311624 249432 311636
rect 248564 311596 249432 311624
rect 248564 311584 248570 311596
rect 249426 311584 249432 311596
rect 249484 311584 249490 311636
rect 249886 311584 249892 311636
rect 249944 311624 249950 311636
rect 250622 311624 250628 311636
rect 249944 311596 250628 311624
rect 249944 311584 249950 311596
rect 250622 311584 250628 311596
rect 250680 311584 250686 311636
rect 223666 311176 223672 311228
rect 223724 311216 223730 311228
rect 224862 311216 224868 311228
rect 223724 311188 224868 311216
rect 223724 311176 223730 311188
rect 224862 311176 224868 311188
rect 224920 311176 224926 311228
rect 247218 309748 247224 309800
rect 247276 309788 247282 309800
rect 248322 309788 248328 309800
rect 247276 309760 248328 309788
rect 247276 309748 247282 309760
rect 248322 309748 248328 309760
rect 248380 309748 248386 309800
rect 251269 309587 251327 309593
rect 251269 309553 251281 309587
rect 251315 309584 251327 309587
rect 251726 309584 251732 309596
rect 251315 309556 251732 309584
rect 251315 309553 251327 309556
rect 251269 309547 251327 309553
rect 251726 309544 251732 309556
rect 251784 309544 251790 309596
rect 77570 309272 77576 309324
rect 77628 309272 77634 309324
rect 77588 309188 77616 309272
rect 193861 309247 193919 309253
rect 193861 309213 193873 309247
rect 193907 309244 193919 309247
rect 193950 309244 193956 309256
rect 193907 309216 193956 309244
rect 193907 309213 193919 309216
rect 193861 309207 193919 309213
rect 193950 309204 193956 309216
rect 194008 309204 194014 309256
rect 70854 309176 70860 309188
rect 70815 309148 70860 309176
rect 70854 309136 70860 309148
rect 70912 309136 70918 309188
rect 77570 309136 77576 309188
rect 77628 309136 77634 309188
rect 78950 309136 78956 309188
rect 79008 309176 79014 309188
rect 79410 309176 79416 309188
rect 79008 309148 79416 309176
rect 79008 309136 79014 309148
rect 79410 309136 79416 309148
rect 79468 309136 79474 309188
rect 84654 309136 84660 309188
rect 84712 309176 84718 309188
rect 85114 309176 85120 309188
rect 84712 309148 85120 309176
rect 84712 309136 84718 309148
rect 85114 309136 85120 309148
rect 85172 309136 85178 309188
rect 147309 309179 147367 309185
rect 147309 309145 147321 309179
rect 147355 309176 147367 309179
rect 151078 309176 151084 309188
rect 147355 309148 151084 309176
rect 147355 309145 147367 309148
rect 147309 309139 147367 309145
rect 151078 309136 151084 309148
rect 151136 309136 151142 309188
rect 162118 309176 162124 309188
rect 162079 309148 162124 309176
rect 162118 309136 162124 309148
rect 162176 309136 162182 309188
rect 197998 309176 198004 309188
rect 197959 309148 198004 309176
rect 197998 309136 198004 309148
rect 198056 309136 198062 309188
rect 204898 309176 204904 309188
rect 204859 309148 204904 309176
rect 204898 309136 204904 309148
rect 204956 309136 204962 309188
rect 251266 309136 251272 309188
rect 251324 309176 251330 309188
rect 251450 309176 251456 309188
rect 251324 309148 251456 309176
rect 251324 309136 251330 309148
rect 251450 309136 251456 309148
rect 251508 309136 251514 309188
rect 259178 309136 259184 309188
rect 259236 309176 259242 309188
rect 259270 309176 259276 309188
rect 259236 309148 259276 309176
rect 259236 309136 259242 309148
rect 259270 309136 259276 309148
rect 259328 309136 259334 309188
rect 270770 309136 270776 309188
rect 270828 309176 270834 309188
rect 271506 309176 271512 309188
rect 270828 309148 271512 309176
rect 270828 309136 270834 309148
rect 271506 309136 271512 309148
rect 271564 309136 271570 309188
rect 245562 309108 245568 309120
rect 245523 309080 245568 309108
rect 245562 309068 245568 309080
rect 245620 309068 245626 309120
rect 254026 309108 254032 309120
rect 253987 309080 254032 309108
rect 254026 309068 254032 309080
rect 254084 309068 254090 309120
rect 264698 309068 264704 309120
rect 264756 309068 264762 309120
rect 324961 309111 325019 309117
rect 324961 309077 324973 309111
rect 325007 309108 325019 309111
rect 325050 309108 325056 309120
rect 325007 309080 325056 309108
rect 325007 309077 325019 309080
rect 324961 309071 325019 309077
rect 325050 309068 325056 309080
rect 325108 309068 325114 309120
rect 264716 309040 264744 309068
rect 264790 309040 264796 309052
rect 264716 309012 264796 309040
rect 264790 309000 264796 309012
rect 264848 309000 264854 309052
rect 94038 307884 94044 307896
rect 93999 307856 94044 307884
rect 94038 307844 94044 307856
rect 94096 307844 94102 307896
rect 70854 307816 70860 307828
rect 70815 307788 70860 307816
rect 70854 307776 70860 307788
rect 70912 307776 70918 307828
rect 73522 307776 73528 307828
rect 73580 307816 73586 307828
rect 73614 307816 73620 307828
rect 73580 307788 73620 307816
rect 73580 307776 73586 307788
rect 73614 307776 73620 307788
rect 73672 307776 73678 307828
rect 92842 307816 92848 307828
rect 92803 307788 92848 307816
rect 92842 307776 92848 307788
rect 92900 307776 92906 307828
rect 193858 307816 193864 307828
rect 193819 307788 193864 307816
rect 193858 307776 193864 307788
rect 193916 307776 193922 307828
rect 236178 307816 236184 307828
rect 236139 307788 236184 307816
rect 236178 307776 236184 307788
rect 236236 307776 236242 307828
rect 238938 307816 238944 307828
rect 238899 307788 238944 307816
rect 238938 307776 238944 307788
rect 238996 307776 239002 307828
rect 94038 307748 94044 307760
rect 93999 307720 94044 307748
rect 94038 307708 94044 307720
rect 94096 307708 94102 307760
rect 247034 307300 247040 307352
rect 247092 307340 247098 307352
rect 248138 307340 248144 307352
rect 247092 307312 248144 307340
rect 247092 307300 247098 307312
rect 248138 307300 248144 307312
rect 248196 307300 248202 307352
rect 255314 307096 255320 307148
rect 255372 307136 255378 307148
rect 256510 307136 256516 307148
rect 255372 307108 256516 307136
rect 255372 307096 255378 307108
rect 256510 307096 256516 307108
rect 256568 307096 256574 307148
rect 224954 307028 224960 307080
rect 225012 307068 225018 307080
rect 226150 307068 226156 307080
rect 225012 307040 226156 307068
rect 225012 307028 225018 307040
rect 226150 307028 226156 307040
rect 226208 307028 226214 307080
rect 230566 307028 230572 307080
rect 230624 307068 230630 307080
rect 231578 307068 231584 307080
rect 230624 307040 231584 307068
rect 230624 307028 230630 307040
rect 231578 307028 231584 307040
rect 231636 307028 231642 307080
rect 231854 307028 231860 307080
rect 231912 307068 231918 307080
rect 233050 307068 233056 307080
rect 231912 307040 233056 307068
rect 231912 307028 231918 307040
rect 233050 307028 233056 307040
rect 233108 307028 233114 307080
rect 233234 307028 233240 307080
rect 233292 307068 233298 307080
rect 234522 307068 234528 307080
rect 233292 307040 234528 307068
rect 233292 307028 233298 307040
rect 234522 307028 234528 307040
rect 234580 307028 234586 307080
rect 234614 307028 234620 307080
rect 234672 307068 234678 307080
rect 235810 307068 235816 307080
rect 234672 307040 235816 307068
rect 234672 307028 234678 307040
rect 235810 307028 235816 307040
rect 235868 307028 235874 307080
rect 235994 307028 236000 307080
rect 236052 307068 236058 307080
rect 237282 307068 237288 307080
rect 236052 307040 237288 307068
rect 236052 307028 236058 307040
rect 237282 307028 237288 307040
rect 237340 307028 237346 307080
rect 237374 307028 237380 307080
rect 237432 307068 237438 307080
rect 238662 307068 238668 307080
rect 237432 307040 238668 307068
rect 237432 307028 237438 307040
rect 238662 307028 238668 307040
rect 238720 307028 238726 307080
rect 238846 307028 238852 307080
rect 238904 307068 238910 307080
rect 239858 307068 239864 307080
rect 238904 307040 239864 307068
rect 238904 307028 238910 307040
rect 239858 307028 239864 307040
rect 239916 307028 239922 307080
rect 240134 307028 240140 307080
rect 240192 307068 240198 307080
rect 241422 307068 241428 307080
rect 240192 307040 241428 307068
rect 240192 307028 240198 307040
rect 241422 307028 241428 307040
rect 241480 307028 241486 307080
rect 241514 307028 241520 307080
rect 241572 307068 241578 307080
rect 242802 307068 242808 307080
rect 241572 307040 242808 307068
rect 241572 307028 241578 307040
rect 242802 307028 242808 307040
rect 242860 307028 242866 307080
rect 244274 307028 244280 307080
rect 244332 307068 244338 307080
rect 245470 307068 245476 307080
rect 244332 307040 245476 307068
rect 244332 307028 244338 307040
rect 245470 307028 245476 307040
rect 245528 307028 245534 307080
rect 245654 307028 245660 307080
rect 245712 307068 245718 307080
rect 246850 307068 246856 307080
rect 245712 307040 246856 307068
rect 245712 307028 245718 307040
rect 246850 307028 246856 307040
rect 246908 307028 246914 307080
rect 248414 307028 248420 307080
rect 248472 307068 248478 307080
rect 249702 307068 249708 307080
rect 248472 307040 249708 307068
rect 248472 307028 248478 307040
rect 249702 307028 249708 307040
rect 249760 307028 249766 307080
rect 249794 307028 249800 307080
rect 249852 307068 249858 307080
rect 251082 307068 251088 307080
rect 249852 307040 251088 307068
rect 249852 307028 249858 307040
rect 251082 307028 251088 307040
rect 251140 307028 251146 307080
rect 252554 307028 252560 307080
rect 252612 307068 252618 307080
rect 253842 307068 253848 307080
rect 252612 307040 253848 307068
rect 252612 307028 252618 307040
rect 253842 307028 253848 307040
rect 253900 307028 253906 307080
rect 253934 307028 253940 307080
rect 253992 307068 253998 307080
rect 255130 307068 255136 307080
rect 253992 307040 255136 307068
rect 253992 307028 253998 307040
rect 255130 307028 255136 307040
rect 255188 307028 255194 307080
rect 255406 307028 255412 307080
rect 255464 307068 255470 307080
rect 256418 307068 256424 307080
rect 255464 307040 256424 307068
rect 255464 307028 255470 307040
rect 256418 307028 256424 307040
rect 256476 307028 256482 307080
rect 256694 307028 256700 307080
rect 256752 307068 256758 307080
rect 257982 307068 257988 307080
rect 256752 307040 257988 307068
rect 256752 307028 256758 307040
rect 257982 307028 257988 307040
rect 258040 307028 258046 307080
rect 259638 307028 259644 307080
rect 259696 307068 259702 307080
rect 260742 307068 260748 307080
rect 259696 307040 260748 307068
rect 259696 307028 259702 307040
rect 260742 307028 260748 307040
rect 260800 307028 260806 307080
rect 262214 307028 262220 307080
rect 262272 307068 262278 307080
rect 263318 307068 263324 307080
rect 262272 307040 263324 307068
rect 262272 307028 262278 307040
rect 263318 307028 263324 307040
rect 263376 307028 263382 307080
rect 267734 307028 267740 307080
rect 267792 307068 267798 307080
rect 268930 307068 268936 307080
rect 267792 307040 268936 307068
rect 267792 307028 267798 307040
rect 268930 307028 268936 307040
rect 268988 307028 268994 307080
rect 270494 307028 270500 307080
rect 270552 307068 270558 307080
rect 271598 307068 271604 307080
rect 270552 307040 271604 307068
rect 270552 307028 270558 307040
rect 271598 307028 271604 307040
rect 271656 307028 271662 307080
rect 230750 306960 230756 307012
rect 230808 307000 230814 307012
rect 231762 307000 231768 307012
rect 230808 306972 231768 307000
rect 230808 306960 230814 306972
rect 231762 306960 231768 306972
rect 231820 306960 231826 307012
rect 238754 306960 238760 307012
rect 238812 307000 238818 307012
rect 240042 307000 240048 307012
rect 238812 306972 240048 307000
rect 238812 306960 238818 306972
rect 240042 306960 240048 306972
rect 240100 306960 240106 307012
rect 255498 306960 255504 307012
rect 255556 307000 255562 307012
rect 256602 307000 256608 307012
rect 255556 306972 256608 307000
rect 255556 306960 255562 306972
rect 256602 306960 256608 306972
rect 256660 306960 256666 307012
rect 259454 306960 259460 307012
rect 259512 307000 259518 307012
rect 260650 307000 260656 307012
rect 259512 306972 260656 307000
rect 259512 306960 259518 306972
rect 260650 306960 260656 306972
rect 260708 306960 260714 307012
rect 262398 306960 262404 307012
rect 262456 307000 262462 307012
rect 263502 307000 263508 307012
rect 262456 306972 263508 307000
rect 262456 306960 262462 306972
rect 263502 306960 263508 306972
rect 263560 306960 263566 307012
rect 266446 306960 266452 307012
rect 266504 307000 266510 307012
rect 267550 307000 267556 307012
rect 266504 306972 267556 307000
rect 266504 306960 266510 306972
rect 267550 306960 267556 306972
rect 267608 306960 267614 307012
rect 251266 306932 251272 306944
rect 251227 306904 251272 306932
rect 251266 306892 251272 306904
rect 251324 306892 251330 306944
rect 242894 306824 242900 306876
rect 242952 306864 242958 306876
rect 243906 306864 243912 306876
rect 242952 306836 243912 306864
rect 242952 306824 242958 306836
rect 243906 306824 243912 306836
rect 243964 306824 243970 306876
rect 236178 306688 236184 306740
rect 236236 306728 236242 306740
rect 237098 306728 237104 306740
rect 236236 306700 237104 306728
rect 236236 306688 236242 306700
rect 237098 306688 237104 306700
rect 237156 306688 237162 306740
rect 266538 306348 266544 306400
rect 266596 306388 266602 306400
rect 267090 306388 267096 306400
rect 266596 306360 267096 306388
rect 266596 306348 266602 306360
rect 267090 306348 267096 306360
rect 267148 306348 267154 306400
rect 262306 306008 262312 306060
rect 262364 306048 262370 306060
rect 263226 306048 263232 306060
rect 262364 306020 263232 306048
rect 262364 306008 262370 306020
rect 263226 306008 263232 306020
rect 263284 306008 263290 306060
rect 269114 305736 269120 305788
rect 269172 305776 269178 305788
rect 270218 305776 270224 305788
rect 269172 305748 270224 305776
rect 269172 305736 269178 305748
rect 270218 305736 270224 305748
rect 270276 305736 270282 305788
rect 267090 303600 267096 303612
rect 267051 303572 267096 303600
rect 267090 303560 267096 303572
rect 267148 303560 267154 303612
rect 70578 302308 70584 302320
rect 70504 302280 70584 302308
rect 70504 302184 70532 302280
rect 70578 302268 70584 302280
rect 70636 302268 70642 302320
rect 233418 302268 233424 302320
rect 233476 302268 233482 302320
rect 259178 302268 259184 302320
rect 259236 302268 259242 302320
rect 105081 302243 105139 302249
rect 105081 302209 105093 302243
rect 105127 302240 105139 302243
rect 105170 302240 105176 302252
rect 105127 302212 105176 302240
rect 105127 302209 105139 302212
rect 105081 302203 105139 302209
rect 105170 302200 105176 302212
rect 105228 302200 105234 302252
rect 106550 302200 106556 302252
rect 106608 302240 106614 302252
rect 106734 302240 106740 302252
rect 106608 302212 106740 302240
rect 106608 302200 106614 302212
rect 106734 302200 106740 302212
rect 106792 302200 106798 302252
rect 211798 302200 211804 302252
rect 211856 302240 211862 302252
rect 211982 302240 211988 302252
rect 211856 302212 211988 302240
rect 211856 302200 211862 302212
rect 211982 302200 211988 302212
rect 212040 302200 212046 302252
rect 232038 302200 232044 302252
rect 232096 302240 232102 302252
rect 233142 302240 233148 302252
rect 232096 302212 233148 302240
rect 232096 302200 232102 302212
rect 233142 302200 233148 302212
rect 233200 302200 233206 302252
rect 233436 302240 233464 302268
rect 234430 302240 234436 302252
rect 233436 302212 234436 302240
rect 234430 302200 234436 302212
rect 234488 302200 234494 302252
rect 238938 302200 238944 302252
rect 238996 302200 239002 302252
rect 70486 302132 70492 302184
rect 70544 302132 70550 302184
rect 237466 302132 237472 302184
rect 237524 302172 237530 302184
rect 238386 302172 238392 302184
rect 237524 302144 238392 302172
rect 237524 302132 237530 302144
rect 238386 302132 238392 302144
rect 238444 302132 238450 302184
rect 238956 302172 238984 302200
rect 259196 302184 259224 302268
rect 239766 302172 239772 302184
rect 238956 302144 239772 302172
rect 239766 302132 239772 302144
rect 239824 302132 239830 302184
rect 259178 302132 259184 302184
rect 259236 302132 259242 302184
rect 265802 302172 265808 302184
rect 265763 302144 265808 302172
rect 265802 302132 265808 302144
rect 265860 302132 265866 302184
rect 259546 302064 259552 302116
rect 259604 302104 259610 302116
rect 260466 302104 260472 302116
rect 259604 302076 260472 302104
rect 259604 302064 259610 302076
rect 260466 302064 260472 302076
rect 260524 302064 260530 302116
rect 92842 299548 92848 299600
rect 92900 299548 92906 299600
rect 70670 299480 70676 299532
rect 70728 299520 70734 299532
rect 70854 299520 70860 299532
rect 70728 299492 70860 299520
rect 70728 299480 70734 299492
rect 70854 299480 70860 299492
rect 70912 299480 70918 299532
rect 92860 299464 92888 299548
rect 234246 299480 234252 299532
rect 234304 299520 234310 299532
rect 234338 299520 234344 299532
rect 234304 299492 234344 299520
rect 234304 299480 234310 299492
rect 234338 299480 234344 299492
rect 234396 299480 234402 299532
rect 245562 299520 245568 299532
rect 245523 299492 245568 299520
rect 245562 299480 245568 299492
rect 245620 299480 245626 299532
rect 250806 299480 250812 299532
rect 250864 299520 250870 299532
rect 250990 299520 250996 299532
rect 250864 299492 250996 299520
rect 250864 299480 250870 299492
rect 250990 299480 250996 299492
rect 251048 299480 251054 299532
rect 254029 299523 254087 299529
rect 254029 299489 254041 299523
rect 254075 299520 254087 299523
rect 255038 299520 255044 299532
rect 254075 299492 255044 299520
rect 254075 299489 254087 299492
rect 254029 299483 254087 299489
rect 255038 299480 255044 299492
rect 255096 299480 255102 299532
rect 255222 299520 255228 299532
rect 255183 299492 255228 299520
rect 255222 299480 255228 299492
rect 255280 299480 255286 299532
rect 266078 299480 266084 299532
rect 266136 299520 266142 299532
rect 266170 299520 266176 299532
rect 266136 299492 266176 299520
rect 266136 299480 266142 299492
rect 266170 299480 266176 299492
rect 266228 299480 266234 299532
rect 267826 299480 267832 299532
rect 267884 299520 267890 299532
rect 268746 299520 268752 299532
rect 267884 299492 268752 299520
rect 267884 299480 267890 299492
rect 268746 299480 268752 299492
rect 268804 299480 268810 299532
rect 324958 299520 324964 299532
rect 324919 299492 324964 299520
rect 324958 299480 324964 299492
rect 325016 299480 325022 299532
rect 70486 299452 70492 299464
rect 70447 299424 70492 299452
rect 70486 299412 70492 299424
rect 70544 299412 70550 299464
rect 73430 299412 73436 299464
rect 73488 299452 73494 299464
rect 73522 299452 73528 299464
rect 73488 299424 73528 299452
rect 73488 299412 73494 299424
rect 73522 299412 73528 299424
rect 73580 299412 73586 299464
rect 92842 299412 92848 299464
rect 92900 299412 92906 299464
rect 151078 299452 151084 299464
rect 151039 299424 151084 299452
rect 151078 299412 151084 299424
rect 151136 299412 151142 299464
rect 227346 299452 227352 299464
rect 227307 299424 227352 299452
rect 227346 299412 227352 299424
rect 227404 299412 227410 299464
rect 251266 299452 251272 299464
rect 251227 299424 251272 299452
rect 251266 299412 251272 299424
rect 251324 299412 251330 299464
rect 267090 299452 267096 299464
rect 267051 299424 267096 299452
rect 267090 299412 267096 299424
rect 267148 299412 267154 299464
rect 271506 299452 271512 299464
rect 271467 299424 271512 299452
rect 271506 299412 271512 299424
rect 271564 299412 271570 299464
rect 89990 298188 89996 298240
rect 90048 298228 90054 298240
rect 90174 298228 90180 298240
rect 90048 298200 90180 298228
rect 90048 298188 90054 298200
rect 90174 298188 90180 298200
rect 90232 298188 90238 298240
rect 94038 298160 94044 298172
rect 93999 298132 94044 298160
rect 94038 298120 94044 298132
rect 94096 298120 94102 298172
rect 105078 298160 105084 298172
rect 105039 298132 105084 298160
rect 105078 298120 105084 298132
rect 105136 298120 105142 298172
rect 255222 298160 255228 298172
rect 255183 298132 255228 298160
rect 255222 298120 255228 298132
rect 255280 298120 255286 298172
rect 70762 298092 70768 298104
rect 70723 298064 70768 298092
rect 70762 298052 70768 298064
rect 70820 298052 70826 298104
rect 73430 298052 73436 298104
rect 73488 298092 73494 298104
rect 73522 298092 73528 298104
rect 73488 298064 73528 298092
rect 73488 298052 73494 298064
rect 73522 298052 73528 298064
rect 73580 298052 73586 298104
rect 193858 298092 193864 298104
rect 193819 298064 193864 298092
rect 193858 298052 193864 298064
rect 193916 298052 193922 298104
rect 242618 298092 242624 298104
rect 242579 298064 242624 298092
rect 242618 298052 242624 298064
rect 242676 298052 242682 298104
rect 243906 298092 243912 298104
rect 243867 298064 243912 298092
rect 243906 298052 243912 298064
rect 243964 298052 243970 298104
rect 246942 298092 246948 298104
rect 246903 298064 246948 298092
rect 246942 298052 246948 298064
rect 247000 298052 247006 298104
rect 248230 298092 248236 298104
rect 248191 298064 248236 298092
rect 248230 298052 248236 298064
rect 248288 298052 248294 298104
rect 255222 298024 255228 298036
rect 255183 297996 255228 298024
rect 255222 297984 255228 297996
rect 255280 297984 255286 298036
rect 259178 297440 259184 297492
rect 259236 297480 259242 297492
rect 259273 297483 259331 297489
rect 259273 297480 259285 297483
rect 259236 297452 259285 297480
rect 259236 297440 259242 297452
rect 259273 297449 259285 297452
rect 259319 297449 259331 297483
rect 259273 297443 259331 297449
rect 268838 297372 268844 297424
rect 268896 297412 268902 297424
rect 269022 297412 269028 297424
rect 268896 297384 269028 297412
rect 268896 297372 268902 297384
rect 269022 297372 269028 297384
rect 269080 297372 269086 297424
rect 251269 297279 251327 297285
rect 251269 297245 251281 297279
rect 251315 297276 251327 297279
rect 252186 297276 252192 297288
rect 251315 297248 252192 297276
rect 251315 297245 251327 297248
rect 251269 297239 251327 297245
rect 252186 297236 252192 297248
rect 252244 297236 252250 297288
rect 234890 296760 234896 296812
rect 234948 296800 234954 296812
rect 235718 296800 235724 296812
rect 234948 296772 235724 296800
rect 234948 296760 234954 296772
rect 235718 296760 235724 296772
rect 235776 296760 235782 296812
rect 72142 296664 72148 296676
rect 72103 296636 72148 296664
rect 72142 296624 72148 296636
rect 72200 296624 72206 296676
rect 235718 296664 235724 296676
rect 235679 296636 235724 296664
rect 235718 296624 235724 296636
rect 235776 296624 235782 296676
rect 244366 296284 244372 296336
rect 244424 296324 244430 296336
rect 245378 296324 245384 296336
rect 244424 296296 245384 296324
rect 244424 296284 244430 296296
rect 245378 296284 245384 296296
rect 245436 296284 245442 296336
rect 249886 296284 249892 296336
rect 249944 296324 249950 296336
rect 250898 296324 250904 296336
rect 249944 296296 250904 296324
rect 249944 296284 249950 296296
rect 250898 296284 250904 296296
rect 250956 296284 250962 296336
rect 245746 294584 245752 294636
rect 245804 294624 245810 294636
rect 246758 294624 246764 294636
rect 245804 294596 246764 294624
rect 245804 294584 245810 294596
rect 246758 294584 246764 294596
rect 246816 294584 246822 294636
rect 247218 294584 247224 294636
rect 247276 294624 247282 294636
rect 248046 294624 248052 294636
rect 247276 294596 248052 294624
rect 247276 294584 247282 294596
rect 248046 294584 248052 294596
rect 248104 294584 248110 294636
rect 248506 294584 248512 294636
rect 248564 294624 248570 294636
rect 249518 294624 249524 294636
rect 248564 294596 249524 294624
rect 248564 294584 248570 294596
rect 249518 294584 249524 294596
rect 249576 294584 249582 294636
rect 252738 294584 252744 294636
rect 252796 294624 252802 294636
rect 253658 294624 253664 294636
rect 252796 294596 253664 294624
rect 252796 294584 252802 294596
rect 253658 294584 253664 294596
rect 253716 294584 253722 294636
rect 271506 293536 271512 293548
rect 271467 293508 271512 293536
rect 271506 293496 271512 293508
rect 271564 293496 271570 293548
rect 265805 292655 265863 292661
rect 265805 292621 265817 292655
rect 265851 292652 265863 292655
rect 265894 292652 265900 292664
rect 265851 292624 265900 292652
rect 265851 292621 265863 292624
rect 265805 292615 265863 292621
rect 265894 292612 265900 292624
rect 265952 292612 265958 292664
rect 265894 292476 265900 292528
rect 265952 292476 265958 292528
rect 105170 292408 105176 292460
rect 105228 292448 105234 292460
rect 105354 292448 105360 292460
rect 105228 292420 105360 292448
rect 105228 292408 105234 292420
rect 105354 292408 105360 292420
rect 105412 292408 105418 292460
rect 265912 292448 265940 292476
rect 265986 292448 265992 292460
rect 265912 292420 265992 292448
rect 265986 292408 265992 292420
rect 266044 292408 266050 292460
rect 78950 289932 78956 289944
rect 78876 289904 78956 289932
rect 78876 289876 78904 289904
rect 78950 289892 78956 289904
rect 79008 289892 79014 289944
rect 70489 289867 70547 289873
rect 70489 289833 70501 289867
rect 70535 289864 70547 289867
rect 70578 289864 70584 289876
rect 70535 289836 70584 289864
rect 70535 289833 70547 289836
rect 70489 289827 70547 289833
rect 70578 289824 70584 289836
rect 70636 289824 70642 289876
rect 77570 289824 77576 289876
rect 77628 289864 77634 289876
rect 77662 289864 77668 289876
rect 77628 289836 77668 289864
rect 77628 289824 77634 289836
rect 77662 289824 77668 289836
rect 77720 289824 77726 289876
rect 78858 289824 78864 289876
rect 78916 289824 78922 289876
rect 81710 289824 81716 289876
rect 81768 289864 81774 289876
rect 81802 289864 81808 289876
rect 81768 289836 81808 289864
rect 81768 289824 81774 289836
rect 81802 289824 81808 289836
rect 81860 289824 81866 289876
rect 151078 289864 151084 289876
rect 151039 289836 151084 289864
rect 151078 289824 151084 289836
rect 151136 289824 151142 289876
rect 227349 289867 227407 289873
rect 227349 289833 227361 289867
rect 227395 289864 227407 289867
rect 227438 289864 227444 289876
rect 227395 289836 227444 289864
rect 227395 289833 227407 289836
rect 227349 289827 227407 289833
rect 227438 289824 227444 289836
rect 227496 289824 227502 289876
rect 249426 289824 249432 289876
rect 249484 289864 249490 289876
rect 249610 289864 249616 289876
rect 249484 289836 249616 289864
rect 249484 289824 249490 289836
rect 249610 289824 249616 289836
rect 249668 289824 249674 289876
rect 250806 289824 250812 289876
rect 250864 289864 250870 289876
rect 250990 289864 250996 289876
rect 250864 289836 250996 289864
rect 250864 289824 250870 289836
rect 250990 289824 250996 289836
rect 251048 289824 251054 289876
rect 259270 289864 259276 289876
rect 259231 289836 259276 289864
rect 259270 289824 259276 289836
rect 259328 289824 259334 289876
rect 324961 289799 325019 289805
rect 324961 289765 324973 289799
rect 325007 289796 325019 289799
rect 325050 289796 325056 289808
rect 325007 289768 325056 289796
rect 325007 289765 325019 289768
rect 324961 289759 325019 289765
rect 325050 289756 325056 289768
rect 325108 289756 325114 289808
rect 70762 288436 70768 288448
rect 70723 288408 70768 288436
rect 70762 288396 70768 288408
rect 70820 288396 70826 288448
rect 94038 288396 94044 288448
rect 94096 288436 94102 288448
rect 94130 288436 94136 288448
rect 94096 288408 94136 288436
rect 94096 288396 94102 288408
rect 94130 288396 94136 288408
rect 94188 288396 94194 288448
rect 193858 288436 193864 288448
rect 193819 288408 193864 288436
rect 193858 288396 193864 288408
rect 193916 288396 193922 288448
rect 242618 288436 242624 288448
rect 242579 288408 242624 288436
rect 242618 288396 242624 288408
rect 242676 288396 242682 288448
rect 243814 288396 243820 288448
rect 243872 288436 243878 288448
rect 243909 288439 243967 288445
rect 243909 288436 243921 288439
rect 243872 288408 243921 288436
rect 243872 288396 243878 288408
rect 243909 288405 243921 288408
rect 243955 288405 243967 288439
rect 246942 288436 246948 288448
rect 246903 288408 246948 288436
rect 243909 288399 243967 288405
rect 246942 288396 246948 288408
rect 247000 288396 247006 288448
rect 248230 288436 248236 288448
rect 248191 288408 248236 288436
rect 248230 288396 248236 288408
rect 248288 288396 248294 288448
rect 255222 288436 255228 288448
rect 255183 288408 255228 288436
rect 255222 288396 255228 288408
rect 255280 288396 255286 288448
rect 72145 288371 72203 288377
rect 72145 288337 72157 288371
rect 72191 288368 72203 288371
rect 72326 288368 72332 288380
rect 72191 288340 72332 288368
rect 72191 288337 72203 288340
rect 72145 288331 72203 288337
rect 72326 288328 72332 288340
rect 72384 288328 72390 288380
rect 267182 287756 267188 287768
rect 267143 287728 267188 287756
rect 267182 287716 267188 287728
rect 267240 287716 267246 287768
rect 268838 287716 268844 287768
rect 268896 287756 268902 287768
rect 269022 287756 269028 287768
rect 268896 287728 269028 287756
rect 268896 287716 268902 287728
rect 269022 287716 269028 287728
rect 269080 287716 269086 287768
rect 235718 287144 235724 287156
rect 235679 287116 235724 287144
rect 235718 287104 235724 287116
rect 235776 287104 235782 287156
rect 90082 287036 90088 287088
rect 90140 287076 90146 287088
rect 90266 287076 90272 287088
rect 90140 287048 90272 287076
rect 90140 287036 90146 287048
rect 90266 287036 90272 287048
rect 90324 287036 90330 287088
rect 233970 287036 233976 287088
rect 234028 287076 234034 287088
rect 234062 287076 234068 287088
rect 234028 287048 234068 287076
rect 234028 287036 234034 287048
rect 234062 287036 234068 287048
rect 234120 287036 234126 287088
rect 264514 284248 264520 284300
rect 264572 284288 264578 284300
rect 264698 284288 264704 284300
rect 264572 284260 264704 284288
rect 264572 284248 264578 284260
rect 264698 284248 264704 284260
rect 264756 284248 264762 284300
rect 77570 282996 77576 283008
rect 77496 282968 77576 282996
rect 70762 282888 70768 282940
rect 70820 282888 70826 282940
rect 70780 282860 70808 282888
rect 77496 282872 77524 282968
rect 77570 282956 77576 282968
rect 77628 282956 77634 283008
rect 105170 282956 105176 283008
rect 105228 282956 105234 283008
rect 78766 282888 78772 282940
rect 78824 282928 78830 282940
rect 78861 282931 78919 282937
rect 78861 282928 78873 282931
rect 78824 282900 78873 282928
rect 78824 282888 78830 282900
rect 78861 282897 78873 282900
rect 78907 282897 78919 282931
rect 78861 282891 78919 282897
rect 70854 282860 70860 282872
rect 70780 282832 70860 282860
rect 70854 282820 70860 282832
rect 70912 282820 70918 282872
rect 77478 282820 77484 282872
rect 77536 282820 77542 282872
rect 105188 282804 105216 282956
rect 106550 282888 106556 282940
rect 106608 282928 106614 282940
rect 106734 282928 106740 282940
rect 106608 282900 106740 282928
rect 106608 282888 106614 282900
rect 106734 282888 106740 282900
rect 106792 282888 106798 282940
rect 211798 282888 211804 282940
rect 211856 282928 211862 282940
rect 211982 282928 211988 282940
rect 211856 282900 211988 282928
rect 211856 282888 211862 282900
rect 211982 282888 211988 282900
rect 212040 282888 212046 282940
rect 227254 282888 227260 282940
rect 227312 282928 227318 282940
rect 227438 282928 227444 282940
rect 227312 282900 227444 282928
rect 227312 282888 227318 282900
rect 227438 282888 227444 282900
rect 227496 282888 227502 282940
rect 267185 282931 267243 282937
rect 267185 282897 267197 282931
rect 267231 282928 267243 282931
rect 267274 282928 267280 282940
rect 267231 282900 267280 282928
rect 267231 282897 267243 282900
rect 267185 282891 267243 282897
rect 267274 282888 267280 282900
rect 267332 282888 267338 282940
rect 105170 282752 105176 282804
rect 105228 282752 105234 282804
rect 324958 280208 324964 280220
rect 324919 280180 324964 280208
rect 324958 280168 324964 280180
rect 325016 280168 325022 280220
rect 105170 280140 105176 280152
rect 105131 280112 105176 280140
rect 105170 280100 105176 280112
rect 105228 280100 105234 280152
rect 106642 280140 106648 280152
rect 106603 280112 106648 280140
rect 106642 280100 106648 280112
rect 106700 280100 106706 280152
rect 151078 280140 151084 280152
rect 151039 280112 151084 280140
rect 151078 280100 151084 280112
rect 151136 280100 151142 280152
rect 73430 278808 73436 278860
rect 73488 278848 73494 278860
rect 73522 278848 73528 278860
rect 73488 278820 73528 278848
rect 73488 278808 73494 278820
rect 73522 278808 73528 278820
rect 73580 278808 73586 278860
rect 243814 278848 243820 278860
rect 243775 278820 243820 278848
rect 243814 278808 243820 278820
rect 243872 278808 243878 278860
rect 78858 278780 78864 278792
rect 78819 278752 78864 278780
rect 78858 278740 78864 278752
rect 78916 278740 78922 278792
rect 81618 278740 81624 278792
rect 81676 278780 81682 278792
rect 81676 278752 81756 278780
rect 81676 278740 81682 278752
rect 81728 278724 81756 278752
rect 81710 278672 81716 278724
rect 81768 278672 81774 278724
rect 268838 278060 268844 278112
rect 268896 278100 268902 278112
rect 269022 278100 269028 278112
rect 268896 278072 269028 278100
rect 268896 278060 268902 278072
rect 269022 278060 269028 278072
rect 269080 278060 269086 278112
rect 72326 277380 72332 277432
rect 72384 277420 72390 277432
rect 72510 277420 72516 277432
rect 72384 277392 72516 277420
rect 72384 277380 72390 277392
rect 72510 277380 72516 277392
rect 72568 277380 72574 277432
rect 94130 277380 94136 277432
rect 94188 277420 94194 277432
rect 94314 277420 94320 277432
rect 94188 277392 94320 277420
rect 94188 277380 94194 277392
rect 94314 277380 94320 277392
rect 94372 277380 94378 277432
rect 243814 277420 243820 277432
rect 243775 277392 243820 277420
rect 243814 277380 243820 277392
rect 243872 277380 243878 277432
rect 81710 275952 81716 276004
rect 81768 275992 81774 276004
rect 81894 275992 81900 276004
rect 81768 275964 81900 275992
rect 81768 275952 81774 275964
rect 81894 275952 81900 275964
rect 81952 275952 81958 276004
rect 264609 274635 264667 274641
rect 264609 274601 264621 274635
rect 264655 274632 264667 274635
rect 264698 274632 264704 274644
rect 264655 274604 264704 274632
rect 264655 274601 264667 274604
rect 264609 274595 264667 274601
rect 264698 274592 264704 274604
rect 264756 274592 264762 274644
rect 89993 273343 90051 273349
rect 89993 273309 90005 273343
rect 90039 273340 90051 273343
rect 90082 273340 90088 273352
rect 90039 273312 90088 273340
rect 90039 273309 90051 273312
rect 89993 273303 90051 273309
rect 90082 273300 90088 273312
rect 90140 273300 90146 273352
rect 106645 273275 106703 273281
rect 106645 273241 106657 273275
rect 106691 273272 106703 273275
rect 106826 273272 106832 273284
rect 106691 273244 106832 273272
rect 106691 273241 106703 273244
rect 106645 273235 106703 273241
rect 106826 273232 106832 273244
rect 106884 273232 106890 273284
rect 268654 273272 268660 273284
rect 268615 273244 268660 273272
rect 268654 273232 268660 273244
rect 268712 273232 268718 273284
rect 105170 273136 105176 273148
rect 105131 273108 105176 273136
rect 105170 273096 105176 273108
rect 105228 273096 105234 273148
rect 70762 270512 70768 270564
rect 70820 270552 70826 270564
rect 70854 270552 70860 270564
rect 70820 270524 70860 270552
rect 70820 270512 70826 270524
rect 70854 270512 70860 270524
rect 70912 270512 70918 270564
rect 151078 270552 151084 270564
rect 151039 270524 151084 270552
rect 151078 270512 151084 270524
rect 151136 270512 151142 270564
rect 77478 270444 77484 270496
rect 77536 270484 77542 270496
rect 77570 270484 77576 270496
rect 77536 270456 77576 270484
rect 77536 270444 77542 270456
rect 77570 270444 77576 270456
rect 77628 270444 77634 270496
rect 78674 270444 78680 270496
rect 78732 270484 78738 270496
rect 78858 270484 78864 270496
rect 78732 270456 78864 270484
rect 78732 270444 78738 270456
rect 78858 270444 78864 270456
rect 78916 270444 78922 270496
rect 105170 270484 105176 270496
rect 105131 270456 105176 270484
rect 105170 270444 105176 270456
rect 105228 270444 105234 270496
rect 106826 270484 106832 270496
rect 106787 270456 106832 270484
rect 106826 270444 106832 270456
rect 106884 270444 106890 270496
rect 242526 270444 242532 270496
rect 242584 270484 242590 270496
rect 242618 270484 242624 270496
rect 242584 270456 242624 270484
rect 242584 270444 242590 270456
rect 242618 270444 242624 270456
rect 242676 270444 242682 270496
rect 249610 270484 249616 270496
rect 249571 270456 249616 270484
rect 249610 270444 249616 270456
rect 249668 270444 249674 270496
rect 250990 270484 250996 270496
rect 250951 270456 250996 270484
rect 250990 270444 250996 270456
rect 251048 270444 251054 270496
rect 252278 270484 252284 270496
rect 252239 270456 252284 270484
rect 252278 270444 252284 270456
rect 252336 270444 252342 270496
rect 259270 270484 259276 270496
rect 259231 270456 259276 270484
rect 259270 270444 259276 270456
rect 259328 270444 259334 270496
rect 324961 270487 325019 270493
rect 324961 270453 324973 270487
rect 325007 270484 325019 270487
rect 325050 270484 325056 270496
rect 325007 270456 325056 270484
rect 325007 270453 325019 270456
rect 324961 270447 325019 270453
rect 325050 270444 325056 270456
rect 325108 270444 325114 270496
rect 234065 270419 234123 270425
rect 234065 270385 234077 270419
rect 234111 270416 234123 270419
rect 234154 270416 234160 270428
rect 234111 270388 234160 270416
rect 234111 270385 234123 270388
rect 234065 270379 234123 270385
rect 234154 270376 234160 270388
rect 234212 270376 234218 270428
rect 243814 269192 243820 269204
rect 243740 269164 243820 269192
rect 92750 269084 92756 269136
rect 92808 269124 92814 269136
rect 92842 269124 92848 269136
rect 92808 269096 92848 269124
rect 92808 269084 92814 269096
rect 92842 269084 92848 269096
rect 92900 269084 92906 269136
rect 193674 269084 193680 269136
rect 193732 269124 193738 269136
rect 193858 269124 193864 269136
rect 193732 269096 193864 269124
rect 193732 269084 193738 269096
rect 193858 269084 193864 269096
rect 193916 269084 193922 269136
rect 243740 269068 243768 269164
rect 243814 269152 243820 269164
rect 243872 269152 243878 269204
rect 255222 269084 255228 269136
rect 255280 269124 255286 269136
rect 255314 269124 255320 269136
rect 255280 269096 255320 269124
rect 255280 269084 255286 269096
rect 255314 269084 255320 269096
rect 255372 269084 255378 269136
rect 243722 269016 243728 269068
rect 243780 269016 243786 269068
rect 268746 268200 268752 268252
rect 268804 268240 268810 268252
rect 269022 268240 269028 268252
rect 268804 268212 269028 268240
rect 268804 268200 268810 268212
rect 269022 268200 269028 268212
rect 269080 268200 269086 268252
rect 72418 267724 72424 267776
rect 72476 267764 72482 267776
rect 72602 267764 72608 267776
rect 72476 267736 72608 267764
rect 72476 267724 72482 267736
rect 72602 267724 72608 267736
rect 72660 267724 72666 267776
rect 73430 267724 73436 267776
rect 73488 267764 73494 267776
rect 73614 267764 73620 267776
rect 73488 267736 73620 267764
rect 73488 267724 73494 267736
rect 73614 267724 73620 267736
rect 73672 267724 73678 267776
rect 89990 267764 89996 267776
rect 89951 267736 89996 267764
rect 89990 267724 89996 267736
rect 90048 267724 90054 267776
rect 268654 267764 268660 267776
rect 268615 267736 268660 267764
rect 268654 267724 268660 267736
rect 268712 267724 268718 267776
rect 264606 264976 264612 264988
rect 264567 264948 264612 264976
rect 264606 264936 264612 264948
rect 264664 264936 264670 264988
rect 70486 264052 70492 264104
rect 70544 264092 70550 264104
rect 70670 264092 70676 264104
rect 70544 264064 70676 264092
rect 70544 264052 70550 264064
rect 70670 264052 70676 264064
rect 70728 264052 70734 264104
rect 70762 263616 70768 263628
rect 70688 263588 70768 263616
rect 70688 263560 70716 263588
rect 70762 263576 70768 263588
rect 70820 263576 70826 263628
rect 73430 263576 73436 263628
rect 73488 263576 73494 263628
rect 84470 263576 84476 263628
rect 84528 263616 84534 263628
rect 84654 263616 84660 263628
rect 84528 263588 84660 263616
rect 84528 263576 84534 263588
rect 84654 263576 84660 263588
rect 84712 263576 84718 263628
rect 211798 263576 211804 263628
rect 211856 263616 211862 263628
rect 211982 263616 211988 263628
rect 211856 263588 211988 263616
rect 211856 263576 211862 263588
rect 211982 263576 211988 263588
rect 212040 263576 212046 263628
rect 227254 263576 227260 263628
rect 227312 263616 227318 263628
rect 227438 263616 227444 263628
rect 227312 263588 227444 263616
rect 227312 263576 227318 263588
rect 227438 263576 227444 263588
rect 227496 263576 227502 263628
rect 70670 263508 70676 263560
rect 70728 263508 70734 263560
rect 73448 263480 73476 263576
rect 73522 263480 73528 263492
rect 73448 263452 73528 263480
rect 73522 263440 73528 263452
rect 73580 263440 73586 263492
rect 105170 263480 105176 263492
rect 105131 263452 105176 263480
rect 105170 263440 105176 263452
rect 105228 263440 105234 263492
rect 92750 260856 92756 260908
rect 92808 260856 92814 260908
rect 106829 260899 106887 260905
rect 106829 260865 106841 260899
rect 106875 260896 106887 260899
rect 106918 260896 106924 260908
rect 106875 260868 106924 260896
rect 106875 260865 106887 260868
rect 106829 260859 106887 260865
rect 106918 260856 106924 260868
rect 106976 260856 106982 260908
rect 234062 260896 234068 260908
rect 234023 260868 234068 260896
rect 234062 260856 234068 260868
rect 234120 260856 234126 260908
rect 249610 260896 249616 260908
rect 249571 260868 249616 260896
rect 249610 260856 249616 260868
rect 249668 260856 249674 260908
rect 250990 260896 250996 260908
rect 250951 260868 250996 260896
rect 250990 260856 250996 260868
rect 251048 260856 251054 260908
rect 252278 260896 252284 260908
rect 252239 260868 252284 260896
rect 252278 260856 252284 260868
rect 252336 260856 252342 260908
rect 259270 260896 259276 260908
rect 259231 260868 259276 260896
rect 259270 260856 259276 260868
rect 259328 260856 259334 260908
rect 324958 260896 324964 260908
rect 324919 260868 324964 260896
rect 324958 260856 324964 260868
rect 325016 260856 325022 260908
rect 89990 260788 89996 260840
rect 90048 260828 90054 260840
rect 90082 260828 90088 260840
rect 90048 260800 90088 260828
rect 90048 260788 90054 260800
rect 90082 260788 90088 260800
rect 90140 260788 90146 260840
rect 92768 260760 92796 260856
rect 105170 260828 105176 260840
rect 105131 260800 105176 260828
rect 105170 260788 105176 260800
rect 105228 260788 105234 260840
rect 151078 260828 151084 260840
rect 151039 260800 151084 260828
rect 151078 260788 151084 260800
rect 151136 260788 151142 260840
rect 92842 260760 92848 260772
rect 92768 260732 92848 260760
rect 92842 260720 92848 260732
rect 92900 260720 92906 260772
rect 70670 259360 70676 259412
rect 70728 259400 70734 259412
rect 70765 259403 70823 259409
rect 70765 259400 70777 259403
rect 70728 259372 70777 259400
rect 70728 259360 70734 259372
rect 70765 259369 70777 259372
rect 70811 259369 70823 259403
rect 70765 259363 70823 259369
rect 268746 258748 268752 258800
rect 268804 258788 268810 258800
rect 269022 258788 269028 258800
rect 268804 258760 269028 258788
rect 268804 258748 268810 258760
rect 269022 258748 269028 258760
rect 269080 258748 269086 258800
rect 106918 254028 106924 254040
rect 106844 254000 106924 254028
rect 89990 253920 89996 253972
rect 90048 253920 90054 253972
rect 70486 253852 70492 253904
rect 70544 253892 70550 253904
rect 70670 253892 70676 253904
rect 70544 253864 70676 253892
rect 70544 253852 70550 253864
rect 70670 253852 70676 253864
rect 70728 253852 70734 253904
rect 90008 253824 90036 253920
rect 106844 253904 106872 254000
rect 106918 253988 106924 254000
rect 106976 253988 106982 254040
rect 106826 253852 106832 253904
rect 106884 253852 106890 253904
rect 90082 253824 90088 253836
rect 90008 253796 90088 253824
rect 90082 253784 90088 253796
rect 90140 253784 90146 253836
rect 105170 253824 105176 253836
rect 105131 253796 105176 253824
rect 105170 253784 105176 253796
rect 105228 253784 105234 253836
rect 73433 252603 73491 252609
rect 73433 252569 73445 252603
rect 73479 252600 73491 252603
rect 73522 252600 73528 252612
rect 73479 252572 73528 252600
rect 73479 252569 73491 252572
rect 73433 252563 73491 252569
rect 73522 252560 73528 252572
rect 73580 252560 73586 252612
rect 94038 251200 94044 251252
rect 94096 251240 94102 251252
rect 94130 251240 94136 251252
rect 94096 251212 94136 251240
rect 94096 251200 94102 251212
rect 94130 251200 94136 251212
rect 94188 251200 94194 251252
rect 151078 251240 151084 251252
rect 151039 251212 151084 251240
rect 151078 251200 151084 251212
rect 151136 251200 151142 251252
rect 234062 251200 234068 251252
rect 234120 251240 234126 251252
rect 234154 251240 234160 251252
rect 234120 251212 234160 251240
rect 234120 251200 234126 251212
rect 234154 251200 234160 251212
rect 234212 251200 234218 251252
rect 324774 251200 324780 251252
rect 324832 251240 324838 251252
rect 324958 251240 324964 251252
rect 324832 251212 324964 251240
rect 324832 251200 324838 251212
rect 324958 251200 324964 251212
rect 325016 251200 325022 251252
rect 105081 251175 105139 251181
rect 105081 251141 105093 251175
rect 105127 251172 105139 251175
rect 105170 251172 105176 251184
rect 105127 251144 105176 251172
rect 105127 251141 105139 251144
rect 105081 251135 105139 251141
rect 105170 251132 105176 251144
rect 105228 251132 105234 251184
rect 252278 251172 252284 251184
rect 252239 251144 252284 251172
rect 252278 251132 252284 251144
rect 252336 251132 252342 251184
rect 324774 251104 324780 251116
rect 324735 251076 324780 251104
rect 324774 251064 324780 251076
rect 324832 251064 324838 251116
rect 81710 250996 81716 251048
rect 81768 250996 81774 251048
rect 81728 250912 81756 250996
rect 81710 250860 81716 250912
rect 81768 250860 81774 250912
rect 72142 249772 72148 249824
rect 72200 249812 72206 249824
rect 72418 249812 72424 249824
rect 72200 249784 72424 249812
rect 72200 249772 72206 249784
rect 72418 249772 72424 249784
rect 72476 249772 72482 249824
rect 92658 249772 92664 249824
rect 92716 249812 92722 249824
rect 92842 249812 92848 249824
rect 92716 249784 92848 249812
rect 92716 249772 92722 249784
rect 92842 249772 92848 249784
rect 92900 249772 92906 249824
rect 193674 249772 193680 249824
rect 193732 249812 193738 249824
rect 193858 249812 193864 249824
rect 193732 249784 193864 249812
rect 193732 249772 193738 249784
rect 193858 249772 193864 249784
rect 193916 249772 193922 249824
rect 243630 249772 243636 249824
rect 243688 249812 243694 249824
rect 243814 249812 243820 249824
rect 243688 249784 243820 249812
rect 243688 249772 243694 249784
rect 243814 249772 243820 249784
rect 243872 249772 243878 249824
rect 246942 249772 246948 249824
rect 247000 249812 247006 249824
rect 247126 249812 247132 249824
rect 247000 249784 247132 249812
rect 247000 249772 247006 249784
rect 247126 249772 247132 249784
rect 247184 249772 247190 249824
rect 78766 248412 78772 248464
rect 78824 248452 78830 248464
rect 78950 248452 78956 248464
rect 78824 248424 78956 248452
rect 78824 248412 78830 248424
rect 78950 248412 78956 248424
rect 79008 248412 79014 248464
rect 77662 244944 77668 244996
rect 77720 244984 77726 244996
rect 77846 244984 77852 244996
rect 77720 244956 77852 244984
rect 77720 244944 77726 244956
rect 77846 244944 77852 244956
rect 77904 244944 77910 244996
rect 94041 244987 94099 244993
rect 94041 244953 94053 244987
rect 94087 244984 94099 244987
rect 94130 244984 94136 244996
rect 94087 244956 94136 244984
rect 94087 244953 94099 244956
rect 94041 244947 94099 244953
rect 94130 244944 94136 244956
rect 94188 244944 94194 244996
rect 268746 244672 268752 244724
rect 268804 244712 268810 244724
rect 269022 244712 269028 244724
rect 268804 244684 269028 244712
rect 268804 244672 268810 244684
rect 269022 244672 269028 244684
rect 269080 244672 269086 244724
rect 70670 244372 70676 244384
rect 70504 244344 70676 244372
rect 70504 244316 70532 244344
rect 70670 244332 70676 244344
rect 70728 244332 70734 244384
rect 70486 244264 70492 244316
rect 70544 244264 70550 244316
rect 84470 244264 84476 244316
rect 84528 244304 84534 244316
rect 84654 244304 84660 244316
rect 84528 244276 84660 244304
rect 84528 244264 84534 244276
rect 84654 244264 84660 244276
rect 84712 244264 84718 244316
rect 211798 244264 211804 244316
rect 211856 244304 211862 244316
rect 211982 244304 211988 244316
rect 211856 244276 211988 244304
rect 211856 244264 211862 244276
rect 211982 244264 211988 244276
rect 212040 244264 212046 244316
rect 227254 244264 227260 244316
rect 227312 244304 227318 244316
rect 227438 244304 227444 244316
rect 227312 244276 227444 244304
rect 227312 244264 227318 244276
rect 227438 244264 227444 244276
rect 227496 244264 227502 244316
rect 268654 244264 268660 244316
rect 268712 244304 268718 244316
rect 268838 244304 268844 244316
rect 268712 244276 268844 244304
rect 268712 244264 268718 244276
rect 268838 244264 268844 244276
rect 268896 244264 268902 244316
rect 324777 241587 324835 241593
rect 324777 241553 324789 241587
rect 324823 241584 324835 241587
rect 324866 241584 324872 241596
rect 324823 241556 324872 241584
rect 324823 241553 324835 241556
rect 324777 241547 324835 241553
rect 324866 241544 324872 241556
rect 324924 241544 324930 241596
rect 70762 241516 70768 241528
rect 70723 241488 70768 241516
rect 70762 241476 70768 241488
rect 70820 241476 70826 241528
rect 73433 241519 73491 241525
rect 73433 241485 73445 241519
rect 73479 241516 73491 241519
rect 73706 241516 73712 241528
rect 73479 241488 73712 241516
rect 73479 241485 73491 241488
rect 73433 241479 73491 241485
rect 73706 241476 73712 241488
rect 73764 241476 73770 241528
rect 81710 241476 81716 241528
rect 81768 241476 81774 241528
rect 105078 241516 105084 241528
rect 105039 241488 105084 241516
rect 105078 241476 105084 241488
rect 105136 241476 105142 241528
rect 252278 241516 252284 241528
rect 252239 241488 252284 241516
rect 252278 241476 252284 241488
rect 252336 241476 252342 241528
rect 81728 241448 81756 241476
rect 81802 241448 81808 241460
rect 81728 241420 81808 241448
rect 81802 241408 81808 241420
rect 81860 241408 81866 241460
rect 324866 241448 324872 241460
rect 324827 241420 324872 241448
rect 324866 241408 324872 241420
rect 324924 241408 324930 241460
rect 72234 240116 72240 240168
rect 72292 240156 72298 240168
rect 72418 240156 72424 240168
rect 72292 240128 72424 240156
rect 72292 240116 72298 240128
rect 72418 240116 72424 240128
rect 72476 240116 72482 240168
rect 78766 240116 78772 240168
rect 78824 240116 78830 240168
rect 234062 240116 234068 240168
rect 234120 240156 234126 240168
rect 234154 240156 234160 240168
rect 234120 240128 234160 240156
rect 234120 240116 234126 240128
rect 234154 240116 234160 240128
rect 234212 240116 234218 240168
rect 242342 240116 242348 240168
rect 242400 240156 242406 240168
rect 242526 240156 242532 240168
rect 242400 240128 242532 240156
rect 242400 240116 242406 240128
rect 242526 240116 242532 240128
rect 242584 240116 242590 240168
rect 255222 240116 255228 240168
rect 255280 240156 255286 240168
rect 255314 240156 255320 240168
rect 255280 240128 255320 240156
rect 255280 240116 255286 240128
rect 255314 240116 255320 240128
rect 255372 240116 255378 240168
rect 78784 240088 78812 240116
rect 78858 240088 78864 240100
rect 78784 240060 78864 240088
rect 78858 240048 78864 240060
rect 78916 240048 78922 240100
rect 268746 239436 268752 239488
rect 268804 239476 268810 239488
rect 269022 239476 269028 239488
rect 268804 239448 269028 239476
rect 268804 239436 268810 239448
rect 269022 239436 269028 239448
rect 269080 239436 269086 239488
rect 81802 234608 81808 234660
rect 81860 234608 81866 234660
rect 95694 234648 95700 234660
rect 95620 234620 95700 234648
rect 70486 234540 70492 234592
rect 70544 234580 70550 234592
rect 70670 234580 70676 234592
rect 70544 234552 70676 234580
rect 70544 234540 70550 234552
rect 70670 234540 70676 234552
rect 70728 234540 70734 234592
rect 70762 234540 70768 234592
rect 70820 234580 70826 234592
rect 70820 234552 70865 234580
rect 70820 234540 70826 234552
rect 81820 234524 81848 234608
rect 95620 234592 95648 234620
rect 95694 234608 95700 234620
rect 95752 234608 95758 234660
rect 105078 234608 105084 234660
rect 105136 234608 105142 234660
rect 234062 234608 234068 234660
rect 234120 234608 234126 234660
rect 324869 234651 324927 234657
rect 324869 234617 324881 234651
rect 324915 234648 324927 234651
rect 325050 234648 325056 234660
rect 324915 234620 325056 234648
rect 324915 234617 324927 234620
rect 324869 234611 324927 234617
rect 325050 234608 325056 234620
rect 325108 234608 325114 234660
rect 95602 234540 95608 234592
rect 95660 234540 95666 234592
rect 81802 234472 81808 234524
rect 81860 234472 81866 234524
rect 105096 234512 105124 234608
rect 105170 234512 105176 234524
rect 105096 234484 105176 234512
rect 105170 234472 105176 234484
rect 105228 234472 105234 234524
rect 234080 234512 234108 234608
rect 234154 234512 234160 234524
rect 234080 234484 234160 234512
rect 234154 234472 234160 234484
rect 234212 234472 234218 234524
rect 70762 231860 70768 231872
rect 70723 231832 70768 231860
rect 70762 231820 70768 231832
rect 70820 231820 70826 231872
rect 72142 231820 72148 231872
rect 72200 231860 72206 231872
rect 72418 231860 72424 231872
rect 72200 231832 72424 231860
rect 72200 231820 72206 231832
rect 72418 231820 72424 231832
rect 72476 231820 72482 231872
rect 73430 231820 73436 231872
rect 73488 231860 73494 231872
rect 73706 231860 73712 231872
rect 73488 231832 73712 231860
rect 73488 231820 73494 231832
rect 73706 231820 73712 231832
rect 73764 231820 73770 231872
rect 94041 231863 94099 231869
rect 94041 231829 94053 231863
rect 94087 231860 94099 231863
rect 94130 231860 94136 231872
rect 94087 231832 94136 231860
rect 94087 231829 94099 231832
rect 94041 231823 94099 231829
rect 94130 231820 94136 231832
rect 94188 231820 94194 231872
rect 150986 231820 150992 231872
rect 151044 231860 151050 231872
rect 151078 231860 151084 231872
rect 151044 231832 151084 231860
rect 151044 231820 151050 231832
rect 151078 231820 151084 231832
rect 151136 231820 151142 231872
rect 89990 230460 89996 230512
rect 90048 230500 90054 230512
rect 90174 230500 90180 230512
rect 90048 230472 90180 230500
rect 90048 230460 90054 230472
rect 90174 230460 90180 230472
rect 90232 230460 90238 230512
rect 90818 230460 90824 230512
rect 90876 230500 90882 230512
rect 90910 230500 90916 230512
rect 90876 230472 90916 230500
rect 90876 230460 90882 230472
rect 90910 230460 90916 230472
rect 90968 230460 90974 230512
rect 193674 230460 193680 230512
rect 193732 230500 193738 230512
rect 193858 230500 193864 230512
rect 193732 230472 193864 230500
rect 193732 230460 193738 230472
rect 193858 230460 193864 230472
rect 193916 230460 193922 230512
rect 243630 230460 243636 230512
rect 243688 230500 243694 230512
rect 243814 230500 243820 230512
rect 243688 230472 243820 230500
rect 243688 230460 243694 230472
rect 243814 230460 243820 230472
rect 243872 230460 243878 230512
rect 246942 230460 246948 230512
rect 247000 230500 247006 230512
rect 247126 230500 247132 230512
rect 247000 230472 247132 230500
rect 247000 230460 247006 230472
rect 247126 230460 247132 230472
rect 247184 230460 247190 230512
rect 250806 230460 250812 230512
rect 250864 230500 250870 230512
rect 250990 230500 250996 230512
rect 250864 230472 250996 230500
rect 250864 230460 250870 230472
rect 250990 230460 250996 230472
rect 251048 230460 251054 230512
rect 252094 230460 252100 230512
rect 252152 230500 252158 230512
rect 252278 230500 252284 230512
rect 252152 230472 252284 230500
rect 252152 230460 252158 230472
rect 252278 230460 252284 230472
rect 252336 230460 252342 230512
rect 255222 230460 255228 230512
rect 255280 230500 255286 230512
rect 255314 230500 255320 230512
rect 255280 230472 255320 230500
rect 255280 230460 255286 230472
rect 255314 230460 255320 230472
rect 255372 230460 255378 230512
rect 259086 230460 259092 230512
rect 259144 230500 259150 230512
rect 259270 230500 259276 230512
rect 259144 230472 259276 230500
rect 259144 230460 259150 230472
rect 259270 230460 259276 230472
rect 259328 230460 259334 230512
rect 265986 230500 265992 230512
rect 265947 230472 265992 230500
rect 265986 230460 265992 230472
rect 266044 230460 266050 230512
rect 106461 230435 106519 230441
rect 106461 230401 106473 230435
rect 106507 230432 106519 230435
rect 106550 230432 106556 230444
rect 106507 230404 106556 230432
rect 106507 230401 106519 230404
rect 106461 230395 106519 230401
rect 106550 230392 106556 230404
rect 106608 230392 106614 230444
rect 268746 229712 268752 229764
rect 268804 229752 268810 229764
rect 269022 229752 269028 229764
rect 268804 229724 269028 229752
rect 268804 229712 268810 229724
rect 269022 229712 269028 229724
rect 269080 229712 269086 229764
rect 78769 229075 78827 229081
rect 78769 229041 78781 229075
rect 78815 229072 78827 229075
rect 78950 229072 78956 229084
rect 78815 229044 78956 229072
rect 78815 229041 78827 229044
rect 78769 229035 78827 229041
rect 78950 229032 78956 229044
rect 79008 229032 79014 229084
rect 255222 229032 255228 229084
rect 255280 229072 255286 229084
rect 255498 229072 255504 229084
rect 255280 229044 255504 229072
rect 255280 229032 255286 229044
rect 255498 229032 255504 229044
rect 255556 229032 255562 229084
rect 77481 225675 77539 225681
rect 77481 225641 77493 225675
rect 77527 225672 77539 225675
rect 77754 225672 77760 225684
rect 77527 225644 77760 225672
rect 77527 225641 77539 225644
rect 77481 225635 77539 225641
rect 77754 225632 77760 225644
rect 77812 225632 77818 225684
rect 70670 225060 70676 225072
rect 70504 225032 70676 225060
rect 70504 225004 70532 225032
rect 70670 225020 70676 225032
rect 70728 225020 70734 225072
rect 94130 225060 94136 225072
rect 94056 225032 94136 225060
rect 70486 224952 70492 225004
rect 70544 224952 70550 225004
rect 84470 224952 84476 225004
rect 84528 224992 84534 225004
rect 84654 224992 84660 225004
rect 84528 224964 84660 224992
rect 84528 224952 84534 224964
rect 84654 224952 84660 224964
rect 84712 224952 84718 225004
rect 94056 224936 94084 225032
rect 94130 225020 94136 225032
rect 94188 225020 94194 225072
rect 234154 225060 234160 225072
rect 234080 225032 234160 225060
rect 105078 224992 105084 225004
rect 105039 224964 105084 224992
rect 105078 224952 105084 224964
rect 105136 224952 105142 225004
rect 211798 224952 211804 225004
rect 211856 224992 211862 225004
rect 211982 224992 211988 225004
rect 211856 224964 211988 224992
rect 211856 224952 211862 224964
rect 211982 224952 211988 224964
rect 212040 224952 212046 225004
rect 227254 224952 227260 225004
rect 227312 224992 227318 225004
rect 227438 224992 227444 225004
rect 227312 224964 227444 224992
rect 227312 224952 227318 224964
rect 227438 224952 227444 224964
rect 227496 224952 227502 225004
rect 234080 224936 234108 225032
rect 234154 225020 234160 225032
rect 234212 225020 234218 225072
rect 268654 224952 268660 225004
rect 268712 224992 268718 225004
rect 268838 224992 268844 225004
rect 268712 224964 268844 224992
rect 268712 224952 268718 224964
rect 268838 224952 268844 224964
rect 268896 224952 268902 225004
rect 94038 224884 94044 224936
rect 94096 224884 94102 224936
rect 234062 224884 234068 224936
rect 234120 224884 234126 224936
rect 268746 224476 268752 224528
rect 268804 224516 268810 224528
rect 269022 224516 269028 224528
rect 268804 224488 269028 224516
rect 268804 224476 268810 224488
rect 269022 224476 269028 224488
rect 269080 224476 269086 224528
rect 72142 222164 72148 222216
rect 72200 222204 72206 222216
rect 72418 222204 72424 222216
rect 72200 222176 72424 222204
rect 72200 222164 72206 222176
rect 72418 222164 72424 222176
rect 72476 222164 72482 222216
rect 81710 222164 81716 222216
rect 81768 222204 81774 222216
rect 81802 222204 81808 222216
rect 81768 222176 81808 222204
rect 81768 222164 81774 222176
rect 81802 222164 81808 222176
rect 81860 222164 81866 222216
rect 105078 222204 105084 222216
rect 105039 222176 105084 222204
rect 105078 222164 105084 222176
rect 105136 222164 105142 222216
rect 324866 222164 324872 222216
rect 324924 222204 324930 222216
rect 325142 222204 325148 222216
rect 324924 222176 325148 222204
rect 324924 222164 324930 222176
rect 325142 222164 325148 222176
rect 325200 222164 325206 222216
rect 106458 220912 106464 220924
rect 106419 220884 106464 220912
rect 106458 220872 106464 220884
rect 106516 220872 106522 220924
rect 90634 220804 90640 220856
rect 90692 220844 90698 220856
rect 91002 220844 91008 220856
rect 90692 220816 91008 220844
rect 90692 220804 90698 220816
rect 91002 220804 91008 220816
rect 91060 220804 91066 220856
rect 242342 220804 242348 220856
rect 242400 220844 242406 220856
rect 242526 220844 242532 220856
rect 242400 220816 242532 220844
rect 242400 220804 242406 220816
rect 242526 220804 242532 220816
rect 242584 220804 242590 220856
rect 106458 220736 106464 220788
rect 106516 220776 106522 220788
rect 106642 220776 106648 220788
rect 106516 220748 106648 220776
rect 106516 220736 106522 220748
rect 106642 220736 106648 220748
rect 106700 220736 106706 220788
rect 91002 220708 91008 220720
rect 90963 220680 91008 220708
rect 91002 220668 91008 220680
rect 91060 220668 91066 220720
rect 78766 219484 78772 219496
rect 78727 219456 78772 219484
rect 78766 219444 78772 219456
rect 78824 219444 78830 219496
rect 265986 218056 265992 218068
rect 265947 218028 265992 218056
rect 265986 218016 265992 218028
rect 266044 218016 266050 218068
rect 77481 217379 77539 217385
rect 77481 217345 77493 217379
rect 77527 217376 77539 217379
rect 77570 217376 77576 217388
rect 77527 217348 77576 217376
rect 77527 217345 77539 217348
rect 77481 217339 77539 217345
rect 77570 217336 77576 217348
rect 77628 217336 77634 217388
rect 233786 216628 233792 216640
rect 233747 216600 233792 216628
rect 233786 216588 233792 216600
rect 233844 216588 233850 216640
rect 325142 215404 325148 215416
rect 325068 215376 325148 215404
rect 95694 215336 95700 215348
rect 95620 215308 95700 215336
rect 95620 215280 95648 215308
rect 95694 215296 95700 215308
rect 95752 215296 95758 215348
rect 105078 215296 105084 215348
rect 105136 215296 105142 215348
rect 70486 215228 70492 215280
rect 70544 215268 70550 215280
rect 70670 215268 70676 215280
rect 70544 215240 70676 215268
rect 70544 215228 70550 215240
rect 70670 215228 70676 215240
rect 70728 215228 70734 215280
rect 70762 215228 70768 215280
rect 70820 215268 70826 215280
rect 70820 215240 70865 215268
rect 70820 215228 70826 215240
rect 95602 215228 95608 215280
rect 95660 215228 95666 215280
rect 105096 215200 105124 215296
rect 325068 215280 325096 215376
rect 325142 215364 325148 215376
rect 325200 215364 325206 215416
rect 325050 215228 325056 215280
rect 325108 215228 325114 215280
rect 105170 215200 105176 215212
rect 105096 215172 105176 215200
rect 105170 215160 105176 215172
rect 105228 215160 105234 215212
rect 70762 212548 70768 212560
rect 70723 212520 70768 212548
rect 70762 212508 70768 212520
rect 70820 212508 70826 212560
rect 72142 212508 72148 212560
rect 72200 212548 72206 212560
rect 72418 212548 72424 212560
rect 72200 212520 72424 212548
rect 72200 212508 72206 212520
rect 72418 212508 72424 212520
rect 72476 212508 72482 212560
rect 73430 212508 73436 212560
rect 73488 212548 73494 212560
rect 73706 212548 73712 212560
rect 73488 212520 73712 212548
rect 73488 212508 73494 212520
rect 73706 212508 73712 212520
rect 73764 212508 73770 212560
rect 94130 212508 94136 212560
rect 94188 212548 94194 212560
rect 94314 212548 94320 212560
rect 94188 212520 94320 212548
rect 94188 212508 94194 212520
rect 94314 212508 94320 212520
rect 94372 212508 94378 212560
rect 150986 212508 150992 212560
rect 151044 212548 151050 212560
rect 151078 212548 151084 212560
rect 151044 212520 151084 212548
rect 151044 212508 151050 212520
rect 151078 212508 151084 212520
rect 151136 212508 151142 212560
rect 91005 212483 91063 212489
rect 91005 212449 91017 212483
rect 91051 212480 91063 212483
rect 91094 212480 91100 212492
rect 91051 212452 91100 212480
rect 91051 212449 91063 212452
rect 91005 212443 91063 212449
rect 91094 212440 91100 212452
rect 91152 212440 91158 212492
rect 78674 211148 78680 211200
rect 78732 211188 78738 211200
rect 78766 211188 78772 211200
rect 78732 211160 78772 211188
rect 78732 211148 78738 211160
rect 78766 211148 78772 211160
rect 78824 211148 78830 211200
rect 243722 211148 243728 211200
rect 243780 211188 243786 211200
rect 243814 211188 243820 211200
rect 243780 211160 243820 211188
rect 243780 211148 243786 211160
rect 243814 211148 243820 211160
rect 243872 211148 243878 211200
rect 255314 211148 255320 211200
rect 255372 211148 255378 211200
rect 91005 211123 91063 211129
rect 91005 211089 91017 211123
rect 91051 211120 91063 211123
rect 91186 211120 91192 211132
rect 91051 211092 91192 211120
rect 91051 211089 91063 211092
rect 91005 211083 91063 211089
rect 91186 211080 91192 211092
rect 91244 211080 91250 211132
rect 242342 211080 242348 211132
rect 242400 211120 242406 211132
rect 242526 211120 242532 211132
rect 242400 211092 242532 211120
rect 242400 211080 242406 211092
rect 242526 211080 242532 211092
rect 242584 211080 242590 211132
rect 255332 211052 255360 211148
rect 255590 211052 255596 211064
rect 255332 211024 255596 211052
rect 255590 211012 255596 211024
rect 255648 211012 255654 211064
rect 268746 210400 268752 210452
rect 268804 210440 268810 210452
rect 269022 210440 269028 210452
rect 268804 210412 269028 210440
rect 268804 210400 268810 210412
rect 269022 210400 269028 210412
rect 269080 210400 269086 210452
rect 235537 209763 235595 209769
rect 235537 209729 235549 209763
rect 235583 209760 235595 209763
rect 235718 209760 235724 209772
rect 235583 209732 235724 209760
rect 235583 209729 235595 209732
rect 235537 209723 235595 209729
rect 235718 209720 235724 209732
rect 235776 209720 235782 209772
rect 233786 208400 233792 208412
rect 233747 208372 233792 208400
rect 233786 208360 233792 208372
rect 233844 208360 233850 208412
rect 255406 206184 255412 206236
rect 255464 206224 255470 206236
rect 255590 206224 255596 206236
rect 255464 206196 255596 206224
rect 255464 206184 255470 206196
rect 255590 206184 255596 206196
rect 255648 206184 255654 206236
rect 70670 205748 70676 205760
rect 70504 205720 70676 205748
rect 70504 205692 70532 205720
rect 70670 205708 70676 205720
rect 70728 205708 70734 205760
rect 94130 205748 94136 205760
rect 94056 205720 94136 205748
rect 70486 205640 70492 205692
rect 70544 205640 70550 205692
rect 77478 205680 77484 205692
rect 77439 205652 77484 205680
rect 77478 205640 77484 205652
rect 77536 205640 77542 205692
rect 84470 205640 84476 205692
rect 84528 205680 84534 205692
rect 84654 205680 84660 205692
rect 84528 205652 84660 205680
rect 84528 205640 84534 205652
rect 84654 205640 84660 205652
rect 84712 205640 84718 205692
rect 89990 205640 89996 205692
rect 90048 205640 90054 205692
rect 90008 205544 90036 205640
rect 94056 205624 94084 205720
rect 94130 205708 94136 205720
rect 94188 205708 94194 205760
rect 105078 205680 105084 205692
rect 105039 205652 105084 205680
rect 105078 205640 105084 205652
rect 105136 205640 105142 205692
rect 211798 205640 211804 205692
rect 211856 205680 211862 205692
rect 211982 205680 211988 205692
rect 211856 205652 211988 205680
rect 211856 205640 211862 205652
rect 211982 205640 211988 205652
rect 212040 205640 212046 205692
rect 227254 205640 227260 205692
rect 227312 205680 227318 205692
rect 227438 205680 227444 205692
rect 227312 205652 227444 205680
rect 227312 205640 227318 205652
rect 227438 205640 227444 205652
rect 227496 205640 227502 205692
rect 268654 205640 268660 205692
rect 268712 205680 268718 205692
rect 268838 205680 268844 205692
rect 268712 205652 268844 205680
rect 268712 205640 268718 205652
rect 268838 205640 268844 205652
rect 268896 205640 268902 205692
rect 94038 205572 94044 205624
rect 94096 205572 94102 205624
rect 90082 205544 90088 205556
rect 90008 205516 90088 205544
rect 90082 205504 90088 205516
rect 90140 205504 90146 205556
rect 233786 203532 233792 203584
rect 233844 203572 233850 203584
rect 234338 203572 234344 203584
rect 233844 203544 234344 203572
rect 233844 203532 233850 203544
rect 234338 203532 234344 203544
rect 234396 203532 234402 203584
rect 72142 202852 72148 202904
rect 72200 202892 72206 202904
rect 72418 202892 72424 202904
rect 72200 202864 72424 202892
rect 72200 202852 72206 202864
rect 72418 202852 72424 202864
rect 72476 202852 72482 202904
rect 77478 202892 77484 202904
rect 77439 202864 77484 202892
rect 77478 202852 77484 202864
rect 77536 202852 77542 202904
rect 105078 202892 105084 202904
rect 105039 202864 105084 202892
rect 105078 202852 105084 202864
rect 105136 202852 105142 202904
rect 106550 202852 106556 202904
rect 106608 202892 106614 202904
rect 106734 202892 106740 202904
rect 106608 202864 106740 202892
rect 106608 202852 106614 202864
rect 106734 202852 106740 202864
rect 106792 202852 106798 202904
rect 324866 202852 324872 202904
rect 324924 202892 324930 202904
rect 325142 202892 325148 202904
rect 324924 202864 325148 202892
rect 324924 202852 324930 202864
rect 325142 202852 325148 202864
rect 325200 202852 325206 202904
rect 91002 202824 91008 202836
rect 90963 202796 91008 202824
rect 91002 202784 91008 202796
rect 91060 202784 91066 202836
rect 94038 202824 94044 202836
rect 93999 202796 94044 202824
rect 94038 202784 94044 202796
rect 94096 202784 94102 202836
rect 193674 201424 193680 201476
rect 193732 201464 193738 201476
rect 193858 201464 193864 201476
rect 193732 201436 193864 201464
rect 193732 201424 193738 201436
rect 193858 201424 193864 201436
rect 193916 201424 193922 201476
rect 246942 201424 246948 201476
rect 247000 201464 247006 201476
rect 247126 201464 247132 201476
rect 247000 201436 247132 201464
rect 247000 201424 247006 201436
rect 247126 201424 247132 201436
rect 247184 201424 247190 201476
rect 252278 201464 252284 201476
rect 252239 201436 252284 201464
rect 252278 201424 252284 201436
rect 252336 201424 252342 201476
rect 268746 200948 268752 201000
rect 268804 200988 268810 201000
rect 269022 200988 269028 201000
rect 268804 200960 269028 200988
rect 268804 200948 268810 200960
rect 269022 200948 269028 200960
rect 269080 200948 269086 201000
rect 235534 200172 235540 200184
rect 235495 200144 235540 200172
rect 235534 200132 235540 200144
rect 235592 200132 235598 200184
rect 325142 196092 325148 196104
rect 325068 196064 325148 196092
rect 81710 195984 81716 196036
rect 81768 195984 81774 196036
rect 95694 196024 95700 196036
rect 95620 195996 95700 196024
rect 70486 195916 70492 195968
rect 70544 195956 70550 195968
rect 70670 195956 70676 195968
rect 70544 195928 70676 195956
rect 70544 195916 70550 195928
rect 70670 195916 70676 195928
rect 70728 195916 70734 195968
rect 70762 195916 70768 195968
rect 70820 195956 70826 195968
rect 81728 195956 81756 195984
rect 95620 195968 95648 195996
rect 95694 195984 95700 195996
rect 95752 195984 95758 196036
rect 105078 195984 105084 196036
rect 105136 195984 105142 196036
rect 106734 195984 106740 196036
rect 106792 195984 106798 196036
rect 81802 195956 81808 195968
rect 70820 195928 70865 195956
rect 81728 195928 81808 195956
rect 70820 195916 70826 195928
rect 81802 195916 81808 195928
rect 81860 195916 81866 195968
rect 95602 195916 95608 195968
rect 95660 195916 95666 195968
rect 105096 195888 105124 195984
rect 106752 195956 106780 195984
rect 325068 195968 325096 196064
rect 325142 196052 325148 196064
rect 325200 196052 325206 196104
rect 106826 195956 106832 195968
rect 106752 195928 106832 195956
rect 106826 195916 106832 195928
rect 106884 195916 106890 195968
rect 325050 195916 325056 195968
rect 325108 195916 325114 195968
rect 105170 195888 105176 195900
rect 105096 195860 105176 195888
rect 105170 195848 105176 195860
rect 105228 195848 105234 195900
rect 92750 193264 92756 193316
rect 92808 193304 92814 193316
rect 92934 193304 92940 193316
rect 92808 193276 92940 193304
rect 92808 193264 92814 193276
rect 92934 193264 92940 193276
rect 92992 193264 92998 193316
rect 70762 193236 70768 193248
rect 70723 193208 70768 193236
rect 70762 193196 70768 193208
rect 70820 193196 70826 193248
rect 72142 193196 72148 193248
rect 72200 193236 72206 193248
rect 72418 193236 72424 193248
rect 72200 193208 72424 193236
rect 72200 193196 72206 193208
rect 72418 193196 72424 193208
rect 72476 193196 72482 193248
rect 73430 193196 73436 193248
rect 73488 193236 73494 193248
rect 73706 193236 73712 193248
rect 73488 193208 73712 193236
rect 73488 193196 73494 193208
rect 73706 193196 73712 193208
rect 73764 193196 73770 193248
rect 94041 193239 94099 193245
rect 94041 193205 94053 193239
rect 94087 193236 94099 193239
rect 94130 193236 94136 193248
rect 94087 193208 94136 193236
rect 94087 193205 94099 193208
rect 94041 193199 94099 193205
rect 94130 193196 94136 193208
rect 94188 193196 94194 193248
rect 150986 193196 150992 193248
rect 151044 193236 151050 193248
rect 151078 193236 151084 193248
rect 151044 193208 151084 193236
rect 151044 193196 151050 193208
rect 151078 193196 151084 193208
rect 151136 193196 151142 193248
rect 264606 192556 264612 192568
rect 264567 192528 264612 192556
rect 264606 192516 264612 192528
rect 264664 192516 264670 192568
rect 243722 191836 243728 191888
rect 243780 191876 243786 191888
rect 243814 191876 243820 191888
rect 243780 191848 243820 191876
rect 243780 191836 243786 191848
rect 243814 191836 243820 191848
rect 243872 191836 243878 191888
rect 252278 191876 252284 191888
rect 252239 191848 252284 191876
rect 252278 191836 252284 191848
rect 252336 191836 252342 191888
rect 72050 191768 72056 191820
rect 72108 191808 72114 191820
rect 72142 191808 72148 191820
rect 72108 191780 72148 191808
rect 72108 191768 72114 191780
rect 72142 191768 72148 191780
rect 72200 191768 72206 191820
rect 73338 191768 73344 191820
rect 73396 191808 73402 191820
rect 73430 191808 73436 191820
rect 73396 191780 73436 191808
rect 73396 191768 73402 191780
rect 73430 191768 73436 191780
rect 73488 191768 73494 191820
rect 242342 191768 242348 191820
rect 242400 191808 242406 191820
rect 242526 191808 242532 191820
rect 242400 191780 242532 191808
rect 242400 191768 242406 191780
rect 242526 191768 242532 191780
rect 242584 191768 242590 191820
rect 268746 191088 268752 191140
rect 268804 191128 268810 191140
rect 269022 191128 269028 191140
rect 268804 191100 269028 191128
rect 268804 191088 268810 191100
rect 269022 191088 269028 191100
rect 269080 191088 269086 191140
rect 255314 190476 255320 190528
rect 255372 190516 255378 190528
rect 255406 190516 255412 190528
rect 255372 190488 255412 190516
rect 255372 190476 255378 190488
rect 255406 190476 255412 190488
rect 255464 190476 255470 190528
rect 260282 190408 260288 190460
rect 260340 190448 260346 190460
rect 260466 190448 260472 190460
rect 260340 190420 260472 190448
rect 260340 190408 260346 190420
rect 260466 190408 260472 190420
rect 260524 190408 260530 190460
rect 70670 186436 70676 186448
rect 70504 186408 70676 186436
rect 70504 186380 70532 186408
rect 70670 186396 70676 186408
rect 70728 186396 70734 186448
rect 77570 186436 77576 186448
rect 77496 186408 77576 186436
rect 70486 186328 70492 186380
rect 70544 186328 70550 186380
rect 77496 186312 77524 186408
rect 77570 186396 77576 186408
rect 77628 186396 77634 186448
rect 267274 186436 267280 186448
rect 267108 186408 267280 186436
rect 267108 186380 267136 186408
rect 267274 186396 267280 186408
rect 267332 186396 267338 186448
rect 78766 186368 78772 186380
rect 78727 186340 78772 186368
rect 78766 186328 78772 186340
rect 78824 186328 78830 186380
rect 84470 186328 84476 186380
rect 84528 186368 84534 186380
rect 84654 186368 84660 186380
rect 84528 186340 84660 186368
rect 84528 186328 84534 186340
rect 84654 186328 84660 186340
rect 84712 186328 84718 186380
rect 105078 186368 105084 186380
rect 105039 186340 105084 186368
rect 105078 186328 105084 186340
rect 105136 186328 105142 186380
rect 211798 186328 211804 186380
rect 211856 186368 211862 186380
rect 211982 186368 211988 186380
rect 211856 186340 211988 186368
rect 211856 186328 211862 186340
rect 211982 186328 211988 186340
rect 212040 186328 212046 186380
rect 227254 186328 227260 186380
rect 227312 186368 227318 186380
rect 227438 186368 227444 186380
rect 227312 186340 227444 186368
rect 227312 186328 227318 186340
rect 227438 186328 227444 186340
rect 227496 186328 227502 186380
rect 267090 186328 267096 186380
rect 267148 186328 267154 186380
rect 268654 186328 268660 186380
rect 268712 186368 268718 186380
rect 268838 186368 268844 186380
rect 268712 186340 268844 186368
rect 268712 186328 268718 186340
rect 268838 186328 268844 186340
rect 268896 186328 268902 186380
rect 77478 186260 77484 186312
rect 77536 186260 77542 186312
rect 264606 185688 264612 185700
rect 264567 185660 264612 185688
rect 264606 185648 264612 185660
rect 264664 185648 264670 185700
rect 204898 183648 204904 183660
rect 204732 183620 204904 183648
rect 204732 183592 204760 183620
rect 204898 183608 204904 183620
rect 204956 183608 204962 183660
rect 78766 183580 78772 183592
rect 78727 183552 78772 183580
rect 78766 183540 78772 183552
rect 78824 183540 78830 183592
rect 91002 183580 91008 183592
rect 90963 183552 91008 183580
rect 91002 183540 91008 183552
rect 91060 183540 91066 183592
rect 105078 183580 105084 183592
rect 105039 183552 105084 183580
rect 105078 183540 105084 183552
rect 105136 183540 105142 183592
rect 106642 183540 106648 183592
rect 106700 183580 106706 183592
rect 106918 183580 106924 183592
rect 106700 183552 106924 183580
rect 106700 183540 106706 183552
rect 106918 183540 106924 183552
rect 106976 183540 106982 183592
rect 204714 183540 204720 183592
rect 204772 183540 204778 183592
rect 324866 183540 324872 183592
rect 324924 183580 324930 183592
rect 325142 183580 325148 183592
rect 324924 183552 325148 183580
rect 324924 183540 324930 183552
rect 325142 183540 325148 183552
rect 325200 183540 325206 183592
rect 77478 183512 77484 183524
rect 77439 183484 77484 183512
rect 77478 183472 77484 183484
rect 77536 183472 77542 183524
rect 193674 182112 193680 182164
rect 193732 182152 193738 182164
rect 193858 182152 193864 182164
rect 193732 182124 193864 182152
rect 193732 182112 193738 182124
rect 193858 182112 193864 182124
rect 193916 182112 193922 182164
rect 246942 182112 246948 182164
rect 247000 182152 247006 182164
rect 247126 182152 247132 182164
rect 247000 182124 247132 182152
rect 247000 182112 247006 182124
rect 247126 182112 247132 182124
rect 247184 182112 247190 182164
rect 250806 182112 250812 182164
rect 250864 182152 250870 182164
rect 250990 182152 250996 182164
rect 250864 182124 250996 182152
rect 250864 182112 250870 182124
rect 250990 182112 250996 182124
rect 251048 182112 251054 182164
rect 252094 182112 252100 182164
rect 252152 182152 252158 182164
rect 252278 182152 252284 182164
rect 252152 182124 252284 182152
rect 252152 182112 252158 182124
rect 252278 182112 252284 182124
rect 252336 182112 252342 182164
rect 259086 182112 259092 182164
rect 259144 182152 259150 182164
rect 259270 182152 259276 182164
rect 259144 182124 259276 182152
rect 259144 182112 259150 182124
rect 259270 182112 259276 182124
rect 259328 182112 259334 182164
rect 268746 181432 268752 181484
rect 268804 181472 268810 181484
rect 269022 181472 269028 181484
rect 268804 181444 269028 181472
rect 268804 181432 268810 181444
rect 269022 181432 269028 181444
rect 269080 181432 269086 181484
rect 265986 180956 265992 181008
rect 266044 180956 266050 181008
rect 266004 180872 266032 180956
rect 91002 180860 91008 180872
rect 90963 180832 91008 180860
rect 91002 180820 91008 180832
rect 91060 180820 91066 180872
rect 265986 180820 265992 180872
rect 266044 180820 266050 180872
rect 235629 180795 235687 180801
rect 235629 180761 235641 180795
rect 235675 180792 235687 180795
rect 235718 180792 235724 180804
rect 235675 180764 235724 180792
rect 235675 180761 235687 180764
rect 235629 180755 235687 180761
rect 235718 180752 235724 180764
rect 235776 180752 235782 180804
rect 265986 179364 265992 179376
rect 265947 179336 265992 179364
rect 265986 179324 265992 179336
rect 266044 179324 266050 179376
rect 267274 179364 267280 179376
rect 267235 179336 267280 179364
rect 267274 179324 267280 179336
rect 267332 179324 267338 179376
rect 91002 178684 91008 178696
rect 90963 178656 91008 178684
rect 91002 178644 91008 178656
rect 91060 178644 91066 178696
rect 325142 176780 325148 176792
rect 325068 176752 325148 176780
rect 95510 176672 95516 176724
rect 95568 176712 95574 176724
rect 95568 176684 95648 176712
rect 95568 176672 95574 176684
rect 95620 176656 95648 176684
rect 105078 176672 105084 176724
rect 105136 176672 105142 176724
rect 70486 176604 70492 176656
rect 70544 176644 70550 176656
rect 70670 176644 70676 176656
rect 70544 176616 70676 176644
rect 70544 176604 70550 176616
rect 70670 176604 70676 176616
rect 70728 176604 70734 176656
rect 70762 176604 70768 176656
rect 70820 176644 70826 176656
rect 70820 176616 70865 176644
rect 70820 176604 70826 176616
rect 95602 176604 95608 176656
rect 95660 176604 95666 176656
rect 105096 176576 105124 176672
rect 325068 176656 325096 176752
rect 325142 176740 325148 176752
rect 325200 176740 325206 176792
rect 325050 176604 325056 176656
rect 325108 176604 325114 176656
rect 105170 176576 105176 176588
rect 105096 176548 105176 176576
rect 105170 176536 105176 176548
rect 105228 176536 105234 176588
rect 72326 174060 72332 174072
rect 72287 174032 72332 174060
rect 72326 174020 72332 174032
rect 72384 174020 72390 174072
rect 89990 173952 89996 174004
rect 90048 173992 90054 174004
rect 90174 173992 90180 174004
rect 90048 173964 90180 173992
rect 90048 173952 90054 173964
rect 90174 173952 90180 173964
rect 90232 173952 90238 174004
rect 70762 173924 70768 173936
rect 70723 173896 70768 173924
rect 70762 173884 70768 173896
rect 70820 173884 70826 173936
rect 73430 173884 73436 173936
rect 73488 173924 73494 173936
rect 73614 173924 73620 173936
rect 73488 173896 73620 173924
rect 73488 173884 73494 173896
rect 73614 173884 73620 173896
rect 73672 173884 73678 173936
rect 77481 173927 77539 173933
rect 77481 173893 77493 173927
rect 77527 173924 77539 173927
rect 77570 173924 77576 173936
rect 77527 173896 77576 173924
rect 77527 173893 77539 173896
rect 77481 173887 77539 173893
rect 77570 173884 77576 173896
rect 77628 173884 77634 173936
rect 78766 173884 78772 173936
rect 78824 173924 78830 173936
rect 78858 173924 78864 173936
rect 78824 173896 78864 173924
rect 78824 173884 78830 173896
rect 78858 173884 78864 173896
rect 78916 173884 78922 173936
rect 81802 173884 81808 173936
rect 81860 173924 81866 173936
rect 81894 173924 81900 173936
rect 81860 173896 81900 173924
rect 81860 173884 81866 173896
rect 81894 173884 81900 173896
rect 81952 173884 81958 173936
rect 94130 173884 94136 173936
rect 94188 173924 94194 173936
rect 94222 173924 94228 173936
rect 94188 173896 94228 173924
rect 94188 173884 94194 173896
rect 94222 173884 94228 173896
rect 94280 173884 94286 173936
rect 106734 173884 106740 173936
rect 106792 173924 106798 173936
rect 106918 173924 106924 173936
rect 106792 173896 106924 173924
rect 106792 173884 106798 173896
rect 106918 173884 106924 173896
rect 106976 173884 106982 173936
rect 150986 173884 150992 173936
rect 151044 173924 151050 173936
rect 151078 173924 151084 173936
rect 151044 173896 151084 173924
rect 151044 173884 151050 173896
rect 151078 173884 151084 173896
rect 151136 173884 151142 173936
rect 204714 173884 204720 173936
rect 204772 173924 204778 173936
rect 204898 173924 204904 173936
rect 204772 173896 204904 173924
rect 204772 173884 204778 173896
rect 204898 173884 204904 173896
rect 204956 173884 204962 173936
rect 211706 173884 211712 173936
rect 211764 173924 211770 173936
rect 211982 173924 211988 173936
rect 211764 173896 211988 173924
rect 211764 173884 211770 173896
rect 211982 173884 211988 173896
rect 212040 173884 212046 173936
rect 227162 173884 227168 173936
rect 227220 173924 227226 173936
rect 227438 173924 227444 173936
rect 227220 173896 227444 173924
rect 227220 173884 227226 173896
rect 227438 173884 227444 173896
rect 227496 173884 227502 173936
rect 243722 172524 243728 172576
rect 243780 172564 243786 172576
rect 243814 172564 243820 172576
rect 243780 172536 243820 172564
rect 243780 172524 243786 172536
rect 243814 172524 243820 172536
rect 243872 172524 243878 172576
rect 73338 172456 73344 172508
rect 73396 172496 73402 172508
rect 73430 172496 73436 172508
rect 73396 172468 73436 172496
rect 73396 172456 73402 172468
rect 73430 172456 73436 172468
rect 73488 172456 73494 172508
rect 94130 172456 94136 172508
rect 94188 172496 94194 172508
rect 94314 172496 94320 172508
rect 94188 172468 94320 172496
rect 94188 172456 94194 172468
rect 94314 172456 94320 172468
rect 94372 172456 94378 172508
rect 242526 172496 242532 172508
rect 242487 172468 242532 172496
rect 242526 172456 242532 172468
rect 242584 172456 242590 172508
rect 243814 172388 243820 172440
rect 243872 172428 243878 172440
rect 243906 172428 243912 172440
rect 243872 172400 243912 172428
rect 243872 172388 243878 172400
rect 243906 172388 243912 172400
rect 243964 172388 243970 172440
rect 268746 171572 268752 171624
rect 268804 171612 268810 171624
rect 269022 171612 269028 171624
rect 268804 171584 269028 171612
rect 268804 171572 268810 171584
rect 269022 171572 269028 171584
rect 269080 171572 269086 171624
rect 72326 171136 72332 171148
rect 72287 171108 72332 171136
rect 72326 171096 72332 171108
rect 72384 171096 72390 171148
rect 91005 171139 91063 171145
rect 91005 171105 91017 171139
rect 91051 171136 91063 171139
rect 91186 171136 91192 171148
rect 91051 171108 91192 171136
rect 91051 171105 91063 171108
rect 91005 171099 91063 171105
rect 91186 171096 91192 171108
rect 91244 171096 91250 171148
rect 235626 171136 235632 171148
rect 235587 171108 235632 171136
rect 235626 171096 235632 171108
rect 235684 171096 235690 171148
rect 255314 171096 255320 171148
rect 255372 171136 255378 171148
rect 255406 171136 255412 171148
rect 255372 171108 255412 171136
rect 255372 171096 255378 171108
rect 255406 171096 255412 171108
rect 255464 171096 255470 171148
rect 265986 169776 265992 169788
rect 265947 169748 265992 169776
rect 265986 169736 265992 169748
rect 266044 169736 266050 169788
rect 267274 169776 267280 169788
rect 267235 169748 267280 169776
rect 267274 169736 267280 169748
rect 267332 169736 267338 169788
rect 264606 169708 264612 169720
rect 264567 169680 264612 169708
rect 264606 169668 264612 169680
rect 264664 169668 264670 169720
rect 104894 169056 104900 169108
rect 104952 169096 104958 169108
rect 105078 169096 105084 169108
rect 104952 169068 105084 169096
rect 104952 169056 104958 169068
rect 105078 169056 105084 169068
rect 105136 169056 105142 169108
rect 77386 167628 77392 167680
rect 77444 167668 77450 167680
rect 77570 167668 77576 167680
rect 77444 167640 77576 167668
rect 77444 167628 77450 167640
rect 77570 167628 77576 167640
rect 77628 167628 77634 167680
rect 78674 167628 78680 167680
rect 78732 167668 78738 167680
rect 78858 167668 78864 167680
rect 78732 167640 78864 167668
rect 78732 167628 78738 167640
rect 78858 167628 78864 167640
rect 78916 167628 78922 167680
rect 81802 167628 81808 167680
rect 81860 167668 81866 167680
rect 81986 167668 81992 167680
rect 81860 167640 81992 167668
rect 81860 167628 81866 167640
rect 81986 167628 81992 167640
rect 82044 167628 82050 167680
rect 70670 167124 70676 167136
rect 70504 167096 70676 167124
rect 70504 167068 70532 167096
rect 70670 167084 70676 167096
rect 70728 167084 70734 167136
rect 70486 167016 70492 167068
rect 70544 167016 70550 167068
rect 84470 167016 84476 167068
rect 84528 167056 84534 167068
rect 84654 167056 84660 167068
rect 84528 167028 84660 167056
rect 84528 167016 84534 167028
rect 84654 167016 84660 167028
rect 84712 167016 84718 167068
rect 211798 167016 211804 167068
rect 211856 167056 211862 167068
rect 211982 167056 211988 167068
rect 211856 167028 211988 167056
rect 211856 167016 211862 167028
rect 211982 167016 211988 167028
rect 212040 167016 212046 167068
rect 227254 167016 227260 167068
rect 227312 167056 227318 167068
rect 227438 167056 227444 167068
rect 227312 167028 227444 167056
rect 227312 167016 227318 167028
rect 227438 167016 227444 167028
rect 227496 167016 227502 167068
rect 324866 166948 324872 167000
rect 324924 166988 324930 167000
rect 325050 166988 325056 167000
rect 324924 166960 325056 166988
rect 324924 166948 324930 166960
rect 325050 166948 325056 166960
rect 325108 166948 325114 167000
rect 106642 164200 106648 164212
rect 106603 164172 106648 164200
rect 106642 164160 106648 164172
rect 106700 164160 106706 164212
rect 151078 164200 151084 164212
rect 151039 164172 151084 164200
rect 151078 164160 151084 164172
rect 151136 164160 151142 164212
rect 211890 164200 211896 164212
rect 211851 164172 211896 164200
rect 211890 164160 211896 164172
rect 211948 164160 211954 164212
rect 227346 164200 227352 164212
rect 227307 164172 227352 164200
rect 227346 164160 227352 164172
rect 227404 164160 227410 164212
rect 204806 164092 204812 164144
rect 204864 164132 204870 164144
rect 204898 164132 204904 164144
rect 204864 164104 204904 164132
rect 204864 164092 204870 164104
rect 204898 164092 204904 164104
rect 204956 164092 204962 164144
rect 242526 162908 242532 162920
rect 242487 162880 242532 162908
rect 242526 162868 242532 162880
rect 242584 162868 242590 162920
rect 193858 162840 193864 162852
rect 193819 162812 193864 162840
rect 193858 162800 193864 162812
rect 193916 162800 193922 162852
rect 234154 162800 234160 162852
rect 234212 162840 234218 162852
rect 234338 162840 234344 162852
rect 234212 162812 234344 162840
rect 234212 162800 234218 162812
rect 234338 162800 234344 162812
rect 234396 162800 234402 162852
rect 250806 162800 250812 162852
rect 250864 162840 250870 162852
rect 250990 162840 250996 162852
rect 250864 162812 250996 162840
rect 250864 162800 250870 162812
rect 250990 162800 250996 162812
rect 251048 162800 251054 162852
rect 252094 162800 252100 162852
rect 252152 162840 252158 162852
rect 252278 162840 252284 162852
rect 252152 162812 252284 162840
rect 252152 162800 252158 162812
rect 252278 162800 252284 162812
rect 252336 162800 252342 162852
rect 259086 162800 259092 162852
rect 259144 162840 259150 162852
rect 259270 162840 259276 162852
rect 259144 162812 259276 162840
rect 259144 162800 259150 162812
rect 259270 162800 259276 162812
rect 259328 162800 259334 162852
rect 268746 162324 268752 162376
rect 268804 162364 268810 162376
rect 269022 162364 269028 162376
rect 268804 162336 269028 162364
rect 268804 162324 268810 162336
rect 269022 162324 269028 162336
rect 269080 162324 269086 162376
rect 81894 161412 81900 161424
rect 81855 161384 81900 161412
rect 81894 161372 81900 161384
rect 81952 161372 81958 161424
rect 234154 161412 234160 161424
rect 234115 161384 234160 161412
rect 234154 161372 234160 161384
rect 234212 161372 234218 161424
rect 243814 161412 243820 161424
rect 243775 161384 243820 161412
rect 243814 161372 243820 161384
rect 243872 161372 243878 161424
rect 264606 160120 264612 160132
rect 264567 160092 264612 160120
rect 264606 160080 264612 160092
rect 264664 160080 264670 160132
rect 265986 160052 265992 160064
rect 265947 160024 265992 160052
rect 265986 160012 265992 160024
rect 266044 160012 266050 160064
rect 267274 160052 267280 160064
rect 267235 160024 267280 160052
rect 267274 160012 267280 160024
rect 267332 160012 267338 160064
rect 70673 157471 70731 157477
rect 70673 157437 70685 157471
rect 70719 157468 70731 157471
rect 70762 157468 70768 157480
rect 70719 157440 70768 157468
rect 70719 157437 70731 157440
rect 70673 157431 70731 157437
rect 70762 157428 70768 157440
rect 70820 157428 70826 157480
rect 89990 157428 89996 157480
rect 90048 157428 90054 157480
rect 325142 157468 325148 157480
rect 325068 157440 325148 157468
rect 90008 157344 90036 157428
rect 105078 157360 105084 157412
rect 105136 157360 105142 157412
rect 70486 157292 70492 157344
rect 70544 157332 70550 157344
rect 70762 157332 70768 157344
rect 70544 157304 70768 157332
rect 70544 157292 70550 157304
rect 70762 157292 70768 157304
rect 70820 157292 70826 157344
rect 89990 157292 89996 157344
rect 90048 157292 90054 157344
rect 105096 157264 105124 157360
rect 106642 157332 106648 157344
rect 106603 157304 106648 157332
rect 106642 157292 106648 157304
rect 106700 157292 106706 157344
rect 211890 157332 211896 157344
rect 211851 157304 211896 157332
rect 211890 157292 211896 157304
rect 211948 157292 211954 157344
rect 227346 157332 227352 157344
rect 227307 157304 227352 157332
rect 227346 157292 227352 157304
rect 227404 157292 227410 157344
rect 325068 157276 325096 157440
rect 325142 157428 325148 157440
rect 325200 157428 325206 157480
rect 105170 157264 105176 157276
rect 105096 157236 105176 157264
rect 105170 157224 105176 157236
rect 105228 157224 105234 157276
rect 325050 157224 325056 157276
rect 325108 157224 325114 157276
rect 94041 156655 94099 156661
rect 94041 156621 94053 156655
rect 94087 156652 94099 156655
rect 94130 156652 94136 156664
rect 94087 156624 94136 156652
rect 94087 156621 94099 156624
rect 94041 156615 94099 156621
rect 94130 156612 94136 156624
rect 94188 156612 94194 156664
rect 70670 154612 70676 154624
rect 70631 154584 70676 154612
rect 70670 154572 70676 154584
rect 70728 154572 70734 154624
rect 73522 154572 73528 154624
rect 73580 154612 73586 154624
rect 73614 154612 73620 154624
rect 73580 154584 73620 154612
rect 73580 154572 73586 154584
rect 73614 154572 73620 154584
rect 73672 154572 73678 154624
rect 151078 154612 151084 154624
rect 151039 154584 151084 154612
rect 151078 154572 151084 154584
rect 151136 154572 151142 154624
rect 325050 154504 325056 154556
rect 325108 154544 325114 154556
rect 325234 154544 325240 154556
rect 325108 154516 325240 154544
rect 325108 154504 325114 154516
rect 325234 154504 325240 154516
rect 325292 154504 325298 154556
rect 193858 153252 193864 153264
rect 193819 153224 193864 153252
rect 193858 153212 193864 153224
rect 193916 153212 193922 153264
rect 73430 153184 73436 153196
rect 73391 153156 73436 153184
rect 73430 153144 73436 153156
rect 73488 153144 73494 153196
rect 77478 153144 77484 153196
rect 77536 153144 77542 153196
rect 78766 153144 78772 153196
rect 78824 153144 78830 153196
rect 242526 153184 242532 153196
rect 242487 153156 242532 153184
rect 242526 153144 242532 153156
rect 242584 153144 242590 153196
rect 77496 153048 77524 153144
rect 77662 153048 77668 153060
rect 77496 153020 77668 153048
rect 77662 153008 77668 153020
rect 77720 153008 77726 153060
rect 78784 153048 78812 153144
rect 78950 153048 78956 153060
rect 78784 153020 78956 153048
rect 78950 153008 78956 153020
rect 79008 153008 79014 153060
rect 268746 152464 268752 152516
rect 268804 152504 268810 152516
rect 269022 152504 269028 152516
rect 268804 152476 269028 152504
rect 268804 152464 268810 152476
rect 269022 152464 269028 152476
rect 269080 152464 269086 152516
rect 72142 151784 72148 151836
rect 72200 151824 72206 151836
rect 72326 151824 72332 151836
rect 72200 151796 72332 151824
rect 72200 151784 72206 151796
rect 72326 151784 72332 151796
rect 72384 151784 72390 151836
rect 234154 151824 234160 151836
rect 234115 151796 234160 151824
rect 234154 151784 234160 151796
rect 234212 151784 234218 151836
rect 243814 151824 243820 151836
rect 243775 151796 243820 151824
rect 243814 151784 243820 151796
rect 243872 151784 243878 151836
rect 264514 150424 264520 150476
rect 264572 150464 264578 150476
rect 264606 150464 264612 150476
rect 264572 150436 264612 150464
rect 264572 150424 264578 150436
rect 264606 150424 264612 150436
rect 264664 150424 264670 150476
rect 265986 150464 265992 150476
rect 265947 150436 265992 150464
rect 265986 150424 265992 150436
rect 266044 150424 266050 150476
rect 267274 150464 267280 150476
rect 267235 150436 267280 150464
rect 267274 150424 267280 150436
rect 267332 150424 267338 150476
rect 105170 147744 105176 147756
rect 105096 147716 105176 147744
rect 70486 147636 70492 147688
rect 70544 147676 70550 147688
rect 70762 147676 70768 147688
rect 70544 147648 70768 147676
rect 70544 147636 70550 147648
rect 70762 147636 70768 147648
rect 70820 147636 70826 147688
rect 84470 147636 84476 147688
rect 84528 147676 84534 147688
rect 84654 147676 84660 147688
rect 84528 147648 84660 147676
rect 84528 147636 84534 147648
rect 84654 147636 84660 147648
rect 84712 147636 84718 147688
rect 105096 147620 105124 147716
rect 105170 147704 105176 147716
rect 105228 147704 105234 147756
rect 106550 147636 106556 147688
rect 106608 147676 106614 147688
rect 106734 147676 106740 147688
rect 106608 147648 106740 147676
rect 106608 147636 106614 147648
rect 106734 147636 106740 147648
rect 106792 147636 106798 147688
rect 211798 147636 211804 147688
rect 211856 147676 211862 147688
rect 211982 147676 211988 147688
rect 211856 147648 211988 147676
rect 211856 147636 211862 147648
rect 211982 147636 211988 147648
rect 212040 147636 212046 147688
rect 227254 147636 227260 147688
rect 227312 147676 227318 147688
rect 227438 147676 227444 147688
rect 227312 147648 227444 147676
rect 227312 147636 227318 147648
rect 227438 147636 227444 147648
rect 227496 147636 227502 147688
rect 268654 147636 268660 147688
rect 268712 147676 268718 147688
rect 268838 147676 268844 147688
rect 268712 147648 268844 147676
rect 268712 147636 268718 147648
rect 268838 147636 268844 147648
rect 268896 147636 268902 147688
rect 105078 147568 105084 147620
rect 105136 147568 105142 147620
rect 94041 146999 94099 147005
rect 94041 146965 94053 146999
rect 94087 146996 94099 146999
rect 94314 146996 94320 147008
rect 94087 146968 94320 146996
rect 94087 146965 94099 146968
rect 94041 146959 94099 146965
rect 94314 146956 94320 146968
rect 94372 146956 94378 147008
rect 234154 144916 234160 144968
rect 234212 144916 234218 144968
rect 73430 144888 73436 144900
rect 73391 144860 73436 144888
rect 73430 144848 73436 144860
rect 73488 144848 73494 144900
rect 106642 144888 106648 144900
rect 106603 144860 106648 144888
rect 106642 144848 106648 144860
rect 106700 144848 106706 144900
rect 151078 144888 151084 144900
rect 151039 144860 151084 144888
rect 151078 144848 151084 144860
rect 151136 144848 151142 144900
rect 211890 144888 211896 144900
rect 211851 144860 211896 144888
rect 211890 144848 211896 144860
rect 211948 144848 211954 144900
rect 227346 144888 227352 144900
rect 227307 144860 227352 144888
rect 227346 144848 227352 144860
rect 227404 144848 227410 144900
rect 81894 144820 81900 144832
rect 81855 144792 81900 144820
rect 81894 144780 81900 144792
rect 81952 144780 81958 144832
rect 204806 144780 204812 144832
rect 204864 144820 204870 144832
rect 204898 144820 204904 144832
rect 204864 144792 204904 144820
rect 204864 144780 204870 144792
rect 204898 144780 204904 144792
rect 204956 144780 204962 144832
rect 234172 144820 234200 144916
rect 234246 144820 234252 144832
rect 234172 144792 234252 144820
rect 234246 144780 234252 144792
rect 234304 144780 234310 144832
rect 242526 143596 242532 143608
rect 242487 143568 242532 143596
rect 242526 143556 242532 143568
rect 242584 143556 242590 143608
rect 243630 143556 243636 143608
rect 243688 143596 243694 143608
rect 243814 143596 243820 143608
rect 243688 143568 243820 143596
rect 243688 143556 243694 143568
rect 243814 143556 243820 143568
rect 243872 143556 243878 143608
rect 72142 143488 72148 143540
rect 72200 143528 72206 143540
rect 72326 143528 72332 143540
rect 72200 143500 72332 143528
rect 72200 143488 72206 143500
rect 72326 143488 72332 143500
rect 72384 143488 72390 143540
rect 81894 143488 81900 143540
rect 81952 143528 81958 143540
rect 82078 143528 82084 143540
rect 81952 143500 82084 143528
rect 81952 143488 81958 143500
rect 82078 143488 82084 143500
rect 82136 143488 82142 143540
rect 105078 143528 105084 143540
rect 105039 143500 105084 143528
rect 105078 143488 105084 143500
rect 105136 143488 105142 143540
rect 193858 143528 193864 143540
rect 193819 143500 193864 143528
rect 193858 143488 193864 143500
rect 193916 143488 193922 143540
rect 246942 143488 246948 143540
rect 247000 143528 247006 143540
rect 247126 143528 247132 143540
rect 247000 143500 247132 143528
rect 247000 143488 247006 143500
rect 247126 143488 247132 143500
rect 247184 143488 247190 143540
rect 248230 143488 248236 143540
rect 248288 143528 248294 143540
rect 248414 143528 248420 143540
rect 248288 143500 248420 143528
rect 248288 143488 248294 143500
rect 248414 143488 248420 143500
rect 248472 143488 248478 143540
rect 249426 143488 249432 143540
rect 249484 143528 249490 143540
rect 249610 143528 249616 143540
rect 249484 143500 249616 143528
rect 249484 143488 249490 143500
rect 249610 143488 249616 143500
rect 249668 143488 249674 143540
rect 250990 143488 250996 143540
rect 251048 143528 251054 143540
rect 251174 143528 251180 143540
rect 251048 143500 251180 143528
rect 251048 143488 251054 143500
rect 251174 143488 251180 143500
rect 251232 143488 251238 143540
rect 252094 143488 252100 143540
rect 252152 143528 252158 143540
rect 252278 143528 252284 143540
rect 252152 143500 252284 143528
rect 252152 143488 252158 143500
rect 252278 143488 252284 143500
rect 252336 143488 252342 143540
rect 259086 143488 259092 143540
rect 259144 143528 259150 143540
rect 259270 143528 259276 143540
rect 259144 143500 259276 143528
rect 259144 143488 259150 143500
rect 259270 143488 259276 143500
rect 259328 143488 259334 143540
rect 264790 143488 264796 143540
rect 264848 143528 264854 143540
rect 264974 143528 264980 143540
rect 264848 143500 264980 143528
rect 264848 143488 264854 143500
rect 264974 143488 264980 143500
rect 265032 143488 265038 143540
rect 73522 143460 73528 143472
rect 73483 143432 73528 143460
rect 73522 143420 73528 143432
rect 73580 143420 73586 143472
rect 268746 142808 268752 142860
rect 268804 142848 268810 142860
rect 269022 142848 269028 142860
rect 268804 142820 269028 142848
rect 268804 142808 268810 142820
rect 269022 142808 269028 142820
rect 269080 142808 269086 142860
rect 234157 142103 234215 142109
rect 234157 142069 234169 142103
rect 234203 142100 234215 142103
rect 234246 142100 234252 142112
rect 234203 142072 234252 142100
rect 234203 142069 234215 142072
rect 234157 142063 234215 142069
rect 234246 142060 234252 142072
rect 234304 142060 234310 142112
rect 264514 140768 264520 140820
rect 264572 140808 264578 140820
rect 264606 140808 264612 140820
rect 264572 140780 264612 140808
rect 264572 140768 264578 140780
rect 264606 140768 264612 140780
rect 264664 140768 264670 140820
rect 265986 140740 265992 140752
rect 265947 140712 265992 140740
rect 265986 140700 265992 140712
rect 266044 140700 266050 140752
rect 267274 140740 267280 140752
rect 267235 140712 267280 140740
rect 267274 140700 267280 140712
rect 267332 140700 267338 140752
rect 324958 137980 324964 138032
rect 325016 137980 325022 138032
rect 105078 137952 105084 137964
rect 105039 137924 105084 137952
rect 105078 137912 105084 137924
rect 105136 137912 105142 137964
rect 106642 137952 106648 137964
rect 106603 137924 106648 137952
rect 106642 137912 106648 137924
rect 106700 137912 106706 137964
rect 211890 137952 211896 137964
rect 211851 137924 211896 137952
rect 211890 137912 211896 137924
rect 211948 137912 211954 137964
rect 227346 137952 227352 137964
rect 227307 137924 227352 137952
rect 227346 137912 227352 137924
rect 227404 137912 227410 137964
rect 324976 137952 325004 137980
rect 325050 137952 325056 137964
rect 324976 137924 325056 137952
rect 325050 137912 325056 137924
rect 325108 137912 325114 137964
rect 151078 135300 151084 135312
rect 151039 135272 151084 135300
rect 151078 135260 151084 135272
rect 151136 135260 151142 135312
rect 325050 135192 325056 135244
rect 325108 135232 325114 135244
rect 325234 135232 325240 135244
rect 325108 135204 325240 135232
rect 325108 135192 325114 135204
rect 325234 135192 325240 135204
rect 325292 135192 325298 135244
rect 91002 133900 91008 133952
rect 91060 133940 91066 133952
rect 91186 133940 91192 133952
rect 91060 133912 91192 133940
rect 91060 133900 91066 133912
rect 91186 133900 91192 133912
rect 91244 133900 91250 133952
rect 193858 133940 193864 133952
rect 193819 133912 193864 133940
rect 193858 133900 193864 133912
rect 193916 133900 193922 133952
rect 243630 133900 243636 133952
rect 243688 133940 243694 133952
rect 243814 133940 243820 133952
rect 243688 133912 243820 133940
rect 243688 133900 243694 133912
rect 243814 133900 243820 133912
rect 243872 133900 243878 133952
rect 72326 133872 72332 133884
rect 72287 133844 72332 133872
rect 72326 133832 72332 133844
rect 72384 133832 72390 133884
rect 242526 133872 242532 133884
rect 242487 133844 242532 133872
rect 242526 133832 242532 133844
rect 242584 133832 242590 133884
rect 243814 133804 243820 133816
rect 243775 133776 243820 133804
rect 243814 133764 243820 133776
rect 243872 133764 243878 133816
rect 268746 133152 268752 133204
rect 268804 133192 268810 133204
rect 269022 133192 269028 133204
rect 268804 133164 269028 133192
rect 268804 133152 268810 133164
rect 269022 133152 269028 133164
rect 269080 133152 269086 133204
rect 73525 131563 73583 131569
rect 73525 131529 73537 131563
rect 73571 131560 73583 131563
rect 73614 131560 73620 131572
rect 73571 131532 73620 131560
rect 73571 131529 73583 131532
rect 73525 131523 73583 131529
rect 73614 131520 73620 131532
rect 73672 131520 73678 131572
rect 264514 131112 264520 131164
rect 264572 131152 264578 131164
rect 264606 131152 264612 131164
rect 264572 131124 264612 131152
rect 264572 131112 264578 131124
rect 264606 131112 264612 131124
rect 264664 131112 264670 131164
rect 265986 131152 265992 131164
rect 265947 131124 265992 131152
rect 265986 131112 265992 131124
rect 266044 131112 266050 131164
rect 267274 131152 267280 131164
rect 267235 131124 267280 131152
rect 267274 131112 267280 131124
rect 267332 131112 267338 131164
rect 70670 128432 70676 128444
rect 70504 128404 70676 128432
rect 70504 128376 70532 128404
rect 70670 128392 70676 128404
rect 70728 128392 70734 128444
rect 70762 128392 70768 128444
rect 70820 128392 70826 128444
rect 105170 128432 105176 128444
rect 105096 128404 105176 128432
rect 70486 128324 70492 128376
rect 70544 128324 70550 128376
rect 70578 128256 70584 128308
rect 70636 128296 70642 128308
rect 70780 128296 70808 128392
rect 84470 128324 84476 128376
rect 84528 128364 84534 128376
rect 84654 128364 84660 128376
rect 84528 128336 84660 128364
rect 84528 128324 84534 128336
rect 84654 128324 84660 128336
rect 84712 128324 84718 128376
rect 105096 128308 105124 128404
rect 105170 128392 105176 128404
rect 105228 128392 105234 128444
rect 211798 128324 211804 128376
rect 211856 128364 211862 128376
rect 211982 128364 211988 128376
rect 211856 128336 211988 128364
rect 211856 128324 211862 128336
rect 211982 128324 211988 128336
rect 212040 128324 212046 128376
rect 227254 128324 227260 128376
rect 227312 128364 227318 128376
rect 227438 128364 227444 128376
rect 227312 128336 227444 128364
rect 227312 128324 227318 128336
rect 227438 128324 227444 128336
rect 227496 128324 227502 128376
rect 268654 128324 268660 128376
rect 268712 128364 268718 128376
rect 268838 128364 268844 128376
rect 268712 128336 268844 128364
rect 268712 128324 268718 128336
rect 268838 128324 268844 128336
rect 268896 128324 268902 128376
rect 70636 128268 70808 128296
rect 70636 128256 70642 128268
rect 105078 128256 105084 128308
rect 105136 128256 105142 128308
rect 70486 125536 70492 125588
rect 70544 125576 70550 125588
rect 70670 125576 70676 125588
rect 70544 125548 70676 125576
rect 70544 125536 70550 125548
rect 70670 125536 70676 125548
rect 70728 125536 70734 125588
rect 90082 125536 90088 125588
rect 90140 125576 90146 125588
rect 90174 125576 90180 125588
rect 90140 125548 90180 125576
rect 90140 125536 90146 125548
rect 90174 125536 90180 125548
rect 90232 125536 90238 125588
rect 92842 125536 92848 125588
rect 92900 125576 92906 125588
rect 92934 125576 92940 125588
rect 92900 125548 92940 125576
rect 92900 125536 92906 125548
rect 92934 125536 92940 125548
rect 92992 125536 92998 125588
rect 151078 125576 151084 125588
rect 151039 125548 151084 125576
rect 151078 125536 151084 125548
rect 151136 125536 151142 125588
rect 211890 125576 211896 125588
rect 211851 125548 211896 125576
rect 211890 125536 211896 125548
rect 211948 125536 211954 125588
rect 227346 125576 227352 125588
rect 227307 125548 227352 125576
rect 227346 125536 227352 125548
rect 227404 125536 227410 125588
rect 70578 125468 70584 125520
rect 70636 125508 70642 125520
rect 70762 125508 70768 125520
rect 70636 125480 70768 125508
rect 70636 125468 70642 125480
rect 70762 125468 70768 125480
rect 70820 125468 70826 125520
rect 72326 124216 72332 124228
rect 72287 124188 72332 124216
rect 72326 124176 72332 124188
rect 72384 124176 72390 124228
rect 106458 124176 106464 124228
rect 106516 124216 106522 124228
rect 106734 124216 106740 124228
rect 106516 124188 106740 124216
rect 106516 124176 106522 124188
rect 106734 124176 106740 124188
rect 106792 124176 106798 124228
rect 234157 124219 234215 124225
rect 234157 124185 234169 124219
rect 234203 124216 234215 124219
rect 234246 124216 234252 124228
rect 234203 124188 234252 124216
rect 234203 124185 234215 124188
rect 234157 124179 234215 124185
rect 234246 124176 234252 124188
rect 234304 124176 234310 124228
rect 242526 124216 242532 124228
rect 242487 124188 242532 124216
rect 242526 124176 242532 124188
rect 242584 124176 242590 124228
rect 243814 124216 243820 124228
rect 243775 124188 243820 124216
rect 243814 124176 243820 124188
rect 243872 124176 243878 124228
rect 70762 124108 70768 124160
rect 70820 124148 70826 124160
rect 70854 124148 70860 124160
rect 70820 124120 70860 124148
rect 70820 124108 70826 124120
rect 70854 124108 70860 124120
rect 70912 124108 70918 124160
rect 91002 124108 91008 124160
rect 91060 124148 91066 124160
rect 91186 124148 91192 124160
rect 91060 124120 91192 124148
rect 91060 124108 91066 124120
rect 91186 124108 91192 124120
rect 91244 124108 91250 124160
rect 105078 124148 105084 124160
rect 105039 124120 105084 124148
rect 105078 124108 105084 124120
rect 105136 124108 105142 124160
rect 193858 124148 193864 124160
rect 193819 124120 193864 124148
rect 193858 124108 193864 124120
rect 193916 124108 193922 124160
rect 252278 124148 252284 124160
rect 252239 124120 252284 124148
rect 252278 124108 252284 124120
rect 252336 124108 252342 124160
rect 255222 124148 255228 124160
rect 255183 124120 255228 124148
rect 255222 124108 255228 124120
rect 255280 124108 255286 124160
rect 106458 124080 106464 124092
rect 106419 124052 106464 124080
rect 106458 124040 106464 124052
rect 106516 124040 106522 124092
rect 268746 123496 268752 123548
rect 268804 123536 268810 123548
rect 269022 123536 269028 123548
rect 268804 123508 269028 123536
rect 268804 123496 268810 123508
rect 269022 123496 269028 123508
rect 269080 123496 269086 123548
rect 243814 122788 243820 122800
rect 243775 122760 243820 122788
rect 243814 122748 243820 122760
rect 243872 122748 243878 122800
rect 268654 122788 268660 122800
rect 268615 122760 268660 122788
rect 268654 122748 268660 122760
rect 268712 122748 268718 122800
rect 264514 121456 264520 121508
rect 264572 121496 264578 121508
rect 264606 121496 264612 121508
rect 264572 121468 264612 121496
rect 264572 121456 264578 121468
rect 264606 121456 264612 121468
rect 264664 121456 264670 121508
rect 265986 121428 265992 121440
rect 265947 121400 265992 121428
rect 265986 121388 265992 121400
rect 266044 121388 266050 121440
rect 267274 121388 267280 121440
rect 267332 121428 267338 121440
rect 267369 121431 267427 121437
rect 267369 121428 267381 121431
rect 267332 121400 267381 121428
rect 267332 121388 267338 121400
rect 267369 121397 267381 121400
rect 267415 121397 267427 121431
rect 267369 121391 267427 121397
rect 234246 119388 234252 119400
rect 234207 119360 234252 119388
rect 234246 119348 234252 119360
rect 234304 119348 234310 119400
rect 95602 118736 95608 118788
rect 95660 118736 95666 118788
rect 95620 118652 95648 118736
rect 324958 118668 324964 118720
rect 325016 118668 325022 118720
rect 95602 118600 95608 118652
rect 95660 118600 95666 118652
rect 211890 118640 211896 118652
rect 211851 118612 211896 118640
rect 211890 118600 211896 118612
rect 211948 118600 211954 118652
rect 227346 118640 227352 118652
rect 227307 118612 227352 118640
rect 227346 118600 227352 118612
rect 227404 118600 227410 118652
rect 324976 118640 325004 118668
rect 325050 118640 325056 118652
rect 324976 118612 325056 118640
rect 325050 118600 325056 118612
rect 325108 118600 325114 118652
rect 94038 118396 94044 118448
rect 94096 118396 94102 118448
rect 94056 118368 94084 118396
rect 94130 118368 94136 118380
rect 94056 118340 94136 118368
rect 94130 118328 94136 118340
rect 94188 118328 94194 118380
rect 151078 115988 151084 116000
rect 151039 115960 151084 115988
rect 151078 115948 151084 115960
rect 151136 115948 151142 116000
rect 204898 115948 204904 116000
rect 204956 115988 204962 116000
rect 205082 115988 205088 116000
rect 204956 115960 205088 115988
rect 204956 115948 204962 115960
rect 205082 115948 205088 115960
rect 205140 115948 205146 116000
rect 78769 115923 78827 115929
rect 78769 115889 78781 115923
rect 78815 115920 78827 115923
rect 78858 115920 78864 115932
rect 78815 115892 78864 115920
rect 78815 115889 78827 115892
rect 78769 115883 78827 115889
rect 78858 115880 78864 115892
rect 78916 115880 78922 115932
rect 89990 115880 89996 115932
rect 90048 115920 90054 115932
rect 90174 115920 90180 115932
rect 90048 115892 90180 115920
rect 90048 115880 90054 115892
rect 90174 115880 90180 115892
rect 90232 115880 90238 115932
rect 92750 115880 92756 115932
rect 92808 115920 92814 115932
rect 92934 115920 92940 115932
rect 92808 115892 92940 115920
rect 92808 115880 92814 115892
rect 92934 115880 92940 115892
rect 92992 115880 92998 115932
rect 325050 115880 325056 115932
rect 325108 115920 325114 115932
rect 325234 115920 325240 115932
rect 325108 115892 325240 115920
rect 325108 115880 325114 115892
rect 325234 115880 325240 115892
rect 325292 115880 325298 115932
rect 106461 114631 106519 114637
rect 106461 114597 106473 114631
rect 106507 114628 106519 114631
rect 106550 114628 106556 114640
rect 106507 114600 106556 114628
rect 106507 114597 106519 114600
rect 106461 114591 106519 114597
rect 106550 114588 106556 114600
rect 106608 114588 106614 114640
rect 234062 114588 234068 114640
rect 234120 114628 234126 114640
rect 234249 114631 234307 114637
rect 234249 114628 234261 114631
rect 234120 114600 234261 114628
rect 234120 114588 234126 114600
rect 234249 114597 234261 114600
rect 234295 114597 234307 114631
rect 234249 114591 234307 114597
rect 72142 114520 72148 114572
rect 72200 114560 72206 114572
rect 72234 114560 72240 114572
rect 72200 114532 72240 114560
rect 72200 114520 72206 114532
rect 72234 114520 72240 114532
rect 72292 114520 72298 114572
rect 73430 114520 73436 114572
rect 73488 114560 73494 114572
rect 73522 114560 73528 114572
rect 73488 114532 73528 114560
rect 73488 114520 73494 114532
rect 73522 114520 73528 114532
rect 73580 114520 73586 114572
rect 105081 114563 105139 114569
rect 105081 114529 105093 114563
rect 105127 114560 105139 114563
rect 105170 114560 105176 114572
rect 105127 114532 105176 114560
rect 105127 114529 105139 114532
rect 105081 114523 105139 114529
rect 105170 114520 105176 114532
rect 105228 114520 105234 114572
rect 193858 114560 193864 114572
rect 193819 114532 193864 114560
rect 193858 114520 193864 114532
rect 193916 114520 193922 114572
rect 252278 114560 252284 114572
rect 252239 114532 252284 114560
rect 252278 114520 252284 114532
rect 252336 114520 252342 114572
rect 259086 114520 259092 114572
rect 259144 114560 259150 114572
rect 259270 114560 259276 114572
rect 259144 114532 259276 114560
rect 259144 114520 259150 114532
rect 259270 114520 259276 114532
rect 259328 114520 259334 114572
rect 90910 114492 90916 114504
rect 90871 114464 90916 114492
rect 90910 114452 90916 114464
rect 90968 114452 90974 114504
rect 234154 114492 234160 114504
rect 234115 114464 234160 114492
rect 234154 114452 234160 114464
rect 234212 114452 234218 114504
rect 242526 114492 242532 114504
rect 242487 114464 242532 114492
rect 242526 114452 242532 114464
rect 242584 114452 242590 114504
rect 268746 113840 268752 113892
rect 268804 113880 268810 113892
rect 269022 113880 269028 113892
rect 268804 113852 269028 113880
rect 268804 113840 268810 113852
rect 269022 113840 269028 113852
rect 269080 113840 269086 113892
rect 243814 113200 243820 113212
rect 243775 113172 243820 113200
rect 243814 113160 243820 113172
rect 243872 113160 243878 113212
rect 268657 113203 268715 113209
rect 268657 113169 268669 113203
rect 268703 113200 268715 113203
rect 268838 113200 268844 113212
rect 268703 113172 268844 113200
rect 268703 113169 268715 113172
rect 268657 113163 268715 113169
rect 268838 113160 268844 113172
rect 268896 113160 268902 113212
rect 264514 111800 264520 111852
rect 264572 111840 264578 111852
rect 264606 111840 264612 111852
rect 264572 111812 264612 111840
rect 264572 111800 264578 111812
rect 264606 111800 264612 111812
rect 264664 111800 264670 111852
rect 265986 111840 265992 111852
rect 265947 111812 265992 111840
rect 265986 111800 265992 111812
rect 266044 111800 266050 111852
rect 267274 111800 267280 111852
rect 267332 111840 267338 111852
rect 267369 111843 267427 111849
rect 267369 111840 267381 111843
rect 267332 111812 267381 111840
rect 267332 111800 267338 111812
rect 267369 111809 267381 111812
rect 267415 111809 267427 111843
rect 267369 111803 267427 111809
rect 264606 111704 264612 111716
rect 264567 111676 264612 111704
rect 264606 111664 264612 111676
rect 264664 111664 264670 111716
rect 70670 109120 70676 109132
rect 70504 109092 70676 109120
rect 70504 109064 70532 109092
rect 70670 109080 70676 109092
rect 70728 109080 70734 109132
rect 77570 109120 77576 109132
rect 77496 109092 77576 109120
rect 70486 109012 70492 109064
rect 70544 109012 70550 109064
rect 77496 108996 77524 109092
rect 77570 109080 77576 109092
rect 77628 109080 77634 109132
rect 81802 109120 81808 109132
rect 81728 109092 81808 109120
rect 81728 108996 81756 109092
rect 81802 109080 81808 109092
rect 81860 109080 81866 109132
rect 105170 109120 105176 109132
rect 105096 109092 105176 109120
rect 84470 109012 84476 109064
rect 84528 109052 84534 109064
rect 84654 109052 84660 109064
rect 84528 109024 84660 109052
rect 84528 109012 84534 109024
rect 84654 109012 84660 109024
rect 84712 109012 84718 109064
rect 105096 108996 105124 109092
rect 105170 109080 105176 109092
rect 105228 109080 105234 109132
rect 106550 109080 106556 109132
rect 106608 109080 106614 109132
rect 106568 108996 106596 109080
rect 211798 109012 211804 109064
rect 211856 109052 211862 109064
rect 211982 109052 211988 109064
rect 211856 109024 211988 109052
rect 211856 109012 211862 109024
rect 211982 109012 211988 109024
rect 212040 109012 212046 109064
rect 227254 109012 227260 109064
rect 227312 109052 227318 109064
rect 227438 109052 227444 109064
rect 227312 109024 227444 109052
rect 227312 109012 227318 109024
rect 227438 109012 227444 109024
rect 227496 109012 227502 109064
rect 268654 109012 268660 109064
rect 268712 109052 268718 109064
rect 268838 109052 268844 109064
rect 268712 109024 268844 109052
rect 268712 109012 268718 109024
rect 268838 109012 268844 109024
rect 268896 109012 268902 109064
rect 77478 108944 77484 108996
rect 77536 108944 77542 108996
rect 81710 108944 81716 108996
rect 81768 108944 81774 108996
rect 105078 108944 105084 108996
rect 105136 108944 105142 108996
rect 106550 108944 106556 108996
rect 106608 108944 106614 108996
rect 268746 108536 268752 108588
rect 268804 108576 268810 108588
rect 269022 108576 269028 108588
rect 268804 108548 269028 108576
rect 268804 108536 268810 108548
rect 269022 108536 269028 108548
rect 269080 108536 269086 108588
rect 78766 106332 78772 106344
rect 78727 106304 78772 106332
rect 78766 106292 78772 106304
rect 78824 106292 78830 106344
rect 204714 106292 204720 106344
rect 204772 106332 204778 106344
rect 204898 106332 204904 106344
rect 204772 106304 204904 106332
rect 204772 106292 204778 106304
rect 204898 106292 204904 106304
rect 204956 106292 204962 106344
rect 255222 106332 255228 106344
rect 255183 106304 255228 106332
rect 255222 106292 255228 106304
rect 255280 106292 255286 106344
rect 72234 106264 72240 106276
rect 72195 106236 72240 106264
rect 72234 106224 72240 106236
rect 72292 106224 72298 106276
rect 73522 106264 73528 106276
rect 73483 106236 73528 106264
rect 73522 106224 73528 106236
rect 73580 106224 73586 106276
rect 151078 106264 151084 106276
rect 151039 106236 151084 106264
rect 151078 106224 151084 106236
rect 151136 106224 151142 106276
rect 211890 106264 211896 106276
rect 211851 106236 211896 106264
rect 211890 106224 211896 106236
rect 211948 106224 211954 106276
rect 227346 106264 227352 106276
rect 227307 106236 227352 106264
rect 227346 106224 227352 106236
rect 227404 106224 227410 106276
rect 243814 104972 243820 104984
rect 243648 104944 243820 104972
rect 243648 104916 243676 104944
rect 243814 104932 243820 104944
rect 243872 104932 243878 104984
rect 90913 104907 90971 104913
rect 90913 104873 90925 104907
rect 90959 104904 90971 104907
rect 91002 104904 91008 104916
rect 90959 104876 91008 104904
rect 90959 104873 90971 104876
rect 90913 104867 90971 104873
rect 91002 104864 91008 104876
rect 91060 104864 91066 104916
rect 234157 104907 234215 104913
rect 234157 104873 234169 104907
rect 234203 104904 234215 104907
rect 234246 104904 234252 104916
rect 234203 104876 234252 104904
rect 234203 104873 234215 104876
rect 234157 104867 234215 104873
rect 234246 104864 234252 104876
rect 234304 104864 234310 104916
rect 242526 104904 242532 104916
rect 242487 104876 242532 104904
rect 242526 104864 242532 104876
rect 242584 104864 242590 104916
rect 243630 104864 243636 104916
rect 243688 104864 243694 104916
rect 70765 104839 70823 104845
rect 70765 104805 70777 104839
rect 70811 104836 70823 104839
rect 70854 104836 70860 104848
rect 70811 104808 70860 104836
rect 70811 104805 70823 104808
rect 70765 104799 70823 104805
rect 70854 104796 70860 104808
rect 70912 104796 70918 104848
rect 94038 104836 94044 104848
rect 93999 104808 94044 104836
rect 94038 104796 94044 104808
rect 94096 104796 94102 104848
rect 105078 104836 105084 104848
rect 105039 104808 105084 104836
rect 105078 104796 105084 104808
rect 105136 104796 105142 104848
rect 193858 104836 193864 104848
rect 193819 104808 193864 104836
rect 193858 104796 193864 104808
rect 193916 104796 193922 104848
rect 246942 104836 246948 104848
rect 246903 104808 246948 104836
rect 246942 104796 246948 104808
rect 247000 104796 247006 104848
rect 252097 104839 252155 104845
rect 252097 104805 252109 104839
rect 252143 104836 252155 104839
rect 252278 104836 252284 104848
rect 252143 104808 252284 104836
rect 252143 104805 252155 104808
rect 252097 104799 252155 104805
rect 252278 104796 252284 104808
rect 252336 104796 252342 104848
rect 255222 104836 255228 104848
rect 255183 104808 255228 104836
rect 255222 104796 255228 104808
rect 255280 104796 255286 104848
rect 259270 104836 259276 104848
rect 259231 104808 259276 104836
rect 259270 104796 259276 104808
rect 259328 104796 259334 104848
rect 106642 103436 106648 103488
rect 106700 103476 106706 103488
rect 268565 103479 268623 103485
rect 106700 103448 106745 103476
rect 106700 103436 106706 103448
rect 268565 103445 268577 103479
rect 268611 103476 268623 103479
rect 268654 103476 268660 103488
rect 268611 103448 268660 103476
rect 268611 103445 268623 103448
rect 268565 103439 268623 103445
rect 268654 103436 268660 103448
rect 268712 103436 268718 103488
rect 264606 102184 264612 102196
rect 264567 102156 264612 102184
rect 264606 102144 264612 102156
rect 264664 102144 264670 102196
rect 265986 102116 265992 102128
rect 265947 102088 265992 102116
rect 265986 102076 265992 102088
rect 266044 102076 266050 102128
rect 267274 102116 267280 102128
rect 267235 102088 267280 102116
rect 267274 102076 267280 102088
rect 267332 102076 267338 102128
rect 324774 101396 324780 101448
rect 324832 101436 324838 101448
rect 324958 101436 324964 101448
rect 324832 101408 324964 101436
rect 324832 101396 324838 101408
rect 324958 101396 324964 101408
rect 325016 101396 325022 101448
rect 234157 100079 234215 100085
rect 234157 100045 234169 100079
rect 234203 100076 234215 100079
rect 234246 100076 234252 100088
rect 234203 100048 234252 100076
rect 234203 100045 234215 100048
rect 234157 100039 234215 100045
rect 234246 100036 234252 100048
rect 234304 100036 234310 100088
rect 211890 99328 211896 99340
rect 211851 99300 211896 99328
rect 211890 99288 211896 99300
rect 211948 99288 211954 99340
rect 227346 99328 227352 99340
rect 227307 99300 227352 99328
rect 227346 99288 227352 99300
rect 227404 99288 227410 99340
rect 72234 96744 72240 96756
rect 72195 96716 72240 96744
rect 72234 96704 72240 96716
rect 72292 96704 72298 96756
rect 151078 96676 151084 96688
rect 151039 96648 151084 96676
rect 151078 96636 151084 96648
rect 151136 96636 151142 96688
rect 204714 96636 204720 96688
rect 204772 96676 204778 96688
rect 204898 96676 204904 96688
rect 204772 96648 204904 96676
rect 204772 96636 204778 96648
rect 204898 96636 204904 96648
rect 204956 96636 204962 96688
rect 235718 96608 235724 96620
rect 235679 96580 235724 96608
rect 235718 96568 235724 96580
rect 235776 96568 235782 96620
rect 70762 95316 70768 95328
rect 70723 95288 70768 95316
rect 70762 95276 70768 95288
rect 70820 95276 70826 95328
rect 70486 95208 70492 95260
rect 70544 95248 70550 95260
rect 70670 95248 70676 95260
rect 70544 95220 70676 95248
rect 70544 95208 70550 95220
rect 70670 95208 70676 95220
rect 70728 95208 70734 95260
rect 73525 95251 73583 95257
rect 73525 95217 73537 95251
rect 73571 95248 73583 95251
rect 73614 95248 73620 95260
rect 73571 95220 73620 95248
rect 73571 95217 73583 95220
rect 73525 95211 73583 95217
rect 73614 95208 73620 95220
rect 73672 95208 73678 95260
rect 91002 95208 91008 95260
rect 91060 95248 91066 95260
rect 91094 95248 91100 95260
rect 91060 95220 91100 95248
rect 91060 95208 91066 95220
rect 91094 95208 91100 95220
rect 91152 95208 91158 95260
rect 94038 95248 94044 95260
rect 93999 95220 94044 95248
rect 94038 95208 94044 95220
rect 94096 95208 94102 95260
rect 105081 95251 105139 95257
rect 105081 95217 105093 95251
rect 105127 95248 105139 95251
rect 105170 95248 105176 95260
rect 105127 95220 105176 95248
rect 105127 95217 105139 95220
rect 105081 95211 105139 95217
rect 105170 95208 105176 95220
rect 105228 95208 105234 95260
rect 193858 95248 193864 95260
rect 193819 95220 193864 95248
rect 193858 95208 193864 95220
rect 193916 95208 193922 95260
rect 234154 95248 234160 95260
rect 234115 95220 234160 95248
rect 234154 95208 234160 95220
rect 234212 95208 234218 95260
rect 243630 95208 243636 95260
rect 243688 95248 243694 95260
rect 243814 95248 243820 95260
rect 243688 95220 243820 95248
rect 243688 95208 243694 95220
rect 243814 95208 243820 95220
rect 243872 95208 243878 95260
rect 246942 95248 246948 95260
rect 246903 95220 246948 95248
rect 246942 95208 246948 95220
rect 247000 95208 247006 95260
rect 252094 95248 252100 95260
rect 252055 95220 252100 95248
rect 252094 95208 252100 95220
rect 252152 95208 252158 95260
rect 259270 95248 259276 95260
rect 259231 95220 259276 95248
rect 259270 95208 259276 95220
rect 259328 95208 259334 95260
rect 70762 95140 70768 95192
rect 70820 95180 70826 95192
rect 70946 95180 70952 95192
rect 70820 95152 70952 95180
rect 70820 95140 70826 95152
rect 70946 95140 70952 95152
rect 71004 95140 71010 95192
rect 242526 95180 242532 95192
rect 242487 95152 242532 95180
rect 242526 95140 242532 95152
rect 242584 95140 242590 95192
rect 268746 94324 268752 94376
rect 268804 94364 268810 94376
rect 269022 94364 269028 94376
rect 268804 94336 269028 94364
rect 268804 94324 268810 94336
rect 269022 94324 269028 94336
rect 269080 94324 269086 94376
rect 106550 93848 106556 93900
rect 106608 93888 106614 93900
rect 106645 93891 106703 93897
rect 106645 93888 106657 93891
rect 106608 93860 106657 93888
rect 106608 93848 106614 93860
rect 106645 93857 106657 93860
rect 106691 93857 106703 93891
rect 268562 93888 268568 93900
rect 268523 93860 268568 93888
rect 106645 93851 106703 93857
rect 268562 93848 268568 93860
rect 268620 93848 268626 93900
rect 78677 93823 78735 93829
rect 78677 93789 78689 93823
rect 78723 93820 78735 93823
rect 78858 93820 78864 93832
rect 78723 93792 78864 93820
rect 78723 93789 78735 93792
rect 78677 93783 78735 93789
rect 78858 93780 78864 93792
rect 78916 93780 78922 93832
rect 264514 92488 264520 92540
rect 264572 92528 264578 92540
rect 264606 92528 264612 92540
rect 264572 92500 264612 92528
rect 264572 92488 264578 92500
rect 264606 92488 264612 92500
rect 264664 92488 264670 92540
rect 265986 92528 265992 92540
rect 265947 92500 265992 92528
rect 265986 92488 265992 92500
rect 266044 92488 266050 92540
rect 267274 92528 267280 92540
rect 267235 92500 267280 92528
rect 267274 92488 267280 92500
rect 267332 92488 267338 92540
rect 264606 92392 264612 92404
rect 264567 92364 264612 92392
rect 264606 92352 264612 92364
rect 264664 92352 264670 92404
rect 234154 91780 234160 91792
rect 234115 91752 234160 91780
rect 234154 91740 234160 91752
rect 234212 91740 234218 91792
rect 70670 89808 70676 89820
rect 70504 89780 70676 89808
rect 70504 89752 70532 89780
rect 70670 89768 70676 89780
rect 70728 89768 70734 89820
rect 105170 89808 105176 89820
rect 105096 89780 105176 89808
rect 70486 89700 70492 89752
rect 70544 89700 70550 89752
rect 84470 89700 84476 89752
rect 84528 89740 84534 89752
rect 84654 89740 84660 89752
rect 84528 89712 84660 89740
rect 84528 89700 84534 89712
rect 84654 89700 84660 89712
rect 84712 89700 84718 89752
rect 105096 89684 105124 89780
rect 105170 89768 105176 89780
rect 105228 89768 105234 89820
rect 106550 89768 106556 89820
rect 106608 89808 106614 89820
rect 106645 89811 106703 89817
rect 106645 89808 106657 89811
rect 106608 89780 106657 89808
rect 106608 89768 106614 89780
rect 106645 89777 106657 89780
rect 106691 89777 106703 89811
rect 106645 89771 106703 89777
rect 211798 89700 211804 89752
rect 211856 89740 211862 89752
rect 211982 89740 211988 89752
rect 211856 89712 211988 89740
rect 211856 89700 211862 89712
rect 211982 89700 211988 89712
rect 212040 89700 212046 89752
rect 227254 89700 227260 89752
rect 227312 89740 227318 89752
rect 227438 89740 227444 89752
rect 227312 89712 227444 89740
rect 227312 89700 227318 89712
rect 227438 89700 227444 89712
rect 227496 89700 227502 89752
rect 105078 89632 105084 89684
rect 105136 89632 105142 89684
rect 234157 87091 234215 87097
rect 234157 87057 234169 87091
rect 234203 87088 234215 87091
rect 234338 87088 234344 87100
rect 234203 87060 234344 87088
rect 234203 87057 234215 87060
rect 234157 87051 234215 87057
rect 234338 87048 234344 87060
rect 234396 87048 234402 87100
rect 204714 86980 204720 87032
rect 204772 87020 204778 87032
rect 204898 87020 204904 87032
rect 204772 86992 204904 87020
rect 204772 86980 204778 86992
rect 204898 86980 204904 86992
rect 204956 86980 204962 87032
rect 235718 87020 235724 87032
rect 235679 86992 235724 87020
rect 235718 86980 235724 86992
rect 235776 86980 235782 87032
rect 255222 87020 255228 87032
rect 255183 86992 255228 87020
rect 255222 86980 255228 86992
rect 255280 86980 255286 87032
rect 151078 86952 151084 86964
rect 151039 86924 151084 86952
rect 151078 86912 151084 86924
rect 151136 86912 151142 86964
rect 211890 86952 211896 86964
rect 211851 86924 211896 86952
rect 211890 86912 211896 86924
rect 211948 86912 211954 86964
rect 227346 86952 227352 86964
rect 227307 86924 227352 86952
rect 227346 86912 227352 86924
rect 227404 86912 227410 86964
rect 89990 86884 89996 86896
rect 89951 86856 89996 86884
rect 89990 86844 89996 86856
rect 90048 86844 90054 86896
rect 92750 86884 92756 86896
rect 92711 86856 92756 86884
rect 92750 86844 92756 86856
rect 92808 86844 92814 86896
rect 106642 85592 106648 85604
rect 106603 85564 106648 85592
rect 106642 85552 106648 85564
rect 106700 85552 106706 85604
rect 242526 85592 242532 85604
rect 242487 85564 242532 85592
rect 242526 85552 242532 85564
rect 242584 85552 242590 85604
rect 72142 85524 72148 85536
rect 72103 85496 72148 85524
rect 72142 85484 72148 85496
rect 72200 85484 72206 85536
rect 73430 85524 73436 85536
rect 73391 85496 73436 85524
rect 73430 85484 73436 85496
rect 73488 85484 73494 85536
rect 77478 85524 77484 85536
rect 77439 85496 77484 85524
rect 77478 85484 77484 85496
rect 77536 85484 77542 85536
rect 81710 85524 81716 85536
rect 81671 85496 81716 85524
rect 81710 85484 81716 85496
rect 81768 85484 81774 85536
rect 94038 85524 94044 85536
rect 93999 85496 94044 85524
rect 94038 85484 94044 85496
rect 94096 85484 94102 85536
rect 105078 85524 105084 85536
rect 105039 85496 105084 85524
rect 105078 85484 105084 85496
rect 105136 85484 105142 85536
rect 193858 85524 193864 85536
rect 193819 85496 193864 85524
rect 193858 85484 193864 85496
rect 193916 85484 193922 85536
rect 204714 85524 204720 85536
rect 204675 85496 204720 85524
rect 204714 85484 204720 85496
rect 204772 85484 204778 85536
rect 234157 85527 234215 85533
rect 234157 85493 234169 85527
rect 234203 85524 234215 85527
rect 234246 85524 234252 85536
rect 234203 85496 234252 85524
rect 234203 85493 234215 85496
rect 234157 85487 234215 85493
rect 234246 85484 234252 85496
rect 234304 85484 234310 85536
rect 246942 85524 246948 85536
rect 246903 85496 246948 85524
rect 246942 85484 246948 85496
rect 247000 85484 247006 85536
rect 252278 85524 252284 85536
rect 252239 85496 252284 85524
rect 252278 85484 252284 85496
rect 252336 85484 252342 85536
rect 255222 85524 255228 85536
rect 255183 85496 255228 85524
rect 255222 85484 255228 85496
rect 255280 85484 255286 85536
rect 259270 85524 259276 85536
rect 259231 85496 259276 85524
rect 259270 85484 259276 85496
rect 259328 85484 259334 85536
rect 268746 84872 268752 84924
rect 268804 84912 268810 84924
rect 269022 84912 269028 84924
rect 268804 84884 269028 84912
rect 268804 84872 268810 84884
rect 269022 84872 269028 84884
rect 269080 84872 269086 84924
rect 78674 84300 78680 84312
rect 78635 84272 78680 84300
rect 78674 84260 78680 84272
rect 78732 84260 78738 84312
rect 78674 84124 78680 84176
rect 78732 84124 78738 84176
rect 105081 84167 105139 84173
rect 105081 84133 105093 84167
rect 105127 84133 105139 84167
rect 105081 84127 105139 84133
rect 78692 84096 78720 84124
rect 78858 84096 78864 84108
rect 78692 84068 78864 84096
rect 78858 84056 78864 84068
rect 78916 84056 78922 84108
rect 104986 84056 104992 84108
rect 105044 84096 105050 84108
rect 105096 84096 105124 84127
rect 105044 84068 105124 84096
rect 105044 84056 105050 84068
rect 264606 82872 264612 82884
rect 264567 82844 264612 82872
rect 264606 82832 264612 82844
rect 264664 82832 264670 82884
rect 78677 82807 78735 82813
rect 78677 82773 78689 82807
rect 78723 82804 78735 82807
rect 78858 82804 78864 82816
rect 78723 82776 78864 82804
rect 78723 82773 78735 82776
rect 78677 82767 78735 82773
rect 78858 82764 78864 82776
rect 78916 82764 78922 82816
rect 265986 82804 265992 82816
rect 265947 82776 265992 82804
rect 265986 82764 265992 82776
rect 266044 82764 266050 82816
rect 267274 82804 267280 82816
rect 267235 82776 267280 82804
rect 267274 82764 267280 82776
rect 267332 82764 267338 82816
rect 94041 80971 94099 80977
rect 94041 80937 94053 80971
rect 94087 80968 94099 80971
rect 94314 80968 94320 80980
rect 94087 80940 94320 80968
rect 94087 80937 94099 80940
rect 94041 80931 94099 80937
rect 94314 80928 94320 80940
rect 94372 80928 94378 80980
rect 324958 80044 324964 80096
rect 325016 80044 325022 80096
rect 324976 79948 325004 80044
rect 325050 79948 325056 79960
rect 324976 79920 325056 79948
rect 325050 79908 325056 79920
rect 325108 79908 325114 79960
rect 89990 77296 89996 77308
rect 89951 77268 89996 77296
rect 89990 77256 89996 77268
rect 90048 77256 90054 77308
rect 92750 77296 92756 77308
rect 92711 77268 92756 77296
rect 92750 77256 92756 77268
rect 92808 77256 92814 77308
rect 151078 77296 151084 77308
rect 151039 77268 151084 77296
rect 151078 77256 151084 77268
rect 151136 77256 151142 77308
rect 211893 77299 211951 77305
rect 211893 77265 211905 77299
rect 211939 77296 211951 77299
rect 211982 77296 211988 77308
rect 211939 77268 211988 77296
rect 211939 77265 211951 77268
rect 211893 77259 211951 77265
rect 211982 77256 211988 77268
rect 212040 77256 212046 77308
rect 227349 77299 227407 77305
rect 227349 77265 227361 77299
rect 227395 77296 227407 77299
rect 227438 77296 227444 77308
rect 227395 77268 227444 77296
rect 227395 77265 227407 77268
rect 227349 77259 227407 77265
rect 227438 77256 227444 77268
rect 227496 77256 227502 77308
rect 93854 77188 93860 77240
rect 93912 77188 93918 77240
rect 93946 77188 93952 77240
rect 94004 77188 94010 77240
rect 235718 77228 235724 77240
rect 235679 77200 235724 77228
rect 235718 77188 235724 77200
rect 235776 77188 235782 77240
rect 324961 77231 325019 77237
rect 324961 77197 324973 77231
rect 325007 77228 325019 77231
rect 325050 77228 325056 77240
rect 325007 77200 325056 77228
rect 325007 77197 325019 77200
rect 324961 77191 325019 77197
rect 325050 77188 325056 77200
rect 325108 77188 325114 77240
rect 93872 77036 93900 77188
rect 93964 77104 93992 77188
rect 93946 77052 93952 77104
rect 94004 77052 94010 77104
rect 93854 76984 93860 77036
rect 93912 76984 93918 77036
rect 72142 75936 72148 75948
rect 72103 75908 72148 75936
rect 72142 75896 72148 75908
rect 72200 75896 72206 75948
rect 73433 75939 73491 75945
rect 73433 75905 73445 75939
rect 73479 75936 73491 75939
rect 73522 75936 73528 75948
rect 73479 75908 73528 75936
rect 73479 75905 73491 75908
rect 73433 75899 73491 75905
rect 73522 75896 73528 75908
rect 73580 75896 73586 75948
rect 77481 75939 77539 75945
rect 77481 75905 77493 75939
rect 77527 75936 77539 75939
rect 77570 75936 77576 75948
rect 77527 75908 77576 75936
rect 77527 75905 77539 75908
rect 77481 75899 77539 75905
rect 77570 75896 77576 75908
rect 77628 75896 77634 75948
rect 81713 75939 81771 75945
rect 81713 75905 81725 75939
rect 81759 75936 81771 75939
rect 81802 75936 81808 75948
rect 81759 75908 81808 75936
rect 81759 75905 81771 75908
rect 81713 75899 81771 75905
rect 81802 75896 81808 75908
rect 81860 75896 81866 75948
rect 193858 75936 193864 75948
rect 193819 75908 193864 75936
rect 193858 75896 193864 75908
rect 193916 75896 193922 75948
rect 204717 75939 204775 75945
rect 204717 75905 204729 75939
rect 204763 75936 204775 75939
rect 204898 75936 204904 75948
rect 204763 75908 204904 75936
rect 204763 75905 204775 75908
rect 204717 75899 204775 75905
rect 204898 75896 204904 75908
rect 204956 75896 204962 75948
rect 234154 75936 234160 75948
rect 234115 75908 234160 75936
rect 234154 75896 234160 75908
rect 234212 75896 234218 75948
rect 243630 75896 243636 75948
rect 243688 75936 243694 75948
rect 243814 75936 243820 75948
rect 243688 75908 243820 75936
rect 243688 75896 243694 75908
rect 243814 75896 243820 75908
rect 243872 75896 243878 75948
rect 246942 75936 246948 75948
rect 246903 75908 246948 75936
rect 246942 75896 246948 75908
rect 247000 75896 247006 75948
rect 252278 75936 252284 75948
rect 252239 75908 252284 75936
rect 252278 75896 252284 75908
rect 252336 75896 252342 75948
rect 255222 75936 255228 75948
rect 255183 75908 255228 75936
rect 255222 75896 255228 75908
rect 255280 75896 255286 75948
rect 259270 75936 259276 75948
rect 259231 75908 259276 75936
rect 259270 75896 259276 75908
rect 259328 75896 259334 75948
rect 106461 75871 106519 75877
rect 106461 75837 106473 75871
rect 106507 75868 106519 75871
rect 106550 75868 106556 75880
rect 106507 75840 106556 75868
rect 106507 75837 106519 75840
rect 106461 75831 106519 75837
rect 106550 75828 106556 75840
rect 106608 75828 106614 75880
rect 211893 75871 211951 75877
rect 211893 75837 211905 75871
rect 211939 75868 211951 75871
rect 211982 75868 211988 75880
rect 211939 75840 211988 75868
rect 211939 75837 211951 75840
rect 211893 75831 211951 75837
rect 211982 75828 211988 75840
rect 212040 75828 212046 75880
rect 242526 75868 242532 75880
rect 242487 75840 242532 75868
rect 242526 75828 242532 75840
rect 242584 75828 242590 75880
rect 268746 75080 268752 75132
rect 268804 75120 268810 75132
rect 269022 75120 269028 75132
rect 268804 75092 269028 75120
rect 268804 75080 268810 75092
rect 269022 75080 269028 75092
rect 269080 75080 269086 75132
rect 104986 74576 104992 74588
rect 104947 74548 104992 74576
rect 104986 74536 104992 74548
rect 105044 74536 105050 74588
rect 94133 74511 94191 74517
rect 94133 74477 94145 74511
rect 94179 74508 94191 74511
rect 94314 74508 94320 74520
rect 94179 74480 94320 74508
rect 94179 74477 94191 74480
rect 94133 74471 94191 74477
rect 94314 74468 94320 74480
rect 94372 74468 94378 74520
rect 264514 73176 264520 73228
rect 264572 73216 264578 73228
rect 264606 73216 264612 73228
rect 264572 73188 264612 73216
rect 264572 73176 264578 73188
rect 264606 73176 264612 73188
rect 264664 73176 264670 73228
rect 265986 73216 265992 73228
rect 265947 73188 265992 73216
rect 265986 73176 265992 73188
rect 266044 73176 266050 73228
rect 267274 73216 267280 73228
rect 267235 73188 267280 73216
rect 267274 73176 267280 73188
rect 267332 73176 267338 73228
rect 72142 72468 72148 72480
rect 72103 72440 72148 72468
rect 72142 72428 72148 72440
rect 72200 72428 72206 72480
rect 70486 71408 70492 71460
rect 70544 71448 70550 71460
rect 70670 71448 70676 71460
rect 70544 71420 70676 71448
rect 70544 71408 70550 71420
rect 70670 71408 70676 71420
rect 70728 71408 70734 71460
rect 70762 70496 70768 70508
rect 70688 70468 70768 70496
rect 70688 70372 70716 70468
rect 70762 70456 70768 70468
rect 70820 70456 70826 70508
rect 77570 70496 77576 70508
rect 77496 70468 77576 70496
rect 77496 70372 77524 70468
rect 77570 70456 77576 70468
rect 77628 70456 77634 70508
rect 81802 70456 81808 70508
rect 81860 70456 81866 70508
rect 81820 70372 81848 70456
rect 268654 70388 268660 70440
rect 268712 70428 268718 70440
rect 268838 70428 268844 70440
rect 268712 70400 268844 70428
rect 268712 70388 268718 70400
rect 268838 70388 268844 70400
rect 268896 70388 268902 70440
rect 70670 70320 70676 70372
rect 70728 70320 70734 70372
rect 77478 70320 77484 70372
rect 77536 70320 77542 70372
rect 81802 70320 81808 70372
rect 81860 70320 81866 70372
rect 211890 70360 211896 70372
rect 211851 70332 211896 70360
rect 211890 70320 211896 70332
rect 211948 70320 211954 70372
rect 72142 67708 72148 67720
rect 72103 67680 72148 67708
rect 72142 67668 72148 67680
rect 72200 67668 72206 67720
rect 234062 67600 234068 67652
rect 234120 67640 234126 67652
rect 234246 67640 234252 67652
rect 234120 67612 234252 67640
rect 234120 67600 234126 67612
rect 234246 67600 234252 67612
rect 234304 67600 234310 67652
rect 235718 67640 235724 67652
rect 235679 67612 235724 67640
rect 235718 67600 235724 67612
rect 235776 67600 235782 67652
rect 324958 67640 324964 67652
rect 324919 67612 324964 67640
rect 324958 67600 324964 67612
rect 325016 67600 325022 67652
rect 70670 67572 70676 67584
rect 70631 67544 70676 67572
rect 70670 67532 70676 67544
rect 70728 67532 70734 67584
rect 89990 67572 89996 67584
rect 89951 67544 89996 67572
rect 89990 67532 89996 67544
rect 90048 67532 90054 67584
rect 92750 67572 92756 67584
rect 92711 67544 92756 67572
rect 92750 67532 92756 67544
rect 92808 67532 92814 67584
rect 151078 67572 151084 67584
rect 151039 67544 151084 67572
rect 151078 67532 151084 67544
rect 151136 67532 151142 67584
rect 70486 67124 70492 67176
rect 70544 67164 70550 67176
rect 70670 67164 70676 67176
rect 70544 67136 70676 67164
rect 70544 67124 70550 67136
rect 70670 67124 70676 67136
rect 70728 67124 70734 67176
rect 91094 66348 91100 66360
rect 91020 66320 91100 66348
rect 91020 66292 91048 66320
rect 91094 66308 91100 66320
rect 91152 66308 91158 66360
rect 106458 66348 106464 66360
rect 106419 66320 106464 66348
rect 106458 66308 106464 66320
rect 106516 66308 106522 66360
rect 84562 66240 84568 66292
rect 84620 66280 84626 66292
rect 84654 66280 84660 66292
rect 84620 66252 84660 66280
rect 84620 66240 84626 66252
rect 84654 66240 84660 66252
rect 84712 66240 84718 66292
rect 91002 66240 91008 66292
rect 91060 66240 91066 66292
rect 104986 66280 104992 66292
rect 104947 66252 104992 66280
rect 104986 66240 104992 66252
rect 105044 66240 105050 66292
rect 242526 66280 242532 66292
rect 242487 66252 242532 66280
rect 242526 66240 242532 66252
rect 242584 66240 242590 66292
rect 72053 66215 72111 66221
rect 72053 66181 72065 66215
rect 72099 66212 72111 66215
rect 72142 66212 72148 66224
rect 72099 66184 72148 66212
rect 72099 66181 72111 66184
rect 72053 66175 72111 66181
rect 72142 66172 72148 66184
rect 72200 66172 72206 66224
rect 77386 66172 77392 66224
rect 77444 66212 77450 66224
rect 77478 66212 77484 66224
rect 77444 66184 77484 66212
rect 77444 66172 77450 66184
rect 77478 66172 77484 66184
rect 77536 66172 77542 66224
rect 106458 66172 106464 66224
rect 106516 66212 106522 66224
rect 106550 66212 106556 66224
rect 106516 66184 106556 66212
rect 106516 66172 106522 66184
rect 106550 66172 106556 66184
rect 106608 66172 106614 66224
rect 193858 66212 193864 66224
rect 193819 66184 193864 66212
rect 193858 66172 193864 66184
rect 193916 66172 193922 66224
rect 204898 66212 204904 66224
rect 204859 66184 204904 66212
rect 204898 66172 204904 66184
rect 204956 66172 204962 66224
rect 234062 66212 234068 66224
rect 234023 66184 234068 66212
rect 234062 66172 234068 66184
rect 234120 66172 234126 66224
rect 246942 66212 246948 66224
rect 246903 66184 246948 66212
rect 246942 66172 246948 66184
rect 247000 66172 247006 66224
rect 252278 66212 252284 66224
rect 252239 66184 252284 66212
rect 252278 66172 252284 66184
rect 252336 66172 252342 66224
rect 255222 66212 255228 66224
rect 255183 66184 255228 66212
rect 255222 66172 255228 66184
rect 255280 66172 255286 66224
rect 259270 66212 259276 66224
rect 259231 66184 259276 66212
rect 259270 66172 259276 66184
rect 259328 66172 259334 66224
rect 262030 66172 262036 66224
rect 262088 66212 262094 66224
rect 262214 66212 262220 66224
rect 262088 66184 262220 66212
rect 262088 66172 262094 66184
rect 262214 66172 262220 66184
rect 262272 66172 262278 66224
rect 268746 65492 268752 65544
rect 268804 65532 268810 65544
rect 269022 65532 269028 65544
rect 268804 65504 269028 65532
rect 268804 65492 268810 65504
rect 269022 65492 269028 65504
rect 269080 65492 269086 65544
rect 78674 64920 78680 64932
rect 78635 64892 78680 64920
rect 78674 64880 78680 64892
rect 78732 64880 78738 64932
rect 94130 64920 94136 64932
rect 94091 64892 94136 64920
rect 94130 64880 94136 64892
rect 94188 64880 94194 64932
rect 104986 64812 104992 64864
rect 105044 64852 105050 64864
rect 105262 64852 105268 64864
rect 105044 64824 105268 64852
rect 105044 64812 105050 64824
rect 105262 64812 105268 64824
rect 105320 64812 105326 64864
rect 267274 63492 267280 63504
rect 267235 63464 267280 63492
rect 267274 63452 267280 63464
rect 267332 63452 267338 63504
rect 78674 61412 78680 61464
rect 78732 61452 78738 61464
rect 78950 61452 78956 61464
rect 78732 61424 78956 61452
rect 78732 61412 78738 61424
rect 78950 61412 78956 61424
rect 79008 61412 79014 61464
rect 94130 60024 94136 60036
rect 94091 59996 94136 60024
rect 94130 59984 94136 59996
rect 94188 59984 94194 60036
rect 89990 58052 89996 58064
rect 89951 58024 89996 58052
rect 89990 58012 89996 58024
rect 90048 58012 90054 58064
rect 92750 58052 92756 58064
rect 92711 58024 92756 58052
rect 92750 58012 92756 58024
rect 92808 58012 92814 58064
rect 70673 57987 70731 57993
rect 70673 57953 70685 57987
rect 70719 57984 70731 57987
rect 70762 57984 70768 57996
rect 70719 57956 70768 57984
rect 70719 57953 70731 57956
rect 70673 57947 70731 57953
rect 70762 57944 70768 57956
rect 70820 57944 70826 57996
rect 151078 57984 151084 57996
rect 151039 57956 151084 57984
rect 151078 57944 151084 57956
rect 151136 57944 151142 57996
rect 211893 57919 211951 57925
rect 211893 57885 211905 57919
rect 211939 57916 211951 57919
rect 211982 57916 211988 57928
rect 211939 57888 211988 57916
rect 211939 57885 211951 57888
rect 211893 57879 211951 57885
rect 211982 57876 211988 57888
rect 212040 57876 212046 57928
rect 227349 57919 227407 57925
rect 227349 57885 227361 57919
rect 227395 57916 227407 57919
rect 227438 57916 227444 57928
rect 227395 57888 227444 57916
rect 227395 57885 227407 57888
rect 227349 57879 227407 57885
rect 227438 57876 227444 57888
rect 227496 57876 227502 57928
rect 235718 57916 235724 57928
rect 235679 57888 235724 57916
rect 235718 57876 235724 57888
rect 235776 57876 235782 57928
rect 234065 57851 234123 57857
rect 234065 57817 234077 57851
rect 234111 57848 234123 57851
rect 234246 57848 234252 57860
rect 234111 57820 234252 57848
rect 234111 57817 234123 57820
rect 234065 57811 234123 57817
rect 234246 57808 234252 57820
rect 234304 57808 234310 57860
rect 90913 56695 90971 56701
rect 90913 56661 90925 56695
rect 90959 56692 90971 56695
rect 91002 56692 91008 56704
rect 90959 56664 91008 56692
rect 90959 56661 90971 56664
rect 90913 56655 90971 56661
rect 91002 56652 91008 56664
rect 91060 56652 91066 56704
rect 72050 56624 72056 56636
rect 72011 56596 72056 56624
rect 72050 56584 72056 56596
rect 72108 56584 72114 56636
rect 193858 56624 193864 56636
rect 193819 56596 193864 56624
rect 193858 56584 193864 56596
rect 193916 56584 193922 56636
rect 204898 56624 204904 56636
rect 204859 56596 204904 56624
rect 204898 56584 204904 56596
rect 204956 56584 204962 56636
rect 243630 56584 243636 56636
rect 243688 56624 243694 56636
rect 243814 56624 243820 56636
rect 243688 56596 243820 56624
rect 243688 56584 243694 56596
rect 243814 56584 243820 56596
rect 243872 56584 243878 56636
rect 246942 56624 246948 56636
rect 246903 56596 246948 56624
rect 246942 56584 246948 56596
rect 247000 56584 247006 56636
rect 252278 56624 252284 56636
rect 252239 56596 252284 56624
rect 252278 56584 252284 56596
rect 252336 56584 252342 56636
rect 255222 56624 255228 56636
rect 255183 56596 255228 56624
rect 255222 56584 255228 56596
rect 255280 56584 255286 56636
rect 259270 56624 259276 56636
rect 259231 56596 259276 56624
rect 259270 56584 259276 56596
rect 259328 56584 259334 56636
rect 96982 56556 96988 56568
rect 96943 56528 96988 56556
rect 96982 56516 96988 56528
rect 97040 56516 97046 56568
rect 242526 56556 242532 56568
rect 242487 56528 242532 56556
rect 242526 56516 242532 56528
rect 242584 56516 242590 56568
rect 268746 55836 268752 55888
rect 268804 55876 268810 55888
rect 269022 55876 269028 55888
rect 268804 55848 269028 55876
rect 268804 55836 268810 55848
rect 269022 55836 269028 55848
rect 269080 55836 269086 55888
rect 90910 55264 90916 55276
rect 90871 55236 90916 55264
rect 90910 55224 90916 55236
rect 90968 55224 90974 55276
rect 267274 53836 267280 53848
rect 267235 53808 267280 53836
rect 267274 53796 267280 53808
rect 267332 53796 267338 53848
rect 264606 53768 264612 53780
rect 264567 53740 264612 53768
rect 264606 53728 264612 53740
rect 264664 53728 264670 53780
rect 70486 53116 70492 53168
rect 70544 53156 70550 53168
rect 70670 53156 70676 53168
rect 70544 53128 70676 53156
rect 70544 53116 70550 53128
rect 70670 53116 70676 53128
rect 70728 53116 70734 53168
rect 81713 51799 81771 51805
rect 81713 51765 81725 51799
rect 81759 51796 81771 51799
rect 81802 51796 81808 51808
rect 81759 51768 81808 51796
rect 81759 51765 81771 51768
rect 81713 51759 81771 51765
rect 81802 51756 81808 51768
rect 81860 51756 81866 51808
rect 70762 51116 70768 51128
rect 70688 51088 70768 51116
rect 70688 51060 70716 51088
rect 70762 51076 70768 51088
rect 70820 51076 70826 51128
rect 70670 51008 70676 51060
rect 70728 51008 70734 51060
rect 106550 51008 106556 51060
rect 106608 51048 106614 51060
rect 106734 51048 106740 51060
rect 106608 51020 106740 51048
rect 106608 51008 106614 51020
rect 106734 51008 106740 51020
rect 106792 51008 106798 51060
rect 227346 51048 227352 51060
rect 227307 51020 227352 51048
rect 227346 51008 227352 51020
rect 227404 51008 227410 51060
rect 211890 50708 211896 50720
rect 211851 50680 211896 50708
rect 211890 50668 211896 50680
rect 211948 50668 211954 50720
rect 94130 50640 94136 50652
rect 94091 50612 94136 50640
rect 94130 50600 94136 50612
rect 94188 50600 94194 50652
rect 262030 49376 262036 49428
rect 262088 49416 262094 49428
rect 262214 49416 262220 49428
rect 262088 49388 262220 49416
rect 262088 49376 262094 49388
rect 262214 49376 262220 49388
rect 262272 49376 262278 49428
rect 73430 48356 73436 48408
rect 73488 48356 73494 48408
rect 72050 48288 72056 48340
rect 72108 48328 72114 48340
rect 72234 48328 72240 48340
rect 72108 48300 72240 48328
rect 72108 48288 72114 48300
rect 72234 48288 72240 48300
rect 72292 48288 72298 48340
rect 73448 48328 73476 48356
rect 73522 48328 73528 48340
rect 73448 48300 73528 48328
rect 73522 48288 73528 48300
rect 73580 48288 73586 48340
rect 78766 48288 78772 48340
rect 78824 48328 78830 48340
rect 78950 48328 78956 48340
rect 78824 48300 78956 48328
rect 78824 48288 78830 48300
rect 78950 48288 78956 48300
rect 79008 48288 79014 48340
rect 84562 48288 84568 48340
rect 84620 48328 84626 48340
rect 84654 48328 84660 48340
rect 84620 48300 84660 48328
rect 84620 48288 84626 48300
rect 84654 48288 84660 48300
rect 84712 48288 84718 48340
rect 92750 48288 92756 48340
rect 92808 48288 92814 48340
rect 234062 48288 234068 48340
rect 234120 48328 234126 48340
rect 234246 48328 234252 48340
rect 234120 48300 234252 48328
rect 234120 48288 234126 48300
rect 234246 48288 234252 48300
rect 234304 48288 234310 48340
rect 235718 48328 235724 48340
rect 235679 48300 235724 48328
rect 235718 48288 235724 48300
rect 235776 48288 235782 48340
rect 92768 48192 92796 48288
rect 151078 48260 151084 48272
rect 151039 48232 151084 48260
rect 151078 48220 151084 48232
rect 151136 48220 151142 48272
rect 324590 48220 324596 48272
rect 324648 48260 324654 48272
rect 324774 48260 324780 48272
rect 324648 48232 324780 48260
rect 324648 48220 324654 48232
rect 324774 48220 324780 48232
rect 324832 48220 324838 48272
rect 92842 48192 92848 48204
rect 92768 48164 92848 48192
rect 92842 48152 92848 48164
rect 92900 48152 92906 48204
rect 96982 47036 96988 47048
rect 96943 47008 96988 47036
rect 96982 46996 96988 47008
rect 97040 46996 97046 47048
rect 90910 46928 90916 46980
rect 90968 46968 90974 46980
rect 91002 46968 91008 46980
rect 90968 46940 91008 46968
rect 90968 46928 90974 46940
rect 91002 46928 91008 46940
rect 91060 46928 91066 46980
rect 104894 46928 104900 46980
rect 104952 46968 104958 46980
rect 105262 46968 105268 46980
rect 104952 46940 105268 46968
rect 104952 46928 104958 46940
rect 105262 46928 105268 46940
rect 105320 46928 105326 46980
rect 242526 46968 242532 46980
rect 242487 46940 242532 46968
rect 242526 46928 242532 46940
rect 242584 46928 242590 46980
rect 72053 46903 72111 46909
rect 72053 46869 72065 46903
rect 72099 46900 72111 46903
rect 72234 46900 72240 46912
rect 72099 46872 72240 46900
rect 72099 46869 72111 46872
rect 72053 46863 72111 46869
rect 72234 46860 72240 46872
rect 72292 46860 72298 46912
rect 73433 46903 73491 46909
rect 73433 46869 73445 46903
rect 73479 46900 73491 46903
rect 73522 46900 73528 46912
rect 73479 46872 73528 46900
rect 73479 46869 73491 46872
rect 73433 46863 73491 46869
rect 73522 46860 73528 46872
rect 73580 46860 73586 46912
rect 96982 46900 96988 46912
rect 96943 46872 96988 46900
rect 96982 46860 96988 46872
rect 97040 46860 97046 46912
rect 193858 46900 193864 46912
rect 193819 46872 193864 46900
rect 193858 46860 193864 46872
rect 193916 46860 193922 46912
rect 204898 46900 204904 46912
rect 204859 46872 204904 46900
rect 204898 46860 204904 46872
rect 204956 46860 204962 46912
rect 234062 46900 234068 46912
rect 234023 46872 234068 46900
rect 234062 46860 234068 46872
rect 234120 46860 234126 46912
rect 246942 46900 246948 46912
rect 246903 46872 246948 46900
rect 246942 46860 246948 46872
rect 247000 46860 247006 46912
rect 250990 46900 250996 46912
rect 250951 46872 250996 46900
rect 250990 46860 250996 46872
rect 251048 46860 251054 46912
rect 252278 46900 252284 46912
rect 252239 46872 252284 46900
rect 252278 46860 252284 46872
rect 252336 46860 252342 46912
rect 255222 46900 255228 46912
rect 255183 46872 255228 46900
rect 255222 46860 255228 46872
rect 255280 46860 255286 46912
rect 259270 46900 259276 46912
rect 259231 46872 259276 46900
rect 259270 46860 259276 46872
rect 259328 46860 259334 46912
rect 324590 46860 324596 46912
rect 324648 46900 324654 46912
rect 324869 46903 324927 46909
rect 324869 46900 324881 46903
rect 324648 46872 324881 46900
rect 324648 46860 324654 46872
rect 324869 46869 324881 46872
rect 324915 46869 324927 46903
rect 324869 46863 324927 46869
rect 91002 46792 91008 46844
rect 91060 46832 91066 46844
rect 91186 46832 91192 46844
rect 91060 46804 91192 46832
rect 91060 46792 91066 46804
rect 91186 46792 91192 46804
rect 91244 46792 91250 46844
rect 268746 46180 268752 46232
rect 268804 46220 268810 46232
rect 269022 46220 269028 46232
rect 268804 46192 269028 46220
rect 268804 46180 268810 46192
rect 269022 46180 269028 46192
rect 269080 46180 269086 46232
rect 264606 44316 264612 44328
rect 264567 44288 264612 44316
rect 264606 44276 264612 44288
rect 264664 44276 264670 44328
rect 267274 44112 267280 44124
rect 267235 44084 267280 44112
rect 267274 44072 267280 44084
rect 267332 44072 267338 44124
rect 70486 41352 70492 41404
rect 70544 41392 70550 41404
rect 70670 41392 70676 41404
rect 70544 41364 70676 41392
rect 70544 41352 70550 41364
rect 70670 41352 70676 41364
rect 70728 41352 70734 41404
rect 70578 41284 70584 41336
rect 70636 41324 70642 41336
rect 70762 41324 70768 41336
rect 70636 41296 70768 41324
rect 70636 41284 70642 41296
rect 70762 41284 70768 41296
rect 70820 41284 70826 41336
rect 89990 41284 89996 41336
rect 90048 41284 90054 41336
rect 104894 41284 104900 41336
rect 104952 41324 104958 41336
rect 105170 41324 105176 41336
rect 104952 41296 105176 41324
rect 104952 41284 104958 41296
rect 105170 41284 105176 41296
rect 105228 41284 105234 41336
rect 90008 41200 90036 41284
rect 89990 41148 89996 41200
rect 90048 41148 90054 41200
rect 77386 38700 77392 38752
rect 77444 38700 77450 38752
rect 77404 38616 77432 38700
rect 78766 38672 78772 38684
rect 78727 38644 78772 38672
rect 78766 38632 78772 38644
rect 78824 38632 78830 38684
rect 81713 38675 81771 38681
rect 81713 38641 81725 38675
rect 81759 38672 81771 38675
rect 81802 38672 81808 38684
rect 81759 38644 81808 38672
rect 81759 38641 81771 38644
rect 81713 38635 81771 38641
rect 81802 38632 81808 38644
rect 81860 38632 81866 38684
rect 151078 38672 151084 38684
rect 151039 38644 151084 38672
rect 151078 38632 151084 38644
rect 151136 38632 151142 38684
rect 234062 38672 234068 38684
rect 234023 38644 234068 38672
rect 234062 38632 234068 38644
rect 234120 38632 234126 38684
rect 77386 38564 77392 38616
rect 77444 38564 77450 38616
rect 106826 38604 106832 38616
rect 106787 38576 106832 38604
rect 106826 38564 106832 38576
rect 106884 38564 106890 38616
rect 211893 38607 211951 38613
rect 211893 38573 211905 38607
rect 211939 38604 211951 38607
rect 211982 38604 211988 38616
rect 211939 38576 211988 38604
rect 211939 38573 211951 38576
rect 211893 38567 211951 38573
rect 211982 38564 211988 38576
rect 212040 38564 212046 38616
rect 235718 38604 235724 38616
rect 235679 38576 235724 38604
rect 235718 38564 235724 38576
rect 235776 38564 235782 38616
rect 324866 38536 324872 38548
rect 324827 38508 324872 38536
rect 324866 38496 324872 38508
rect 324924 38496 324930 38548
rect 72050 37312 72056 37324
rect 72011 37284 72056 37312
rect 72050 37272 72056 37284
rect 72108 37272 72114 37324
rect 73430 37312 73436 37324
rect 73391 37284 73436 37312
rect 73430 37272 73436 37284
rect 73488 37272 73494 37324
rect 78766 37312 78772 37324
rect 78727 37284 78772 37312
rect 78766 37272 78772 37284
rect 78824 37272 78830 37324
rect 96982 37312 96988 37324
rect 96943 37284 96988 37312
rect 96982 37272 96988 37284
rect 97040 37272 97046 37324
rect 204898 37312 204904 37324
rect 204859 37284 204904 37312
rect 204898 37272 204904 37284
rect 204956 37272 204962 37324
rect 243630 37272 243636 37324
rect 243688 37312 243694 37324
rect 243814 37312 243820 37324
rect 243688 37284 243820 37312
rect 243688 37272 243694 37284
rect 243814 37272 243820 37284
rect 243872 37272 243878 37324
rect 246942 37312 246948 37324
rect 246903 37284 246948 37312
rect 246942 37272 246948 37284
rect 247000 37272 247006 37324
rect 250990 37312 250996 37324
rect 250951 37284 250996 37312
rect 250990 37272 250996 37284
rect 251048 37272 251054 37324
rect 252278 37312 252284 37324
rect 252239 37284 252284 37312
rect 252278 37272 252284 37284
rect 252336 37272 252342 37324
rect 255222 37312 255228 37324
rect 255183 37284 255228 37312
rect 255222 37272 255228 37284
rect 255280 37272 255286 37324
rect 259270 37312 259276 37324
rect 259231 37284 259276 37312
rect 259270 37272 259276 37284
rect 259328 37272 259334 37324
rect 242526 37244 242532 37256
rect 242487 37216 242532 37244
rect 242526 37204 242532 37216
rect 242584 37204 242590 37256
rect 73430 36292 73436 36304
rect 73391 36264 73436 36292
rect 73430 36252 73436 36264
rect 73488 36252 73494 36304
rect 267277 35819 267335 35825
rect 267277 35785 267289 35819
rect 267323 35816 267335 35819
rect 267366 35816 267372 35828
rect 267323 35788 267372 35816
rect 267323 35785 267335 35788
rect 267277 35779 267335 35785
rect 267366 35776 267372 35788
rect 267424 35776 267430 35828
rect 70486 33804 70492 33856
rect 70544 33844 70550 33856
rect 70670 33844 70676 33856
rect 70544 33816 70676 33844
rect 70544 33804 70550 33816
rect 70670 33804 70676 33816
rect 70728 33804 70734 33856
rect 262030 33232 262036 33244
rect 261864 33204 262036 33232
rect 261864 33164 261892 33204
rect 262030 33192 262036 33204
rect 262088 33192 262094 33244
rect 264422 33192 264428 33244
rect 264480 33232 264486 33244
rect 264606 33232 264612 33244
rect 264480 33204 264612 33232
rect 264480 33192 264486 33204
rect 264606 33192 264612 33204
rect 264664 33192 264670 33244
rect 261941 33167 261999 33173
rect 261941 33164 261953 33167
rect 261864 33136 261953 33164
rect 261941 33133 261953 33136
rect 261987 33133 261999 33167
rect 261941 33127 261999 33133
rect 268746 32172 268752 32224
rect 268804 32212 268810 32224
rect 269022 32212 269028 32224
rect 268804 32184 269028 32212
rect 268804 32172 268810 32184
rect 269022 32172 269028 32184
rect 269080 32172 269086 32224
rect 70762 31804 70768 31816
rect 70688 31776 70768 31804
rect 70688 31748 70716 31776
rect 70762 31764 70768 31776
rect 70820 31764 70826 31816
rect 94130 31764 94136 31816
rect 94188 31764 94194 31816
rect 105170 31804 105176 31816
rect 105096 31776 105176 31804
rect 70670 31696 70676 31748
rect 70728 31696 70734 31748
rect 94148 31612 94176 31764
rect 105096 31748 105124 31776
rect 105170 31764 105176 31776
rect 105228 31764 105234 31816
rect 324866 31764 324872 31816
rect 324924 31764 324930 31816
rect 105078 31696 105084 31748
rect 105136 31696 105142 31748
rect 227254 31696 227260 31748
rect 227312 31736 227318 31748
rect 227438 31736 227444 31748
rect 227312 31708 227444 31736
rect 227312 31696 227318 31708
rect 227438 31696 227444 31708
rect 227496 31696 227502 31748
rect 324884 31680 324912 31764
rect 324866 31628 324872 31680
rect 324924 31628 324930 31680
rect 94130 31560 94136 31612
rect 94188 31560 94194 31612
rect 106826 31600 106832 31612
rect 106787 31572 106832 31600
rect 106826 31560 106832 31572
rect 106884 31560 106890 31612
rect 261941 29699 261999 29705
rect 261941 29665 261953 29699
rect 261987 29696 261999 29699
rect 262030 29696 262036 29708
rect 261987 29668 262036 29696
rect 261987 29665 261999 29668
rect 261941 29659 261999 29665
rect 262030 29656 262036 29668
rect 262088 29656 262094 29708
rect 84654 29084 84660 29096
rect 84580 29056 84660 29084
rect 84580 29028 84608 29056
rect 84654 29044 84660 29056
rect 84712 29044 84718 29096
rect 72050 28976 72056 29028
rect 72108 29016 72114 29028
rect 72234 29016 72240 29028
rect 72108 28988 72240 29016
rect 72108 28976 72114 28988
rect 72234 28976 72240 28988
rect 72292 28976 72298 29028
rect 73433 29019 73491 29025
rect 73433 28985 73445 29019
rect 73479 29016 73491 29019
rect 73522 29016 73528 29028
rect 73479 28988 73528 29016
rect 73479 28985 73491 28988
rect 73433 28979 73491 28985
rect 73522 28976 73528 28988
rect 73580 28976 73586 29028
rect 84562 28976 84568 29028
rect 84620 28976 84626 29028
rect 91002 28976 91008 29028
rect 91060 29016 91066 29028
rect 91186 29016 91192 29028
rect 91060 28988 91192 29016
rect 91060 28976 91066 28988
rect 91186 28976 91192 28988
rect 91244 28976 91250 29028
rect 193861 29019 193919 29025
rect 193861 28985 193873 29019
rect 193907 29016 193919 29019
rect 193950 29016 193956 29028
rect 193907 28988 193956 29016
rect 193907 28985 193919 28988
rect 193861 28979 193919 28985
rect 193950 28976 193956 28988
rect 194008 28976 194014 29028
rect 211890 29016 211896 29028
rect 211851 28988 211896 29016
rect 211890 28976 211896 28988
rect 211948 28976 211954 29028
rect 235718 29016 235724 29028
rect 235679 28988 235724 29016
rect 235718 28976 235724 28988
rect 235776 28976 235782 29028
rect 89990 28948 89996 28960
rect 89951 28920 89996 28948
rect 89990 28908 89996 28920
rect 90048 28908 90054 28960
rect 96982 28948 96988 28960
rect 96943 28920 96988 28948
rect 96982 28908 96988 28920
rect 97040 28908 97046 28960
rect 151078 28948 151084 28960
rect 151039 28920 151084 28948
rect 151078 28908 151084 28920
rect 151136 28908 151142 28960
rect 92842 27724 92848 27736
rect 92768 27696 92848 27724
rect 92768 27668 92796 27696
rect 92842 27684 92848 27696
rect 92900 27684 92906 27736
rect 92750 27616 92756 27668
rect 92808 27616 92814 27668
rect 242526 27656 242532 27668
rect 242487 27628 242532 27656
rect 242526 27616 242532 27628
rect 242584 27616 242590 27668
rect 77478 27588 77484 27600
rect 77439 27560 77484 27588
rect 77478 27548 77484 27560
rect 77536 27548 77542 27600
rect 78861 27591 78919 27597
rect 78861 27557 78873 27591
rect 78907 27588 78919 27591
rect 78950 27588 78956 27600
rect 78907 27560 78956 27588
rect 78907 27557 78919 27560
rect 78861 27551 78919 27557
rect 78950 27548 78956 27560
rect 79008 27548 79014 27600
rect 91002 27548 91008 27600
rect 91060 27588 91066 27600
rect 91097 27591 91155 27597
rect 91097 27588 91109 27591
rect 91060 27560 91109 27588
rect 91060 27548 91066 27560
rect 91097 27557 91109 27560
rect 91143 27557 91155 27591
rect 204898 27588 204904 27600
rect 204859 27560 204904 27588
rect 91097 27551 91155 27557
rect 204898 27548 204904 27560
rect 204956 27548 204962 27600
rect 248230 27588 248236 27600
rect 248191 27560 248236 27588
rect 248230 27548 248236 27560
rect 248288 27548 248294 27600
rect 249610 27588 249616 27600
rect 249571 27560 249616 27588
rect 249610 27548 249616 27560
rect 249668 27548 249674 27600
rect 255222 27588 255228 27600
rect 255183 27560 255228 27588
rect 255222 27548 255228 27560
rect 255280 27548 255286 27600
rect 268746 26868 268752 26920
rect 268804 26908 268810 26920
rect 269022 26908 269028 26920
rect 268804 26880 269028 26908
rect 268804 26868 268810 26880
rect 269022 26868 269028 26880
rect 269080 26868 269086 26920
rect 260377 26231 260435 26237
rect 260377 26197 260389 26231
rect 260423 26228 260435 26231
rect 260466 26228 260472 26240
rect 260423 26200 260472 26228
rect 260423 26197 260435 26200
rect 260377 26191 260435 26197
rect 260466 26188 260472 26200
rect 260524 26188 260530 26240
rect 264422 24828 264428 24880
rect 264480 24868 264486 24880
rect 264698 24868 264704 24880
rect 264480 24840 264704 24868
rect 264480 24828 264486 24840
rect 264698 24828 264704 24840
rect 264756 24828 264762 24880
rect 262030 23332 262036 23384
rect 262088 23372 262094 23384
rect 262214 23372 262220 23384
rect 262088 23344 262220 23372
rect 262088 23332 262094 23344
rect 262214 23332 262220 23344
rect 262272 23332 262278 23384
rect 259178 22760 259184 22772
rect 259139 22732 259184 22760
rect 259178 22720 259184 22732
rect 259236 22720 259242 22772
rect 70486 22652 70492 22704
rect 70544 22692 70550 22704
rect 70670 22692 70676 22704
rect 70544 22664 70676 22692
rect 70544 22652 70550 22664
rect 70670 22652 70676 22664
rect 70728 22652 70734 22704
rect 72234 22148 72240 22160
rect 72160 22120 72240 22148
rect 72160 22092 72188 22120
rect 72234 22108 72240 22120
rect 72292 22108 72298 22160
rect 72142 22040 72148 22092
rect 72200 22040 72206 22092
rect 96982 21944 96988 21956
rect 96943 21916 96988 21944
rect 96982 21904 96988 21916
rect 97040 21904 97046 21956
rect 250806 19864 250812 19916
rect 250864 19904 250870 19916
rect 250990 19904 250996 19916
rect 250864 19876 250996 19904
rect 250864 19864 250870 19876
rect 250990 19864 250996 19876
rect 251048 19864 251054 19916
rect 89990 19360 89996 19372
rect 89951 19332 89996 19360
rect 89990 19320 89996 19332
rect 90048 19320 90054 19372
rect 151078 19360 151084 19372
rect 151039 19332 151084 19360
rect 151078 19320 151084 19332
rect 151136 19320 151142 19372
rect 193766 19292 193772 19304
rect 193727 19264 193772 19292
rect 193766 19252 193772 19264
rect 193824 19252 193830 19304
rect 227346 19292 227352 19304
rect 227307 19264 227352 19292
rect 227346 19252 227352 19264
rect 227404 19252 227410 19304
rect 234338 19252 234344 19304
rect 234396 19292 234402 19304
rect 234614 19292 234620 19304
rect 234396 19264 234620 19292
rect 234396 19252 234402 19264
rect 234614 19252 234620 19264
rect 234672 19252 234678 19304
rect 235718 19292 235724 19304
rect 235679 19264 235724 19292
rect 235718 19252 235724 19264
rect 235776 19252 235782 19304
rect 245286 19252 245292 19304
rect 245344 19292 245350 19304
rect 245562 19292 245568 19304
rect 245344 19264 245568 19292
rect 245344 19252 245350 19264
rect 245562 19252 245568 19264
rect 245620 19252 245626 19304
rect 77478 18000 77484 18012
rect 77439 17972 77484 18000
rect 77478 17960 77484 17972
rect 77536 17960 77542 18012
rect 78858 18000 78864 18012
rect 78819 17972 78864 18000
rect 78858 17960 78864 17972
rect 78916 17960 78922 18012
rect 91002 17960 91008 18012
rect 91060 18000 91066 18012
rect 91097 18003 91155 18009
rect 91097 18000 91109 18003
rect 91060 17972 91109 18000
rect 91060 17960 91066 17972
rect 91097 17969 91109 17972
rect 91143 17969 91155 18003
rect 204898 18000 204904 18012
rect 204859 17972 204904 18000
rect 91097 17963 91155 17969
rect 204898 17960 204904 17972
rect 204956 17960 204962 18012
rect 243722 17960 243728 18012
rect 243780 18000 243786 18012
rect 243814 18000 243820 18012
rect 243780 17972 243820 18000
rect 243780 17960 243786 17972
rect 243814 17960 243820 17972
rect 243872 17960 243878 18012
rect 248230 18000 248236 18012
rect 248191 17972 248236 18000
rect 248230 17960 248236 17972
rect 248288 17960 248294 18012
rect 249610 18000 249616 18012
rect 249571 17972 249616 18000
rect 249610 17960 249616 17972
rect 249668 17960 249674 18012
rect 255222 18000 255228 18012
rect 255183 17972 255228 18000
rect 255222 17960 255228 17972
rect 255280 17960 255286 18012
rect 73341 17935 73399 17941
rect 73341 17901 73353 17935
rect 73387 17932 73399 17935
rect 73430 17932 73436 17944
rect 73387 17904 73436 17932
rect 73387 17901 73399 17904
rect 73341 17895 73399 17901
rect 73430 17892 73436 17904
rect 73488 17892 73494 17944
rect 268746 17212 268752 17264
rect 268804 17252 268810 17264
rect 269022 17252 269028 17264
rect 268804 17224 269028 17252
rect 268804 17212 268810 17224
rect 269022 17212 269028 17224
rect 269080 17212 269086 17264
rect 248230 17076 248236 17128
rect 248288 17116 248294 17128
rect 248414 17116 248420 17128
rect 248288 17088 248420 17116
rect 248288 17076 248294 17088
rect 248414 17076 248420 17088
rect 248472 17076 248478 17128
rect 219066 16532 219072 16584
rect 219124 16572 219130 16584
rect 219342 16572 219348 16584
rect 219124 16544 219348 16572
rect 219124 16532 219130 16544
rect 219342 16532 219348 16544
rect 219400 16532 219406 16584
rect 169478 16396 169484 16448
rect 169536 16436 169542 16448
rect 285674 16436 285680 16448
rect 169536 16408 285680 16436
rect 169536 16396 169542 16408
rect 285674 16396 285680 16408
rect 285732 16396 285738 16448
rect 170858 16328 170864 16380
rect 170916 16368 170922 16380
rect 288434 16368 288440 16380
rect 170916 16340 288440 16368
rect 170916 16328 170922 16340
rect 288434 16328 288440 16340
rect 288492 16328 288498 16380
rect 172146 16260 172152 16312
rect 172204 16300 172210 16312
rect 292574 16300 292580 16312
rect 172204 16272 292580 16300
rect 172204 16260 172210 16272
rect 292574 16260 292580 16272
rect 292632 16260 292638 16312
rect 173618 16192 173624 16244
rect 173676 16232 173682 16244
rect 296714 16232 296720 16244
rect 173676 16204 296720 16232
rect 173676 16192 173682 16204
rect 296714 16192 296720 16204
rect 296772 16192 296778 16244
rect 176286 16124 176292 16176
rect 176344 16164 176350 16176
rect 303614 16164 303620 16176
rect 176344 16136 303620 16164
rect 176344 16124 176350 16136
rect 303614 16124 303620 16136
rect 303672 16124 303678 16176
rect 206738 16056 206744 16108
rect 206796 16096 206802 16108
rect 391934 16096 391940 16108
rect 206796 16068 391940 16096
rect 206796 16056 206802 16068
rect 391934 16056 391940 16068
rect 391992 16056 391998 16108
rect 212258 15988 212264 16040
rect 212316 16028 212322 16040
rect 407114 16028 407120 16040
rect 212316 16000 407120 16028
rect 212316 15988 212322 16000
rect 407114 15988 407120 16000
rect 407172 15988 407178 16040
rect 216306 15920 216312 15972
rect 216364 15960 216370 15972
rect 420914 15960 420920 15972
rect 216364 15932 420920 15960
rect 216364 15920 216370 15932
rect 420914 15920 420920 15932
rect 420972 15920 420978 15972
rect 235721 15895 235779 15901
rect 235721 15861 235733 15895
rect 235767 15892 235779 15895
rect 477494 15892 477500 15904
rect 235767 15864 477500 15892
rect 235767 15861 235779 15864
rect 235721 15855 235779 15861
rect 477494 15852 477500 15864
rect 477552 15852 477558 15904
rect 202782 15104 202788 15156
rect 202840 15144 202846 15156
rect 379514 15144 379520 15156
rect 202840 15116 379520 15144
rect 202840 15104 202846 15116
rect 379514 15104 379520 15116
rect 379572 15104 379578 15156
rect 204070 15036 204076 15088
rect 204128 15076 204134 15088
rect 382366 15076 382372 15088
rect 204128 15048 382372 15076
rect 204128 15036 204134 15048
rect 382366 15036 382372 15048
rect 382424 15036 382430 15088
rect 202690 14968 202696 15020
rect 202748 15008 202754 15020
rect 380894 15008 380900 15020
rect 202748 14980 380900 15008
rect 202748 14968 202754 14980
rect 380894 14968 380900 14980
rect 380952 14968 380958 15020
rect 203886 14900 203892 14952
rect 203944 14940 203950 14952
rect 383654 14940 383660 14952
rect 203944 14912 383660 14940
rect 203944 14900 203950 14912
rect 383654 14900 383660 14912
rect 383712 14900 383718 14952
rect 205450 14832 205456 14884
rect 205508 14872 205514 14884
rect 387794 14872 387800 14884
rect 205508 14844 387800 14872
rect 205508 14832 205514 14844
rect 387794 14832 387800 14844
rect 387852 14832 387858 14884
rect 203978 14764 203984 14816
rect 204036 14804 204042 14816
rect 386414 14804 386420 14816
rect 204036 14776 386420 14804
rect 204036 14764 204042 14776
rect 386414 14764 386420 14776
rect 386472 14764 386478 14816
rect 206830 14696 206836 14748
rect 206888 14736 206894 14748
rect 390554 14736 390560 14748
rect 206888 14708 390560 14736
rect 206888 14696 206894 14708
rect 390554 14696 390560 14708
rect 390612 14696 390618 14748
rect 237098 14628 237104 14680
rect 237156 14668 237162 14680
rect 478874 14668 478880 14680
rect 237156 14640 478880 14668
rect 237156 14628 237162 14640
rect 478874 14628 478880 14640
rect 478932 14628 478938 14680
rect 238570 14560 238576 14612
rect 238628 14600 238634 14612
rect 484394 14600 484400 14612
rect 238628 14572 484400 14600
rect 238628 14560 238634 14572
rect 484394 14560 484400 14572
rect 484452 14560 484458 14612
rect 238386 14492 238392 14544
rect 238444 14532 238450 14544
rect 485774 14532 485780 14544
rect 238444 14504 485780 14532
rect 238444 14492 238450 14504
rect 485774 14492 485780 14504
rect 485832 14492 485838 14544
rect 239674 14424 239680 14476
rect 239732 14464 239738 14476
rect 487154 14464 487160 14476
rect 239732 14436 487160 14464
rect 239732 14424 239738 14436
rect 487154 14424 487160 14436
rect 487212 14424 487218 14476
rect 201218 14356 201224 14408
rect 201276 14396 201282 14408
rect 375374 14396 375380 14408
rect 201276 14368 375380 14396
rect 201276 14356 201282 14368
rect 375374 14356 375380 14368
rect 375432 14356 375438 14408
rect 170950 14288 170956 14340
rect 171008 14328 171014 14340
rect 287054 14328 287060 14340
rect 171008 14300 287060 14328
rect 171008 14288 171014 14300
rect 287054 14288 287060 14300
rect 287112 14288 287118 14340
rect 169570 14220 169576 14272
rect 169628 14260 169634 14272
rect 284294 14260 284300 14272
rect 169628 14232 284300 14260
rect 169628 14220 169634 14232
rect 284294 14220 284300 14232
rect 284352 14220 284358 14272
rect 168190 14152 168196 14204
rect 168248 14192 168254 14204
rect 282914 14192 282920 14204
rect 168248 14164 282920 14192
rect 168248 14152 168254 14164
rect 282914 14152 282920 14164
rect 282972 14152 282978 14204
rect 168006 14084 168012 14136
rect 168064 14124 168070 14136
rect 281534 14124 281540 14136
rect 168064 14096 281540 14124
rect 168064 14084 168070 14096
rect 281534 14084 281540 14096
rect 281592 14084 281598 14136
rect 166718 14016 166724 14068
rect 166776 14056 166782 14068
rect 278866 14056 278872 14068
rect 166776 14028 278872 14056
rect 166776 14016 166782 14028
rect 278866 14016 278872 14028
rect 278924 14016 278930 14068
rect 168282 13948 168288 14000
rect 168340 13988 168346 14000
rect 280154 13988 280160 14000
rect 168340 13960 280160 13988
rect 168340 13948 168346 13960
rect 280154 13948 280160 13960
rect 280212 13948 280218 14000
rect 168098 13880 168104 13932
rect 168156 13920 168162 13932
rect 278774 13920 278780 13932
rect 168156 13892 278780 13920
rect 168156 13880 168162 13892
rect 278774 13880 278780 13892
rect 278832 13880 278838 13932
rect 166810 13812 166816 13864
rect 166868 13852 166874 13864
rect 277394 13852 277400 13864
rect 166868 13824 277400 13852
rect 166868 13812 166874 13824
rect 277394 13812 277400 13824
rect 277452 13812 277458 13864
rect 248138 13744 248144 13796
rect 248196 13784 248202 13796
rect 510614 13784 510620 13796
rect 248196 13756 510620 13784
rect 248196 13744 248202 13756
rect 510614 13744 510620 13756
rect 510672 13744 510678 13796
rect 248046 13676 248052 13728
rect 248104 13716 248110 13728
rect 513374 13716 513380 13728
rect 248104 13688 513380 13716
rect 248104 13676 248110 13688
rect 513374 13676 513380 13688
rect 513432 13676 513438 13728
rect 249518 13608 249524 13660
rect 249576 13648 249582 13660
rect 517514 13648 517520 13660
rect 249576 13620 517520 13648
rect 249576 13608 249582 13620
rect 517514 13608 517520 13620
rect 517572 13608 517578 13660
rect 250898 13540 250904 13592
rect 250956 13580 250962 13592
rect 520274 13580 520280 13592
rect 250956 13552 520280 13580
rect 250956 13540 250962 13552
rect 520274 13540 520280 13552
rect 520332 13540 520338 13592
rect 252186 13472 252192 13524
rect 252244 13512 252250 13524
rect 524414 13512 524420 13524
rect 252244 13484 524420 13512
rect 252244 13472 252250 13484
rect 524414 13472 524420 13484
rect 524472 13472 524478 13524
rect 253658 13404 253664 13456
rect 253716 13444 253722 13456
rect 528554 13444 528560 13456
rect 253716 13416 528560 13444
rect 253716 13404 253722 13416
rect 528554 13404 528560 13416
rect 528612 13404 528618 13456
rect 255038 13336 255044 13388
rect 255096 13376 255102 13388
rect 531314 13376 531320 13388
rect 255096 13348 531320 13376
rect 255096 13336 255102 13348
rect 531314 13336 531320 13348
rect 531372 13336 531378 13388
rect 256326 13268 256332 13320
rect 256384 13308 256390 13320
rect 535454 13308 535460 13320
rect 256384 13280 535460 13308
rect 256384 13268 256390 13280
rect 535454 13268 535460 13280
rect 535512 13268 535518 13320
rect 257798 13200 257804 13252
rect 257856 13240 257862 13252
rect 538214 13240 538220 13252
rect 257856 13212 538220 13240
rect 257856 13200 257862 13212
rect 538214 13200 538220 13212
rect 538272 13200 538278 13252
rect 259181 13175 259239 13181
rect 259181 13141 259193 13175
rect 259227 13172 259239 13175
rect 542354 13172 542360 13184
rect 259227 13144 542360 13172
rect 259227 13141 259239 13144
rect 259181 13135 259239 13141
rect 542354 13132 542360 13144
rect 542412 13132 542418 13184
rect 255130 13104 255136 13116
rect 255091 13076 255136 13104
rect 255130 13064 255136 13076
rect 255188 13064 255194 13116
rect 260377 13107 260435 13113
rect 260377 13073 260389 13107
rect 260423 13104 260435 13107
rect 546494 13104 546500 13116
rect 260423 13076 546500 13104
rect 260423 13073 260435 13076
rect 260377 13067 260435 13073
rect 546494 13064 546500 13076
rect 546552 13064 546558 13116
rect 246758 12996 246764 13048
rect 246816 13036 246822 13048
rect 506474 13036 506480 13048
rect 246816 13008 506480 13036
rect 246816 12996 246822 13008
rect 506474 12996 506480 13008
rect 506532 12996 506538 13048
rect 245378 12928 245384 12980
rect 245436 12968 245442 12980
rect 502334 12968 502340 12980
rect 245436 12940 502340 12968
rect 245436 12928 245442 12940
rect 502334 12928 502340 12940
rect 502392 12928 502398 12980
rect 243814 12860 243820 12912
rect 243872 12900 243878 12912
rect 499574 12900 499580 12912
rect 243872 12872 499580 12900
rect 243872 12860 243878 12872
rect 499574 12860 499580 12872
rect 499632 12860 499638 12912
rect 242434 12792 242440 12844
rect 242492 12832 242498 12844
rect 495434 12832 495440 12844
rect 242492 12804 495440 12832
rect 242492 12792 242498 12804
rect 495434 12792 495440 12804
rect 495492 12792 495498 12844
rect 241146 12724 241152 12776
rect 241204 12764 241210 12776
rect 492674 12764 492680 12776
rect 241204 12736 492680 12764
rect 241204 12724 241210 12736
rect 492674 12724 492680 12736
rect 492732 12724 492738 12776
rect 240042 12656 240048 12708
rect 240100 12696 240106 12708
rect 488534 12696 488540 12708
rect 240100 12668 488540 12696
rect 240100 12656 240106 12668
rect 488534 12656 488540 12668
rect 488592 12656 488598 12708
rect 239950 12588 239956 12640
rect 240008 12628 240014 12640
rect 485866 12628 485872 12640
rect 240008 12600 485872 12628
rect 240008 12588 240014 12600
rect 485866 12588 485872 12600
rect 485924 12588 485930 12640
rect 70670 12560 70676 12572
rect 70504 12532 70676 12560
rect 70504 12504 70532 12532
rect 70670 12520 70676 12532
rect 70728 12520 70734 12572
rect 238662 12520 238668 12572
rect 238720 12560 238726 12572
rect 483014 12560 483020 12572
rect 238720 12532 483020 12560
rect 238720 12520 238726 12532
rect 483014 12520 483020 12532
rect 483072 12520 483078 12572
rect 70486 12452 70492 12504
rect 70544 12452 70550 12504
rect 91002 12492 91008 12504
rect 90928 12464 91008 12492
rect 90928 12436 90956 12464
rect 91002 12452 91008 12464
rect 91060 12452 91066 12504
rect 94130 12452 94136 12504
rect 94188 12452 94194 12504
rect 165338 12452 165344 12504
rect 165396 12492 165402 12504
rect 271874 12492 271880 12504
rect 165396 12464 271880 12492
rect 165396 12452 165402 12464
rect 271874 12452 271880 12464
rect 271932 12452 271938 12504
rect 90910 12384 90916 12436
rect 90968 12384 90974 12436
rect 94148 12356 94176 12452
rect 193766 12424 193772 12436
rect 193727 12396 193772 12424
rect 193766 12384 193772 12396
rect 193824 12384 193830 12436
rect 217870 12384 217876 12436
rect 217928 12424 217934 12436
rect 423674 12424 423680 12436
rect 217928 12396 423680 12424
rect 217928 12384 217934 12396
rect 423674 12384 423680 12396
rect 423732 12384 423738 12436
rect 94222 12356 94228 12368
rect 94148 12328 94228 12356
rect 94222 12316 94228 12328
rect 94280 12316 94286 12368
rect 219158 12316 219164 12368
rect 219216 12356 219222 12368
rect 426434 12356 426440 12368
rect 219216 12328 426440 12356
rect 219216 12316 219222 12328
rect 426434 12316 426440 12328
rect 426492 12316 426498 12368
rect 220538 12248 220544 12300
rect 220596 12288 220602 12300
rect 430574 12288 430580 12300
rect 220596 12260 430580 12288
rect 220596 12248 220602 12260
rect 430574 12248 430580 12260
rect 430632 12248 430638 12300
rect 220630 12180 220636 12232
rect 220688 12220 220694 12232
rect 433334 12220 433340 12232
rect 220688 12192 433340 12220
rect 220688 12180 220694 12192
rect 433334 12180 433340 12192
rect 433392 12180 433398 12232
rect 221918 12112 221924 12164
rect 221976 12152 221982 12164
rect 437474 12152 437480 12164
rect 221976 12124 437480 12152
rect 221976 12112 221982 12124
rect 437474 12112 437480 12124
rect 437532 12112 437538 12164
rect 223390 12044 223396 12096
rect 223448 12084 223454 12096
rect 441614 12084 441620 12096
rect 223448 12056 441620 12084
rect 223448 12044 223454 12056
rect 441614 12044 441620 12056
rect 441672 12044 441678 12096
rect 224678 11976 224684 12028
rect 224736 12016 224742 12028
rect 444374 12016 444380 12028
rect 224736 11988 444380 12016
rect 224736 11976 224742 11988
rect 444374 11976 444380 11988
rect 444432 11976 444438 12028
rect 226058 11908 226064 11960
rect 226116 11948 226122 11960
rect 448514 11948 448520 11960
rect 226116 11920 448520 11948
rect 226116 11908 226122 11920
rect 448514 11908 448520 11920
rect 448572 11908 448578 11960
rect 227349 11883 227407 11889
rect 227349 11849 227361 11883
rect 227395 11880 227407 11883
rect 451274 11880 451280 11892
rect 227395 11852 451280 11880
rect 227395 11849 227407 11852
rect 227349 11843 227407 11849
rect 451274 11840 451280 11852
rect 451332 11840 451338 11892
rect 228818 11772 228824 11824
rect 228876 11812 228882 11824
rect 455414 11812 455420 11824
rect 228876 11784 455420 11812
rect 228876 11772 228882 11784
rect 455414 11772 455420 11784
rect 455472 11772 455478 11824
rect 230290 11704 230296 11756
rect 230348 11744 230354 11756
rect 459646 11744 459652 11756
rect 230348 11716 459652 11744
rect 230348 11704 230354 11716
rect 459646 11704 459652 11716
rect 459704 11704 459710 11756
rect 216398 11636 216404 11688
rect 216456 11676 216462 11688
rect 419534 11676 419540 11688
rect 216456 11648 419540 11676
rect 216456 11636 216462 11648
rect 419534 11636 419540 11648
rect 419592 11636 419598 11688
rect 215110 11568 215116 11620
rect 215168 11608 215174 11620
rect 416866 11608 416872 11620
rect 215168 11580 416872 11608
rect 215168 11568 215174 11580
rect 416866 11568 416872 11580
rect 416924 11568 416930 11620
rect 213638 11500 213644 11552
rect 213696 11540 213702 11552
rect 412634 11540 412640 11552
rect 213696 11512 412640 11540
rect 213696 11500 213702 11512
rect 412634 11500 412640 11512
rect 412692 11500 412698 11552
rect 212350 11432 212356 11484
rect 212408 11472 212414 11484
rect 408494 11472 408500 11484
rect 212408 11444 408500 11472
rect 212408 11432 212414 11444
rect 408494 11432 408500 11444
rect 408552 11432 408558 11484
rect 210970 11364 210976 11416
rect 211028 11404 211034 11416
rect 405734 11404 405740 11416
rect 211028 11376 405740 11404
rect 211028 11364 211034 11376
rect 405734 11364 405740 11376
rect 405792 11364 405798 11416
rect 209590 11296 209596 11348
rect 209648 11336 209654 11348
rect 401594 11336 401600 11348
rect 209648 11308 401600 11336
rect 209648 11296 209654 11308
rect 401594 11296 401600 11308
rect 401652 11296 401658 11348
rect 208026 11228 208032 11280
rect 208084 11268 208090 11280
rect 398834 11268 398840 11280
rect 208084 11240 398840 11268
rect 208084 11228 208090 11240
rect 398834 11228 398840 11240
rect 398892 11228 398898 11280
rect 208118 11160 208124 11212
rect 208176 11200 208182 11212
rect 394694 11200 394700 11212
rect 208176 11172 394700 11200
rect 208176 11160 208182 11172
rect 394694 11160 394700 11172
rect 394752 11160 394758 11212
rect 165430 11092 165436 11144
rect 165488 11132 165494 11144
rect 274634 11132 274640 11144
rect 165488 11104 274640 11132
rect 165488 11092 165494 11104
rect 274634 11092 274640 11104
rect 274692 11092 274698 11144
rect 253658 11024 253664 11076
rect 253716 11064 253722 11076
rect 253842 11064 253848 11076
rect 253716 11036 253848 11064
rect 253716 11024 253722 11036
rect 253842 11024 253848 11036
rect 253900 11024 253906 11076
rect 255130 11064 255136 11076
rect 255091 11036 255136 11064
rect 255130 11024 255136 11036
rect 255188 11024 255194 11076
rect 183370 10956 183376 11008
rect 183428 10996 183434 11008
rect 322934 10996 322940 11008
rect 183428 10968 322940 10996
rect 183428 10956 183434 10968
rect 322934 10956 322940 10968
rect 322992 10956 322998 11008
rect 184658 10888 184664 10940
rect 184716 10928 184722 10940
rect 327074 10928 327080 10940
rect 184716 10900 327080 10928
rect 184716 10888 184722 10900
rect 327074 10888 327080 10900
rect 327132 10888 327138 10940
rect 184566 10820 184572 10872
rect 184624 10860 184630 10872
rect 331306 10860 331312 10872
rect 184624 10832 331312 10860
rect 184624 10820 184630 10832
rect 331306 10820 331312 10832
rect 331364 10820 331370 10872
rect 186130 10752 186136 10804
rect 186188 10792 186194 10804
rect 333974 10792 333980 10804
rect 186188 10764 333980 10792
rect 186188 10752 186194 10764
rect 333974 10752 333980 10764
rect 334032 10752 334038 10804
rect 187418 10684 187424 10736
rect 187476 10724 187482 10736
rect 338114 10724 338120 10736
rect 187476 10696 338120 10724
rect 187476 10684 187482 10696
rect 338114 10684 338120 10696
rect 338172 10684 338178 10736
rect 188798 10616 188804 10668
rect 188856 10656 188862 10668
rect 340874 10656 340880 10668
rect 188856 10628 340880 10656
rect 188856 10616 188862 10628
rect 340874 10616 340880 10628
rect 340932 10616 340938 10668
rect 190270 10548 190276 10600
rect 190328 10588 190334 10600
rect 345014 10588 345020 10600
rect 190328 10560 345020 10588
rect 190328 10548 190334 10560
rect 345014 10548 345020 10560
rect 345072 10548 345078 10600
rect 191558 10480 191564 10532
rect 191616 10520 191622 10532
rect 347774 10520 347780 10532
rect 191616 10492 347780 10520
rect 191616 10480 191622 10492
rect 347774 10480 347780 10492
rect 347832 10480 347838 10532
rect 192938 10412 192944 10464
rect 192996 10452 193002 10464
rect 351914 10452 351920 10464
rect 192996 10424 351920 10452
rect 192996 10412 193002 10424
rect 351914 10412 351920 10424
rect 351972 10412 351978 10464
rect 194318 10344 194324 10396
rect 194376 10384 194382 10396
rect 356146 10384 356152 10396
rect 194376 10356 356152 10384
rect 194376 10344 194382 10356
rect 356146 10344 356152 10356
rect 356204 10344 356210 10396
rect 195790 10276 195796 10328
rect 195848 10316 195854 10328
rect 358814 10316 358820 10328
rect 195848 10288 358820 10316
rect 195848 10276 195854 10288
rect 358814 10276 358820 10288
rect 358872 10276 358878 10328
rect 181898 10208 181904 10260
rect 181956 10248 181962 10260
rect 320174 10248 320180 10260
rect 181956 10220 320180 10248
rect 181956 10208 181962 10220
rect 320174 10208 320180 10220
rect 320232 10208 320238 10260
rect 180518 10140 180524 10192
rect 180576 10180 180582 10192
rect 316034 10180 316040 10192
rect 180576 10152 316040 10180
rect 180576 10140 180582 10152
rect 316034 10140 316040 10152
rect 316092 10140 316098 10192
rect 179138 10072 179144 10124
rect 179196 10112 179202 10124
rect 313366 10112 313372 10124
rect 179196 10084 313372 10112
rect 179196 10072 179202 10084
rect 313366 10072 313372 10084
rect 313424 10072 313430 10124
rect 177850 10004 177856 10056
rect 177908 10044 177914 10056
rect 309134 10044 309140 10056
rect 177908 10016 309140 10044
rect 177908 10004 177914 10016
rect 309134 10004 309140 10016
rect 309192 10004 309198 10056
rect 176378 9936 176384 9988
rect 176436 9976 176442 9988
rect 304994 9976 305000 9988
rect 176436 9948 305000 9976
rect 176436 9936 176442 9948
rect 304994 9936 305000 9948
rect 305052 9936 305058 9988
rect 174998 9868 175004 9920
rect 175056 9908 175062 9920
rect 302234 9908 302240 9920
rect 175056 9880 302240 9908
rect 175056 9868 175062 9880
rect 302234 9868 302240 9880
rect 302292 9868 302298 9920
rect 173710 9800 173716 9852
rect 173768 9840 173774 9852
rect 298094 9840 298100 9852
rect 173768 9812 298100 9840
rect 173768 9800 173774 9812
rect 298094 9800 298100 9812
rect 298152 9800 298158 9852
rect 162118 9772 162124 9784
rect 161952 9744 162124 9772
rect 161952 9716 161980 9744
rect 162118 9732 162124 9744
rect 162176 9732 162182 9784
rect 172330 9732 172336 9784
rect 172388 9772 172394 9784
rect 295334 9772 295340 9784
rect 172388 9744 295340 9772
rect 172388 9732 172394 9744
rect 295334 9732 295340 9744
rect 295392 9732 295398 9784
rect 161934 9664 161940 9716
rect 161992 9664 161998 9716
rect 172238 9664 172244 9716
rect 172296 9704 172302 9716
rect 291194 9704 291200 9716
rect 172296 9676 291200 9704
rect 172296 9664 172302 9676
rect 291194 9664 291200 9676
rect 291252 9664 291258 9716
rect 90910 9596 90916 9648
rect 90968 9596 90974 9648
rect 94222 9636 94228 9648
rect 94183 9608 94228 9636
rect 94222 9596 94228 9608
rect 94280 9596 94286 9648
rect 154390 9596 154396 9648
rect 154448 9636 154454 9648
rect 238849 9639 238907 9645
rect 238849 9636 238861 9639
rect 154448 9608 238861 9636
rect 154448 9596 154454 9608
rect 238849 9605 238861 9608
rect 238895 9605 238907 9639
rect 238849 9599 238907 9605
rect 239401 9639 239459 9645
rect 239401 9605 239413 9639
rect 239447 9636 239459 9639
rect 250346 9636 250352 9648
rect 239447 9608 250352 9636
rect 239447 9605 239459 9608
rect 239401 9599 239459 9605
rect 250346 9596 250352 9608
rect 250404 9596 250410 9648
rect 250898 9596 250904 9648
rect 250956 9636 250962 9648
rect 520366 9636 520372 9648
rect 250956 9608 520372 9636
rect 250956 9596 250962 9608
rect 520366 9596 520372 9608
rect 520424 9596 520430 9648
rect 90928 9512 90956 9596
rect 155770 9528 155776 9580
rect 155828 9568 155834 9580
rect 239309 9571 239367 9577
rect 239309 9568 239321 9571
rect 155828 9540 239321 9568
rect 155828 9528 155834 9540
rect 239309 9537 239321 9540
rect 239355 9537 239367 9571
rect 246758 9568 246764 9580
rect 239309 9531 239367 9537
rect 239416 9540 246764 9568
rect 90910 9460 90916 9512
rect 90968 9460 90974 9512
rect 155678 9460 155684 9512
rect 155736 9500 155742 9512
rect 239416 9500 239444 9540
rect 246758 9528 246764 9540
rect 246816 9528 246822 9580
rect 246868 9540 249748 9568
rect 155736 9472 239444 9500
rect 239493 9503 239551 9509
rect 155736 9460 155742 9472
rect 239493 9469 239505 9503
rect 239539 9500 239551 9503
rect 244829 9503 244887 9509
rect 244829 9500 244841 9503
rect 239539 9472 244841 9500
rect 239539 9469 239551 9472
rect 239493 9463 239551 9469
rect 244829 9469 244841 9472
rect 244875 9469 244887 9503
rect 245562 9500 245568 9512
rect 244829 9463 244887 9469
rect 244936 9472 245568 9500
rect 157058 9392 157064 9444
rect 157116 9432 157122 9444
rect 239217 9435 239275 9441
rect 239217 9432 239229 9435
rect 157116 9404 239229 9432
rect 157116 9392 157122 9404
rect 239217 9401 239229 9404
rect 239263 9401 239275 9435
rect 239217 9395 239275 9401
rect 239309 9435 239367 9441
rect 239309 9401 239321 9435
rect 239355 9432 239367 9435
rect 244936 9432 244964 9472
rect 245562 9460 245568 9472
rect 245620 9460 245626 9512
rect 246669 9503 246727 9509
rect 246669 9469 246681 9503
rect 246715 9500 246727 9503
rect 246868 9500 246896 9540
rect 246715 9472 246896 9500
rect 246715 9469 246727 9472
rect 246669 9463 246727 9469
rect 239355 9404 244964 9432
rect 239355 9401 239367 9404
rect 239309 9395 239367 9401
rect 245470 9392 245476 9444
rect 245528 9432 245534 9444
rect 249429 9435 249487 9441
rect 249429 9432 249441 9435
rect 245528 9404 249441 9432
rect 245528 9392 245534 9404
rect 249429 9401 249441 9404
rect 249475 9401 249487 9435
rect 249720 9432 249748 9540
rect 252186 9528 252192 9580
rect 252244 9568 252250 9580
rect 523862 9568 523868 9580
rect 252244 9540 523868 9568
rect 252244 9528 252250 9540
rect 523862 9528 523868 9540
rect 523920 9528 523926 9580
rect 253750 9460 253756 9512
rect 253808 9500 253814 9512
rect 527450 9500 527456 9512
rect 253808 9472 527456 9500
rect 253808 9460 253814 9472
rect 527450 9460 527456 9472
rect 527508 9460 527514 9512
rect 253842 9432 253848 9444
rect 249720 9404 253848 9432
rect 249429 9395 249487 9401
rect 253842 9392 253848 9404
rect 253900 9392 253906 9444
rect 256418 9392 256424 9444
rect 256476 9432 256482 9444
rect 258997 9435 259055 9441
rect 256476 9404 258948 9432
rect 256476 9392 256482 9404
rect 156966 9324 156972 9376
rect 157024 9364 157030 9376
rect 239401 9367 239459 9373
rect 239401 9364 239413 9367
rect 157024 9336 239413 9364
rect 157024 9324 157030 9336
rect 239401 9333 239413 9336
rect 239447 9333 239459 9367
rect 239401 9327 239459 9333
rect 243998 9324 244004 9376
rect 244056 9364 244062 9376
rect 249153 9367 249211 9373
rect 249153 9364 249165 9367
rect 244056 9336 249165 9364
rect 244056 9324 244062 9336
rect 249153 9333 249165 9336
rect 249199 9333 249211 9367
rect 249153 9327 249211 9333
rect 249245 9367 249303 9373
rect 249245 9333 249257 9367
rect 249291 9364 249303 9367
rect 249291 9336 249472 9364
rect 249291 9333 249303 9336
rect 249245 9327 249303 9333
rect 158530 9256 158536 9308
rect 158588 9296 158594 9308
rect 246669 9299 246727 9305
rect 246669 9296 246681 9299
rect 158588 9268 246681 9296
rect 158588 9256 158594 9268
rect 246669 9265 246681 9268
rect 246715 9265 246727 9299
rect 246669 9259 246727 9265
rect 246850 9256 246856 9308
rect 246908 9296 246914 9308
rect 249337 9299 249395 9305
rect 249337 9296 249349 9299
rect 246908 9268 249349 9296
rect 246908 9256 246914 9268
rect 249337 9265 249349 9268
rect 249383 9265 249395 9299
rect 249444 9296 249472 9336
rect 249518 9324 249524 9376
rect 249576 9364 249582 9376
rect 258721 9367 258779 9373
rect 258721 9364 258733 9367
rect 249576 9336 258733 9364
rect 249576 9324 249582 9336
rect 258721 9333 258733 9336
rect 258767 9333 258779 9367
rect 258920 9364 258948 9404
rect 258997 9401 259009 9435
rect 259043 9432 259055 9435
rect 531038 9432 531044 9444
rect 259043 9404 531044 9432
rect 259043 9401 259055 9404
rect 258997 9395 259055 9401
rect 531038 9392 531044 9404
rect 531096 9392 531102 9444
rect 534534 9364 534540 9376
rect 258920 9336 534540 9364
rect 258721 9327 258779 9333
rect 534534 9324 534540 9336
rect 534592 9324 534598 9376
rect 252646 9296 252652 9308
rect 249444 9268 252652 9296
rect 249337 9259 249395 9265
rect 252646 9256 252652 9268
rect 252704 9256 252710 9308
rect 254949 9299 255007 9305
rect 254949 9265 254961 9299
rect 254995 9296 255007 9299
rect 254995 9268 256372 9296
rect 254995 9265 255007 9268
rect 254949 9259 255007 9265
rect 158438 9188 158444 9240
rect 158496 9228 158502 9240
rect 248969 9231 249027 9237
rect 248969 9228 248981 9231
rect 158496 9200 248981 9228
rect 158496 9188 158502 9200
rect 248969 9197 248981 9200
rect 249015 9197 249027 9231
rect 256234 9228 256240 9240
rect 248969 9191 249027 9197
rect 249076 9200 256240 9228
rect 159910 9120 159916 9172
rect 159968 9160 159974 9172
rect 249076 9160 249104 9200
rect 256234 9188 256240 9200
rect 256292 9188 256298 9240
rect 256344 9228 256372 9268
rect 256510 9256 256516 9308
rect 256568 9296 256574 9308
rect 538122 9296 538128 9308
rect 256568 9268 538128 9296
rect 256568 9256 256574 9268
rect 538122 9256 538128 9268
rect 538180 9256 538186 9308
rect 257798 9228 257804 9240
rect 256344 9200 257804 9228
rect 257798 9188 257804 9200
rect 257856 9188 257862 9240
rect 257890 9188 257896 9240
rect 257948 9228 257954 9240
rect 541710 9228 541716 9240
rect 257948 9200 541716 9228
rect 257948 9188 257954 9200
rect 541710 9188 541716 9200
rect 541768 9188 541774 9240
rect 255041 9163 255099 9169
rect 255041 9160 255053 9163
rect 159968 9132 249104 9160
rect 249168 9132 255053 9160
rect 159968 9120 159974 9132
rect 159818 9052 159824 9104
rect 159876 9092 159882 9104
rect 249168 9092 249196 9132
rect 255041 9129 255053 9132
rect 255087 9129 255099 9163
rect 255041 9123 255099 9129
rect 255130 9120 255136 9172
rect 255188 9160 255194 9172
rect 258997 9163 259055 9169
rect 258997 9160 259009 9163
rect 255188 9132 259009 9160
rect 255188 9120 255194 9132
rect 258997 9129 259009 9132
rect 259043 9129 259055 9163
rect 258997 9123 259055 9129
rect 259089 9163 259147 9169
rect 259089 9129 259101 9163
rect 259135 9160 259147 9163
rect 259822 9160 259828 9172
rect 259135 9132 259828 9160
rect 259135 9129 259147 9132
rect 259089 9123 259147 9129
rect 259822 9120 259828 9132
rect 259880 9120 259886 9172
rect 260650 9120 260656 9172
rect 260708 9160 260714 9172
rect 548886 9160 548892 9172
rect 260708 9132 548892 9160
rect 260708 9120 260714 9132
rect 548886 9120 548892 9132
rect 548944 9120 548950 9172
rect 159876 9064 249196 9092
rect 249245 9095 249303 9101
rect 159876 9052 159882 9064
rect 249245 9061 249257 9095
rect 249291 9092 249303 9095
rect 267366 9092 267372 9104
rect 249291 9064 267372 9092
rect 249291 9061 249303 9064
rect 249245 9055 249303 9061
rect 267366 9052 267372 9064
rect 267424 9052 267430 9104
rect 267458 9052 267464 9104
rect 267516 9092 267522 9104
rect 566734 9092 566740 9104
rect 267516 9064 566740 9092
rect 267516 9052 267522 9064
rect 566734 9052 566740 9064
rect 566792 9052 566798 9104
rect 162670 8984 162676 9036
rect 162728 9024 162734 9036
rect 266998 9024 267004 9036
rect 162728 8996 267004 9024
rect 162728 8984 162734 8996
rect 266998 8984 267004 8996
rect 267056 8984 267062 9036
rect 267550 8984 267556 9036
rect 267608 9024 267614 9036
rect 570230 9024 570236 9036
rect 267608 8996 570236 9024
rect 267608 8984 267614 8996
rect 570230 8984 570236 8996
rect 570288 8984 570294 9036
rect 153010 8916 153016 8968
rect 153068 8956 153074 8968
rect 161293 8959 161351 8965
rect 161293 8956 161305 8959
rect 153068 8928 161305 8956
rect 153068 8916 153074 8928
rect 161293 8925 161305 8928
rect 161339 8925 161351 8959
rect 161293 8919 161351 8925
rect 164050 8916 164056 8968
rect 164108 8956 164114 8968
rect 270494 8956 270500 8968
rect 164108 8928 270500 8956
rect 164108 8916 164114 8928
rect 270494 8916 270500 8928
rect 270552 8916 270558 8968
rect 271690 8916 271696 8968
rect 271748 8956 271754 8968
rect 581086 8956 581092 8968
rect 271748 8928 581092 8956
rect 271748 8916 271754 8928
rect 581086 8916 581092 8928
rect 581144 8916 581150 8968
rect 154298 8848 154304 8900
rect 154356 8888 154362 8900
rect 239217 8891 239275 8897
rect 154356 8860 238616 8888
rect 154356 8848 154362 8860
rect 161293 8823 161351 8829
rect 161293 8789 161305 8823
rect 161339 8820 161351 8823
rect 166997 8823 167055 8829
rect 166997 8820 167009 8823
rect 161339 8792 167009 8820
rect 161339 8789 161351 8792
rect 161293 8783 161351 8789
rect 166997 8789 167009 8792
rect 167043 8789 167055 8823
rect 166997 8783 167055 8789
rect 176565 8823 176623 8829
rect 176565 8789 176577 8823
rect 176611 8820 176623 8823
rect 186317 8823 186375 8829
rect 186317 8820 186329 8823
rect 176611 8792 186329 8820
rect 176611 8789 176623 8792
rect 176565 8783 176623 8789
rect 186317 8789 186329 8792
rect 186363 8789 186375 8823
rect 186317 8783 186375 8789
rect 195885 8823 195943 8829
rect 195885 8789 195897 8823
rect 195931 8820 195943 8823
rect 205634 8820 205640 8832
rect 195931 8792 205640 8820
rect 195931 8789 195943 8792
rect 195885 8783 195943 8789
rect 205634 8780 205640 8792
rect 205692 8780 205698 8832
rect 215110 8780 215116 8832
rect 215168 8820 215174 8832
rect 224954 8820 224960 8832
rect 215168 8792 224960 8820
rect 215168 8780 215174 8792
rect 224954 8780 224960 8792
rect 225012 8780 225018 8832
rect 152918 8712 152924 8764
rect 152976 8752 152982 8764
rect 238386 8752 238392 8764
rect 152976 8724 238392 8752
rect 152976 8712 152982 8724
rect 238386 8712 238392 8724
rect 238444 8712 238450 8764
rect 238588 8752 238616 8860
rect 239217 8857 239229 8891
rect 239263 8888 239275 8891
rect 248782 8888 248788 8900
rect 239263 8860 248788 8888
rect 239263 8857 239275 8860
rect 239217 8851 239275 8857
rect 248782 8848 248788 8860
rect 248840 8848 248846 8900
rect 248969 8891 249027 8897
rect 248969 8857 248981 8891
rect 249015 8888 249027 8891
rect 254949 8891 255007 8897
rect 254949 8888 254961 8891
rect 249015 8860 254961 8888
rect 249015 8857 249027 8860
rect 248969 8851 249027 8857
rect 254949 8857 254961 8860
rect 254995 8857 255007 8891
rect 254949 8851 255007 8857
rect 255041 8891 255099 8897
rect 255041 8857 255053 8891
rect 255087 8888 255099 8891
rect 258629 8891 258687 8897
rect 258629 8888 258641 8891
rect 255087 8860 258641 8888
rect 255087 8857 255099 8860
rect 255041 8851 255099 8857
rect 258629 8857 258641 8860
rect 258675 8857 258687 8891
rect 258629 8851 258687 8857
rect 258721 8891 258779 8897
rect 258721 8857 258733 8891
rect 258767 8888 258779 8891
rect 516778 8888 516784 8900
rect 258767 8860 516784 8888
rect 258767 8857 258779 8860
rect 258721 8851 258779 8857
rect 516778 8848 516784 8860
rect 516836 8848 516842 8900
rect 242710 8780 242716 8832
rect 242768 8820 242774 8832
rect 249061 8823 249119 8829
rect 249061 8820 249073 8823
rect 242768 8792 249073 8820
rect 242768 8780 242774 8792
rect 249061 8789 249073 8792
rect 249107 8789 249119 8823
rect 513190 8820 513196 8832
rect 249061 8783 249119 8789
rect 249168 8792 513196 8820
rect 241974 8752 241980 8764
rect 238588 8724 241980 8752
rect 241974 8712 241980 8724
rect 242032 8712 242038 8764
rect 244829 8755 244887 8761
rect 244829 8721 244841 8755
rect 244875 8752 244887 8755
rect 248138 8752 248144 8764
rect 244875 8724 248144 8752
rect 244875 8721 244887 8724
rect 244829 8715 244887 8721
rect 248138 8712 248144 8724
rect 248196 8712 248202 8764
rect 248414 8712 248420 8764
rect 248472 8752 248478 8764
rect 249168 8752 249196 8792
rect 513190 8780 513196 8792
rect 513248 8780 513254 8832
rect 248472 8724 249196 8752
rect 249337 8755 249395 8761
rect 248472 8712 248478 8724
rect 249337 8721 249349 8755
rect 249383 8752 249395 8755
rect 509602 8752 509608 8764
rect 249383 8724 509608 8752
rect 249383 8721 249395 8724
rect 249337 8715 249395 8721
rect 509602 8712 509608 8724
rect 509660 8712 509666 8764
rect 152826 8644 152832 8696
rect 152884 8684 152890 8696
rect 235994 8684 236000 8696
rect 152884 8656 236000 8684
rect 152884 8644 152890 8656
rect 235994 8644 236000 8656
rect 236052 8644 236058 8696
rect 238849 8687 238907 8693
rect 238849 8653 238861 8687
rect 238895 8684 238907 8687
rect 243170 8684 243176 8696
rect 238895 8656 243176 8684
rect 238895 8653 238907 8656
rect 238849 8647 238907 8653
rect 243170 8644 243176 8656
rect 243228 8644 243234 8696
rect 249245 8687 249303 8693
rect 249245 8684 249257 8687
rect 246316 8656 249257 8684
rect 166997 8619 167055 8625
rect 166997 8585 167009 8619
rect 167043 8616 167055 8619
rect 176565 8619 176623 8625
rect 176565 8616 176577 8619
rect 167043 8588 176577 8616
rect 167043 8585 167055 8588
rect 166997 8579 167055 8585
rect 176565 8585 176577 8588
rect 176611 8585 176623 8619
rect 193217 8619 193275 8625
rect 193217 8616 193229 8619
rect 176565 8579 176623 8585
rect 181456 8588 193229 8616
rect 176470 8440 176476 8492
rect 176528 8480 176534 8492
rect 181456 8480 181484 8588
rect 193217 8585 193229 8588
rect 193263 8585 193275 8619
rect 193217 8579 193275 8585
rect 197170 8576 197176 8628
rect 197228 8616 197234 8628
rect 246316 8616 246344 8656
rect 249245 8653 249257 8656
rect 249291 8653 249303 8687
rect 249245 8647 249303 8653
rect 249429 8687 249487 8693
rect 249429 8653 249441 8687
rect 249475 8684 249487 8687
rect 506014 8684 506020 8696
rect 249475 8656 506020 8684
rect 249475 8653 249487 8656
rect 249429 8647 249487 8653
rect 506014 8644 506020 8656
rect 506072 8644 506078 8696
rect 197228 8588 246344 8616
rect 197228 8576 197234 8588
rect 249334 8576 249340 8628
rect 249392 8616 249398 8628
rect 502426 8616 502432 8628
rect 249392 8588 502432 8616
rect 249392 8576 249398 8588
rect 502426 8576 502432 8588
rect 502484 8576 502490 8628
rect 181990 8508 181996 8560
rect 182048 8548 182054 8560
rect 239493 8551 239551 8557
rect 239493 8548 239505 8551
rect 182048 8520 239505 8548
rect 182048 8508 182054 8520
rect 239493 8517 239505 8520
rect 239539 8517 239551 8551
rect 242894 8548 242900 8560
rect 239493 8511 239551 8517
rect 239692 8520 242900 8548
rect 195793 8483 195851 8489
rect 195793 8480 195805 8483
rect 176528 8452 181484 8480
rect 190380 8452 195805 8480
rect 176528 8440 176534 8452
rect 186317 8415 186375 8421
rect 186317 8381 186329 8415
rect 186363 8412 186375 8415
rect 190380 8412 190408 8452
rect 195793 8449 195805 8452
rect 195839 8449 195851 8483
rect 195793 8443 195851 8449
rect 196069 8483 196127 8489
rect 196069 8449 196081 8483
rect 196115 8480 196127 8483
rect 215113 8483 215171 8489
rect 215113 8480 215125 8483
rect 196115 8452 215125 8480
rect 196115 8449 196127 8452
rect 196069 8443 196127 8449
rect 215113 8449 215125 8452
rect 215159 8449 215171 8483
rect 215113 8443 215171 8449
rect 215389 8483 215447 8489
rect 215389 8449 215401 8483
rect 215435 8480 215447 8483
rect 215435 8452 234568 8480
rect 215435 8449 215447 8452
rect 215389 8443 215447 8449
rect 186363 8384 190408 8412
rect 186363 8381 186375 8384
rect 186317 8375 186375 8381
rect 191650 8372 191656 8424
rect 191708 8412 191714 8424
rect 197173 8415 197231 8421
rect 197173 8412 197185 8415
rect 191708 8384 197185 8412
rect 191708 8372 191714 8384
rect 197173 8381 197185 8384
rect 197219 8381 197231 8415
rect 197173 8375 197231 8381
rect 202877 8415 202935 8421
rect 202877 8381 202889 8415
rect 202923 8412 202935 8415
rect 205545 8415 205603 8421
rect 205545 8412 205557 8415
rect 202923 8384 205557 8412
rect 202923 8381 202935 8384
rect 202877 8375 202935 8381
rect 205545 8381 205557 8384
rect 205591 8381 205603 8415
rect 205545 8375 205603 8381
rect 205637 8415 205695 8421
rect 205637 8381 205649 8415
rect 205683 8412 205695 8415
rect 215205 8415 215263 8421
rect 215205 8412 215217 8415
rect 205683 8384 215217 8412
rect 205683 8381 205695 8384
rect 205637 8375 205695 8381
rect 215205 8381 215217 8384
rect 215251 8381 215263 8415
rect 215205 8375 215263 8381
rect 215297 8415 215355 8421
rect 215297 8381 215309 8415
rect 215343 8412 215355 8415
rect 234430 8412 234436 8424
rect 215343 8384 234436 8412
rect 215343 8381 215355 8384
rect 215297 8375 215355 8381
rect 234430 8372 234436 8384
rect 234488 8372 234494 8424
rect 234540 8412 234568 8452
rect 239692 8412 239720 8520
rect 242894 8508 242900 8520
rect 242952 8508 242958 8560
rect 249153 8551 249211 8557
rect 249153 8517 249165 8551
rect 249199 8548 249211 8551
rect 498930 8548 498936 8560
rect 249199 8520 498936 8548
rect 249199 8517 249211 8520
rect 249153 8511 249211 8517
rect 498930 8508 498936 8520
rect 498988 8508 498994 8560
rect 239766 8440 239772 8492
rect 239824 8480 239830 8492
rect 248969 8483 249027 8489
rect 248969 8480 248981 8483
rect 239824 8452 248981 8480
rect 239824 8440 239830 8452
rect 248969 8449 248981 8452
rect 249015 8449 249027 8483
rect 248969 8443 249027 8449
rect 249061 8483 249119 8489
rect 249061 8449 249073 8483
rect 249107 8480 249119 8483
rect 495342 8480 495348 8492
rect 249107 8452 495348 8480
rect 249107 8449 249119 8452
rect 249061 8443 249119 8449
rect 495342 8440 495348 8452
rect 495400 8440 495406 8492
rect 234540 8384 239720 8412
rect 241330 8372 241336 8424
rect 241388 8412 241394 8424
rect 491754 8412 491760 8424
rect 241388 8384 491760 8412
rect 241388 8372 241394 8384
rect 491754 8372 491760 8384
rect 491812 8372 491818 8424
rect 73338 8344 73344 8356
rect 73299 8316 73344 8344
rect 73338 8304 73344 8316
rect 73396 8304 73402 8356
rect 165522 8304 165528 8356
rect 165580 8344 165586 8356
rect 205453 8347 205511 8353
rect 205453 8344 205465 8347
rect 165580 8316 205465 8344
rect 165580 8304 165586 8316
rect 205453 8313 205465 8316
rect 205499 8313 205511 8347
rect 205453 8307 205511 8313
rect 205729 8347 205787 8353
rect 205729 8313 205741 8347
rect 205775 8344 205787 8347
rect 274082 8344 274088 8356
rect 205775 8316 274088 8344
rect 205775 8313 205787 8316
rect 205729 8307 205787 8313
rect 274082 8304 274088 8316
rect 274140 8304 274146 8356
rect 193217 8279 193275 8285
rect 193217 8245 193229 8279
rect 193263 8276 193275 8279
rect 196069 8279 196127 8285
rect 196069 8276 196081 8279
rect 193263 8248 196081 8276
rect 193263 8245 193275 8248
rect 193217 8239 193275 8245
rect 196069 8245 196081 8248
rect 196115 8245 196127 8279
rect 196069 8239 196127 8245
rect 216490 8236 216496 8288
rect 216548 8276 216554 8288
rect 419166 8276 419172 8288
rect 216548 8248 419172 8276
rect 216548 8236 216554 8248
rect 419166 8236 419172 8248
rect 419224 8236 419230 8288
rect 197173 8211 197231 8217
rect 197173 8177 197185 8211
rect 197219 8208 197231 8211
rect 202877 8211 202935 8217
rect 202877 8208 202889 8211
rect 197219 8180 202889 8208
rect 197219 8177 197231 8180
rect 197173 8171 197231 8177
rect 202877 8177 202889 8180
rect 202923 8177 202935 8211
rect 202877 8171 202935 8177
rect 216582 8168 216588 8220
rect 216640 8208 216646 8220
rect 422754 8208 422760 8220
rect 216640 8180 422760 8208
rect 216640 8168 216646 8180
rect 422754 8168 422760 8180
rect 422812 8168 422818 8220
rect 217962 8100 217968 8152
rect 218020 8140 218026 8152
rect 426342 8140 426348 8152
rect 218020 8112 426348 8140
rect 218020 8100 218026 8112
rect 426342 8100 426348 8112
rect 426400 8100 426406 8152
rect 215205 8075 215263 8081
rect 215205 8041 215217 8075
rect 215251 8072 215263 8075
rect 215297 8075 215355 8081
rect 215297 8072 215309 8075
rect 215251 8044 215309 8072
rect 215251 8041 215263 8044
rect 215205 8035 215263 8041
rect 215297 8041 215309 8044
rect 215343 8041 215355 8075
rect 215297 8035 215355 8041
rect 219250 8032 219256 8084
rect 219308 8072 219314 8084
rect 429930 8072 429936 8084
rect 219308 8044 429936 8072
rect 219308 8032 219314 8044
rect 429930 8032 429936 8044
rect 429988 8032 429994 8084
rect 140498 7964 140504 8016
rect 140556 8004 140562 8016
rect 202690 8004 202696 8016
rect 140556 7976 202696 8004
rect 140556 7964 140562 7976
rect 202690 7964 202696 7976
rect 202748 7964 202754 8016
rect 215113 8007 215171 8013
rect 215113 7973 215125 8007
rect 215159 8004 215171 8007
rect 215389 8007 215447 8013
rect 215389 8004 215401 8007
rect 215159 7976 215401 8004
rect 215159 7973 215171 7976
rect 215113 7967 215171 7973
rect 215389 7973 215401 7976
rect 215435 7973 215447 8007
rect 215389 7967 215447 7973
rect 220722 7964 220728 8016
rect 220780 8004 220786 8016
rect 433518 8004 433524 8016
rect 220780 7976 433524 8004
rect 220780 7964 220786 7976
rect 433518 7964 433524 7976
rect 433576 7964 433582 8016
rect 141970 7896 141976 7948
rect 142028 7936 142034 7948
rect 206278 7936 206284 7948
rect 142028 7908 206284 7936
rect 142028 7896 142034 7908
rect 206278 7896 206284 7908
rect 206336 7896 206342 7948
rect 218698 7896 218704 7948
rect 218756 7936 218762 7948
rect 219250 7936 219256 7948
rect 218756 7908 219256 7936
rect 218756 7896 218762 7908
rect 219250 7896 219256 7908
rect 219308 7896 219314 7948
rect 222010 7896 222016 7948
rect 222068 7936 222074 7948
rect 437014 7936 437020 7948
rect 222068 7908 437020 7936
rect 222068 7896 222074 7908
rect 437014 7896 437020 7908
rect 437072 7896 437078 7948
rect 143350 7828 143356 7880
rect 143408 7868 143414 7880
rect 209866 7868 209872 7880
rect 143408 7840 209872 7868
rect 143408 7828 143414 7840
rect 209866 7828 209872 7840
rect 209924 7828 209930 7880
rect 223482 7828 223488 7880
rect 223540 7868 223546 7880
rect 440602 7868 440608 7880
rect 223540 7840 440608 7868
rect 223540 7828 223546 7840
rect 440602 7828 440608 7840
rect 440660 7828 440666 7880
rect 144546 7760 144552 7812
rect 144604 7800 144610 7812
rect 213454 7800 213460 7812
rect 144604 7772 213460 7800
rect 144604 7760 144610 7772
rect 213454 7760 213460 7772
rect 213512 7760 213518 7812
rect 224770 7760 224776 7812
rect 224828 7800 224834 7812
rect 444190 7800 444196 7812
rect 224828 7772 444196 7800
rect 224828 7760 224834 7772
rect 444190 7760 444196 7772
rect 444248 7760 444254 7812
rect 146110 7692 146116 7744
rect 146168 7732 146174 7744
rect 217042 7732 217048 7744
rect 146168 7704 217048 7732
rect 146168 7692 146174 7704
rect 217042 7692 217048 7704
rect 217100 7692 217106 7744
rect 226150 7692 226156 7744
rect 226208 7732 226214 7744
rect 447778 7732 447784 7744
rect 226208 7704 447784 7732
rect 226208 7692 226214 7704
rect 447778 7692 447784 7704
rect 447836 7692 447842 7744
rect 147490 7624 147496 7676
rect 147548 7664 147554 7676
rect 220538 7664 220544 7676
rect 147548 7636 220544 7664
rect 147548 7624 147554 7636
rect 220538 7624 220544 7636
rect 220596 7624 220602 7676
rect 227622 7624 227628 7676
rect 227680 7664 227686 7676
rect 451366 7664 451372 7676
rect 227680 7636 451372 7664
rect 227680 7624 227686 7636
rect 451366 7624 451372 7636
rect 451424 7624 451430 7676
rect 148778 7556 148784 7608
rect 148836 7596 148842 7608
rect 224126 7596 224132 7608
rect 148836 7568 224132 7596
rect 148836 7556 148842 7568
rect 224126 7556 224132 7568
rect 224184 7556 224190 7608
rect 227530 7556 227536 7608
rect 227588 7596 227594 7608
rect 454862 7596 454868 7608
rect 227588 7568 454868 7596
rect 227588 7556 227594 7568
rect 454862 7556 454868 7568
rect 454920 7556 454926 7608
rect 215202 7488 215208 7540
rect 215260 7528 215266 7540
rect 415670 7528 415676 7540
rect 215260 7500 415676 7528
rect 215260 7488 215266 7500
rect 415670 7488 415676 7500
rect 415728 7488 415734 7540
rect 156598 7420 156604 7472
rect 156656 7460 156662 7472
rect 161201 7463 161259 7469
rect 161201 7460 161213 7463
rect 156656 7432 161213 7460
rect 156656 7420 156662 7432
rect 161201 7429 161213 7432
rect 161247 7429 161259 7463
rect 161201 7423 161259 7429
rect 213730 7420 213736 7472
rect 213788 7460 213794 7472
rect 412082 7460 412088 7472
rect 213788 7432 412088 7460
rect 213788 7420 213794 7432
rect 412082 7420 412088 7432
rect 412140 7420 412146 7472
rect 212442 7352 212448 7404
rect 212500 7392 212506 7404
rect 408586 7392 408592 7404
rect 212500 7364 408592 7392
rect 212500 7352 212506 7364
rect 408586 7352 408592 7364
rect 408644 7352 408650 7404
rect 211062 7284 211068 7336
rect 211120 7324 211126 7336
rect 404906 7324 404912 7336
rect 211120 7296 404912 7324
rect 211120 7284 211126 7296
rect 404906 7284 404912 7296
rect 404964 7284 404970 7336
rect 209682 7216 209688 7268
rect 209740 7256 209746 7268
rect 401318 7256 401324 7268
rect 209740 7228 401324 7256
rect 209740 7216 209746 7228
rect 401318 7216 401324 7228
rect 401376 7216 401382 7268
rect 208210 7148 208216 7200
rect 208268 7188 208274 7200
rect 397822 7188 397828 7200
rect 208268 7160 397828 7188
rect 208268 7148 208274 7160
rect 397822 7148 397828 7160
rect 397880 7148 397886 7200
rect 206922 7080 206928 7132
rect 206980 7120 206986 7132
rect 394234 7120 394240 7132
rect 206980 7092 394240 7120
rect 206980 7080 206986 7092
rect 394234 7080 394240 7092
rect 394292 7080 394298 7132
rect 197998 7012 198004 7064
rect 198056 7052 198062 7064
rect 201589 7055 201647 7061
rect 201589 7052 201601 7055
rect 198056 7024 201601 7052
rect 198056 7012 198062 7024
rect 201589 7021 201601 7024
rect 201635 7021 201647 7055
rect 201589 7015 201647 7021
rect 204806 7012 204812 7064
rect 204864 7052 204870 7064
rect 205177 7055 205235 7061
rect 205177 7052 205189 7055
rect 204864 7024 205189 7052
rect 204864 7012 204870 7024
rect 205177 7021 205189 7024
rect 205223 7021 205235 7055
rect 205177 7015 205235 7021
rect 205542 7012 205548 7064
rect 205600 7052 205606 7064
rect 390646 7052 390652 7064
rect 205600 7024 390652 7052
rect 205600 7012 205606 7024
rect 390646 7012 390652 7024
rect 390704 7012 390710 7064
rect 161290 6944 161296 6996
rect 161348 6984 161354 6996
rect 263410 6984 263416 6996
rect 161348 6956 263416 6984
rect 161348 6944 161354 6956
rect 263410 6944 263416 6956
rect 263468 6944 263474 6996
rect 241422 6916 241428 6928
rect 241383 6888 241428 6916
rect 241422 6876 241428 6888
rect 241480 6876 241486 6928
rect 248322 6876 248328 6928
rect 248380 6916 248386 6928
rect 249613 6919 249671 6925
rect 249613 6916 249625 6919
rect 248380 6888 249625 6916
rect 248380 6876 248386 6888
rect 249613 6885 249625 6888
rect 249659 6885 249671 6919
rect 249613 6879 249671 6885
rect 180610 6808 180616 6860
rect 180668 6848 180674 6860
rect 319254 6848 319260 6860
rect 180668 6820 319260 6848
rect 180668 6808 180674 6820
rect 319254 6808 319260 6820
rect 319312 6808 319318 6860
rect 182082 6740 182088 6792
rect 182140 6780 182146 6792
rect 322842 6780 322848 6792
rect 182140 6752 322848 6780
rect 182140 6740 182146 6752
rect 322842 6740 322848 6752
rect 322900 6740 322906 6792
rect 183462 6672 183468 6724
rect 183520 6712 183526 6724
rect 326430 6712 326436 6724
rect 183520 6684 326436 6712
rect 183520 6672 183526 6684
rect 326430 6672 326436 6684
rect 326488 6672 326494 6724
rect 161934 6604 161940 6656
rect 161992 6644 161998 6656
rect 162121 6647 162179 6653
rect 162121 6644 162133 6647
rect 161992 6616 162133 6644
rect 161992 6604 161998 6616
rect 162121 6613 162133 6616
rect 162167 6613 162179 6647
rect 162121 6607 162179 6613
rect 184750 6604 184756 6656
rect 184808 6644 184814 6656
rect 330018 6644 330024 6656
rect 184808 6616 330024 6644
rect 184808 6604 184814 6616
rect 330018 6604 330024 6616
rect 330076 6604 330082 6656
rect 129458 6536 129464 6588
rect 129516 6576 129522 6588
rect 170582 6576 170588 6588
rect 129516 6548 170588 6576
rect 129516 6536 129522 6548
rect 170582 6536 170588 6548
rect 170640 6536 170646 6588
rect 186222 6536 186228 6588
rect 186280 6576 186286 6588
rect 333606 6576 333612 6588
rect 186280 6548 333612 6576
rect 186280 6536 186286 6548
rect 333606 6536 333612 6548
rect 333664 6536 333670 6588
rect 130838 6468 130844 6520
rect 130896 6508 130902 6520
rect 174170 6508 174176 6520
rect 130896 6480 174176 6508
rect 130896 6468 130902 6480
rect 174170 6468 174176 6480
rect 174228 6468 174234 6520
rect 187510 6468 187516 6520
rect 187568 6508 187574 6520
rect 337102 6508 337108 6520
rect 187568 6480 337108 6508
rect 187568 6468 187574 6480
rect 337102 6468 337108 6480
rect 337160 6468 337166 6520
rect 132218 6400 132224 6452
rect 132276 6440 132282 6452
rect 177758 6440 177764 6452
rect 132276 6412 177764 6440
rect 132276 6400 132282 6412
rect 177758 6400 177764 6412
rect 177816 6400 177822 6452
rect 188890 6400 188896 6452
rect 188948 6440 188954 6452
rect 340690 6440 340696 6452
rect 188948 6412 340696 6440
rect 188948 6400 188954 6412
rect 340690 6400 340696 6412
rect 340748 6400 340754 6452
rect 133782 6332 133788 6384
rect 133840 6372 133846 6384
rect 181346 6372 181352 6384
rect 133840 6344 181352 6372
rect 133840 6332 133846 6344
rect 181346 6332 181352 6344
rect 181404 6332 181410 6384
rect 190362 6332 190368 6384
rect 190420 6372 190426 6384
rect 344278 6372 344284 6384
rect 190420 6344 344284 6372
rect 190420 6332 190426 6344
rect 344278 6332 344284 6344
rect 344336 6332 344342 6384
rect 135162 6264 135168 6316
rect 135220 6304 135226 6316
rect 184842 6304 184848 6316
rect 135220 6276 184848 6304
rect 135220 6264 135226 6276
rect 184842 6264 184848 6276
rect 184900 6264 184906 6316
rect 191742 6264 191748 6316
rect 191800 6304 191806 6316
rect 347866 6304 347872 6316
rect 191800 6276 347872 6304
rect 191800 6264 191806 6276
rect 347866 6264 347872 6276
rect 347924 6264 347930 6316
rect 136542 6196 136548 6248
rect 136600 6236 136606 6248
rect 188430 6236 188436 6248
rect 136600 6208 188436 6236
rect 136600 6196 136606 6208
rect 188430 6196 188436 6208
rect 188488 6196 188494 6248
rect 193030 6196 193036 6248
rect 193088 6236 193094 6248
rect 351362 6236 351368 6248
rect 193088 6208 351368 6236
rect 193088 6196 193094 6208
rect 351362 6196 351368 6208
rect 351420 6196 351426 6248
rect 136450 6128 136456 6180
rect 136508 6168 136514 6180
rect 192018 6168 192024 6180
rect 136508 6140 192024 6168
rect 136508 6128 136514 6140
rect 192018 6128 192024 6140
rect 192076 6128 192082 6180
rect 193122 6128 193128 6180
rect 193180 6168 193186 6180
rect 354950 6168 354956 6180
rect 193180 6140 354956 6168
rect 193180 6128 193186 6140
rect 354950 6128 354956 6140
rect 355008 6128 355014 6180
rect 180702 6060 180708 6112
rect 180760 6100 180766 6112
rect 315758 6100 315764 6112
rect 180760 6072 315764 6100
rect 180760 6060 180766 6072
rect 315758 6060 315764 6072
rect 315816 6060 315822 6112
rect 179230 5992 179236 6044
rect 179288 6032 179294 6044
rect 312170 6032 312176 6044
rect 179288 6004 312176 6032
rect 179288 5992 179294 6004
rect 312170 5992 312176 6004
rect 312228 5992 312234 6044
rect 177942 5924 177948 5976
rect 178000 5964 178006 5976
rect 308582 5964 308588 5976
rect 178000 5936 308588 5964
rect 178000 5924 178006 5936
rect 308582 5924 308588 5936
rect 308640 5924 308646 5976
rect 176562 5856 176568 5908
rect 176620 5896 176626 5908
rect 305086 5896 305092 5908
rect 176620 5868 305092 5896
rect 176620 5856 176626 5868
rect 305086 5856 305092 5868
rect 305144 5856 305150 5908
rect 175090 5788 175096 5840
rect 175148 5828 175154 5840
rect 301406 5828 301412 5840
rect 175148 5800 301412 5828
rect 175148 5788 175154 5800
rect 301406 5788 301412 5800
rect 301464 5788 301470 5840
rect 173802 5720 173808 5772
rect 173860 5760 173866 5772
rect 297910 5760 297916 5772
rect 173860 5732 297916 5760
rect 173860 5720 173866 5732
rect 297910 5720 297916 5732
rect 297968 5720 297974 5772
rect 172422 5652 172428 5704
rect 172480 5692 172486 5704
rect 294322 5692 294328 5704
rect 172480 5664 294328 5692
rect 172480 5652 172486 5664
rect 294322 5652 294328 5664
rect 294380 5652 294386 5704
rect 171042 5584 171048 5636
rect 171100 5624 171106 5636
rect 290734 5624 290740 5636
rect 171100 5596 290740 5624
rect 171100 5584 171106 5596
rect 290734 5584 290740 5596
rect 290792 5584 290798 5636
rect 157150 5516 157156 5568
rect 157208 5556 157214 5568
rect 157337 5559 157395 5565
rect 157337 5556 157349 5559
rect 157208 5528 157349 5556
rect 157208 5516 157214 5528
rect 157337 5525 157349 5528
rect 157383 5525 157395 5559
rect 157337 5519 157395 5525
rect 169662 5516 169668 5568
rect 169720 5556 169726 5568
rect 286962 5556 286968 5568
rect 169720 5528 286968 5556
rect 169720 5516 169726 5528
rect 286962 5516 286968 5528
rect 287020 5516 287026 5568
rect 287054 5516 287060 5568
rect 287112 5556 287118 5568
rect 288342 5556 288348 5568
rect 287112 5528 288348 5556
rect 287112 5516 287118 5528
rect 288342 5516 288348 5528
rect 288400 5516 288406 5568
rect 367738 5516 367744 5568
rect 367796 5556 367802 5568
rect 368198 5556 368204 5568
rect 367796 5528 368204 5556
rect 367796 5516 367802 5528
rect 368198 5516 368204 5528
rect 368256 5516 368262 5568
rect 148962 5448 148968 5500
rect 149020 5488 149026 5500
rect 226518 5488 226524 5500
rect 149020 5460 226524 5488
rect 149020 5448 149026 5460
rect 226518 5448 226524 5460
rect 226576 5448 226582 5500
rect 245378 5448 245384 5500
rect 245436 5488 245442 5500
rect 249429 5491 249487 5497
rect 249429 5488 249441 5491
rect 245436 5460 249441 5488
rect 245436 5448 245442 5460
rect 249429 5457 249441 5460
rect 249475 5457 249487 5491
rect 249429 5451 249487 5457
rect 252370 5448 252376 5500
rect 252428 5488 252434 5500
rect 526254 5488 526260 5500
rect 252428 5460 526260 5488
rect 252428 5448 252434 5460
rect 526254 5448 526260 5460
rect 526312 5448 526318 5500
rect 148870 5380 148876 5432
rect 148928 5420 148934 5432
rect 227714 5420 227720 5432
rect 148928 5392 227720 5420
rect 148928 5380 148934 5392
rect 227714 5380 227720 5392
rect 227772 5380 227778 5432
rect 253658 5380 253664 5432
rect 253716 5420 253722 5432
rect 529842 5420 529848 5432
rect 253716 5392 529848 5420
rect 253716 5380 253722 5392
rect 529842 5380 529848 5392
rect 529900 5380 529906 5432
rect 150250 5312 150256 5364
rect 150308 5352 150314 5364
rect 230106 5352 230112 5364
rect 150308 5324 230112 5352
rect 150308 5312 150314 5324
rect 230106 5312 230112 5324
rect 230164 5312 230170 5364
rect 249702 5312 249708 5364
rect 249760 5352 249766 5364
rect 258721 5355 258779 5361
rect 258721 5352 258733 5355
rect 249760 5324 258733 5352
rect 249760 5312 249766 5324
rect 258721 5321 258733 5324
rect 258767 5321 258779 5355
rect 258721 5315 258779 5321
rect 258813 5355 258871 5361
rect 258813 5321 258825 5355
rect 258859 5352 258871 5355
rect 533430 5352 533436 5364
rect 258859 5324 533436 5352
rect 258859 5321 258871 5324
rect 258813 5315 258871 5321
rect 533430 5312 533436 5324
rect 533488 5312 533494 5364
rect 58802 5244 58808 5296
rect 58860 5284 58866 5296
rect 89806 5284 89812 5296
rect 58860 5256 89812 5284
rect 58860 5244 58866 5256
rect 89806 5244 89812 5256
rect 89864 5244 89870 5296
rect 150342 5244 150348 5296
rect 150400 5284 150406 5296
rect 231302 5284 231308 5296
rect 150400 5256 231308 5284
rect 150400 5244 150406 5256
rect 231302 5244 231308 5256
rect 231360 5244 231366 5296
rect 256602 5244 256608 5296
rect 256660 5284 256666 5296
rect 536926 5284 536932 5296
rect 256660 5256 536932 5284
rect 256660 5244 256666 5256
rect 536926 5244 536932 5256
rect 536984 5244 536990 5296
rect 55214 5176 55220 5228
rect 55272 5216 55278 5228
rect 88426 5216 88432 5228
rect 55272 5188 88432 5216
rect 55272 5176 55278 5188
rect 88426 5176 88432 5188
rect 88484 5176 88490 5228
rect 151630 5176 151636 5228
rect 151688 5216 151694 5228
rect 233694 5216 233700 5228
rect 151688 5188 233700 5216
rect 151688 5176 151694 5188
rect 233694 5176 233700 5188
rect 233752 5176 233758 5228
rect 257982 5176 257988 5228
rect 258040 5216 258046 5228
rect 540514 5216 540520 5228
rect 258040 5188 540520 5216
rect 258040 5176 258046 5188
rect 540514 5176 540520 5188
rect 540572 5176 540578 5228
rect 51626 5108 51632 5160
rect 51684 5148 51690 5160
rect 87046 5148 87052 5160
rect 51684 5120 87052 5148
rect 51684 5108 51690 5120
rect 87046 5108 87052 5120
rect 87104 5108 87110 5160
rect 151722 5108 151728 5160
rect 151780 5148 151786 5160
rect 234798 5148 234804 5160
rect 151780 5120 234804 5148
rect 151780 5108 151786 5120
rect 234798 5108 234804 5120
rect 234856 5108 234862 5160
rect 247865 5151 247923 5157
rect 247865 5117 247877 5151
rect 247911 5148 247923 5151
rect 251450 5148 251456 5160
rect 247911 5120 251456 5148
rect 247911 5117 247923 5120
rect 247865 5111 247923 5117
rect 251450 5108 251456 5120
rect 251508 5108 251514 5160
rect 255130 5108 255136 5160
rect 255188 5148 255194 5160
rect 258813 5151 258871 5157
rect 258813 5148 258825 5151
rect 255188 5120 258825 5148
rect 255188 5108 255194 5120
rect 258813 5117 258825 5120
rect 258859 5117 258871 5151
rect 258813 5111 258871 5117
rect 260742 5108 260748 5160
rect 260800 5148 260806 5160
rect 268473 5151 268531 5157
rect 260800 5120 268424 5148
rect 260800 5108 260806 5120
rect 48222 5040 48228 5092
rect 48280 5080 48286 5092
rect 85666 5080 85672 5092
rect 48280 5052 85672 5080
rect 48280 5040 48286 5052
rect 85666 5040 85672 5052
rect 85724 5040 85730 5092
rect 116946 5040 116952 5092
rect 117004 5080 117010 5092
rect 117222 5080 117228 5092
rect 117004 5052 117228 5080
rect 117004 5040 117010 5052
rect 117222 5040 117228 5052
rect 117280 5040 117286 5092
rect 153102 5040 153108 5092
rect 153160 5080 153166 5092
rect 237190 5080 237196 5092
rect 153160 5052 237196 5080
rect 153160 5040 153166 5052
rect 237190 5040 237196 5052
rect 237248 5040 237254 5092
rect 242802 5040 242808 5092
rect 242860 5080 242866 5092
rect 248877 5083 248935 5089
rect 248877 5080 248889 5083
rect 242860 5052 248889 5080
rect 242860 5040 242866 5052
rect 248877 5049 248889 5052
rect 248923 5049 248935 5083
rect 248877 5043 248935 5049
rect 254857 5083 254915 5089
rect 254857 5049 254869 5083
rect 254903 5080 254915 5083
rect 264606 5080 264612 5092
rect 254903 5052 264612 5080
rect 254903 5049 254915 5052
rect 254857 5043 254915 5049
rect 264606 5040 264612 5052
rect 264664 5040 264670 5092
rect 264882 5040 264888 5092
rect 264940 5080 264946 5092
rect 268396 5080 268424 5120
rect 268473 5117 268485 5151
rect 268519 5148 268531 5151
rect 544102 5148 544108 5160
rect 268519 5120 544108 5148
rect 268519 5117 268531 5120
rect 268473 5111 268531 5117
rect 544102 5108 544108 5120
rect 544160 5108 544166 5160
rect 547690 5080 547696 5092
rect 264940 5052 268240 5080
rect 268396 5052 547696 5080
rect 264940 5040 264946 5052
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 72142 5012 72148 5024
rect 7708 4984 72148 5012
rect 7708 4972 7714 4984
rect 72142 4972 72148 4984
rect 72200 4972 72206 5024
rect 154482 4972 154488 5024
rect 154540 5012 154546 5024
rect 240778 5012 240784 5024
rect 154540 4984 240784 5012
rect 154540 4972 154546 4984
rect 240778 4972 240784 4984
rect 240836 4972 240842 5024
rect 244182 4972 244188 5024
rect 244240 5012 244246 5024
rect 249337 5015 249395 5021
rect 249337 5012 249349 5015
rect 244240 4984 249349 5012
rect 244240 4972 244246 4984
rect 249337 4981 249349 4984
rect 249383 4981 249395 5015
rect 249337 4975 249395 4981
rect 252462 4972 252468 5024
rect 252520 5012 252526 5024
rect 255041 5015 255099 5021
rect 255041 5012 255053 5015
rect 252520 4984 255053 5012
rect 252520 4972 252526 4984
rect 255041 4981 255053 4984
rect 255087 4981 255099 5015
rect 255041 4975 255099 4981
rect 257433 5015 257491 5021
rect 257433 4981 257445 5015
rect 257479 5012 257491 5015
rect 261018 5012 261024 5024
rect 257479 4984 261024 5012
rect 257479 4981 257491 4984
rect 257433 4975 257491 4981
rect 261018 4972 261024 4984
rect 261076 4972 261082 5024
rect 262122 4972 262128 5024
rect 262180 5012 262186 5024
rect 268013 5015 268071 5021
rect 268013 5012 268025 5015
rect 262180 4984 268025 5012
rect 262180 4972 262186 4984
rect 268013 4981 268025 4984
rect 268059 4981 268071 5015
rect 268013 4975 268071 4981
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 70762 4944 70768 4956
rect 2924 4916 70768 4944
rect 2924 4904 2930 4916
rect 70762 4904 70768 4916
rect 70820 4904 70826 4956
rect 155862 4904 155868 4956
rect 155920 4944 155926 4956
rect 244366 4944 244372 4956
rect 155920 4916 244372 4944
rect 155920 4904 155926 4916
rect 244366 4904 244372 4916
rect 244424 4904 244430 4956
rect 257525 4947 257583 4953
rect 257525 4944 257537 4947
rect 248800 4916 257537 4944
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 69014 4876 69020 4888
rect 624 4848 69020 4876
rect 624 4836 630 4848
rect 69014 4836 69020 4848
rect 69072 4836 69078 4888
rect 157242 4836 157248 4888
rect 157300 4876 157306 4888
rect 247954 4876 247960 4888
rect 157300 4848 247960 4876
rect 157300 4836 157306 4848
rect 247954 4836 247960 4848
rect 248012 4836 248018 4888
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 70486 4808 70492 4820
rect 1728 4780 70492 4808
rect 1728 4768 1734 4780
rect 70486 4768 70492 4780
rect 70544 4768 70550 4820
rect 157337 4811 157395 4817
rect 157337 4777 157349 4811
rect 157383 4808 157395 4811
rect 171781 4811 171839 4817
rect 171781 4808 171793 4811
rect 157383 4780 171793 4808
rect 157383 4777 157395 4780
rect 157337 4771 157395 4777
rect 171781 4777 171793 4780
rect 171827 4777 171839 4811
rect 171781 4771 171839 4777
rect 181441 4811 181499 4817
rect 181441 4777 181453 4811
rect 181487 4808 181499 4811
rect 195885 4811 195943 4817
rect 195885 4808 195897 4811
rect 181487 4780 195897 4808
rect 181487 4777 181499 4780
rect 181441 4771 181499 4777
rect 195885 4777 195897 4780
rect 195931 4777 195943 4811
rect 195885 4771 195943 4777
rect 195977 4811 196035 4817
rect 195977 4777 195989 4811
rect 196023 4808 196035 4811
rect 215110 4808 215116 4820
rect 196023 4780 215116 4808
rect 196023 4777 196035 4780
rect 195977 4771 196035 4777
rect 215110 4768 215116 4780
rect 215168 4768 215174 4820
rect 215205 4811 215263 4817
rect 215205 4777 215217 4811
rect 215251 4808 215263 4811
rect 215389 4811 215447 4817
rect 215389 4808 215401 4811
rect 215251 4780 215401 4808
rect 215251 4777 215263 4780
rect 215205 4771 215263 4777
rect 215389 4777 215401 4780
rect 215435 4777 215447 4811
rect 215389 4771 215447 4777
rect 215570 4768 215576 4820
rect 215628 4808 215634 4820
rect 229557 4811 229615 4817
rect 229557 4808 229569 4811
rect 215628 4780 229569 4808
rect 215628 4768 215634 4780
rect 229557 4777 229569 4780
rect 229603 4777 229615 4811
rect 229557 4771 229615 4777
rect 229741 4811 229799 4817
rect 229741 4777 229753 4811
rect 229787 4808 229799 4811
rect 229787 4780 239076 4808
rect 229787 4777 229799 4780
rect 229741 4771 229799 4777
rect 147582 4700 147588 4752
rect 147640 4740 147646 4752
rect 215297 4743 215355 4749
rect 215297 4740 215309 4743
rect 147640 4712 215309 4740
rect 147640 4700 147646 4712
rect 215297 4709 215309 4712
rect 215343 4709 215355 4743
rect 215297 4703 215355 4709
rect 215481 4743 215539 4749
rect 215481 4709 215493 4743
rect 215527 4740 215539 4743
rect 219345 4743 219403 4749
rect 215527 4712 219204 4740
rect 215527 4709 215539 4712
rect 215481 4703 215539 4709
rect 146202 4632 146208 4684
rect 146260 4672 146266 4684
rect 218974 4672 218980 4684
rect 146260 4644 218980 4672
rect 146260 4632 146266 4644
rect 218974 4632 218980 4644
rect 219032 4632 219038 4684
rect 219176 4681 219204 4712
rect 219345 4709 219357 4743
rect 219391 4740 219403 4743
rect 223025 4743 223083 4749
rect 223025 4740 223037 4743
rect 219391 4712 223037 4740
rect 219391 4709 219403 4712
rect 219345 4703 219403 4709
rect 223025 4709 223037 4712
rect 223071 4709 223083 4743
rect 223025 4703 223083 4709
rect 225064 4712 229876 4740
rect 219161 4675 219219 4681
rect 219161 4641 219173 4675
rect 219207 4641 219219 4675
rect 219161 4635 219219 4641
rect 219250 4632 219256 4684
rect 219308 4672 219314 4684
rect 225064 4672 225092 4712
rect 219308 4644 225092 4672
rect 219308 4632 219314 4644
rect 144730 4564 144736 4616
rect 144788 4604 144794 4616
rect 215846 4604 215852 4616
rect 144788 4576 215852 4604
rect 144788 4564 144794 4576
rect 215846 4564 215852 4576
rect 215904 4564 215910 4616
rect 222930 4604 222936 4616
rect 215956 4576 222936 4604
rect 144638 4496 144644 4548
rect 144696 4536 144702 4548
rect 212258 4536 212264 4548
rect 144696 4508 212264 4536
rect 144696 4496 144702 4508
rect 212258 4496 212264 4508
rect 212316 4496 212322 4548
rect 212353 4539 212411 4545
rect 212353 4505 212365 4539
rect 212399 4536 212411 4539
rect 215110 4536 215116 4548
rect 212399 4508 215116 4536
rect 212399 4505 212411 4508
rect 212353 4499 212411 4505
rect 215110 4496 215116 4508
rect 215168 4496 215174 4548
rect 215389 4539 215447 4545
rect 215389 4505 215401 4539
rect 215435 4536 215447 4539
rect 215956 4536 215984 4576
rect 222930 4564 222936 4576
rect 222988 4564 222994 4616
rect 223025 4607 223083 4613
rect 223025 4573 223037 4607
rect 223071 4604 223083 4607
rect 229741 4607 229799 4613
rect 229741 4604 229753 4607
rect 223071 4576 229753 4604
rect 223071 4573 223083 4576
rect 223025 4567 223083 4573
rect 229741 4573 229753 4576
rect 229787 4573 229799 4607
rect 229741 4567 229799 4573
rect 215435 4508 215984 4536
rect 215435 4505 215447 4508
rect 215389 4499 215447 4505
rect 216030 4496 216036 4548
rect 216088 4536 216094 4548
rect 219069 4539 219127 4545
rect 219069 4536 219081 4539
rect 216088 4508 219081 4536
rect 216088 4496 216094 4508
rect 219069 4505 219081 4508
rect 219115 4505 219127 4539
rect 219069 4499 219127 4505
rect 219161 4539 219219 4545
rect 219161 4505 219173 4539
rect 219207 4536 219219 4539
rect 229649 4539 229707 4545
rect 229649 4536 229661 4539
rect 219207 4508 229661 4536
rect 219207 4505 219219 4508
rect 219161 4499 219219 4505
rect 229649 4505 229661 4508
rect 229695 4505 229707 4539
rect 229848 4536 229876 4712
rect 239048 4604 239076 4780
rect 239125 4743 239183 4749
rect 239125 4709 239137 4743
rect 239171 4740 239183 4743
rect 247865 4743 247923 4749
rect 247865 4740 247877 4743
rect 239171 4712 247877 4740
rect 239171 4709 239183 4712
rect 239125 4703 239183 4709
rect 247865 4709 247877 4712
rect 247911 4709 247923 4743
rect 247865 4703 247923 4709
rect 239217 4675 239275 4681
rect 239217 4641 239229 4675
rect 239263 4672 239275 4675
rect 248800 4672 248828 4916
rect 257525 4913 257537 4916
rect 257571 4913 257583 4947
rect 257525 4907 257583 4913
rect 258261 4947 258319 4953
rect 258261 4913 258273 4947
rect 258307 4944 258319 4947
rect 268102 4944 268108 4956
rect 258307 4916 268108 4944
rect 258307 4913 258319 4916
rect 258261 4907 258319 4913
rect 268102 4904 268108 4916
rect 268160 4904 268166 4956
rect 268212 4944 268240 5052
rect 547690 5040 547696 5052
rect 547748 5040 547754 5092
rect 268289 5015 268347 5021
rect 268289 4981 268301 5015
rect 268335 5012 268347 5015
rect 551186 5012 551192 5024
rect 268335 4984 551192 5012
rect 268335 4981 268347 4984
rect 268289 4975 268347 4981
rect 551186 4972 551192 4984
rect 551244 4972 551250 5024
rect 561950 4944 561956 4956
rect 268212 4916 561956 4944
rect 561950 4904 561956 4916
rect 562008 4904 562014 4956
rect 258077 4879 258135 4885
rect 258077 4876 258089 4879
rect 239263 4644 248828 4672
rect 248892 4848 258089 4876
rect 239263 4641 239275 4644
rect 239217 4635 239275 4641
rect 248892 4604 248920 4848
rect 258077 4845 258089 4848
rect 258123 4845 258135 4879
rect 258077 4839 258135 4845
rect 259270 4836 259276 4888
rect 259328 4876 259334 4888
rect 268473 4879 268531 4885
rect 268473 4876 268485 4879
rect 259328 4848 268485 4876
rect 259328 4836 259334 4848
rect 268473 4845 268485 4848
rect 268519 4845 268531 4879
rect 268473 4839 268531 4845
rect 268746 4836 268752 4888
rect 268804 4876 268810 4888
rect 572622 4876 572628 4888
rect 268804 4848 572628 4876
rect 268804 4836 268810 4848
rect 572622 4836 572628 4848
rect 572680 4836 572686 4888
rect 254857 4811 254915 4817
rect 254857 4808 254869 4811
rect 239048 4576 248920 4604
rect 248984 4780 254869 4808
rect 234617 4539 234675 4545
rect 229848 4508 234568 4536
rect 229649 4499 229707 4505
rect 143442 4428 143448 4480
rect 143500 4468 143506 4480
rect 208670 4468 208676 4480
rect 143500 4440 208676 4468
rect 143500 4428 143506 4440
rect 208670 4428 208676 4440
rect 208728 4428 208734 4480
rect 209038 4428 209044 4480
rect 209096 4468 209102 4480
rect 211709 4471 211767 4477
rect 211709 4468 211721 4471
rect 209096 4440 211721 4468
rect 209096 4428 209102 4440
rect 211709 4437 211721 4440
rect 211755 4437 211767 4471
rect 211709 4431 211767 4437
rect 211798 4428 211804 4480
rect 211856 4468 211862 4480
rect 215205 4471 215263 4477
rect 215205 4468 215217 4471
rect 211856 4440 215217 4468
rect 211856 4428 211862 4440
rect 215205 4437 215217 4440
rect 215251 4437 215263 4471
rect 215205 4431 215263 4437
rect 215294 4428 215300 4480
rect 215352 4468 215358 4480
rect 225877 4471 225935 4477
rect 225877 4468 225889 4471
rect 215352 4440 225889 4468
rect 215352 4428 215358 4440
rect 225877 4437 225889 4440
rect 225923 4437 225935 4471
rect 225877 4431 225935 4437
rect 229557 4471 229615 4477
rect 229557 4437 229569 4471
rect 229603 4468 229615 4471
rect 234433 4471 234491 4477
rect 234433 4468 234445 4471
rect 229603 4440 234445 4468
rect 229603 4437 229615 4440
rect 229557 4431 229615 4437
rect 234433 4437 234445 4440
rect 234479 4437 234491 4471
rect 234540 4468 234568 4508
rect 234617 4505 234629 4539
rect 234663 4536 234675 4539
rect 239125 4539 239183 4545
rect 239125 4536 239137 4539
rect 234663 4508 239137 4536
rect 234663 4505 234675 4508
rect 234617 4499 234675 4505
rect 239125 4505 239137 4508
rect 239171 4505 239183 4539
rect 239125 4499 239183 4505
rect 239401 4539 239459 4545
rect 239401 4505 239413 4539
rect 239447 4536 239459 4539
rect 248984 4536 249012 4780
rect 254857 4777 254869 4780
rect 254903 4777 254915 4811
rect 257433 4811 257491 4817
rect 257433 4808 257445 4811
rect 254857 4771 254915 4777
rect 254964 4780 257445 4808
rect 249058 4700 249064 4752
rect 249116 4740 249122 4752
rect 254964 4740 254992 4780
rect 257433 4777 257445 4780
rect 257479 4777 257491 4811
rect 257433 4771 257491 4777
rect 257525 4811 257583 4817
rect 257525 4777 257537 4811
rect 257571 4808 257583 4811
rect 271690 4808 271696 4820
rect 257571 4780 271696 4808
rect 257571 4777 257583 4780
rect 257525 4771 257583 4777
rect 271690 4768 271696 4780
rect 271748 4768 271754 4820
rect 271782 4768 271788 4820
rect 271840 4808 271846 4820
rect 579798 4808 579804 4820
rect 271840 4780 579804 4808
rect 271840 4768 271846 4780
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 249116 4712 254992 4740
rect 255041 4743 255099 4749
rect 249116 4700 249122 4712
rect 255041 4709 255053 4743
rect 255087 4740 255099 4743
rect 522666 4740 522672 4752
rect 255087 4712 522672 4740
rect 255087 4709 255099 4712
rect 255041 4703 255099 4709
rect 522666 4700 522672 4712
rect 522724 4700 522730 4752
rect 251082 4632 251088 4684
rect 251140 4672 251146 4684
rect 519078 4672 519084 4684
rect 251140 4644 519084 4672
rect 251140 4632 251146 4644
rect 519078 4632 519084 4644
rect 519136 4632 519142 4684
rect 257430 4604 257436 4616
rect 239447 4508 249012 4536
rect 249076 4576 257436 4604
rect 239447 4505 239459 4508
rect 239401 4499 239459 4505
rect 239217 4471 239275 4477
rect 239217 4468 239229 4471
rect 234540 4440 239229 4468
rect 234433 4431 234491 4437
rect 239217 4437 239229 4440
rect 239263 4437 239275 4471
rect 244182 4468 244188 4480
rect 239217 4431 239275 4437
rect 239324 4440 244188 4468
rect 142062 4360 142068 4412
rect 142120 4400 142126 4412
rect 205082 4400 205088 4412
rect 142120 4372 205088 4400
rect 142120 4360 142126 4372
rect 205082 4360 205088 4372
rect 205140 4360 205146 4412
rect 205177 4403 205235 4409
rect 205177 4369 205189 4403
rect 205223 4400 205235 4403
rect 231854 4400 231860 4412
rect 205223 4372 231860 4400
rect 205223 4369 205235 4372
rect 205177 4363 205235 4369
rect 231854 4360 231860 4372
rect 231912 4360 231918 4412
rect 231949 4403 232007 4409
rect 231949 4369 231961 4403
rect 231995 4400 232007 4403
rect 232593 4403 232651 4409
rect 232593 4400 232605 4403
rect 231995 4372 232605 4400
rect 231995 4369 232007 4372
rect 231949 4363 232007 4369
rect 232593 4369 232605 4372
rect 232639 4369 232651 4403
rect 232593 4363 232651 4369
rect 232685 4403 232743 4409
rect 232685 4369 232697 4403
rect 232731 4400 232743 4403
rect 239324 4400 239352 4440
rect 244182 4428 244188 4440
rect 244240 4428 244246 4480
rect 244093 4403 244151 4409
rect 244093 4400 244105 4403
rect 232731 4372 239352 4400
rect 239416 4372 244105 4400
rect 232731 4369 232743 4372
rect 232685 4363 232743 4369
rect 140590 4292 140596 4344
rect 140648 4332 140654 4344
rect 201494 4332 201500 4344
rect 140648 4304 201500 4332
rect 140648 4292 140654 4304
rect 201494 4292 201500 4304
rect 201552 4292 201558 4344
rect 201589 4335 201647 4341
rect 201589 4301 201601 4335
rect 201635 4332 201647 4335
rect 204809 4335 204867 4341
rect 204809 4332 204821 4335
rect 201635 4304 204821 4332
rect 201635 4301 201647 4304
rect 201589 4295 201647 4301
rect 204809 4301 204821 4304
rect 204855 4301 204867 4335
rect 232498 4332 232504 4344
rect 204809 4295 204867 4301
rect 205284 4304 232504 4332
rect 132497 4267 132555 4273
rect 132497 4233 132509 4267
rect 132543 4264 132555 4267
rect 132543 4236 136312 4264
rect 132543 4233 132555 4236
rect 132497 4227 132555 4233
rect 127897 4199 127955 4205
rect 127897 4196 127909 4199
rect 127544 4168 127909 4196
rect 36170 4088 36176 4140
rect 36228 4128 36234 4140
rect 81526 4128 81532 4140
rect 36228 4100 81532 4128
rect 36228 4088 36234 4100
rect 81526 4088 81532 4100
rect 81584 4088 81590 4140
rect 81621 4131 81679 4137
rect 81621 4097 81633 4131
rect 81667 4128 81679 4131
rect 81667 4100 81940 4128
rect 81667 4097 81679 4100
rect 81621 4091 81679 4097
rect 34974 4020 34980 4072
rect 35032 4060 35038 4072
rect 81802 4060 81808 4072
rect 35032 4032 81808 4060
rect 35032 4020 35038 4032
rect 81802 4020 81808 4032
rect 81860 4020 81866 4072
rect 81912 4060 81940 4100
rect 82630 4088 82636 4140
rect 82688 4128 82694 4140
rect 84838 4128 84844 4140
rect 82688 4100 84844 4128
rect 82688 4088 82694 4100
rect 84838 4088 84844 4100
rect 84896 4088 84902 4140
rect 87322 4088 87328 4140
rect 87380 4128 87386 4140
rect 88242 4128 88248 4140
rect 87380 4100 88248 4128
rect 87380 4088 87386 4100
rect 88242 4088 88248 4100
rect 88300 4088 88306 4140
rect 89714 4088 89720 4140
rect 89772 4128 89778 4140
rect 91738 4128 91744 4140
rect 89772 4100 91744 4128
rect 89772 4088 89778 4100
rect 91738 4088 91744 4100
rect 91796 4088 91802 4140
rect 93302 4088 93308 4140
rect 93360 4128 93366 4140
rect 93762 4128 93768 4140
rect 93360 4100 93768 4128
rect 93360 4088 93366 4100
rect 93762 4088 93768 4100
rect 93820 4088 93826 4140
rect 94498 4088 94504 4140
rect 94556 4128 94562 4140
rect 95878 4128 95884 4140
rect 94556 4100 95884 4128
rect 94556 4088 94562 4100
rect 95878 4088 95884 4100
rect 95936 4088 95942 4140
rect 96890 4088 96896 4140
rect 96948 4128 96954 4140
rect 97902 4128 97908 4140
rect 96948 4100 97908 4128
rect 96948 4088 96954 4100
rect 97902 4088 97908 4100
rect 97960 4088 97966 4140
rect 102778 4088 102784 4140
rect 102836 4128 102842 4140
rect 103422 4128 103428 4140
rect 102836 4100 103428 4128
rect 102836 4088 102842 4100
rect 103422 4088 103428 4100
rect 103480 4088 103486 4140
rect 105170 4088 105176 4140
rect 105228 4128 105234 4140
rect 106274 4128 106280 4140
rect 105228 4100 106280 4128
rect 105228 4088 105234 4100
rect 106274 4088 106280 4100
rect 106332 4088 106338 4140
rect 106826 4088 106832 4140
rect 106884 4128 106890 4140
rect 107562 4128 107568 4140
rect 106884 4100 107568 4128
rect 106884 4088 106890 4100
rect 107562 4088 107568 4100
rect 107620 4088 107626 4140
rect 107838 4088 107844 4140
rect 107896 4128 107902 4140
rect 108758 4128 108764 4140
rect 107896 4100 108764 4128
rect 107896 4088 107902 4100
rect 108758 4088 108764 4100
rect 108816 4088 108822 4140
rect 125318 4088 125324 4140
rect 125376 4128 125382 4140
rect 127544 4128 127572 4168
rect 127897 4165 127909 4168
rect 127943 4165 127955 4199
rect 127897 4159 127955 4165
rect 134518 4156 134524 4208
rect 134576 4196 134582 4208
rect 136177 4199 136235 4205
rect 136177 4196 136189 4199
rect 134576 4168 136189 4196
rect 134576 4156 134582 4168
rect 136177 4165 136189 4168
rect 136223 4165 136235 4199
rect 136284 4196 136312 4236
rect 139302 4224 139308 4276
rect 139360 4264 139366 4276
rect 197998 4264 198004 4276
rect 139360 4236 198004 4264
rect 139360 4224 139366 4236
rect 197998 4224 198004 4236
rect 198056 4224 198062 4276
rect 202138 4224 202144 4276
rect 202196 4264 202202 4276
rect 205284 4264 205312 4304
rect 232498 4292 232504 4304
rect 232556 4292 232562 4344
rect 202196 4236 205312 4264
rect 205361 4267 205419 4273
rect 202196 4224 202202 4236
rect 205361 4233 205373 4267
rect 205407 4264 205419 4267
rect 225877 4267 225935 4273
rect 205407 4236 225828 4264
rect 205407 4233 205419 4236
rect 205361 4227 205419 4233
rect 157337 4199 157395 4205
rect 157337 4196 157349 4199
rect 136284 4168 145696 4196
rect 136177 4159 136235 4165
rect 145558 4128 145564 4140
rect 125376 4100 127572 4128
rect 127636 4100 145564 4128
rect 125376 4088 125382 4100
rect 84378 4060 84384 4072
rect 81912 4032 84384 4060
rect 84378 4020 84384 4032
rect 84436 4020 84442 4072
rect 86126 4020 86132 4072
rect 86184 4060 86190 4072
rect 89070 4060 89076 4072
rect 86184 4032 89076 4060
rect 86184 4020 86190 4032
rect 89070 4020 89076 4032
rect 89128 4020 89134 4072
rect 89165 4063 89223 4069
rect 89165 4029 89177 4063
rect 89211 4060 89223 4063
rect 91557 4063 91615 4069
rect 91557 4060 91569 4063
rect 89211 4032 91569 4060
rect 89211 4029 89223 4032
rect 89165 4023 89223 4029
rect 91557 4029 91569 4032
rect 91603 4029 91615 4063
rect 91557 4023 91615 4029
rect 91649 4063 91707 4069
rect 91649 4029 91661 4063
rect 91695 4060 91707 4063
rect 96706 4060 96712 4072
rect 91695 4032 96712 4060
rect 91695 4029 91707 4032
rect 91649 4023 91707 4029
rect 96706 4020 96712 4032
rect 96764 4020 96770 4072
rect 101582 4020 101588 4072
rect 101640 4060 101646 4072
rect 104986 4060 104992 4072
rect 101640 4032 104992 4060
rect 101640 4020 101646 4032
rect 104986 4020 104992 4032
rect 105044 4020 105050 4072
rect 114278 4020 114284 4072
rect 114336 4060 114342 4072
rect 127526 4060 127532 4072
rect 114336 4032 127532 4060
rect 114336 4020 114342 4032
rect 127526 4020 127532 4032
rect 127584 4020 127590 4072
rect 30282 3952 30288 4004
rect 30340 3992 30346 4004
rect 80330 3992 80336 4004
rect 30340 3964 80336 3992
rect 30340 3952 30346 3964
rect 80330 3952 80336 3964
rect 80388 3952 80394 4004
rect 81434 3952 81440 4004
rect 81492 3992 81498 4004
rect 88978 3992 88984 4004
rect 81492 3964 88984 3992
rect 81492 3952 81498 3964
rect 88978 3952 88984 3964
rect 89036 3952 89042 4004
rect 89257 3995 89315 4001
rect 89257 3961 89269 3995
rect 89303 3992 89315 3995
rect 96614 3992 96620 4004
rect 89303 3964 96620 3992
rect 89303 3961 89315 3964
rect 89257 3955 89315 3961
rect 96614 3952 96620 3964
rect 96672 3952 96678 4004
rect 110322 3952 110328 4004
rect 110380 3992 110386 4004
rect 114738 3992 114744 4004
rect 110380 3964 114744 3992
rect 110380 3952 110386 3964
rect 114738 3952 114744 3964
rect 114796 3952 114802 4004
rect 115658 3952 115664 4004
rect 115716 3992 115722 4004
rect 127437 3995 127495 4001
rect 127437 3992 127449 3995
rect 115716 3964 127449 3992
rect 115716 3952 115722 3964
rect 127437 3961 127449 3964
rect 127483 3961 127495 3995
rect 127437 3955 127495 3961
rect 27890 3884 27896 3936
rect 27948 3924 27954 3936
rect 70673 3927 70731 3933
rect 70673 3924 70685 3927
rect 27948 3896 70685 3924
rect 27948 3884 27954 3896
rect 70673 3893 70685 3896
rect 70719 3893 70731 3927
rect 70673 3887 70731 3893
rect 71866 3884 71872 3936
rect 71924 3924 71930 3936
rect 79965 3927 80023 3933
rect 79965 3924 79977 3927
rect 71924 3896 79977 3924
rect 71924 3884 71930 3896
rect 79965 3893 79977 3896
rect 80011 3893 80023 3927
rect 79965 3887 80023 3893
rect 80054 3884 80060 3936
rect 80112 3924 80118 3936
rect 81621 3927 81679 3933
rect 81621 3924 81633 3927
rect 80112 3896 81633 3924
rect 80112 3884 80118 3896
rect 81621 3893 81633 3896
rect 81667 3893 81679 3927
rect 96982 3924 96988 3936
rect 81621 3887 81679 3893
rect 81820 3896 96988 3924
rect 20714 3816 20720 3868
rect 20772 3856 20778 3868
rect 76006 3856 76012 3868
rect 20772 3828 76012 3856
rect 20772 3816 20778 3828
rect 76006 3816 76012 3828
rect 76064 3816 76070 3868
rect 78858 3856 78864 3868
rect 76116 3828 78864 3856
rect 21910 3748 21916 3800
rect 21968 3788 21974 3800
rect 70489 3791 70547 3797
rect 70489 3788 70501 3791
rect 21968 3760 70501 3788
rect 21968 3748 21974 3760
rect 70489 3757 70501 3760
rect 70535 3757 70547 3791
rect 73154 3788 73160 3800
rect 70489 3751 70547 3757
rect 70596 3760 73160 3788
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 70596 3720 70624 3760
rect 73154 3748 73160 3760
rect 73212 3748 73218 3800
rect 76116 3788 76144 3828
rect 78858 3816 78864 3828
rect 78916 3816 78922 3868
rect 79042 3816 79048 3868
rect 79100 3856 79106 3868
rect 81820 3856 81848 3896
rect 96982 3884 96988 3896
rect 97040 3884 97046 3936
rect 100478 3884 100484 3936
rect 100536 3924 100542 3936
rect 103698 3924 103704 3936
rect 100536 3896 103704 3924
rect 100536 3884 100542 3896
rect 103698 3884 103704 3896
rect 103756 3884 103762 3936
rect 121362 3884 121368 3936
rect 121420 3924 121426 3936
rect 127636 3924 127664 4100
rect 145558 4088 145564 4100
rect 145616 4088 145622 4140
rect 145668 4128 145696 4168
rect 157168 4168 157349 4196
rect 153657 4131 153715 4137
rect 153657 4128 153669 4131
rect 145668 4100 153669 4128
rect 153657 4097 153669 4100
rect 153703 4097 153715 4131
rect 153657 4091 153715 4097
rect 153933 4131 153991 4137
rect 153933 4097 153945 4131
rect 153979 4128 153991 4131
rect 157168 4128 157196 4168
rect 157337 4165 157349 4168
rect 157383 4165 157395 4199
rect 157337 4159 157395 4165
rect 171781 4199 171839 4205
rect 171781 4165 171793 4199
rect 171827 4196 171839 4199
rect 181441 4199 181499 4205
rect 181441 4196 181453 4199
rect 171827 4168 181453 4196
rect 171827 4165 171839 4168
rect 171781 4159 171839 4165
rect 181441 4165 181453 4168
rect 181487 4165 181499 4199
rect 181441 4159 181499 4165
rect 193858 4156 193864 4208
rect 193916 4196 193922 4208
rect 225322 4196 225328 4208
rect 193916 4168 225328 4196
rect 193916 4156 193922 4168
rect 225322 4156 225328 4168
rect 225380 4156 225386 4208
rect 225800 4196 225828 4236
rect 225877 4233 225889 4267
rect 225923 4264 225935 4267
rect 231857 4267 231915 4273
rect 231857 4264 231869 4267
rect 225923 4236 231869 4264
rect 225923 4233 225935 4236
rect 225877 4227 225935 4233
rect 231857 4233 231869 4236
rect 231903 4233 231915 4267
rect 231857 4227 231915 4233
rect 231946 4224 231952 4276
rect 232004 4264 232010 4276
rect 239416 4264 239444 4372
rect 244093 4369 244105 4372
rect 244139 4369 244151 4403
rect 244093 4363 244151 4369
rect 244369 4403 244427 4409
rect 244369 4369 244381 4403
rect 244415 4400 244427 4403
rect 249076 4400 249104 4576
rect 257430 4564 257436 4576
rect 257488 4564 257494 4616
rect 258721 4607 258779 4613
rect 258721 4573 258733 4607
rect 258767 4604 258779 4607
rect 515582 4604 515588 4616
rect 258767 4576 515588 4604
rect 258767 4573 258779 4576
rect 258721 4567 258779 4573
rect 515582 4564 515588 4576
rect 515640 4564 515646 4616
rect 249613 4539 249671 4545
rect 249613 4505 249625 4539
rect 249659 4536 249671 4539
rect 511994 4536 512000 4548
rect 249659 4508 512000 4536
rect 249659 4505 249671 4508
rect 249613 4499 249671 4505
rect 511994 4496 512000 4508
rect 512052 4496 512058 4548
rect 249242 4428 249248 4480
rect 249300 4468 249306 4480
rect 508406 4468 508412 4480
rect 249300 4440 508412 4468
rect 249300 4428 249306 4440
rect 508406 4428 508412 4440
rect 508464 4428 508470 4480
rect 244415 4372 249104 4400
rect 249429 4403 249487 4409
rect 244415 4369 244427 4372
rect 244369 4363 244427 4369
rect 249429 4369 249441 4403
rect 249475 4400 249487 4403
rect 504818 4400 504824 4412
rect 249475 4372 504824 4400
rect 249475 4369 249487 4372
rect 249429 4363 249487 4369
rect 504818 4360 504824 4372
rect 504876 4360 504882 4412
rect 249337 4335 249395 4341
rect 249337 4301 249349 4335
rect 249383 4332 249395 4335
rect 501230 4332 501236 4344
rect 249383 4304 501236 4332
rect 249383 4301 249395 4304
rect 249337 4295 249395 4301
rect 501230 4292 501236 4304
rect 501288 4292 501294 4344
rect 232004 4236 239444 4264
rect 248877 4267 248935 4273
rect 232004 4224 232010 4236
rect 248877 4233 248889 4267
rect 248923 4264 248935 4267
rect 497734 4264 497740 4276
rect 248923 4236 497740 4264
rect 248923 4233 248935 4236
rect 248877 4227 248935 4233
rect 497734 4224 497740 4236
rect 497792 4224 497798 4276
rect 228910 4196 228916 4208
rect 225800 4168 228916 4196
rect 228910 4156 228916 4168
rect 228968 4156 228974 4208
rect 229649 4199 229707 4205
rect 229649 4165 229661 4199
rect 229695 4196 229707 4199
rect 239401 4199 239459 4205
rect 239401 4196 239413 4199
rect 229695 4168 239413 4196
rect 229695 4165 229707 4168
rect 229649 4159 229707 4165
rect 239401 4165 239413 4168
rect 239447 4165 239459 4199
rect 239401 4159 239459 4165
rect 241425 4199 241483 4205
rect 241425 4165 241437 4199
rect 241471 4196 241483 4199
rect 494146 4196 494152 4208
rect 241471 4168 494152 4196
rect 241471 4165 241483 4168
rect 241425 4159 241483 4165
rect 494146 4156 494152 4168
rect 494204 4156 494210 4208
rect 153979 4100 157196 4128
rect 157245 4131 157303 4137
rect 153979 4097 153991 4100
rect 153933 4091 153991 4097
rect 157245 4097 157257 4131
rect 157291 4128 157303 4131
rect 183738 4128 183744 4140
rect 157291 4100 183744 4128
rect 157291 4097 157303 4100
rect 157245 4091 157303 4097
rect 183738 4088 183744 4100
rect 183796 4088 183802 4140
rect 184750 4088 184756 4140
rect 184808 4128 184814 4140
rect 328822 4128 328828 4140
rect 184808 4100 328828 4128
rect 184808 4088 184814 4100
rect 328822 4088 328828 4100
rect 328880 4088 328886 4140
rect 340141 4131 340199 4137
rect 340141 4097 340153 4131
rect 340187 4128 340199 4131
rect 345014 4128 345020 4140
rect 340187 4100 345020 4128
rect 340187 4097 340199 4100
rect 340141 4091 340199 4097
rect 345014 4088 345020 4100
rect 345072 4088 345078 4140
rect 354582 4088 354588 4140
rect 354640 4128 354646 4140
rect 368014 4128 368020 4140
rect 354640 4100 368020 4128
rect 354640 4088 354646 4100
rect 368014 4088 368020 4100
rect 368072 4088 368078 4140
rect 368198 4088 368204 4140
rect 368256 4128 368262 4140
rect 369029 4131 369087 4137
rect 369029 4128 369041 4131
rect 368256 4100 369041 4128
rect 368256 4088 368262 4100
rect 369029 4097 369041 4100
rect 369075 4097 369087 4131
rect 369029 4091 369087 4097
rect 369118 4088 369124 4140
rect 369176 4128 369182 4140
rect 446582 4128 446588 4140
rect 369176 4100 446588 4128
rect 369176 4088 369182 4100
rect 446582 4088 446588 4100
rect 446640 4088 446646 4140
rect 128170 4020 128176 4072
rect 128228 4060 128234 4072
rect 132497 4063 132555 4069
rect 132497 4060 132509 4063
rect 128228 4032 132509 4060
rect 128228 4020 128234 4032
rect 132497 4029 132509 4032
rect 132543 4029 132555 4063
rect 132497 4023 132555 4029
rect 148318 4020 148324 4072
rect 148376 4060 148382 4072
rect 153013 4063 153071 4069
rect 153013 4060 153025 4063
rect 148376 4032 153025 4060
rect 148376 4020 148382 4032
rect 153013 4029 153025 4032
rect 153059 4029 153071 4063
rect 153013 4023 153071 4029
rect 153838 4020 153844 4072
rect 153896 4060 153902 4072
rect 156322 4060 156328 4072
rect 153896 4032 156328 4060
rect 153896 4020 153902 4032
rect 156322 4020 156328 4032
rect 156380 4020 156386 4072
rect 157337 4063 157395 4069
rect 157337 4029 157349 4063
rect 157383 4060 157395 4063
rect 164694 4060 164700 4072
rect 157383 4032 164700 4060
rect 157383 4029 157395 4032
rect 157337 4023 157395 4029
rect 164694 4020 164700 4032
rect 164752 4020 164758 4072
rect 164789 4063 164847 4069
rect 164789 4029 164801 4063
rect 164835 4060 164847 4063
rect 186038 4060 186044 4072
rect 164835 4032 186044 4060
rect 164835 4029 164847 4032
rect 164789 4023 164847 4029
rect 186038 4020 186044 4032
rect 186096 4020 186102 4072
rect 187602 4020 187608 4072
rect 187660 4060 187666 4072
rect 335906 4060 335912 4072
rect 187660 4032 335912 4060
rect 187660 4020 187666 4032
rect 335906 4020 335912 4032
rect 335964 4020 335970 4072
rect 335998 4020 336004 4072
rect 336056 4060 336062 4072
rect 364886 4060 364892 4072
rect 336056 4032 364892 4060
rect 336056 4020 336062 4032
rect 364886 4020 364892 4032
rect 364944 4020 364950 4072
rect 364978 4020 364984 4072
rect 365036 4060 365042 4072
rect 453666 4060 453672 4072
rect 365036 4032 453672 4060
rect 365036 4020 365042 4032
rect 453666 4020 453672 4032
rect 453724 4020 453730 4072
rect 127805 3995 127863 4001
rect 127805 3961 127817 3995
rect 127851 3992 127863 3995
rect 128998 3992 129004 4004
rect 127851 3964 129004 3992
rect 127851 3961 127863 3964
rect 127805 3955 127863 3961
rect 128998 3952 129004 3964
rect 129056 3952 129062 4004
rect 129642 3952 129648 4004
rect 129700 3992 129706 4004
rect 169386 3992 169392 4004
rect 129700 3964 169392 3992
rect 129700 3952 129706 3964
rect 169386 3952 169392 3964
rect 169444 3952 169450 4004
rect 195885 3995 195943 4001
rect 195885 3961 195897 3995
rect 195931 3992 195943 3995
rect 195977 3995 196035 4001
rect 195977 3992 195989 3995
rect 195931 3964 195989 3992
rect 195931 3961 195943 3964
rect 195885 3955 195943 3961
rect 195977 3961 195989 3964
rect 196023 3961 196035 3995
rect 195977 3955 196035 3961
rect 331858 3952 331864 4004
rect 331916 3992 331922 4004
rect 340141 3995 340199 4001
rect 340141 3992 340153 3995
rect 331916 3964 340153 3992
rect 331916 3952 331922 3964
rect 340141 3961 340153 3964
rect 340187 3961 340199 3995
rect 340141 3955 340199 3961
rect 340230 3952 340236 4004
rect 340288 3992 340294 4004
rect 382274 3992 382280 4004
rect 340288 3964 382280 3992
rect 340288 3952 340294 3964
rect 382274 3952 382280 3964
rect 382332 3952 382338 4004
rect 121420 3896 127664 3924
rect 127713 3927 127771 3933
rect 121420 3884 121426 3896
rect 127713 3893 127725 3927
rect 127759 3924 127771 3927
rect 149238 3924 149244 3936
rect 127759 3896 149244 3924
rect 127759 3893 127771 3896
rect 127713 3887 127771 3893
rect 149238 3884 149244 3896
rect 149296 3884 149302 3936
rect 151170 3884 151176 3936
rect 151228 3924 151234 3936
rect 155126 3924 155132 3936
rect 151228 3896 155132 3924
rect 151228 3884 151234 3896
rect 155126 3884 155132 3896
rect 155184 3884 155190 3936
rect 155221 3927 155279 3933
rect 155221 3893 155233 3927
rect 155267 3924 155279 3927
rect 190822 3924 190828 3936
rect 155267 3896 190828 3924
rect 155267 3893 155279 3896
rect 155221 3887 155279 3893
rect 190822 3884 190828 3896
rect 190880 3884 190886 3936
rect 194502 3884 194508 3936
rect 194560 3924 194566 3936
rect 357342 3924 357348 3936
rect 194560 3896 357348 3924
rect 194560 3884 194566 3896
rect 357342 3884 357348 3896
rect 357400 3884 357406 3936
rect 357805 3927 357863 3933
rect 357805 3893 357817 3927
rect 357851 3924 357863 3927
rect 360930 3924 360936 3936
rect 357851 3896 360936 3924
rect 357851 3893 357863 3896
rect 357805 3887 357863 3893
rect 360930 3884 360936 3896
rect 360988 3884 360994 3936
rect 361022 3884 361028 3936
rect 361080 3924 361086 3936
rect 369118 3924 369124 3936
rect 361080 3896 369124 3924
rect 361080 3884 361086 3896
rect 369118 3884 369124 3896
rect 369176 3884 369182 3936
rect 369213 3927 369271 3933
rect 369213 3893 369225 3927
rect 369259 3924 369271 3927
rect 369259 3896 371740 3924
rect 369259 3893 369271 3896
rect 369213 3887 369271 3893
rect 79100 3828 81848 3856
rect 82449 3859 82507 3865
rect 79100 3816 79106 3828
rect 82449 3825 82461 3859
rect 82495 3856 82507 3859
rect 95694 3856 95700 3868
rect 82495 3828 95700 3856
rect 82495 3825 82507 3828
rect 82449 3819 82507 3825
rect 95694 3816 95700 3828
rect 95752 3816 95758 3868
rect 111610 3816 111616 3868
rect 111668 3856 111674 3868
rect 119430 3856 119436 3868
rect 111668 3828 119436 3856
rect 111668 3816 111674 3828
rect 119430 3816 119436 3828
rect 119488 3816 119494 3868
rect 122650 3816 122656 3868
rect 122708 3856 122714 3868
rect 151538 3856 151544 3868
rect 122708 3828 151544 3856
rect 122708 3816 122714 3828
rect 151538 3816 151544 3828
rect 151596 3816 151602 3868
rect 152458 3816 152464 3868
rect 152516 3856 152522 3868
rect 194410 3856 194416 3868
rect 152516 3828 194416 3856
rect 152516 3816 152522 3828
rect 194410 3816 194416 3828
rect 194468 3816 194474 3868
rect 200022 3816 200028 3868
rect 200080 3856 200086 3868
rect 371602 3856 371608 3868
rect 200080 3828 371608 3856
rect 200080 3816 200086 3828
rect 371602 3816 371608 3828
rect 371660 3816 371666 3868
rect 371712 3856 371740 3896
rect 371878 3884 371884 3936
rect 371936 3924 371942 3936
rect 467926 3924 467932 3936
rect 371936 3896 467932 3924
rect 371936 3884 371942 3896
rect 467926 3884 467932 3896
rect 467984 3884 467990 3936
rect 378689 3859 378747 3865
rect 378689 3856 378701 3859
rect 371712 3828 378701 3856
rect 378689 3825 378701 3828
rect 378735 3825 378747 3859
rect 378689 3819 378747 3825
rect 378873 3859 378931 3865
rect 378873 3825 378885 3859
rect 378919 3856 378931 3859
rect 482278 3856 482284 3868
rect 378919 3828 482284 3856
rect 378919 3825 378931 3828
rect 378873 3819 378931 3825
rect 482278 3816 482284 3828
rect 482336 3816 482342 3868
rect 73264 3760 76144 3788
rect 76193 3791 76251 3797
rect 12492 3692 70624 3720
rect 70673 3723 70731 3729
rect 12492 3680 12498 3692
rect 70673 3689 70685 3723
rect 70719 3720 70731 3723
rect 73264 3720 73292 3760
rect 76193 3757 76205 3791
rect 76239 3788 76251 3791
rect 77478 3788 77484 3800
rect 76239 3760 77484 3788
rect 76239 3757 76251 3760
rect 76193 3751 76251 3757
rect 77478 3748 77484 3760
rect 77536 3748 77542 3800
rect 77846 3748 77852 3800
rect 77904 3788 77910 3800
rect 91649 3791 91707 3797
rect 91649 3788 91661 3791
rect 77904 3760 91661 3788
rect 77904 3748 77910 3760
rect 91649 3757 91661 3760
rect 91695 3757 91707 3791
rect 93946 3788 93952 3800
rect 91649 3751 91707 3757
rect 91848 3760 93952 3788
rect 70719 3692 73292 3720
rect 73709 3723 73767 3729
rect 70719 3689 70731 3692
rect 70673 3683 70731 3689
rect 73709 3689 73721 3723
rect 73755 3720 73767 3723
rect 79873 3723 79931 3729
rect 79873 3720 79885 3723
rect 73755 3692 79885 3720
rect 73755 3689 73767 3692
rect 73709 3683 73767 3689
rect 79873 3689 79885 3692
rect 79919 3689 79931 3723
rect 79873 3683 79931 3689
rect 79965 3723 80023 3729
rect 79965 3689 79977 3723
rect 80011 3720 80023 3723
rect 91848 3720 91876 3760
rect 93946 3748 93952 3760
rect 94004 3748 94010 3800
rect 115842 3748 115848 3800
rect 115900 3788 115906 3800
rect 130194 3788 130200 3800
rect 115900 3760 130200 3788
rect 115900 3748 115906 3760
rect 130194 3748 130200 3760
rect 130252 3748 130258 3800
rect 131022 3748 131028 3800
rect 131080 3788 131086 3800
rect 172974 3788 172980 3800
rect 131080 3760 172980 3788
rect 131080 3748 131086 3760
rect 172974 3748 172980 3760
rect 173032 3748 173038 3800
rect 201402 3748 201408 3800
rect 201460 3788 201466 3800
rect 378778 3788 378784 3800
rect 201460 3760 378784 3788
rect 201460 3748 201466 3760
rect 378778 3748 378784 3760
rect 378836 3748 378842 3800
rect 382366 3748 382372 3800
rect 382424 3788 382430 3800
rect 383562 3788 383568 3800
rect 382424 3760 383568 3788
rect 382424 3748 382430 3760
rect 383562 3748 383568 3760
rect 383620 3748 383626 3800
rect 80011 3692 91876 3720
rect 80011 3689 80023 3692
rect 79965 3683 80023 3689
rect 92106 3680 92112 3732
rect 92164 3720 92170 3732
rect 100110 3720 100116 3732
rect 92164 3692 100116 3720
rect 92164 3680 92170 3692
rect 100110 3680 100116 3692
rect 100168 3680 100174 3732
rect 115750 3680 115756 3732
rect 115808 3720 115814 3732
rect 131390 3720 131396 3732
rect 115808 3692 131396 3720
rect 115808 3680 115814 3692
rect 131390 3680 131396 3692
rect 131448 3680 131454 3732
rect 132402 3680 132408 3732
rect 132460 3720 132466 3732
rect 176562 3720 176568 3732
rect 132460 3692 176568 3720
rect 132460 3680 132466 3692
rect 176562 3680 176568 3692
rect 176620 3680 176626 3732
rect 179322 3680 179328 3732
rect 179380 3720 179386 3732
rect 180245 3723 180303 3729
rect 180245 3720 180257 3723
rect 179380 3692 180257 3720
rect 179380 3680 179386 3692
rect 180245 3689 180257 3692
rect 180291 3689 180303 3723
rect 180245 3683 180303 3689
rect 204162 3680 204168 3732
rect 204220 3720 204226 3732
rect 385862 3720 385868 3732
rect 204220 3692 385868 3720
rect 204220 3680 204226 3692
rect 385862 3680 385868 3692
rect 385920 3680 385926 3732
rect 390554 3680 390560 3732
rect 390612 3720 390618 3732
rect 391842 3720 391848 3732
rect 390612 3692 391848 3720
rect 390612 3680 390618 3692
rect 391842 3680 391848 3692
rect 391900 3680 391906 3732
rect 11238 3612 11244 3664
rect 11296 3652 11302 3664
rect 70305 3655 70363 3661
rect 70305 3652 70317 3655
rect 11296 3624 70317 3652
rect 11296 3612 11302 3624
rect 70305 3621 70317 3624
rect 70351 3621 70363 3655
rect 70305 3615 70363 3621
rect 70397 3655 70455 3661
rect 70397 3621 70409 3655
rect 70443 3652 70455 3655
rect 73246 3652 73252 3664
rect 70443 3624 73252 3652
rect 70443 3621 70455 3624
rect 70397 3615 70455 3621
rect 73246 3612 73252 3624
rect 73304 3612 73310 3664
rect 75454 3612 75460 3664
rect 75512 3652 75518 3664
rect 95234 3652 95240 3664
rect 75512 3624 95240 3652
rect 75512 3612 75518 3624
rect 95234 3612 95240 3624
rect 95292 3612 95298 3664
rect 98086 3612 98092 3664
rect 98144 3652 98150 3664
rect 102594 3652 102600 3664
rect 98144 3624 102600 3652
rect 98144 3612 98150 3624
rect 102594 3612 102600 3624
rect 102652 3612 102658 3664
rect 111150 3612 111156 3664
rect 111208 3652 111214 3664
rect 111208 3624 112484 3652
rect 111208 3612 111214 3624
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 71774 3584 71780 3596
rect 8904 3556 71780 3584
rect 8904 3544 8910 3556
rect 71774 3544 71780 3556
rect 71832 3544 71838 3596
rect 74258 3544 74264 3596
rect 74316 3584 74322 3596
rect 95418 3584 95424 3596
rect 74316 3556 95424 3584
rect 74316 3544 74322 3556
rect 95418 3544 95424 3556
rect 95476 3544 95482 3596
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 71958 3516 71964 3528
rect 6512 3488 71964 3516
rect 6512 3476 6518 3488
rect 71958 3476 71964 3488
rect 72016 3476 72022 3528
rect 73062 3476 73068 3528
rect 73120 3516 73126 3528
rect 95326 3516 95332 3528
rect 73120 3488 95332 3516
rect 73120 3476 73126 3488
rect 95326 3476 95332 3488
rect 95384 3476 95390 3528
rect 99282 3476 99288 3528
rect 99340 3516 99346 3528
rect 100018 3516 100024 3528
rect 99340 3488 100024 3516
rect 99340 3476 99346 3488
rect 100018 3476 100024 3488
rect 100076 3476 100082 3528
rect 103974 3476 103980 3528
rect 104032 3516 104038 3528
rect 104802 3516 104808 3528
rect 104032 3488 104808 3516
rect 104032 3476 104038 3488
rect 104802 3476 104808 3488
rect 104860 3476 104866 3528
rect 111058 3476 111064 3528
rect 111116 3516 111122 3528
rect 112346 3516 112352 3528
rect 111116 3488 112352 3516
rect 111116 3476 111122 3488
rect 112346 3476 112352 3488
rect 112404 3476 112410 3528
rect 112456 3516 112484 3624
rect 113082 3612 113088 3664
rect 113140 3652 113146 3664
rect 123018 3652 123024 3664
rect 113140 3624 123024 3652
rect 113140 3612 113146 3624
rect 123018 3612 123024 3624
rect 123076 3612 123082 3664
rect 127713 3655 127771 3661
rect 127713 3652 127725 3655
rect 123404 3624 127725 3652
rect 113818 3544 113824 3596
rect 113876 3584 113882 3596
rect 117130 3584 117136 3596
rect 113876 3556 117136 3584
rect 113876 3544 113882 3556
rect 117130 3544 117136 3556
rect 117188 3544 117194 3596
rect 123205 3587 123263 3593
rect 123205 3584 123217 3587
rect 118344 3556 123217 3584
rect 115934 3516 115940 3528
rect 112456 3488 115940 3516
rect 115934 3476 115940 3488
rect 115992 3476 115998 3528
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 70394 3448 70400 3460
rect 4120 3420 70400 3448
rect 4120 3408 4126 3420
rect 70394 3408 70400 3420
rect 70452 3408 70458 3460
rect 70489 3451 70547 3457
rect 70489 3417 70501 3451
rect 70535 3448 70547 3451
rect 71501 3451 71559 3457
rect 71501 3448 71513 3451
rect 70535 3420 71513 3448
rect 70535 3417 70547 3420
rect 70489 3411 70547 3417
rect 71501 3417 71513 3420
rect 71547 3417 71559 3451
rect 75181 3451 75239 3457
rect 75181 3448 75193 3451
rect 71501 3411 71559 3417
rect 71608 3420 75193 3448
rect 16022 3340 16028 3392
rect 16080 3380 16086 3392
rect 16482 3380 16488 3392
rect 16080 3352 16488 3380
rect 16080 3340 16086 3352
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 17862 3380 17868 3392
rect 17276 3352 17868 3380
rect 17276 3340 17282 3352
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 24302 3340 24308 3392
rect 24360 3380 24366 3392
rect 24762 3380 24768 3392
rect 24360 3352 24768 3380
rect 24360 3340 24366 3352
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 25498 3340 25504 3392
rect 25556 3380 25562 3392
rect 26142 3380 26148 3392
rect 25556 3352 26148 3380
rect 25556 3340 25562 3352
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 26694 3340 26700 3392
rect 26752 3380 26758 3392
rect 27522 3380 27528 3392
rect 26752 3352 27528 3380
rect 26752 3340 26758 3352
rect 27522 3340 27528 3352
rect 27580 3340 27586 3392
rect 33870 3340 33876 3392
rect 33928 3380 33934 3392
rect 34422 3380 34428 3392
rect 33928 3352 34428 3380
rect 33928 3340 33934 3352
rect 34422 3340 34428 3352
rect 34480 3340 34486 3392
rect 45373 3383 45431 3389
rect 45373 3349 45385 3383
rect 45419 3380 45431 3383
rect 55217 3383 55275 3389
rect 55217 3380 55229 3383
rect 45419 3352 55229 3380
rect 45419 3349 45431 3352
rect 45373 3343 45431 3349
rect 55217 3349 55229 3352
rect 55263 3349 55275 3383
rect 55217 3343 55275 3349
rect 64785 3383 64843 3389
rect 64785 3349 64797 3383
rect 64831 3380 64843 3383
rect 71608 3380 71636 3420
rect 75181 3417 75193 3420
rect 75227 3417 75239 3451
rect 75181 3411 75239 3417
rect 75273 3451 75331 3457
rect 75273 3417 75285 3451
rect 75319 3448 75331 3451
rect 76193 3451 76251 3457
rect 76193 3448 76205 3451
rect 75319 3420 76205 3448
rect 75319 3417 75331 3420
rect 75273 3411 75331 3417
rect 76193 3417 76205 3420
rect 76239 3417 76251 3451
rect 76193 3411 76251 3417
rect 76650 3408 76656 3460
rect 76708 3448 76714 3460
rect 79965 3451 80023 3457
rect 76708 3420 79916 3448
rect 76708 3408 76714 3420
rect 79778 3380 79784 3392
rect 64831 3352 71636 3380
rect 71700 3352 79784 3380
rect 64831 3349 64843 3352
rect 64785 3343 64843 3349
rect 45465 3315 45523 3321
rect 45465 3281 45477 3315
rect 45511 3312 45523 3315
rect 55309 3315 55367 3321
rect 55309 3312 55321 3315
rect 45511 3284 55321 3312
rect 45511 3281 45523 3284
rect 45465 3275 45523 3281
rect 55309 3281 55321 3284
rect 55355 3281 55367 3315
rect 55309 3275 55367 3281
rect 64601 3315 64659 3321
rect 64601 3281 64613 3315
rect 64647 3312 64659 3315
rect 71700 3312 71728 3352
rect 79778 3340 79784 3352
rect 79836 3340 79842 3392
rect 79888 3380 79916 3420
rect 79965 3417 79977 3451
rect 80011 3448 80023 3451
rect 93854 3448 93860 3460
rect 80011 3420 93860 3448
rect 80011 3417 80023 3420
rect 79965 3411 80023 3417
rect 93854 3408 93860 3420
rect 93912 3408 93918 3460
rect 95694 3408 95700 3460
rect 95752 3448 95758 3460
rect 96522 3448 96528 3460
rect 95752 3420 96528 3448
rect 95752 3408 95758 3420
rect 96522 3408 96528 3420
rect 96580 3408 96586 3460
rect 110230 3408 110236 3460
rect 110288 3448 110294 3460
rect 110288 3420 111288 3448
rect 110288 3408 110294 3420
rect 82449 3383 82507 3389
rect 82449 3380 82461 3383
rect 79888 3352 82461 3380
rect 82449 3349 82461 3352
rect 82495 3349 82507 3383
rect 82449 3343 82507 3349
rect 82538 3340 82544 3392
rect 82596 3380 82602 3392
rect 88426 3380 88432 3392
rect 82596 3352 88432 3380
rect 82596 3340 82602 3352
rect 88426 3340 88432 3352
rect 88484 3340 88490 3392
rect 88518 3340 88524 3392
rect 88576 3380 88582 3392
rect 91465 3383 91523 3389
rect 91465 3380 91477 3383
rect 88576 3352 91477 3380
rect 88576 3340 88582 3352
rect 91465 3349 91477 3352
rect 91511 3349 91523 3383
rect 91465 3343 91523 3349
rect 91557 3383 91615 3389
rect 91557 3349 91569 3383
rect 91603 3380 91615 3383
rect 98270 3380 98276 3392
rect 91603 3352 98276 3380
rect 91603 3349 91615 3352
rect 91557 3343 91615 3349
rect 98270 3340 98276 3352
rect 98328 3340 98334 3392
rect 108942 3340 108948 3392
rect 109000 3380 109006 3392
rect 111150 3380 111156 3392
rect 109000 3352 111156 3380
rect 109000 3340 109006 3352
rect 111150 3340 111156 3352
rect 111208 3340 111214 3392
rect 111260 3380 111288 3420
rect 111702 3408 111708 3460
rect 111760 3448 111766 3460
rect 118234 3448 118240 3460
rect 111760 3420 118240 3448
rect 111760 3408 111766 3420
rect 118234 3408 118240 3420
rect 118292 3408 118298 3460
rect 113542 3380 113548 3392
rect 111260 3352 113548 3380
rect 113542 3340 113548 3352
rect 113600 3340 113606 3392
rect 114370 3340 114376 3392
rect 114428 3380 114434 3392
rect 118344 3380 118372 3556
rect 123205 3553 123217 3556
rect 123251 3553 123263 3587
rect 123205 3547 123263 3553
rect 122558 3476 122564 3528
rect 122616 3516 122622 3528
rect 123404 3516 123432 3624
rect 127713 3621 127725 3624
rect 127759 3621 127771 3655
rect 127713 3615 127771 3621
rect 127805 3655 127863 3661
rect 127805 3621 127817 3655
rect 127851 3652 127863 3655
rect 153930 3652 153936 3664
rect 127851 3624 153936 3652
rect 127851 3621 127863 3624
rect 127805 3615 127863 3621
rect 153930 3612 153936 3624
rect 153988 3612 153994 3664
rect 155218 3612 155224 3664
rect 155276 3652 155282 3664
rect 199194 3652 199200 3664
rect 155276 3624 199200 3652
rect 155276 3612 155282 3624
rect 199194 3612 199200 3624
rect 199252 3612 199258 3664
rect 208302 3612 208308 3664
rect 208360 3652 208366 3664
rect 396626 3652 396632 3664
rect 208360 3624 396632 3652
rect 208360 3612 208366 3624
rect 396626 3612 396632 3624
rect 396684 3612 396690 3664
rect 408494 3612 408500 3664
rect 408552 3652 408558 3664
rect 409690 3652 409696 3664
rect 408552 3624 409696 3652
rect 408552 3612 408558 3624
rect 409690 3612 409696 3624
rect 409748 3612 409754 3664
rect 123573 3587 123631 3593
rect 123573 3553 123585 3587
rect 123619 3584 123631 3587
rect 126606 3584 126612 3596
rect 123619 3556 126612 3584
rect 123619 3553 123631 3556
rect 123573 3547 123631 3553
rect 126606 3544 126612 3556
rect 126664 3544 126670 3596
rect 126882 3544 126888 3596
rect 126940 3584 126946 3596
rect 162302 3584 162308 3596
rect 126940 3556 162308 3584
rect 126940 3544 126946 3556
rect 162302 3544 162308 3556
rect 162360 3544 162366 3596
rect 162397 3587 162455 3593
rect 162397 3553 162409 3587
rect 162443 3584 162455 3587
rect 164786 3584 164792 3596
rect 162443 3556 164792 3584
rect 162443 3553 162455 3556
rect 162397 3547 162455 3553
rect 164786 3544 164792 3556
rect 164844 3544 164850 3596
rect 164878 3544 164884 3596
rect 164936 3584 164942 3596
rect 167086 3584 167092 3596
rect 164936 3556 167092 3584
rect 164936 3544 164942 3556
rect 167086 3544 167092 3556
rect 167144 3544 167150 3596
rect 167638 3544 167644 3596
rect 167696 3584 167702 3596
rect 168282 3584 168288 3596
rect 167696 3556 168288 3584
rect 167696 3544 167702 3556
rect 168282 3544 168288 3556
rect 168340 3544 168346 3596
rect 169021 3587 169079 3593
rect 169021 3553 169033 3587
rect 169067 3584 169079 3587
rect 211062 3584 211068 3596
rect 169067 3556 211068 3584
rect 169067 3553 169079 3556
rect 169021 3547 169079 3553
rect 211062 3544 211068 3556
rect 211120 3544 211126 3596
rect 213822 3544 213828 3596
rect 213880 3584 213886 3596
rect 414474 3584 414480 3596
rect 213880 3556 414480 3584
rect 213880 3544 213886 3556
rect 414474 3544 414480 3556
rect 414532 3544 414538 3596
rect 477494 3544 477500 3596
rect 477552 3584 477558 3596
rect 478690 3584 478696 3596
rect 477552 3556 478696 3584
rect 477552 3544 477558 3556
rect 478690 3544 478696 3556
rect 478748 3544 478754 3596
rect 122616 3488 123432 3516
rect 122616 3476 122622 3488
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124214 3516 124220 3528
rect 123536 3488 124220 3516
rect 123536 3476 123542 3488
rect 124214 3476 124220 3488
rect 124272 3476 124278 3528
rect 124306 3476 124312 3528
rect 124364 3516 124370 3528
rect 127529 3519 127587 3525
rect 127529 3516 127541 3519
rect 124364 3488 127541 3516
rect 124364 3476 124370 3488
rect 127529 3485 127541 3488
rect 127575 3485 127587 3519
rect 127529 3479 127587 3485
rect 127621 3519 127679 3525
rect 127621 3485 127633 3519
rect 127667 3516 127679 3519
rect 132957 3519 133015 3525
rect 132957 3516 132969 3519
rect 127667 3488 132969 3516
rect 127667 3485 127679 3488
rect 127621 3479 127679 3485
rect 132957 3485 132969 3488
rect 133003 3485 133015 3519
rect 132957 3479 133015 3485
rect 133230 3476 133236 3528
rect 133288 3516 133294 3528
rect 136082 3516 136088 3528
rect 133288 3488 136088 3516
rect 133288 3476 133294 3488
rect 136082 3476 136088 3488
rect 136140 3476 136146 3528
rect 136177 3519 136235 3525
rect 136177 3485 136189 3519
rect 136223 3516 136235 3519
rect 138661 3519 138719 3525
rect 138661 3516 138673 3519
rect 136223 3488 138673 3516
rect 136223 3485 136235 3488
rect 136177 3479 136235 3485
rect 138661 3485 138673 3488
rect 138707 3485 138719 3519
rect 138661 3479 138719 3485
rect 141418 3476 141424 3528
rect 141476 3516 141482 3528
rect 144454 3516 144460 3528
rect 141476 3488 144460 3516
rect 141476 3476 141482 3488
rect 144454 3476 144460 3488
rect 144512 3476 144518 3528
rect 145650 3476 145656 3528
rect 145708 3516 145714 3528
rect 148042 3516 148048 3528
rect 145708 3488 148048 3516
rect 145708 3476 145714 3488
rect 148042 3476 148048 3488
rect 148100 3476 148106 3528
rect 148873 3519 148931 3525
rect 148873 3485 148885 3519
rect 148919 3516 148931 3519
rect 193214 3516 193220 3528
rect 148919 3488 193220 3516
rect 148919 3485 148931 3488
rect 148873 3479 148931 3485
rect 193214 3476 193220 3488
rect 193272 3476 193278 3528
rect 219158 3476 219164 3528
rect 219216 3516 219222 3528
rect 428734 3516 428740 3528
rect 219216 3488 428740 3516
rect 219216 3476 219222 3488
rect 428734 3476 428740 3488
rect 428792 3476 428798 3528
rect 433334 3476 433340 3528
rect 433392 3516 433398 3528
rect 434622 3516 434628 3528
rect 433392 3488 434628 3516
rect 433392 3476 433398 3488
rect 434622 3476 434628 3488
rect 434680 3476 434686 3528
rect 451274 3476 451280 3528
rect 451332 3516 451338 3528
rect 452470 3516 452476 3528
rect 451332 3488 452476 3516
rect 451332 3476 451338 3488
rect 452470 3476 452476 3488
rect 452528 3476 452534 3528
rect 502334 3476 502340 3528
rect 502392 3516 502398 3528
rect 503622 3516 503628 3528
rect 502392 3488 503628 3516
rect 502392 3476 502398 3488
rect 503622 3476 503628 3488
rect 503680 3476 503686 3528
rect 520274 3476 520280 3528
rect 520332 3516 520338 3528
rect 521470 3516 521476 3528
rect 520332 3488 521476 3516
rect 520332 3476 520338 3488
rect 521470 3476 521476 3488
rect 521528 3476 521534 3528
rect 563054 3476 563060 3528
rect 563112 3516 563118 3528
rect 564342 3516 564348 3528
rect 563112 3488 564348 3516
rect 563112 3476 563118 3488
rect 564342 3476 564348 3488
rect 564400 3476 564406 3528
rect 580994 3476 581000 3528
rect 581052 3516 581058 3528
rect 582190 3516 582196 3528
rect 581052 3488 582196 3516
rect 581052 3476 581058 3488
rect 582190 3476 582196 3488
rect 582248 3476 582254 3528
rect 118602 3408 118608 3460
rect 118660 3448 118666 3460
rect 133049 3451 133107 3457
rect 133049 3448 133061 3451
rect 118660 3420 133061 3448
rect 118660 3408 118666 3420
rect 133049 3417 133061 3420
rect 133095 3417 133107 3451
rect 133049 3411 133107 3417
rect 133138 3408 133144 3460
rect 133196 3448 133202 3460
rect 139670 3448 139676 3460
rect 133196 3420 139676 3448
rect 133196 3408 133202 3420
rect 139670 3408 139676 3420
rect 139728 3408 139734 3460
rect 140682 3408 140688 3460
rect 140740 3448 140746 3460
rect 200390 3448 200396 3460
rect 140740 3420 200396 3448
rect 140740 3408 140746 3420
rect 200390 3408 200396 3420
rect 200448 3408 200454 3460
rect 222102 3408 222108 3460
rect 222160 3448 222166 3460
rect 435818 3448 435824 3460
rect 222160 3420 435824 3448
rect 222160 3408 222166 3420
rect 435818 3408 435824 3420
rect 435876 3408 435882 3460
rect 114428 3352 118372 3380
rect 114428 3340 114434 3352
rect 118510 3340 118516 3392
rect 118568 3380 118574 3392
rect 122009 3383 122067 3389
rect 118568 3352 121960 3380
rect 118568 3340 118574 3352
rect 84470 3312 84476 3324
rect 64647 3284 71728 3312
rect 71792 3284 84476 3312
rect 64647 3281 64659 3284
rect 64601 3275 64659 3281
rect 45738 3204 45744 3256
rect 45796 3244 45802 3256
rect 46842 3244 46848 3256
rect 45796 3216 46848 3244
rect 45796 3204 45802 3216
rect 46842 3204 46848 3216
rect 46900 3204 46906 3256
rect 46934 3204 46940 3256
rect 46992 3244 46998 3256
rect 48130 3244 48136 3256
rect 46992 3216 48136 3244
rect 46992 3204 46998 3216
rect 48130 3204 48136 3216
rect 48188 3204 48194 3256
rect 50522 3204 50528 3256
rect 50580 3244 50586 3256
rect 50982 3244 50988 3256
rect 50580 3216 50988 3244
rect 50580 3204 50586 3216
rect 50982 3204 50988 3216
rect 51040 3204 51046 3256
rect 64693 3247 64751 3253
rect 64693 3213 64705 3247
rect 64739 3244 64751 3247
rect 71792 3244 71820 3284
rect 84470 3272 84476 3284
rect 84528 3272 84534 3324
rect 84930 3272 84936 3324
rect 84988 3312 84994 3324
rect 93118 3312 93124 3324
rect 84988 3284 93124 3312
rect 84988 3272 84994 3284
rect 93118 3272 93124 3284
rect 93176 3272 93182 3324
rect 116578 3272 116584 3324
rect 116636 3312 116642 3324
rect 121822 3312 121828 3324
rect 116636 3284 121828 3312
rect 116636 3272 116642 3284
rect 121822 3272 121828 3284
rect 121880 3272 121886 3324
rect 121932 3312 121960 3352
rect 122009 3349 122021 3383
rect 122055 3380 122067 3383
rect 125410 3380 125416 3392
rect 122055 3352 125416 3380
rect 122055 3349 122067 3352
rect 122009 3343 122067 3349
rect 125410 3340 125416 3352
rect 125468 3340 125474 3392
rect 125502 3340 125508 3392
rect 125560 3380 125566 3392
rect 127897 3383 127955 3389
rect 125560 3352 127756 3380
rect 125560 3340 125566 3352
rect 127621 3315 127679 3321
rect 127621 3312 127633 3315
rect 121932 3284 127633 3312
rect 127621 3281 127633 3284
rect 127667 3281 127679 3315
rect 127728 3312 127756 3352
rect 127897 3349 127909 3383
rect 127943 3380 127955 3383
rect 149057 3383 149115 3389
rect 149057 3380 149069 3383
rect 127943 3352 149069 3380
rect 127943 3349 127955 3352
rect 127897 3343 127955 3349
rect 149057 3349 149069 3352
rect 149103 3349 149115 3383
rect 149057 3343 149115 3349
rect 151262 3340 151268 3392
rect 151320 3380 151326 3392
rect 155221 3383 155279 3389
rect 155221 3380 155233 3383
rect 151320 3352 155233 3380
rect 151320 3340 151326 3352
rect 155221 3349 155233 3352
rect 155267 3349 155279 3383
rect 155221 3343 155279 3349
rect 159358 3340 159364 3392
rect 159416 3380 159422 3392
rect 164789 3383 164847 3389
rect 164789 3380 164801 3383
rect 159416 3352 164801 3380
rect 159416 3340 159422 3352
rect 164789 3349 164801 3352
rect 164835 3349 164847 3383
rect 164789 3343 164847 3349
rect 164878 3340 164884 3392
rect 164936 3380 164942 3392
rect 182542 3380 182548 3392
rect 164936 3352 182548 3380
rect 164936 3340 164942 3352
rect 182542 3340 182548 3352
rect 182600 3340 182606 3392
rect 278774 3340 278780 3392
rect 278832 3380 278838 3392
rect 280062 3380 280068 3392
rect 278832 3352 280068 3380
rect 278832 3340 278838 3352
rect 280062 3340 280068 3352
rect 280120 3340 280126 3392
rect 300118 3340 300124 3392
rect 300176 3380 300182 3392
rect 300176 3352 300440 3380
rect 300176 3340 300182 3352
rect 157518 3312 157524 3324
rect 127728 3284 157524 3312
rect 127621 3275 127679 3281
rect 157518 3272 157524 3284
rect 157576 3272 157582 3324
rect 157978 3272 157984 3324
rect 158036 3312 158042 3324
rect 158036 3284 158852 3312
rect 158036 3272 158042 3284
rect 64739 3216 71820 3244
rect 71869 3247 71927 3253
rect 64739 3213 64751 3216
rect 64693 3207 64751 3213
rect 71869 3213 71881 3247
rect 71915 3244 71927 3247
rect 75089 3247 75147 3253
rect 75089 3244 75101 3247
rect 71915 3216 75101 3244
rect 71915 3213 71927 3216
rect 71869 3207 71927 3213
rect 75089 3213 75101 3216
rect 75135 3213 75147 3247
rect 75089 3207 75147 3213
rect 75181 3247 75239 3253
rect 75181 3213 75193 3247
rect 75227 3244 75239 3247
rect 82998 3244 83004 3256
rect 75227 3216 83004 3244
rect 75227 3213 75239 3216
rect 75181 3207 75239 3213
rect 82998 3204 83004 3216
rect 83056 3204 83062 3256
rect 83826 3204 83832 3256
rect 83884 3244 83890 3256
rect 89165 3247 89223 3253
rect 89165 3244 89177 3247
rect 83884 3216 89177 3244
rect 83884 3204 83890 3216
rect 89165 3213 89177 3216
rect 89211 3213 89223 3247
rect 89165 3207 89223 3213
rect 91465 3247 91523 3253
rect 91465 3213 91477 3247
rect 91511 3244 91523 3247
rect 97258 3244 97264 3256
rect 91511 3216 97264 3244
rect 91511 3213 91523 3216
rect 91465 3207 91523 3213
rect 97258 3204 97264 3216
rect 97316 3204 97322 3256
rect 108850 3204 108856 3256
rect 108908 3244 108914 3256
rect 109954 3244 109960 3256
rect 108908 3216 109960 3244
rect 108908 3204 108914 3216
rect 109954 3204 109960 3216
rect 110012 3204 110018 3256
rect 124030 3204 124036 3256
rect 124088 3244 124094 3256
rect 127805 3247 127863 3253
rect 127805 3244 127817 3247
rect 124088 3216 127817 3244
rect 124088 3204 124094 3216
rect 127805 3213 127817 3216
rect 127851 3213 127863 3247
rect 127805 3207 127863 3213
rect 127897 3247 127955 3253
rect 127897 3213 127909 3247
rect 127943 3244 127955 3247
rect 148965 3247 149023 3253
rect 148965 3244 148977 3247
rect 127943 3216 148977 3244
rect 127943 3213 127955 3216
rect 127897 3207 127955 3213
rect 148965 3213 148977 3216
rect 149011 3213 149023 3247
rect 148965 3207 149023 3213
rect 149057 3247 149115 3253
rect 149057 3213 149069 3247
rect 149103 3244 149115 3247
rect 158714 3244 158720 3256
rect 149103 3216 158720 3244
rect 149103 3213 149115 3216
rect 149057 3207 149115 3213
rect 158714 3204 158720 3216
rect 158772 3204 158778 3256
rect 158824 3244 158852 3284
rect 159450 3272 159456 3324
rect 159508 3312 159514 3324
rect 162029 3315 162087 3321
rect 162029 3312 162041 3315
rect 159508 3284 162041 3312
rect 159508 3272 159514 3284
rect 162029 3281 162041 3284
rect 162075 3281 162087 3315
rect 162029 3275 162087 3281
rect 162121 3315 162179 3321
rect 162121 3281 162133 3315
rect 162167 3312 162179 3315
rect 170125 3315 170183 3321
rect 162167 3284 170076 3312
rect 162167 3281 162179 3284
rect 162121 3275 162179 3281
rect 162397 3247 162455 3253
rect 162397 3244 162409 3247
rect 158824 3216 162409 3244
rect 162397 3213 162409 3216
rect 162443 3213 162455 3247
rect 162397 3207 162455 3213
rect 162489 3247 162547 3253
rect 162489 3213 162501 3247
rect 162535 3244 162547 3247
rect 163409 3247 163467 3253
rect 163409 3244 163421 3247
rect 162535 3216 163421 3244
rect 162535 3213 162547 3216
rect 162489 3207 162547 3213
rect 163409 3213 163421 3216
rect 163455 3213 163467 3247
rect 163409 3207 163467 3213
rect 163498 3204 163504 3256
rect 163556 3244 163562 3256
rect 169021 3247 169079 3253
rect 169021 3244 169033 3247
rect 163556 3216 169033 3244
rect 163556 3204 163562 3216
rect 169021 3213 169033 3216
rect 169067 3213 169079 3247
rect 169021 3207 169079 3213
rect 44542 3136 44548 3188
rect 44600 3176 44606 3188
rect 44600 3148 45784 3176
rect 44600 3136 44606 3148
rect 43346 3068 43352 3120
rect 43404 3108 43410 3120
rect 45465 3111 45523 3117
rect 45465 3108 45477 3111
rect 43404 3080 45477 3108
rect 43404 3068 43410 3080
rect 45465 3077 45477 3080
rect 45511 3077 45523 3111
rect 45756 3108 45784 3148
rect 54018 3136 54024 3188
rect 54076 3176 54082 3188
rect 80146 3176 80152 3188
rect 54076 3148 80152 3176
rect 54076 3136 54082 3148
rect 80146 3136 80152 3148
rect 80204 3136 80210 3188
rect 80238 3136 80244 3188
rect 80296 3176 80302 3188
rect 89257 3179 89315 3185
rect 89257 3176 89269 3179
rect 80296 3148 89269 3176
rect 80296 3136 80302 3148
rect 89257 3145 89269 3148
rect 89303 3145 89315 3179
rect 89257 3139 89315 3145
rect 114462 3136 114468 3188
rect 114520 3176 114526 3188
rect 122009 3179 122067 3185
rect 122009 3176 122021 3179
rect 114520 3148 122021 3176
rect 114520 3136 114526 3148
rect 122009 3145 122021 3148
rect 122055 3145 122067 3179
rect 122009 3139 122067 3145
rect 122742 3136 122748 3188
rect 122800 3176 122806 3188
rect 150434 3176 150440 3188
rect 122800 3148 150440 3176
rect 122800 3136 122806 3148
rect 150434 3136 150440 3148
rect 150492 3136 150498 3188
rect 153013 3179 153071 3185
rect 153013 3145 153025 3179
rect 153059 3176 153071 3179
rect 157245 3179 157303 3185
rect 157245 3176 157257 3179
rect 153059 3148 157257 3176
rect 153059 3145 153071 3148
rect 153013 3139 153071 3145
rect 157245 3145 157257 3148
rect 157291 3145 157303 3179
rect 157245 3139 157303 3145
rect 158625 3179 158683 3185
rect 158625 3145 158637 3179
rect 158671 3176 158683 3179
rect 161106 3176 161112 3188
rect 158671 3148 161112 3176
rect 158671 3145 158683 3148
rect 158625 3139 158683 3145
rect 161106 3136 161112 3148
rect 161164 3136 161170 3188
rect 161201 3179 161259 3185
rect 161201 3145 161213 3179
rect 161247 3176 161259 3179
rect 168190 3176 168196 3188
rect 161247 3148 168196 3176
rect 161247 3145 161259 3148
rect 161201 3139 161259 3145
rect 168190 3136 168196 3148
rect 168248 3136 168254 3188
rect 168282 3136 168288 3188
rect 168340 3176 168346 3188
rect 169941 3179 169999 3185
rect 169941 3176 169953 3179
rect 168340 3148 169953 3176
rect 168340 3136 168346 3148
rect 169941 3145 169953 3148
rect 169987 3145 169999 3179
rect 170048 3176 170076 3284
rect 170125 3281 170137 3315
rect 170171 3312 170183 3315
rect 170171 3284 171916 3312
rect 170171 3281 170183 3284
rect 170125 3275 170183 3281
rect 171888 3244 171916 3284
rect 175182 3272 175188 3324
rect 175240 3312 175246 3324
rect 300302 3312 300308 3324
rect 175240 3284 300308 3312
rect 175240 3272 175246 3284
rect 300302 3272 300308 3284
rect 300360 3272 300366 3324
rect 300412 3312 300440 3352
rect 304994 3340 305000 3392
rect 305052 3380 305058 3392
rect 306190 3380 306196 3392
rect 305052 3352 306196 3380
rect 305052 3340 305058 3352
rect 306190 3340 306196 3352
rect 306248 3340 306254 3392
rect 307018 3340 307024 3392
rect 307076 3380 307082 3392
rect 314749 3383 314807 3389
rect 314749 3380 314761 3383
rect 307076 3352 314761 3380
rect 307076 3340 307082 3352
rect 314749 3349 314761 3352
rect 314795 3349 314807 3383
rect 314749 3343 314807 3349
rect 329098 3340 329104 3392
rect 329156 3380 329162 3392
rect 357805 3383 357863 3389
rect 357805 3380 357817 3383
rect 329156 3352 357817 3380
rect 329156 3340 329162 3352
rect 357805 3349 357817 3352
rect 357851 3349 357863 3383
rect 359553 3383 359611 3389
rect 359553 3380 359565 3383
rect 357805 3343 357863 3349
rect 359292 3352 359565 3380
rect 310974 3312 310980 3324
rect 300412 3284 310980 3312
rect 310974 3272 310980 3284
rect 311032 3272 311038 3324
rect 311158 3272 311164 3324
rect 311216 3312 311222 3324
rect 325234 3312 325240 3324
rect 311216 3284 325240 3312
rect 311216 3272 311222 3284
rect 325234 3272 325240 3284
rect 325292 3272 325298 3324
rect 325326 3272 325332 3324
rect 325384 3312 325390 3324
rect 347685 3315 347743 3321
rect 347685 3312 347697 3315
rect 325384 3284 347697 3312
rect 325384 3272 325390 3284
rect 347685 3281 347697 3284
rect 347731 3281 347743 3315
rect 347685 3275 347743 3281
rect 347774 3272 347780 3324
rect 347832 3312 347838 3324
rect 349062 3312 349068 3324
rect 347832 3284 349068 3312
rect 347832 3272 347838 3284
rect 349062 3272 349068 3284
rect 349120 3272 349126 3324
rect 349157 3315 349215 3321
rect 349157 3281 349169 3315
rect 349203 3312 349215 3315
rect 359292 3312 359320 3352
rect 359553 3349 359565 3352
rect 359599 3349 359611 3383
rect 359553 3343 359611 3349
rect 359642 3340 359648 3392
rect 359700 3380 359706 3392
rect 439406 3380 439412 3392
rect 359700 3352 439412 3380
rect 359700 3340 359706 3352
rect 439406 3340 439412 3352
rect 439464 3340 439470 3392
rect 349203 3284 359320 3312
rect 359369 3315 359427 3321
rect 349203 3281 349215 3284
rect 349157 3275 349215 3281
rect 359369 3281 359381 3315
rect 359415 3312 359427 3315
rect 432322 3312 432328 3324
rect 359415 3284 432328 3312
rect 359415 3281 359427 3284
rect 359369 3275 359427 3281
rect 432322 3272 432328 3284
rect 432380 3272 432386 3324
rect 221734 3244 221740 3256
rect 171888 3216 221740 3244
rect 221734 3204 221740 3216
rect 221792 3204 221798 3256
rect 276658 3204 276664 3256
rect 276716 3244 276722 3256
rect 400214 3244 400220 3256
rect 276716 3216 400220 3244
rect 276716 3204 276722 3216
rect 400214 3204 400220 3216
rect 400272 3204 400278 3256
rect 203886 3176 203892 3188
rect 170048 3148 203892 3176
rect 169941 3139 169999 3145
rect 203886 3136 203892 3148
rect 203944 3136 203950 3188
rect 267366 3136 267372 3188
rect 267424 3176 267430 3188
rect 364518 3176 364524 3188
rect 267424 3148 364524 3176
rect 267424 3136 267430 3148
rect 364518 3136 364524 3148
rect 364576 3136 364582 3188
rect 365714 3136 365720 3188
rect 365772 3176 365778 3188
rect 366910 3176 366916 3188
rect 365772 3148 366916 3176
rect 365772 3136 365778 3148
rect 366910 3136 366916 3148
rect 366968 3136 366974 3188
rect 367002 3136 367008 3188
rect 367060 3176 367066 3188
rect 375190 3176 375196 3188
rect 367060 3148 375196 3176
rect 367060 3136 367066 3148
rect 375190 3136 375196 3148
rect 375248 3136 375254 3188
rect 375282 3136 375288 3188
rect 375340 3176 375346 3188
rect 378597 3179 378655 3185
rect 378597 3176 378609 3179
rect 375340 3148 378609 3176
rect 375340 3136 375346 3148
rect 378597 3145 378609 3148
rect 378643 3145 378655 3179
rect 378597 3139 378655 3145
rect 378689 3179 378747 3185
rect 378689 3145 378701 3179
rect 378735 3176 378747 3179
rect 460842 3176 460848 3188
rect 378735 3148 460848 3176
rect 378735 3145 378747 3148
rect 378689 3139 378747 3145
rect 460842 3136 460848 3148
rect 460900 3136 460906 3188
rect 62301 3111 62359 3117
rect 62301 3108 62313 3111
rect 45756 3080 62313 3108
rect 45465 3071 45523 3077
rect 62301 3077 62313 3080
rect 62347 3077 62359 3111
rect 62301 3071 62359 3077
rect 62390 3068 62396 3120
rect 62448 3108 62454 3120
rect 63402 3108 63408 3120
rect 62448 3080 63408 3108
rect 62448 3068 62454 3080
rect 63402 3068 63408 3080
rect 63460 3068 63466 3120
rect 91278 3108 91284 3120
rect 63512 3080 91284 3108
rect 37366 3000 37372 3052
rect 37424 3040 37430 3052
rect 45373 3043 45431 3049
rect 45373 3040 45385 3043
rect 37424 3012 45385 3040
rect 37424 3000 37430 3012
rect 45373 3009 45385 3012
rect 45419 3009 45431 3043
rect 45373 3003 45431 3009
rect 55309 3043 55367 3049
rect 55309 3009 55321 3043
rect 55355 3040 55367 3043
rect 61105 3043 61163 3049
rect 61105 3040 61117 3043
rect 55355 3012 61117 3040
rect 55355 3009 55367 3012
rect 55309 3003 55367 3009
rect 61105 3009 61117 3012
rect 61151 3009 61163 3043
rect 61105 3003 61163 3009
rect 61194 3000 61200 3052
rect 61252 3040 61258 3052
rect 63512 3040 63540 3080
rect 91278 3068 91284 3080
rect 91336 3068 91342 3120
rect 119890 3068 119896 3120
rect 119948 3108 119954 3120
rect 142062 3108 142068 3120
rect 119948 3080 142068 3108
rect 119948 3068 119954 3080
rect 142062 3068 142068 3080
rect 142120 3068 142126 3120
rect 145466 3068 145472 3120
rect 145524 3108 145530 3120
rect 151817 3111 151875 3117
rect 151817 3108 151829 3111
rect 145524 3080 151829 3108
rect 145524 3068 145530 3080
rect 151817 3077 151829 3080
rect 151863 3077 151875 3111
rect 151817 3071 151875 3077
rect 153838 3068 153844 3120
rect 153896 3108 153902 3120
rect 195606 3108 195612 3120
rect 153896 3080 195612 3108
rect 153896 3068 153902 3080
rect 195606 3068 195612 3080
rect 195664 3068 195670 3120
rect 257798 3068 257804 3120
rect 257856 3108 257862 3120
rect 350258 3108 350264 3120
rect 257856 3080 350264 3108
rect 257856 3068 257862 3080
rect 350258 3068 350264 3080
rect 350316 3068 350322 3120
rect 350353 3111 350411 3117
rect 350353 3077 350365 3111
rect 350399 3108 350411 3111
rect 353849 3111 353907 3117
rect 353849 3108 353861 3111
rect 350399 3080 353861 3108
rect 350399 3077 350411 3080
rect 350353 3071 350411 3077
rect 353849 3077 353861 3080
rect 353895 3077 353907 3111
rect 353849 3071 353907 3077
rect 353938 3068 353944 3120
rect 353996 3108 354002 3120
rect 359369 3111 359427 3117
rect 359369 3108 359381 3111
rect 353996 3080 359381 3108
rect 353996 3068 354002 3080
rect 359369 3077 359381 3080
rect 359415 3077 359427 3111
rect 425146 3108 425152 3120
rect 359369 3071 359427 3077
rect 359476 3080 425152 3108
rect 61252 3012 63540 3040
rect 61252 3000 61258 3012
rect 63586 3000 63592 3052
rect 63644 3040 63650 3052
rect 64690 3040 64696 3052
rect 63644 3012 64696 3040
rect 63644 3000 63650 3012
rect 64690 3000 64696 3012
rect 64748 3000 64754 3052
rect 89990 3040 89996 3052
rect 64892 3012 89996 3040
rect 59998 2932 60004 2984
rect 60056 2972 60062 2984
rect 64892 2972 64920 3012
rect 89990 3000 89996 3012
rect 90048 3000 90054 3052
rect 117038 3000 117044 3052
rect 117096 3040 117102 3052
rect 134886 3040 134892 3052
rect 117096 3012 134892 3040
rect 117096 3000 117102 3012
rect 134886 3000 134892 3012
rect 134944 3000 134950 3052
rect 135898 3000 135904 3052
rect 135956 3040 135962 3052
rect 137373 3043 137431 3049
rect 137373 3040 137385 3043
rect 135956 3012 137385 3040
rect 135956 3000 135962 3012
rect 137373 3009 137385 3012
rect 137419 3009 137431 3043
rect 137373 3003 137431 3009
rect 137922 3000 137928 3052
rect 137980 3040 137986 3052
rect 138661 3043 138719 3049
rect 137980 3012 138612 3040
rect 137980 3000 137986 3012
rect 60056 2944 64920 2972
rect 60056 2932 60062 2944
rect 67174 2932 67180 2984
rect 67232 2972 67238 2984
rect 92750 2972 92756 2984
rect 67232 2944 92756 2972
rect 67232 2932 67238 2944
rect 92750 2932 92756 2944
rect 92808 2932 92814 2984
rect 117222 2932 117228 2984
rect 117280 2972 117286 2984
rect 132586 2972 132592 2984
rect 117280 2944 132592 2972
rect 117280 2932 117286 2944
rect 132586 2932 132592 2944
rect 132644 2932 132650 2984
rect 133049 2975 133107 2981
rect 133049 2941 133061 2975
rect 133095 2972 133107 2975
rect 138474 2972 138480 2984
rect 133095 2944 138480 2972
rect 133095 2941 133107 2944
rect 133049 2935 133107 2941
rect 138474 2932 138480 2944
rect 138532 2932 138538 2984
rect 138584 2972 138612 3012
rect 138661 3009 138673 3043
rect 138707 3040 138719 3043
rect 143258 3040 143264 3052
rect 138707 3012 143264 3040
rect 138707 3009 138719 3012
rect 138661 3003 138719 3009
rect 143258 3000 143264 3012
rect 143316 3000 143322 3052
rect 148873 3043 148931 3049
rect 148873 3040 148885 3043
rect 146864 3012 148885 3040
rect 146864 2972 146892 3012
rect 148873 3009 148885 3012
rect 148919 3009 148931 3043
rect 148873 3003 148931 3009
rect 148965 3043 149023 3049
rect 148965 3009 148977 3043
rect 149011 3040 149023 3043
rect 152734 3040 152740 3052
rect 149011 3012 152740 3040
rect 149011 3009 149023 3012
rect 148965 3003 149023 3009
rect 152734 3000 152740 3012
rect 152792 3000 152798 3052
rect 153194 3000 153200 3052
rect 153252 3040 153258 3052
rect 187234 3040 187240 3052
rect 153252 3012 187240 3040
rect 153252 3000 153258 3012
rect 187234 3000 187240 3012
rect 187292 3000 187298 3052
rect 188982 3000 188988 3052
rect 189040 3040 189046 3052
rect 189721 3043 189779 3049
rect 189721 3040 189733 3043
rect 189040 3012 189733 3040
rect 189040 3000 189046 3012
rect 189721 3009 189733 3012
rect 189767 3009 189779 3043
rect 189721 3003 189779 3009
rect 249794 3000 249800 3052
rect 249852 3040 249858 3052
rect 321646 3040 321652 3052
rect 249852 3012 321652 3040
rect 249852 3000 249858 3012
rect 321646 3000 321652 3012
rect 321704 3000 321710 3052
rect 322198 3000 322204 3052
rect 322256 3040 322262 3052
rect 346670 3040 346676 3052
rect 322256 3012 346676 3040
rect 322256 3000 322262 3012
rect 346670 3000 346676 3012
rect 346728 3000 346734 3052
rect 347685 3043 347743 3049
rect 347685 3009 347697 3043
rect 347731 3040 347743 3043
rect 353754 3040 353760 3052
rect 347731 3012 353760 3040
rect 347731 3009 347743 3012
rect 347685 3003 347743 3009
rect 353754 3000 353760 3012
rect 353812 3000 353818 3052
rect 359476 3040 359504 3080
rect 425146 3068 425152 3080
rect 425204 3068 425210 3120
rect 353864 3012 359504 3040
rect 359553 3043 359611 3049
rect 138584 2944 146892 2972
rect 157242 2932 157248 2984
rect 157300 2972 157306 2984
rect 158625 2975 158683 2981
rect 158625 2972 158637 2975
rect 157300 2944 158637 2972
rect 157300 2932 157306 2944
rect 158625 2941 158637 2944
rect 158671 2941 158683 2975
rect 158625 2935 158683 2941
rect 158809 2975 158867 2981
rect 158809 2941 158821 2975
rect 158855 2972 158867 2975
rect 163498 2972 163504 2984
rect 158855 2944 163504 2972
rect 158855 2941 158867 2944
rect 158809 2935 158867 2941
rect 163498 2932 163504 2944
rect 163556 2932 163562 2984
rect 163590 2932 163596 2984
rect 163648 2972 163654 2984
rect 196802 2972 196808 2984
rect 163648 2944 196808 2972
rect 163648 2932 163654 2944
rect 196802 2932 196808 2944
rect 196860 2932 196866 2984
rect 242894 2932 242900 2984
rect 242952 2972 242958 2984
rect 307386 2972 307392 2984
rect 242952 2944 307392 2972
rect 242952 2932 242958 2944
rect 307386 2932 307392 2944
rect 307444 2932 307450 2984
rect 313918 2932 313924 2984
rect 313976 2972 313982 2984
rect 314749 2975 314807 2981
rect 313976 2944 314700 2972
rect 313976 2932 313982 2944
rect 52822 2864 52828 2916
rect 52880 2904 52886 2916
rect 69382 2904 69388 2916
rect 52880 2876 69388 2904
rect 52880 2864 52886 2876
rect 69382 2864 69388 2876
rect 69440 2864 69446 2916
rect 69474 2864 69480 2916
rect 69532 2904 69538 2916
rect 94225 2907 94283 2913
rect 94225 2904 94237 2907
rect 69532 2876 94237 2904
rect 69532 2864 69538 2876
rect 94225 2873 94237 2876
rect 94271 2873 94283 2907
rect 94225 2867 94283 2873
rect 119982 2864 119988 2916
rect 120040 2904 120046 2916
rect 140866 2904 140872 2916
rect 120040 2876 140872 2904
rect 120040 2864 120046 2876
rect 140866 2864 140872 2876
rect 140924 2864 140930 2916
rect 151722 2904 151728 2916
rect 149624 2876 151728 2904
rect 55217 2839 55275 2845
rect 55217 2805 55229 2839
rect 55263 2836 55275 2839
rect 64785 2839 64843 2845
rect 64785 2836 64797 2839
rect 55263 2808 64797 2836
rect 55263 2805 55275 2808
rect 55217 2799 55275 2805
rect 64785 2805 64797 2808
rect 64831 2805 64843 2839
rect 64785 2799 64843 2805
rect 65978 2796 65984 2848
rect 66036 2836 66042 2848
rect 68186 2836 68192 2848
rect 66036 2808 68192 2836
rect 66036 2796 66042 2808
rect 68186 2796 68192 2808
rect 68244 2796 68250 2848
rect 68278 2796 68284 2848
rect 68336 2836 68342 2848
rect 92566 2836 92572 2848
rect 68336 2808 92572 2836
rect 68336 2796 68342 2808
rect 92566 2796 92572 2808
rect 92624 2796 92630 2848
rect 116946 2796 116952 2848
rect 117004 2836 117010 2848
rect 133782 2836 133788 2848
rect 117004 2808 133788 2836
rect 117004 2796 117010 2808
rect 133782 2796 133788 2808
rect 133840 2796 133846 2848
rect 137278 2836 137284 2848
rect 133892 2808 137284 2836
rect 62301 2771 62359 2777
rect 62301 2737 62313 2771
rect 62347 2768 62359 2771
rect 64693 2771 64751 2777
rect 64693 2768 64705 2771
rect 62347 2740 64705 2768
rect 62347 2737 62359 2740
rect 62301 2731 62359 2737
rect 64693 2737 64705 2740
rect 64739 2737 64751 2771
rect 64693 2731 64751 2737
rect 132957 2771 133015 2777
rect 132957 2737 132969 2771
rect 133003 2768 133015 2771
rect 133892 2768 133920 2808
rect 137278 2796 137284 2808
rect 137336 2796 137342 2848
rect 137373 2839 137431 2845
rect 137373 2805 137385 2839
rect 137419 2836 137431 2839
rect 149624 2836 149652 2876
rect 151722 2864 151728 2876
rect 151780 2864 151786 2916
rect 151817 2907 151875 2913
rect 151817 2873 151829 2907
rect 151863 2904 151875 2907
rect 180150 2904 180156 2916
rect 151863 2876 180156 2904
rect 151863 2873 151875 2876
rect 151817 2867 151875 2873
rect 180150 2864 180156 2876
rect 180208 2864 180214 2916
rect 180245 2907 180303 2913
rect 180245 2873 180257 2907
rect 180291 2904 180303 2907
rect 314562 2904 314568 2916
rect 180291 2876 314568 2904
rect 180291 2873 180303 2876
rect 180245 2867 180303 2873
rect 314562 2864 314568 2876
rect 314620 2864 314626 2916
rect 314672 2904 314700 2944
rect 314749 2941 314761 2975
rect 314795 2972 314807 2975
rect 318058 2972 318064 2984
rect 314795 2944 318064 2972
rect 314795 2941 314807 2944
rect 314749 2935 314807 2941
rect 318058 2932 318064 2944
rect 318116 2932 318122 2984
rect 318150 2932 318156 2984
rect 318208 2972 318214 2984
rect 339494 2972 339500 2984
rect 318208 2944 339500 2972
rect 318208 2932 318214 2944
rect 339494 2932 339500 2944
rect 339552 2932 339558 2984
rect 345658 2932 345664 2984
rect 345716 2972 345722 2984
rect 348329 2975 348387 2981
rect 348329 2972 348341 2975
rect 345716 2944 348341 2972
rect 345716 2932 345722 2944
rect 348329 2941 348341 2944
rect 348375 2941 348387 2975
rect 348329 2935 348387 2941
rect 348418 2932 348424 2984
rect 348476 2972 348482 2984
rect 349157 2975 349215 2981
rect 349157 2972 349169 2975
rect 348476 2944 349169 2972
rect 348476 2932 348482 2944
rect 349157 2941 349169 2944
rect 349203 2941 349215 2975
rect 349157 2935 349215 2941
rect 349798 2932 349804 2984
rect 349856 2972 349862 2984
rect 353864 2972 353892 3012
rect 359553 3009 359565 3043
rect 359599 3040 359611 3043
rect 417970 3040 417976 3052
rect 359599 3012 417976 3040
rect 359599 3009 359611 3012
rect 359553 3003 359611 3009
rect 417970 3000 417976 3012
rect 418028 3000 418034 3052
rect 410886 2972 410892 2984
rect 349856 2944 353892 2972
rect 353956 2944 410892 2972
rect 349856 2932 349862 2944
rect 332410 2904 332416 2916
rect 314672 2876 332416 2904
rect 332410 2864 332416 2876
rect 332468 2864 332474 2916
rect 342898 2864 342904 2916
rect 342956 2904 342962 2916
rect 342956 2876 343220 2904
rect 342956 2864 342962 2876
rect 137419 2808 149652 2836
rect 137419 2805 137431 2808
rect 137373 2799 137431 2805
rect 149698 2796 149704 2848
rect 149756 2836 149762 2848
rect 153933 2839 153991 2845
rect 153933 2836 153945 2839
rect 149756 2808 153945 2836
rect 149756 2796 149762 2808
rect 153933 2805 153945 2808
rect 153979 2805 153991 2839
rect 153933 2799 153991 2805
rect 155236 2808 156552 2836
rect 133003 2740 133920 2768
rect 154025 2771 154083 2777
rect 133003 2737 133015 2740
rect 132957 2731 133015 2737
rect 154025 2737 154037 2771
rect 154071 2768 154083 2771
rect 155236 2768 155264 2808
rect 154071 2740 155264 2768
rect 156524 2768 156552 2808
rect 160738 2796 160744 2848
rect 160796 2836 160802 2848
rect 163590 2836 163596 2848
rect 160796 2808 163596 2836
rect 160796 2796 160802 2808
rect 163590 2796 163596 2808
rect 163648 2796 163654 2848
rect 163685 2839 163743 2845
rect 163685 2805 163697 2839
rect 163731 2836 163743 2839
rect 189626 2836 189632 2848
rect 163731 2808 189632 2836
rect 163731 2805 163743 2808
rect 163685 2799 163743 2805
rect 189626 2796 189632 2808
rect 189684 2796 189690 2848
rect 189721 2839 189779 2845
rect 189721 2805 189733 2839
rect 189767 2836 189779 2839
rect 343082 2836 343088 2848
rect 189767 2808 343088 2836
rect 189767 2805 189779 2808
rect 189721 2799 189779 2805
rect 343082 2796 343088 2808
rect 343140 2796 343146 2848
rect 343192 2836 343220 2876
rect 347038 2864 347044 2916
rect 347096 2904 347102 2916
rect 353956 2904 353984 2944
rect 410886 2932 410892 2944
rect 410944 2932 410950 2984
rect 347096 2876 353984 2904
rect 354033 2907 354091 2913
rect 347096 2864 347102 2876
rect 354033 2873 354045 2907
rect 354079 2904 354091 2907
rect 403710 2904 403716 2916
rect 354079 2876 403716 2904
rect 354079 2873 354091 2876
rect 354033 2867 354091 2873
rect 403710 2864 403716 2876
rect 403768 2864 403774 2916
rect 389450 2836 389456 2848
rect 343192 2808 389456 2836
rect 389450 2796 389456 2808
rect 389508 2796 389514 2848
rect 158809 2771 158867 2777
rect 158809 2768 158821 2771
rect 156524 2740 158821 2768
rect 154071 2737 154083 2740
rect 154025 2731 154083 2737
rect 158809 2737 158821 2740
rect 158855 2737 158867 2771
rect 158809 2731 158867 2737
rect 348329 2771 348387 2777
rect 348329 2737 348341 2771
rect 348375 2768 348387 2771
rect 350353 2771 350411 2777
rect 350353 2768 350365 2771
rect 348375 2740 350365 2768
rect 348375 2737 348387 2740
rect 348329 2731 348387 2737
rect 350353 2737 350365 2740
rect 350399 2737 350411 2771
rect 350353 2731 350411 2737
rect 61105 2703 61163 2709
rect 61105 2669 61117 2703
rect 61151 2700 61163 2703
rect 64601 2703 64659 2709
rect 64601 2700 64613 2703
rect 61151 2672 64613 2700
rect 61151 2669 61163 2672
rect 61105 2663 61163 2669
rect 64601 2669 64613 2672
rect 64647 2669 64659 2703
rect 64601 2663 64659 2669
rect 70670 960 70676 1012
rect 70728 1000 70734 1012
rect 73709 1003 73767 1009
rect 73709 1000 73721 1003
rect 70728 972 73721 1000
rect 70728 960 70734 972
rect 73709 969 73721 972
rect 73755 969 73767 1003
rect 73709 963 73767 969
rect 146570 552 146576 604
rect 146628 592 146634 604
rect 146846 592 146852 604
rect 146628 564 146852 592
rect 146628 552 146634 564
rect 146846 552 146852 564
rect 146904 552 146910 604
rect 271874 552 271880 604
rect 271932 592 271938 604
rect 272886 592 272892 604
rect 271932 564 272892 592
rect 271932 552 271938 564
rect 272886 552 272892 564
rect 272944 552 272950 604
rect 274634 552 274640 604
rect 274692 592 274698 604
rect 275278 592 275284 604
rect 274692 564 275284 592
rect 274692 552 274698 564
rect 275278 552 275284 564
rect 275336 552 275342 604
rect 277394 552 277400 604
rect 277452 592 277458 604
rect 277670 592 277676 604
rect 277452 564 277676 592
rect 277452 552 277458 564
rect 277670 552 277676 564
rect 277728 552 277734 604
rect 280154 552 280160 604
rect 280212 592 280218 604
rect 281258 592 281264 604
rect 280212 564 281264 592
rect 280212 552 280218 564
rect 281258 552 281264 564
rect 281316 552 281322 604
rect 281534 552 281540 604
rect 281592 592 281598 604
rect 282454 592 282460 604
rect 281592 564 282460 592
rect 281592 552 281598 564
rect 282454 552 282460 564
rect 282512 552 282518 604
rect 282914 552 282920 604
rect 282972 592 282978 604
rect 283650 592 283656 604
rect 282972 564 283656 592
rect 282972 552 282978 564
rect 283650 552 283656 564
rect 283708 552 283714 604
rect 285674 552 285680 604
rect 285732 592 285738 604
rect 285950 592 285956 604
rect 285732 564 285956 592
rect 285732 552 285738 564
rect 285950 552 285956 564
rect 286008 552 286014 604
rect 288434 552 288440 604
rect 288492 592 288498 604
rect 289538 592 289544 604
rect 288492 564 289544 592
rect 288492 552 288498 564
rect 289538 552 289544 564
rect 289596 552 289602 604
rect 291194 552 291200 604
rect 291252 592 291258 604
rect 291930 592 291936 604
rect 291252 564 291936 592
rect 291252 552 291258 564
rect 291930 552 291936 564
rect 291988 552 291994 604
rect 292574 552 292580 604
rect 292632 592 292638 604
rect 293126 592 293132 604
rect 292632 564 293132 592
rect 292632 552 292638 564
rect 293126 552 293132 564
rect 293184 552 293190 604
rect 295334 552 295340 604
rect 295392 592 295398 604
rect 295518 592 295524 604
rect 295392 564 295524 592
rect 295392 552 295398 564
rect 295518 552 295524 564
rect 295576 552 295582 604
rect 298094 552 298100 604
rect 298152 592 298158 604
rect 299106 592 299112 604
rect 298152 564 299112 592
rect 298152 552 298158 564
rect 299106 552 299112 564
rect 299164 552 299170 604
rect 303614 552 303620 604
rect 303672 592 303678 604
rect 303798 592 303804 604
rect 303672 564 303804 592
rect 303672 552 303678 564
rect 303798 552 303804 564
rect 303856 552 303862 604
rect 309134 552 309140 604
rect 309192 592 309198 604
rect 309778 592 309784 604
rect 309192 564 309784 592
rect 309192 552 309198 564
rect 309778 552 309784 564
rect 309836 552 309842 604
rect 316034 552 316040 604
rect 316092 592 316098 604
rect 316954 592 316960 604
rect 316092 564 316960 592
rect 316092 552 316098 564
rect 316954 552 316960 564
rect 317012 552 317018 604
rect 322934 552 322940 604
rect 322992 592 322998 604
rect 324038 592 324044 604
rect 322992 564 324044 592
rect 322992 552 322998 564
rect 324038 552 324044 564
rect 324096 552 324102 604
rect 327074 552 327080 604
rect 327132 592 327138 604
rect 327626 592 327632 604
rect 327132 564 327632 592
rect 327132 552 327138 564
rect 327626 552 327632 564
rect 327684 552 327690 604
rect 333974 552 333980 604
rect 334032 592 334038 604
rect 334710 592 334716 604
rect 334032 564 334716 592
rect 334032 552 334038 564
rect 334710 552 334716 564
rect 334768 552 334774 604
rect 340874 552 340880 604
rect 340932 592 340938 604
rect 341886 592 341892 604
rect 340932 564 341892 592
rect 340932 552 340938 564
rect 341886 552 341892 564
rect 341944 552 341950 604
rect 351914 552 351920 604
rect 351972 592 351978 604
rect 352558 592 352564 604
rect 351972 564 352564 592
rect 351972 552 351978 564
rect 352558 552 352564 564
rect 352616 552 352622 604
rect 358814 552 358820 604
rect 358872 592 358878 604
rect 359734 592 359740 604
rect 358872 564 359740 592
rect 358872 552 358878 564
rect 359734 552 359740 564
rect 359792 552 359798 604
rect 369854 552 369860 604
rect 369912 592 369918 604
rect 370406 592 370412 604
rect 369912 564 370412 592
rect 369912 552 369918 564
rect 370406 552 370412 564
rect 370464 552 370470 604
rect 375374 552 375380 604
rect 375432 592 375438 604
rect 376386 592 376392 604
rect 375432 564 376392 592
rect 375432 552 375438 564
rect 376386 552 376392 564
rect 376444 552 376450 604
rect 376754 552 376760 604
rect 376812 592 376818 604
rect 377582 592 377588 604
rect 376812 564 377588 592
rect 376812 552 376818 564
rect 377582 552 377588 564
rect 377640 552 377646 604
rect 379514 552 379520 604
rect 379572 592 379578 604
rect 379974 592 379980 604
rect 379572 564 379980 592
rect 379572 552 379578 564
rect 379974 552 379980 564
rect 380032 552 380038 604
rect 394694 552 394700 604
rect 394752 592 394758 604
rect 395430 592 395436 604
rect 394752 564 395436 592
rect 394752 552 394758 564
rect 395430 552 395436 564
rect 395488 552 395494 604
rect 401594 552 401600 604
rect 401652 592 401658 604
rect 402514 592 402520 604
rect 401652 564 402520 592
rect 401652 552 401658 564
rect 402514 552 402520 564
rect 402572 552 402578 604
rect 405734 552 405740 604
rect 405792 592 405798 604
rect 406102 592 406108 604
rect 405792 564 406108 592
rect 405792 552 405798 564
rect 406102 552 406108 564
rect 406160 552 406166 604
rect 412634 552 412640 604
rect 412692 592 412698 604
rect 413278 592 413284 604
rect 412692 564 413284 592
rect 412692 552 412698 564
rect 413278 552 413284 564
rect 413336 552 413342 604
rect 419534 552 419540 604
rect 419592 592 419598 604
rect 420362 592 420368 604
rect 419592 564 420368 592
rect 419592 552 419598 564
rect 420362 552 420368 564
rect 420420 552 420426 604
rect 420914 552 420920 604
rect 420972 592 420978 604
rect 421558 592 421564 604
rect 420972 564 421564 592
rect 420972 552 420978 564
rect 421558 552 421564 564
rect 421616 552 421622 604
rect 423674 552 423680 604
rect 423732 592 423738 604
rect 423950 592 423956 604
rect 423732 564 423956 592
rect 423732 552 423738 564
rect 423950 552 423956 564
rect 424008 552 424014 604
rect 426434 552 426440 604
rect 426492 592 426498 604
rect 427538 592 427544 604
rect 426492 564 427544 592
rect 426492 552 426498 564
rect 427538 552 427544 564
rect 427596 552 427602 604
rect 430574 552 430580 604
rect 430632 592 430638 604
rect 431126 592 431132 604
rect 430632 564 431132 592
rect 430632 552 430638 564
rect 431126 552 431132 564
rect 431184 552 431190 604
rect 437474 552 437480 604
rect 437532 592 437538 604
rect 438210 592 438216 604
rect 437532 564 438216 592
rect 437532 552 437538 564
rect 438210 552 438216 564
rect 438268 552 438274 604
rect 455414 552 455420 604
rect 455472 592 455478 604
rect 456058 592 456064 604
rect 455472 564 456064 592
rect 455472 552 455478 564
rect 456058 552 456064 564
rect 456116 552 456122 604
rect 462314 552 462320 604
rect 462372 592 462378 604
rect 463234 592 463240 604
rect 462372 564 463240 592
rect 462372 552 462378 564
rect 463234 552 463240 564
rect 463292 552 463298 604
rect 466454 552 466460 604
rect 466512 592 466518 604
rect 466822 592 466828 604
rect 466512 564 466828 592
rect 466512 552 466518 564
rect 466822 552 466828 564
rect 466880 552 466886 604
rect 469214 552 469220 604
rect 469272 592 469278 604
rect 470318 592 470324 604
rect 469272 564 470324 592
rect 469272 552 469278 564
rect 470318 552 470324 564
rect 470376 552 470382 604
rect 478874 552 478880 604
rect 478932 592 478938 604
rect 479886 592 479892 604
rect 478932 564 479892 592
rect 478932 552 478938 564
rect 479886 552 479892 564
rect 479944 552 479950 604
rect 489914 552 489920 604
rect 489972 592 489978 604
rect 490558 592 490564 604
rect 489972 564 490564 592
rect 489972 552 489978 564
rect 490558 552 490564 564
rect 490616 552 490622 604
rect 495434 552 495440 604
rect 495492 592 495498 604
rect 496538 592 496544 604
rect 495492 564 496544 592
rect 495492 552 495498 564
rect 496538 552 496544 564
rect 496596 552 496602 604
rect 499574 552 499580 604
rect 499632 592 499638 604
rect 500126 592 500132 604
rect 499632 564 500132 592
rect 499632 552 499638 564
rect 500126 552 500132 564
rect 500184 552 500190 604
rect 506474 552 506480 604
rect 506532 592 506538 604
rect 507210 592 507216 604
rect 506532 564 507216 592
rect 506532 552 506538 564
rect 507210 552 507216 564
rect 507268 552 507274 604
rect 510614 552 510620 604
rect 510672 592 510678 604
rect 510798 592 510804 604
rect 510672 564 510804 592
rect 510672 552 510678 564
rect 510798 552 510804 564
rect 510856 552 510862 604
rect 513374 552 513380 604
rect 513432 592 513438 604
rect 514386 592 514392 604
rect 513432 564 514392 592
rect 513432 552 513438 564
rect 514386 552 514392 564
rect 514444 552 514450 604
rect 524414 552 524420 604
rect 524472 592 524478 604
rect 525058 592 525064 604
rect 524472 564 525064 592
rect 524472 552 524478 564
rect 525058 552 525064 564
rect 525116 552 525122 604
rect 531314 552 531320 604
rect 531372 592 531378 604
rect 532234 592 532240 604
rect 531372 564 532240 592
rect 531372 552 531378 564
rect 532234 552 532240 564
rect 532292 552 532298 604
rect 538214 552 538220 604
rect 538272 592 538278 604
rect 539318 592 539324 604
rect 538272 564 539324 592
rect 538272 552 538278 564
rect 539318 552 539324 564
rect 539376 552 539382 604
rect 542354 552 542360 604
rect 542412 592 542418 604
rect 542906 592 542912 604
rect 542412 564 542912 592
rect 542412 552 542418 564
rect 542906 552 542912 564
rect 542964 552 542970 604
rect 549254 552 549260 604
rect 549312 592 549318 604
rect 550082 592 550088 604
rect 549312 564 550088 592
rect 549312 552 549318 564
rect 550082 552 550088 564
rect 550140 552 550146 604
rect 556154 552 556160 604
rect 556212 592 556218 604
rect 557166 592 557172 604
rect 556212 564 557172 592
rect 556212 552 556218 564
rect 557166 552 557172 564
rect 557224 552 557230 604
rect 576854 552 576860 604
rect 576912 592 576918 604
rect 577406 592 577412 604
rect 576912 564 577412 592
rect 576912 552 576918 564
rect 577406 552 577412 564
rect 577464 552 577470 604
<< via1 >>
rect 156604 655528 156656 655580
rect 187700 655528 187752 655580
rect 95148 568488 95200 568540
rect 103152 568488 103204 568540
rect 119436 568488 119488 568540
rect 128452 568488 128504 568540
rect 132408 568488 132460 568540
rect 209596 568488 209648 568540
rect 110328 568420 110380 568472
rect 135904 568420 135956 568472
rect 117964 568352 118016 568404
rect 137284 568352 137336 568404
rect 98368 568284 98420 568336
rect 107752 568284 107804 568336
rect 117136 568284 117188 568336
rect 121000 568284 121052 568336
rect 140044 568284 140096 568336
rect 217140 568284 217192 568336
rect 225880 568284 225932 568336
rect 234620 568284 234672 568336
rect 100668 568216 100720 568268
rect 109040 568216 109092 568268
rect 97908 568148 97960 568200
rect 106648 568148 106700 568200
rect 115848 568148 115900 568200
rect 93768 568080 93820 568132
rect 101772 568080 101824 568132
rect 110696 568080 110748 568132
rect 103152 568012 103204 568064
rect 112260 568012 112312 568064
rect 96528 567944 96580 567996
rect 105268 567944 105320 567996
rect 114744 567944 114796 567996
rect 124312 568216 124364 568268
rect 117136 568148 117188 568200
rect 126612 568216 126664 568268
rect 144920 568216 144972 568268
rect 215576 568216 215628 568268
rect 224776 568216 224828 568268
rect 233240 568216 233292 568268
rect 128452 568148 128504 568200
rect 149060 568148 149112 568200
rect 209596 568148 209648 568200
rect 218980 568148 219032 568200
rect 228364 568148 228416 568200
rect 237380 568148 237432 568200
rect 102048 567876 102100 567928
rect 109868 567876 109920 567928
rect 94872 567808 94924 567860
rect 104072 567808 104124 567860
rect 113640 567808 113692 567860
rect 123484 568080 123536 568132
rect 124128 568080 124180 568132
rect 146944 568080 146996 568132
rect 217876 568080 217928 568132
rect 227168 568080 227220 568132
rect 236000 568080 236052 568132
rect 120080 568012 120132 568064
rect 144184 568012 144236 568064
rect 202236 568012 202288 568064
rect 211896 568012 211948 568064
rect 221464 568012 221516 568064
rect 230480 568012 230532 568064
rect 119252 567944 119304 567996
rect 142896 567944 142948 567996
rect 203708 567944 203760 567996
rect 213092 567944 213144 567996
rect 222384 567944 222436 567996
rect 231860 567944 231912 567996
rect 125508 567876 125560 567928
rect 152464 567876 152516 567928
rect 204812 567876 204864 567928
rect 214104 567876 214156 567928
rect 223672 567876 223724 567928
rect 231952 567876 232004 567928
rect 118056 567808 118108 567860
rect 142804 567808 142856 567860
rect 208308 567808 208360 567860
rect 217140 567808 217192 567860
rect 220084 567808 220136 567860
rect 229376 567808 229428 567860
rect 238760 567808 238812 567860
rect 102968 567740 103020 567792
rect 156696 567740 156748 567792
rect 85488 567672 85540 567724
rect 91100 567672 91152 567724
rect 100668 567672 100720 567724
rect 156788 567672 156840 567724
rect 97908 567604 97960 567656
rect 155224 567604 155276 567656
rect 95148 567536 95200 567588
rect 153844 567536 153896 567588
rect 194416 567536 194468 567588
rect 252192 567536 252244 567588
rect 110328 567468 110380 567520
rect 138664 567468 138716 567520
rect 124864 567400 124916 567452
rect 81348 567332 81400 567384
rect 88340 567332 88392 567384
rect 120632 567332 120684 567384
rect 127624 567400 127676 567452
rect 128268 567400 128320 567452
rect 207020 567400 207072 567452
rect 208308 567400 208360 567452
rect 82728 567264 82780 567316
rect 89996 567264 90048 567316
rect 118332 567264 118384 567316
rect 125416 567332 125468 567384
rect 204812 567332 204864 567384
rect 209044 567332 209096 567384
rect 217876 567332 217928 567384
rect 121276 567264 121328 567316
rect 202236 567264 202288 567316
rect 210424 567264 210476 567316
rect 220084 567264 220136 567316
rect 78128 567196 78180 567248
rect 86960 567196 87012 567248
rect 110696 567196 110748 567248
rect 120724 567196 120776 567248
rect 122656 567196 122708 567248
rect 203708 567196 203760 567248
rect 206284 567196 206336 567248
rect 215576 567196 215628 567248
rect 252560 557540 252612 557592
rect 257988 557472 258040 557524
rect 258080 551624 258132 551676
rect 259736 551624 259788 551676
rect 259736 549176 259788 549228
rect 261484 549176 261536 549228
rect 261484 540948 261536 541000
rect 263600 540880 263652 540932
rect 263600 538840 263652 538892
rect 272064 538840 272116 538892
rect 272064 534556 272116 534608
rect 273904 534556 273956 534608
rect 111708 525716 111760 525768
rect 181444 525716 181496 525768
rect 119988 525648 120040 525700
rect 194784 525648 194836 525700
rect 128176 525580 128228 525632
rect 208124 525580 208176 525632
rect 101404 525512 101456 525564
rect 188344 525512 188396 525564
rect 99472 525444 99524 525496
rect 188436 525444 188488 525496
rect 97632 525376 97684 525428
rect 188528 525376 188580 525428
rect 95700 525308 95752 525360
rect 188620 525308 188672 525360
rect 93768 525240 93820 525292
rect 188712 525240 188764 525292
rect 91836 525172 91888 525224
rect 188804 525172 188856 525224
rect 86132 525104 86184 525156
rect 188896 525104 188948 525156
rect 89996 525036 90048 525088
rect 195980 525036 196032 525088
rect 108948 524968 109000 525020
rect 175740 524968 175792 525020
rect 107568 524900 107620 524952
rect 173808 524900 173860 524952
rect 104808 524832 104860 524884
rect 170036 524832 170088 524884
rect 106188 524764 106240 524816
rect 171968 524764 172020 524816
rect 93676 524696 93728 524748
rect 150992 524696 151044 524748
rect 74724 524356 74776 524408
rect 75828 524356 75880 524408
rect 80428 524356 80480 524408
rect 81348 524356 81400 524408
rect 84292 524356 84344 524408
rect 85488 524356 85540 524408
rect 95056 524356 95108 524408
rect 152832 524356 152884 524408
rect 153844 524356 153896 524408
rect 154764 524356 154816 524408
rect 155224 524356 155276 524408
rect 158536 524356 158588 524408
rect 99196 524288 99248 524340
rect 96436 524220 96488 524272
rect 156420 524288 156472 524340
rect 156696 524288 156748 524340
rect 156788 524220 156840 524272
rect 162400 524356 162452 524408
rect 208308 524356 208360 524408
rect 219532 524356 219584 524408
rect 229008 524356 229060 524408
rect 253848 524356 253900 524408
rect 166172 524288 166224 524340
rect 211068 524288 211120 524340
rect 223396 524288 223448 524340
rect 227628 524288 227680 524340
rect 252008 524288 252060 524340
rect 209688 524220 209740 524272
rect 221464 524220 221516 524272
rect 231768 524220 231820 524272
rect 257712 524220 257764 524272
rect 101956 524152 102008 524204
rect 164332 524152 164384 524204
rect 212448 524152 212500 524204
rect 227168 524152 227220 524204
rect 230388 524152 230440 524204
rect 255780 524152 255832 524204
rect 78864 524084 78916 524136
rect 88064 524084 88116 524136
rect 103336 524084 103388 524136
rect 168104 524084 168156 524136
rect 225328 524084 225380 524136
rect 233148 524084 233200 524136
rect 259552 524084 259604 524136
rect 78772 524016 78824 524068
rect 78680 523948 78732 524000
rect 120448 524016 120500 524068
rect 121276 524016 121328 524068
rect 185308 524016 185360 524068
rect 204168 524016 204220 524068
rect 213828 524016 213880 524068
rect 213920 524016 213972 524068
rect 229100 524016 229152 524068
rect 234528 524016 234580 524068
rect 263416 524016 263468 524068
rect 78312 523880 78364 523932
rect 109040 523948 109092 524000
rect 118516 523948 118568 524000
rect 191012 523948 191064 524000
rect 205548 523948 205600 524000
rect 215760 523948 215812 524000
rect 216588 523948 216640 524000
rect 232872 523948 232924 524000
rect 235908 523948 235960 524000
rect 261484 523948 261536 524000
rect 110972 523880 111024 523932
rect 114468 523880 114520 523932
rect 122748 523880 122800 523932
rect 198648 523880 198700 523932
rect 202788 523880 202840 523932
rect 211988 523880 212040 523932
rect 215208 523880 215260 523932
rect 231032 523880 231084 523932
rect 233056 523880 233108 523932
rect 78404 523812 78456 523864
rect 114744 523812 114796 523864
rect 124312 523812 124364 523864
rect 125416 523812 125468 523864
rect 133788 523812 133840 523864
rect 210424 523812 210476 523864
rect 210976 523812 211028 523864
rect 217968 523812 218020 523864
rect 234804 523812 234856 523864
rect 237288 523880 237340 523932
rect 267188 523880 267240 523932
rect 78496 523744 78548 523796
rect 116676 523744 116728 523796
rect 130016 523744 130068 523796
rect 209044 523744 209096 523796
rect 219348 523744 219400 523796
rect 238300 523744 238352 523796
rect 78588 523676 78640 523728
rect 118516 523676 118568 523728
rect 126152 523676 126204 523728
rect 206284 523676 206336 523728
rect 206928 523676 206980 523728
rect 217692 523676 217744 523728
rect 217876 523676 217928 523728
rect 236736 523676 236788 523728
rect 238668 523812 238720 523864
rect 240048 523812 240100 523864
rect 265348 523812 265400 523864
rect 269120 523744 269172 523796
rect 273904 523744 273956 523796
rect 275376 523744 275428 523796
rect 271052 523676 271104 523728
rect 78220 523608 78272 523660
rect 107108 523608 107160 523660
rect 123484 523608 123536 523660
rect 139492 523608 139544 523660
rect 140044 523608 140096 523660
rect 196716 523608 196768 523660
rect 226248 523608 226300 523660
rect 250076 523608 250128 523660
rect 103336 523540 103388 523592
rect 155960 523540 156012 523592
rect 160468 523540 160520 523592
rect 226156 523540 226208 523592
rect 248144 523540 248196 523592
rect 86776 523472 86828 523524
rect 105176 523472 105228 523524
rect 112812 523472 112864 523524
rect 127624 523472 127676 523524
rect 147128 523472 147180 523524
rect 124864 523404 124916 523456
rect 143356 523404 143408 523456
rect 146944 523404 146996 523456
rect 200488 523472 200540 523524
rect 223488 523472 223540 523524
rect 244372 523472 244424 523524
rect 125048 523336 125100 523388
rect 141424 523336 141476 523388
rect 144184 523336 144236 523388
rect 192852 523404 192904 523456
rect 224868 523404 224920 523456
rect 246212 523404 246264 523456
rect 189080 523336 189132 523388
rect 222108 523336 222160 523388
rect 242440 523336 242492 523388
rect 120724 523268 120776 523320
rect 135720 523268 135772 523320
rect 137284 523268 137336 523320
rect 183376 523268 183428 523320
rect 220728 523268 220780 523320
rect 240508 523268 240560 523320
rect 122104 523200 122156 523252
rect 137652 523200 137704 523252
rect 142896 523200 142948 523252
rect 187148 523200 187200 523252
rect 135904 523132 135956 523184
rect 177672 523132 177724 523184
rect 138664 523064 138716 523116
rect 179512 523064 179564 523116
rect 142804 522996 142856 523048
rect 275376 518984 275428 519036
rect 278780 518984 278832 519036
rect 274272 518916 274324 518968
rect 301504 518916 301556 518968
rect 278780 517012 278832 517064
rect 280068 517012 280120 517064
rect 280068 516808 280120 516860
rect 320180 516808 320232 516860
rect 273904 516740 273956 516792
rect 337752 516740 337804 516792
rect 338396 516740 338448 516792
rect 340880 516740 340932 516792
rect 275376 516672 275428 516724
rect 398840 516672 398892 516724
rect 275468 516604 275520 516656
rect 400220 516604 400272 516656
rect 274364 516536 274416 516588
rect 401600 516536 401652 516588
rect 274456 516468 274508 516520
rect 403348 516468 403400 516520
rect 274548 516400 274600 516452
rect 404360 516400 404412 516452
rect 406016 516400 406068 516452
rect 273812 516332 273864 516384
rect 273628 514768 273680 514820
rect 298744 514768 298796 514820
rect 275284 511980 275336 512032
rect 320180 511980 320232 512032
rect 273536 510620 273588 510672
rect 297364 510620 297416 510672
rect 279424 509260 279476 509312
rect 320364 509260 320416 509312
rect 302884 507832 302936 507884
rect 320180 507832 320232 507884
rect 273720 506540 273772 506592
rect 294604 506540 294656 506592
rect 275560 506472 275612 506524
rect 319812 506472 319864 506524
rect 273536 505180 273588 505232
rect 291844 505180 291896 505232
rect 275652 505112 275704 505164
rect 320180 505112 320232 505164
rect 276664 503684 276716 503736
rect 319996 503684 320048 503736
rect 320272 502528 320324 502580
rect 276756 502460 276808 502512
rect 273628 501032 273680 501084
rect 290464 501032 290516 501084
rect 276848 500964 276900 501016
rect 319812 500964 319864 501016
rect 273720 499604 273772 499656
rect 287704 499604 287756 499656
rect 276940 499536 276992 499588
rect 320180 499536 320232 499588
rect 277032 498176 277084 498228
rect 319812 498176 319864 498228
rect 273720 496884 273772 496936
rect 286324 496884 286376 496936
rect 278596 496816 278648 496868
rect 320180 496816 320232 496868
rect 273720 495592 273772 495644
rect 284944 495592 284996 495644
rect 279516 495524 279568 495576
rect 319812 495524 319864 495576
rect 275744 495456 275796 495508
rect 319996 495456 320048 495508
rect 320640 495499 320692 495508
rect 320640 495465 320649 495499
rect 320649 495465 320683 495499
rect 320683 495465 320692 495499
rect 320640 495456 320692 495465
rect 273628 494096 273680 494148
rect 278044 494096 278096 494148
rect 275836 494028 275888 494080
rect 319812 494028 319864 494080
rect 275928 492668 275980 492720
rect 320180 492668 320232 492720
rect 320732 492328 320784 492380
rect 320824 492328 320876 492380
rect 320732 492124 320784 492176
rect 320824 492124 320876 492176
rect 273628 491376 273680 491428
rect 283564 491376 283616 491428
rect 275192 491308 275244 491360
rect 319812 491308 319864 491360
rect 320640 490943 320692 490952
rect 320640 490909 320649 490943
rect 320649 490909 320683 490943
rect 320683 490909 320692 490943
rect 320640 490900 320692 490909
rect 273444 489948 273496 490000
rect 280804 489948 280856 490000
rect 275100 489880 275152 489932
rect 320180 489880 320232 489932
rect 320640 489923 320692 489932
rect 320640 489889 320649 489923
rect 320649 489889 320683 489923
rect 320683 489889 320692 489923
rect 320640 489880 320692 489889
rect 320088 489812 320140 489864
rect 320732 489812 320784 489864
rect 320824 489855 320876 489864
rect 320824 489821 320833 489855
rect 320833 489821 320867 489855
rect 320867 489821 320876 489855
rect 320824 489812 320876 489821
rect 320824 489404 320876 489456
rect 273628 488656 273680 488708
rect 278136 488656 278188 488708
rect 275008 488588 275060 488640
rect 319812 488588 319864 488640
rect 274916 488520 274968 488572
rect 319720 488520 319772 488572
rect 320456 487228 320508 487280
rect 274824 487160 274876 487212
rect 320180 487160 320232 487212
rect 320548 486208 320600 486260
rect 320640 486208 320692 486260
rect 320548 486004 320600 486056
rect 320640 486004 320692 486056
rect 273536 485868 273588 485920
rect 278228 485868 278280 485920
rect 274732 485800 274784 485852
rect 319812 485800 319864 485852
rect 273628 484440 273680 484492
rect 278320 484440 278372 484492
rect 274640 484372 274692 484424
rect 320180 484372 320232 484424
rect 277216 483012 277268 483064
rect 319812 483012 319864 483064
rect 320456 482851 320508 482860
rect 320456 482817 320465 482851
rect 320465 482817 320499 482851
rect 320499 482817 320508 482851
rect 320456 482808 320508 482817
rect 320456 482672 320508 482724
rect 320640 482672 320692 482724
rect 320824 482672 320876 482724
rect 320548 482332 320600 482384
rect 273628 481720 273680 481772
rect 278412 481720 278464 481772
rect 277308 481652 277360 481704
rect 320180 481652 320232 481704
rect 320272 480428 320324 480480
rect 320824 480428 320876 480480
rect 273628 480292 273680 480344
rect 278504 480292 278556 480344
rect 320272 480292 320324 480344
rect 276572 480224 276624 480276
rect 319812 480224 319864 480276
rect 320824 479451 320876 479460
rect 320824 479417 320833 479451
rect 320833 479417 320867 479451
rect 320867 479417 320876 479451
rect 320824 479408 320876 479417
rect 320180 479272 320232 479324
rect 320824 479272 320876 479324
rect 320640 478932 320692 478984
rect 273628 478864 273680 478916
rect 315304 478864 315356 478916
rect 320456 476960 320508 477012
rect 320640 476960 320692 477012
rect 320180 476824 320232 476876
rect 320272 476620 320324 476672
rect 273628 476076 273680 476128
rect 312544 476076 312596 476128
rect 320732 476051 320784 476060
rect 320732 476017 320741 476051
rect 320741 476017 320775 476051
rect 320775 476017 320784 476051
rect 320732 476008 320784 476017
rect 320640 475872 320692 475924
rect 320456 475804 320508 475856
rect 320824 475779 320876 475788
rect 320824 475745 320833 475779
rect 320833 475745 320867 475779
rect 320867 475745 320876 475779
rect 320824 475736 320876 475745
rect 273628 474784 273680 474836
rect 309784 474784 309836 474836
rect 276480 474716 276532 474768
rect 320180 474716 320232 474768
rect 273536 473968 273588 474020
rect 320364 473968 320416 474020
rect 273628 473356 273680 473408
rect 308404 473356 308456 473408
rect 273444 471996 273496 472048
rect 320180 471996 320232 472048
rect 273536 470636 273588 470688
rect 305644 470636 305696 470688
rect 273352 470568 273404 470620
rect 320272 470568 320324 470620
rect 320272 470432 320324 470484
rect 273536 469276 273588 469328
rect 304264 469276 304316 469328
rect 276388 469208 276440 469260
rect 320364 469208 320416 469260
rect 276296 467916 276348 467968
rect 320456 467916 320508 467968
rect 276204 467848 276256 467900
rect 320272 467848 320324 467900
rect 320548 467780 320600 467832
rect 320272 467712 320324 467764
rect 320732 467712 320784 467764
rect 320088 467644 320140 467696
rect 320548 467644 320600 467696
rect 320364 467619 320416 467628
rect 320364 467585 320373 467619
rect 320373 467585 320407 467619
rect 320407 467585 320416 467619
rect 320364 467576 320416 467585
rect 320640 467508 320692 467560
rect 320732 467372 320784 467424
rect 273536 466488 273588 466540
rect 302976 466488 303028 466540
rect 276112 466420 276164 466472
rect 320180 466420 320232 466472
rect 276020 465060 276072 465112
rect 320180 465060 320232 465112
rect 273260 463700 273312 463752
rect 277124 463700 277176 463752
rect 273260 460912 273312 460964
rect 278688 460912 278740 460964
rect 273260 460028 273312 460080
rect 276020 460028 276072 460080
rect 273260 458124 273312 458176
rect 276112 458124 276164 458176
rect 320456 457444 320508 457496
rect 320640 457444 320692 457496
rect 320824 457308 320876 457360
rect 320180 457104 320232 457156
rect 320364 456943 320416 456952
rect 320364 456909 320373 456943
rect 320373 456909 320407 456943
rect 320407 456909 320416 456943
rect 320364 456900 320416 456909
rect 320732 456900 320784 456952
rect 320364 456671 320416 456680
rect 320364 456637 320373 456671
rect 320373 456637 320407 456671
rect 320407 456637 320416 456671
rect 320364 456628 320416 456637
rect 320456 456628 320508 456680
rect 320640 456492 320692 456544
rect 273260 456220 273312 456272
rect 276204 456220 276256 456272
rect 273260 454316 273312 454368
rect 276296 454316 276348 454368
rect 273260 452412 273312 452464
rect 276388 452412 276440 452464
rect 320180 452319 320232 452328
rect 320180 452285 320189 452319
rect 320189 452285 320223 452319
rect 320223 452285 320232 452319
rect 320180 452276 320232 452285
rect 320640 449871 320692 449880
rect 320640 449837 320649 449871
rect 320649 449837 320683 449871
rect 320683 449837 320692 449871
rect 320640 449828 320692 449837
rect 320364 447355 320416 447364
rect 320364 447321 320373 447355
rect 320373 447321 320407 447355
rect 320407 447321 320416 447355
rect 320364 447312 320416 447321
rect 320456 447312 320508 447364
rect 320548 447312 320600 447364
rect 320456 447176 320508 447228
rect 320548 447176 320600 447228
rect 320640 447108 320692 447160
rect 273444 447040 273496 447092
rect 320364 447015 320416 447024
rect 320364 446981 320373 447015
rect 320373 446981 320407 447015
rect 320407 446981 320416 447015
rect 320364 446972 320416 446981
rect 320824 446904 320876 446956
rect 320732 446836 320784 446888
rect 320824 446768 320876 446820
rect 273444 444796 273496 444848
rect 276480 444796 276532 444848
rect 273444 442892 273496 442944
rect 276572 442892 276624 442944
rect 320548 442416 320600 442468
rect 320732 442416 320784 442468
rect 320548 442144 320600 442196
rect 320456 442008 320508 442060
rect 273444 441260 273496 441312
rect 277308 441260 277360 441312
rect 273444 439696 273496 439748
rect 277216 439696 277268 439748
rect 273260 433372 273312 433424
rect 274824 433372 274876 433424
rect 320272 431944 320324 431996
rect 320824 431944 320876 431996
rect 273260 431468 273312 431520
rect 274916 431468 274968 431520
rect 273260 429564 273312 429616
rect 275008 429564 275060 429616
rect 320272 427728 320324 427780
rect 320824 427728 320876 427780
rect 273260 427660 273312 427712
rect 275100 427660 275152 427712
rect 273260 425756 273312 425808
rect 275192 425756 275244 425808
rect 273444 423988 273496 424040
rect 275928 423988 275980 424040
rect 273444 422016 273496 422068
rect 275836 422016 275888 422068
rect 273444 420044 273496 420096
rect 275744 420044 275796 420096
rect 273444 418072 273496 418124
rect 279516 418072 279568 418124
rect 273444 416236 273496 416288
rect 278596 416236 278648 416288
rect 273444 414332 273496 414384
rect 277032 414332 277084 414384
rect 273444 412428 273496 412480
rect 276940 412428 276992 412480
rect 273444 410524 273496 410576
rect 276848 410524 276900 410576
rect 273444 408620 273496 408672
rect 276756 408620 276808 408672
rect 273444 406716 273496 406768
rect 276664 406716 276716 406768
rect 273444 402908 273496 402960
rect 275652 402908 275704 402960
rect 273444 401004 273496 401056
rect 275560 401004 275612 401056
rect 273444 400120 273496 400172
rect 320732 400120 320784 400172
rect 320180 398828 320232 398880
rect 320824 398828 320876 398880
rect 273444 397400 273496 397452
rect 320640 397400 320692 397452
rect 273260 396788 273312 396840
rect 338672 396788 338724 396840
rect 275744 396720 275796 396772
rect 397460 396720 397512 396772
rect 275928 396652 275980 396704
rect 398840 396652 398892 396704
rect 275192 396584 275244 396636
rect 400220 396584 400272 396636
rect 275100 396516 275152 396568
rect 401600 396516 401652 396568
rect 275008 396448 275060 396500
rect 403348 396448 403400 396500
rect 274916 396380 274968 396432
rect 404360 396380 404412 396432
rect 406016 396380 406068 396432
rect 274824 396312 274876 396364
rect 273444 395972 273496 396024
rect 320548 395972 320600 396024
rect 273444 394612 273496 394664
rect 320456 394612 320508 394664
rect 275836 392028 275888 392080
rect 320180 392028 320232 392080
rect 275560 391960 275612 392012
rect 320272 391960 320324 392012
rect 273444 391892 273496 391944
rect 320364 391892 320416 391944
rect 275652 390532 275704 390584
rect 320088 390532 320140 390584
rect 273536 390464 273588 390516
rect 320180 390464 320232 390516
rect 273444 389172 273496 389224
rect 320272 389172 320324 389224
rect 273352 388016 273404 388068
rect 273536 388016 273588 388068
rect 320180 387812 320232 387864
rect 273628 387744 273680 387796
rect 320824 387744 320876 387796
rect 278688 387676 278740 387728
rect 320364 387676 320416 387728
rect 273628 387540 273680 387592
rect 277124 386316 277176 386368
rect 320272 386316 320324 386368
rect 273352 384956 273404 385008
rect 320180 384956 320232 385008
rect 302976 384888 303028 384940
rect 320364 384888 320416 384940
rect 304264 383596 304316 383648
rect 320180 383596 320232 383648
rect 273352 383528 273404 383580
rect 273444 383324 273496 383376
rect 305644 382168 305696 382220
rect 320548 382168 320600 382220
rect 320640 381352 320692 381404
rect 308404 380808 308456 380860
rect 320180 380808 320232 380860
rect 320824 380307 320876 380316
rect 320824 380273 320833 380307
rect 320833 380273 320867 380307
rect 320867 380273 320876 380307
rect 320824 380264 320876 380273
rect 273536 380196 273588 380248
rect 320088 380196 320140 380248
rect 273628 380128 273680 380180
rect 320456 380128 320508 380180
rect 320640 379763 320692 379772
rect 320640 379729 320649 379763
rect 320649 379729 320683 379763
rect 320683 379729 320692 379763
rect 320640 379720 320692 379729
rect 320732 379559 320784 379568
rect 320732 379525 320741 379559
rect 320741 379525 320775 379559
rect 320775 379525 320784 379559
rect 320732 379516 320784 379525
rect 309784 379448 309836 379500
rect 320272 379448 320324 379500
rect 273536 378904 273588 378956
rect 274456 378904 274508 378956
rect 274640 378836 274692 378888
rect 320364 378836 320416 378888
rect 274456 378768 274508 378820
rect 320824 378768 320876 378820
rect 320548 378292 320600 378344
rect 315304 376796 315356 376848
rect 319996 376796 320048 376848
rect 312544 376728 312596 376780
rect 319812 376728 319864 376780
rect 278596 376660 278648 376712
rect 320364 376524 320416 376576
rect 274456 375980 274508 376032
rect 320548 375980 320600 376032
rect 278412 375300 278464 375352
rect 320272 375300 320324 375352
rect 273628 374620 273680 374672
rect 273812 374620 273864 374672
rect 274456 374620 274508 374672
rect 273536 374484 273588 374536
rect 273812 374484 273864 374536
rect 320548 374416 320600 374468
rect 320640 374212 320692 374264
rect 278320 373940 278372 373992
rect 320180 373940 320232 373992
rect 320088 372963 320140 372972
rect 320088 372929 320097 372963
rect 320097 372929 320131 372963
rect 320131 372929 320140 372963
rect 320088 372920 320140 372929
rect 278228 372512 278280 372564
rect 320364 372444 320416 372496
rect 274456 371832 274508 371884
rect 319904 371832 319956 371884
rect 320548 371832 320600 371884
rect 320824 371603 320876 371612
rect 320824 371569 320833 371603
rect 320833 371569 320867 371603
rect 320867 371569 320876 371603
rect 320824 371560 320876 371569
rect 278136 371152 278188 371204
rect 320272 371152 320324 371204
rect 320824 371016 320876 371068
rect 274456 370472 274508 370524
rect 319996 370472 320048 370524
rect 320640 370472 320692 370524
rect 320824 370515 320876 370524
rect 320824 370481 320833 370515
rect 320833 370481 320867 370515
rect 320867 370481 320876 370515
rect 320824 370472 320876 370481
rect 320640 370268 320692 370320
rect 280804 369792 280856 369844
rect 320180 369792 320232 369844
rect 283564 369724 283616 369776
rect 319812 369724 319864 369776
rect 319996 369452 320048 369504
rect 320640 369452 320692 369504
rect 319904 369044 319956 369096
rect 320364 369044 320416 369096
rect 320456 368568 320508 368620
rect 278044 368432 278096 368484
rect 320456 368432 320508 368484
rect 320272 367863 320324 367872
rect 320272 367829 320281 367863
rect 320281 367829 320315 367863
rect 320315 367829 320324 367863
rect 320272 367820 320324 367829
rect 284944 366868 284996 366920
rect 318800 366256 318852 366308
rect 320364 365780 320416 365832
rect 320180 365712 320232 365764
rect 286324 365644 286376 365696
rect 320364 365644 320416 365696
rect 287704 364284 287756 364336
rect 320272 364284 320324 364336
rect 319996 363740 320048 363792
rect 273720 362856 273772 362908
rect 320456 362856 320508 362908
rect 290464 362788 290516 362840
rect 319812 362788 319864 362840
rect 320088 362652 320140 362704
rect 273536 361020 273588 361072
rect 275468 361020 275520 361072
rect 320272 360884 320324 360936
rect 320732 360884 320784 360936
rect 320824 360272 320876 360324
rect 320456 360204 320508 360256
rect 320272 360179 320324 360188
rect 320272 360145 320281 360179
rect 320281 360145 320315 360179
rect 320315 360145 320324 360179
rect 320272 360136 320324 360145
rect 320272 360000 320324 360052
rect 320732 360000 320784 360052
rect 320732 359864 320784 359916
rect 319996 359796 320048 359848
rect 320824 359796 320876 359848
rect 273812 359660 273864 359712
rect 275376 359660 275428 359712
rect 320180 356872 320232 356924
rect 320364 356872 320416 356924
rect 291844 355988 291896 356040
rect 320180 355988 320232 356040
rect 274364 355920 274416 355972
rect 275284 355920 275336 355972
rect 320640 355852 320692 355904
rect 294604 354628 294656 354680
rect 320180 354628 320232 354680
rect 273812 353404 273864 353456
rect 274824 353404 274876 353456
rect 274272 353200 274324 353252
rect 320180 353200 320232 353252
rect 297364 351840 297416 351892
rect 320272 351840 320324 351892
rect 274180 350412 274232 350464
rect 320272 350412 320324 350464
rect 273536 349596 273588 349648
rect 275008 349596 275060 349648
rect 274088 349052 274140 349104
rect 320180 349052 320232 349104
rect 298744 348984 298796 349036
rect 320364 348984 320416 349036
rect 273536 347692 273588 347744
rect 275100 347692 275152 347744
rect 301504 347692 301556 347744
rect 320180 347692 320232 347744
rect 273996 346332 274048 346384
rect 320180 346332 320232 346384
rect 273536 345856 273588 345908
rect 275192 345856 275244 345908
rect 273628 343952 273680 344004
rect 275928 343952 275980 344004
rect 273536 342116 273588 342168
rect 275744 342116 275796 342168
rect 273536 340076 273588 340128
rect 275836 340076 275888 340128
rect 273812 335248 273864 335300
rect 302884 335248 302936 335300
rect 274272 332460 274324 332512
rect 279424 332460 279476 332512
rect 273352 331304 273404 331356
rect 273536 331304 273588 331356
rect 273352 331168 273404 331220
rect 319444 331168 319496 331220
rect 273996 329740 274048 329792
rect 316684 329740 316736 329792
rect 273536 323280 273588 323332
rect 275652 323280 275704 323332
rect 273444 321240 273496 321292
rect 275560 321240 275612 321292
rect 230664 320152 230716 320204
rect 231492 320152 231544 320204
rect 235632 320152 235684 320204
rect 240692 320152 240744 320204
rect 241336 320152 241388 320204
rect 241888 320152 241940 320204
rect 242716 320152 242768 320204
rect 244280 320152 244332 320204
rect 245108 320152 245160 320204
rect 245660 320152 245712 320204
rect 246396 320152 246448 320204
rect 247132 320152 247184 320204
rect 248052 320152 248104 320204
rect 253020 320152 253072 320204
rect 253756 320152 253808 320204
rect 255964 320152 256016 320204
rect 256332 320152 256384 320204
rect 260840 320152 260892 320204
rect 261576 320152 261628 320204
rect 263600 320152 263652 320204
rect 264060 320152 264112 320204
rect 266636 320152 266688 320204
rect 267464 320152 267516 320204
rect 269120 320152 269172 320204
rect 269856 320152 269908 320204
rect 235448 319880 235500 319932
rect 251456 319404 251508 319456
rect 251640 319404 251692 319456
rect 267372 319404 267424 319456
rect 267556 319404 267608 319456
rect 271696 319404 271748 319456
rect 271880 319404 271932 319456
rect 142068 318792 142120 318844
rect 150808 318792 150860 318844
rect 49608 318724 49660 318776
rect 87052 318724 87104 318776
rect 118424 318724 118476 318776
rect 133144 318724 133196 318776
rect 135720 318724 135772 318776
rect 159456 318724 159508 318776
rect 164240 318724 164292 318776
rect 167000 318724 167052 318776
rect 46848 318656 46900 318708
rect 85856 318656 85908 318708
rect 126612 318656 126664 318708
rect 145656 318656 145708 318708
rect 148140 318656 148192 318708
rect 164148 318656 164200 318708
rect 39948 318588 40000 318640
rect 83740 318588 83792 318640
rect 91008 318588 91060 318640
rect 101496 318588 101548 318640
rect 117136 318588 117188 318640
rect 133236 318588 133288 318640
rect 134524 318588 134576 318640
rect 159364 318588 159416 318640
rect 162952 318588 163004 318640
rect 164056 318588 164108 318640
rect 41328 318520 41380 318572
rect 84200 318520 84252 318572
rect 93124 318520 93176 318572
rect 99472 318520 99524 318572
rect 127900 318520 127952 318572
rect 164884 318520 164936 318572
rect 185216 318520 185268 318572
rect 192668 318724 192720 318776
rect 204996 318724 205048 318776
rect 208676 318724 208728 318776
rect 214932 318724 214984 318776
rect 220176 318724 220228 318776
rect 237656 318792 237708 318844
rect 238024 318792 238076 318844
rect 240508 318792 240560 318844
rect 240876 318792 240928 318844
rect 241612 318792 241664 318844
rect 242072 318792 242124 318844
rect 245016 318792 245068 318844
rect 245568 318792 245620 318844
rect 245752 318792 245804 318844
rect 245844 318792 245896 318844
rect 256424 318792 256476 318844
rect 256608 318792 256660 318844
rect 261576 318792 261628 318844
rect 261668 318792 261720 318844
rect 269212 318792 269264 318844
rect 269396 318792 269448 318844
rect 353944 318724 353996 318776
rect 197544 318656 197596 318708
rect 202144 318656 202196 318708
rect 202696 318656 202748 318708
rect 214472 318656 214524 318708
rect 215116 318656 215168 318708
rect 222292 318656 222344 318708
rect 356704 318656 356756 318708
rect 195060 318588 195112 318640
rect 329104 318588 329156 318640
rect 38568 318452 38620 318504
rect 34428 318384 34480 318436
rect 81716 318452 81768 318504
rect 93768 318452 93820 318504
rect 102324 318452 102376 318504
rect 132132 318452 132184 318504
rect 132408 318452 132460 318504
rect 133512 318452 133564 318504
rect 157984 318452 158036 318504
rect 161664 318452 161716 318504
rect 331864 318520 331916 318572
rect 215944 318452 215996 318504
rect 217324 318452 217376 318504
rect 348424 318452 348476 318504
rect 78864 318384 78916 318436
rect 33048 318316 33100 318368
rect 81348 318384 81400 318436
rect 88984 318384 89036 318436
rect 98184 318384 98236 318436
rect 123760 318384 123812 318436
rect 147404 318384 147456 318436
rect 149704 318384 149756 318436
rect 149796 318384 149848 318436
rect 150256 318384 150308 318436
rect 159272 318384 159324 318436
rect 91744 318316 91796 318368
rect 101128 318316 101180 318368
rect 124220 318316 124272 318368
rect 149336 318316 149388 318368
rect 153844 318316 153896 318368
rect 154304 318316 154356 318368
rect 160468 318316 160520 318368
rect 209044 318384 209096 318436
rect 209964 318384 210016 318436
rect 202512 318316 202564 318368
rect 212448 318384 212500 318436
rect 347044 318384 347096 318436
rect 345664 318316 345716 318368
rect 27528 318248 27580 318300
rect 79232 318248 79284 318300
rect 89076 318248 89128 318300
rect 99840 318248 99892 318300
rect 108948 318248 109000 318300
rect 111064 318248 111116 318300
rect 120080 318248 120132 318300
rect 140688 318248 140740 318300
rect 31668 318180 31720 318232
rect 26148 318112 26200 318164
rect 24768 318044 24820 318096
rect 78404 318112 78456 318164
rect 80888 318112 80940 318164
rect 88248 318112 88300 318164
rect 100300 318180 100352 318232
rect 113088 318180 113140 318232
rect 123484 318180 123536 318232
rect 128268 318180 128320 318232
rect 97264 318112 97316 318164
rect 100668 318112 100720 318164
rect 110144 318112 110196 318164
rect 111156 318112 111208 318164
rect 112260 318112 112312 318164
rect 116584 318112 116636 318164
rect 121276 318112 121328 318164
rect 83372 318044 83424 318096
rect 48136 317976 48188 318028
rect 86224 318044 86276 318096
rect 111800 318044 111852 318096
rect 92848 317976 92900 318028
rect 110972 317976 111024 318028
rect 111708 317976 111760 318028
rect 112628 317976 112680 318028
rect 113088 317976 113140 318028
rect 50988 317908 51040 317960
rect 87512 317908 87564 317960
rect 109316 317908 109368 317960
rect 110236 317908 110288 317960
rect 113916 318044 113968 318096
rect 114376 318044 114428 318096
rect 114744 318044 114796 318096
rect 115664 318044 115716 318096
rect 116308 318044 116360 318096
rect 117228 318044 117280 318096
rect 119252 318044 119304 318096
rect 119896 318044 119948 318096
rect 121736 318044 121788 318096
rect 122564 318044 122616 318096
rect 152464 318248 152516 318300
rect 200028 318248 200080 318300
rect 336004 318248 336056 318300
rect 163964 318180 164016 318232
rect 218704 318180 218756 318232
rect 224776 318180 224828 318232
rect 360844 318180 360896 318232
rect 147864 318112 147916 318164
rect 150900 318112 150952 318164
rect 156604 318112 156656 318164
rect 113456 317976 113508 318028
rect 114468 317976 114520 318028
rect 115940 317976 115992 318028
rect 117136 317976 117188 318028
rect 118792 317976 118844 318028
rect 119988 317976 120040 318028
rect 120908 317976 120960 318028
rect 120264 317908 120316 317960
rect 56416 317840 56468 317892
rect 89536 317840 89588 317892
rect 96528 317840 96580 317892
rect 103152 317840 103204 317892
rect 115112 317840 115164 317892
rect 115848 317840 115900 317892
rect 119620 317840 119672 317892
rect 122932 317908 122984 317960
rect 124128 317908 124180 317960
rect 124588 317908 124640 317960
rect 125508 317908 125560 317960
rect 126244 317908 126296 317960
rect 126888 317908 126940 317960
rect 127440 317908 127492 317960
rect 128268 317908 128320 317960
rect 128728 317908 128780 317960
rect 129648 317908 129700 317960
rect 129924 317908 129976 317960
rect 131028 317908 131080 317960
rect 132868 317976 132920 318028
rect 133788 317976 133840 318028
rect 135352 317976 135404 318028
rect 136548 317976 136600 318028
rect 137008 317976 137060 318028
rect 137928 317976 137980 318028
rect 145656 318044 145708 318096
rect 146852 318044 146904 318096
rect 146576 317976 146628 318028
rect 125876 317840 125928 317892
rect 131212 317840 131264 317892
rect 132408 317840 132460 317892
rect 57888 317772 57940 317824
rect 64788 317704 64840 317756
rect 84936 317772 84988 317824
rect 89996 317704 90048 317756
rect 96344 317772 96396 317824
rect 102784 317772 102836 317824
rect 122104 317772 122156 317824
rect 122748 317772 122800 317824
rect 129096 317772 129148 317824
rect 129464 317772 129516 317824
rect 130384 317772 130436 317824
rect 130844 317772 130896 317824
rect 131580 317772 131632 317824
rect 132224 317772 132276 317824
rect 98644 317704 98696 317756
rect 123392 317704 123444 317756
rect 124036 317704 124088 317756
rect 127072 317704 127124 317756
rect 128176 317704 128228 317756
rect 63408 317636 63460 317688
rect 91652 317636 91704 317688
rect 97908 317636 97960 317688
rect 103612 317636 103664 317688
rect 132132 317636 132184 317688
rect 134524 317908 134576 317960
rect 141424 317908 141476 317960
rect 136180 317840 136232 317892
rect 153844 317908 153896 317960
rect 134064 317772 134116 317824
rect 135168 317772 135220 317824
rect 137376 317772 137428 317824
rect 148324 317772 148376 317824
rect 134892 317704 134944 317756
rect 145564 317704 145616 317756
rect 147680 317704 147732 317756
rect 148784 317704 148836 317756
rect 167644 317840 167696 317892
rect 211988 318112 212040 318164
rect 215300 318112 215352 318164
rect 216496 318112 216548 318164
rect 218612 318112 218664 318164
rect 219348 318112 219400 318164
rect 220268 318112 220320 318164
rect 220728 318112 220780 318164
rect 221096 318112 221148 318164
rect 222108 318112 222160 318164
rect 342904 318112 342956 318164
rect 207848 318044 207900 318096
rect 208308 318044 208360 318096
rect 340144 318044 340196 318096
rect 202144 317976 202196 318028
rect 203340 317976 203392 318028
rect 203892 317976 203944 318028
rect 206192 317976 206244 318028
rect 206652 317976 206704 318028
rect 207480 317976 207532 318028
rect 208216 317976 208268 318028
rect 211620 317976 211672 318028
rect 212448 317976 212500 318028
rect 213276 317976 213328 318028
rect 213644 317976 213696 318028
rect 214104 317976 214156 318028
rect 215208 317976 215260 318028
rect 215760 317976 215812 318028
rect 216404 317976 216456 318028
rect 216956 317976 217008 318028
rect 217876 317976 217928 318028
rect 218152 317976 218204 318028
rect 219164 317976 219216 318028
rect 219440 317976 219492 318028
rect 220544 317976 220596 318028
rect 221464 317976 221516 318028
rect 222016 317976 222068 318028
rect 222752 317976 222804 318028
rect 223488 317976 223540 318028
rect 223948 317976 224000 318028
rect 224776 317976 224828 318028
rect 226432 317976 226484 318028
rect 227628 317976 227680 318028
rect 228088 317976 228140 318028
rect 228824 317976 228876 318028
rect 229284 317976 229336 318028
rect 230296 317976 230348 318028
rect 231860 317976 231912 318028
rect 233056 317976 233108 318028
rect 233332 317976 233384 318028
rect 234252 317976 234304 318028
rect 349804 317976 349856 318028
rect 190184 317908 190236 317960
rect 322204 317908 322256 317960
rect 325056 317840 325108 317892
rect 160744 317772 160796 317824
rect 182732 317772 182784 317824
rect 193772 317772 193824 317824
rect 155224 317704 155276 317756
rect 177764 317704 177816 317756
rect 187700 317704 187752 317756
rect 318064 317772 318116 317824
rect 196348 317704 196400 317756
rect 197176 317704 197228 317756
rect 198832 317704 198884 317756
rect 200028 317704 200080 317756
rect 202972 317704 203024 317756
rect 204076 317704 204128 317756
rect 92480 317568 92532 317620
rect 100024 317568 100076 317620
rect 104348 317568 104400 317620
rect 117596 317568 117648 317620
rect 118516 317568 118568 317620
rect 120448 317568 120500 317620
rect 121368 317568 121420 317620
rect 135904 317636 135956 317688
rect 138204 317636 138256 317688
rect 139400 317568 139452 317620
rect 140688 317568 140740 317620
rect 144368 317568 144420 317620
rect 144828 317568 144880 317620
rect 158076 317636 158128 317688
rect 180248 317636 180300 317688
rect 151084 317568 151136 317620
rect 64696 317500 64748 317552
rect 92020 317500 92072 317552
rect 103428 317500 103480 317552
rect 105636 317500 105688 317552
rect 137744 317500 137796 317552
rect 153936 317568 153988 317620
rect 166172 317568 166224 317620
rect 171600 317568 171652 317620
rect 172152 317568 172204 317620
rect 183928 317568 183980 317620
rect 184848 317568 184900 317620
rect 186412 317636 186464 317688
rect 187608 317636 187660 317688
rect 189724 317636 189776 317688
rect 190276 317636 190328 317688
rect 191012 317636 191064 317688
rect 191564 317636 191616 317688
rect 191840 317636 191892 317688
rect 193036 317636 193088 317688
rect 193864 317636 193916 317688
rect 194508 317636 194560 317688
rect 194692 317636 194744 317688
rect 195796 317636 195848 317688
rect 313924 317636 313976 317688
rect 307024 317568 307076 317620
rect 311164 317568 311216 317620
rect 152188 317500 152240 317552
rect 153108 317500 153160 317552
rect 154672 317500 154724 317552
rect 155868 317500 155920 317552
rect 155960 317500 156012 317552
rect 157248 317500 157300 317552
rect 158812 317500 158864 317552
rect 159916 317500 159968 317552
rect 163780 317500 163832 317552
rect 164056 317500 164108 317552
rect 164976 317500 165028 317552
rect 165528 317500 165580 317552
rect 165804 317500 165856 317552
rect 166908 317500 166960 317552
rect 167460 317500 167512 317552
rect 168288 317500 168340 317552
rect 171968 317500 172020 317552
rect 172428 317500 172480 317552
rect 173256 317500 173308 317552
rect 173808 317500 173860 317552
rect 174084 317500 174136 317552
rect 175188 317500 175240 317552
rect 175740 317500 175792 317552
rect 176568 317500 176620 317552
rect 177396 317500 177448 317552
rect 177856 317500 177908 317552
rect 178592 317500 178644 317552
rect 179052 317500 179104 317552
rect 179420 317500 179472 317552
rect 180708 317500 180760 317552
rect 183560 317500 183612 317552
rect 184664 317500 184716 317552
rect 300124 317500 300176 317552
rect 68284 317432 68336 317484
rect 69664 317432 69716 317484
rect 88340 317432 88392 317484
rect 100116 317432 100168 317484
rect 101956 317432 102008 317484
rect 102784 317432 102836 317484
rect 103980 317432 104032 317484
rect 104808 317432 104860 317484
rect 106004 317432 106056 317484
rect 108120 317432 108172 317484
rect 108856 317432 108908 317484
rect 110604 317432 110656 317484
rect 113824 317432 113876 317484
rect 133696 317432 133748 317484
rect 138572 317432 138624 317484
rect 139308 317432 139360 317484
rect 139860 317432 139912 317484
rect 140596 317432 140648 317484
rect 141056 317432 141108 317484
rect 142068 317432 142120 317484
rect 142344 317432 142396 317484
rect 143448 317432 143500 317484
rect 143540 317432 143592 317484
rect 144644 317432 144696 317484
rect 145196 317432 145248 317484
rect 146116 317432 146168 317484
rect 146484 317432 146536 317484
rect 147404 317432 147456 317484
rect 93032 317364 93084 317416
rect 94044 317407 94096 317416
rect 94044 317373 94053 317407
rect 94053 317373 94087 317407
rect 94087 317373 94096 317407
rect 94044 317364 94096 317373
rect 139216 317364 139268 317416
rect 148508 317432 148560 317484
rect 148968 317432 149020 317484
rect 151820 317432 151872 317484
rect 152648 317432 152700 317484
rect 153476 317432 153528 317484
rect 154488 317432 154540 317484
rect 155132 317432 155184 317484
rect 155776 317432 155828 317484
rect 156328 317432 156380 317484
rect 157064 317432 157116 317484
rect 159640 317432 159692 317484
rect 160008 317432 160060 317484
rect 160836 317432 160888 317484
rect 161388 317432 161440 317484
rect 162124 317432 162176 317484
rect 162768 317432 162820 317484
rect 163320 317432 163372 317484
rect 164148 317432 164200 317484
rect 164608 317432 164660 317484
rect 165344 317432 165396 317484
rect 166264 317432 166316 317484
rect 166816 317432 166868 317484
rect 167092 317432 167144 317484
rect 168104 317432 168156 317484
rect 168748 317432 168800 317484
rect 169576 317432 169628 317484
rect 169944 317432 169996 317484
rect 170956 317432 171008 317484
rect 171232 317432 171284 317484
rect 172244 317432 172296 317484
rect 172796 317432 172848 317484
rect 173624 317432 173676 317484
rect 174452 317432 174504 317484
rect 175096 317432 175148 317484
rect 175280 317432 175332 317484
rect 176292 317432 176344 317484
rect 176936 317432 176988 317484
rect 177948 317432 178000 317484
rect 178224 317432 178276 317484
rect 179144 317432 179196 317484
rect 179880 317432 179932 317484
rect 180524 317432 180576 317484
rect 181076 317432 181128 317484
rect 181628 317432 181680 317484
rect 182364 317432 182416 317484
rect 183192 317432 183244 317484
rect 184388 317432 184440 317484
rect 184756 317432 184808 317484
rect 185584 317432 185636 317484
rect 186228 317432 186280 317484
rect 186872 317432 186924 317484
rect 187516 317432 187568 317484
rect 188068 317432 188120 317484
rect 188896 317432 188948 317484
rect 189356 317432 189408 317484
rect 190368 317432 190420 317484
rect 190552 317432 190604 317484
rect 191748 317432 191800 317484
rect 192208 317432 192260 317484
rect 192944 317432 192996 317484
rect 193496 317432 193548 317484
rect 194324 317432 194376 317484
rect 195520 317432 195572 317484
rect 195888 317432 195940 317484
rect 196716 317432 196768 317484
rect 197268 317432 197320 317484
rect 198004 317432 198056 317484
rect 198648 317432 198700 317484
rect 199200 317432 199252 317484
rect 199936 317432 199988 317484
rect 200488 317432 200540 317484
rect 201224 317432 201276 317484
rect 201684 317432 201736 317484
rect 202788 317432 202840 317484
rect 203800 317432 203852 317484
rect 204168 317432 204220 317484
rect 204628 317432 204680 317484
rect 205456 317432 205508 317484
rect 205824 317432 205876 317484
rect 206744 317432 206796 317484
rect 207020 317432 207072 317484
rect 208032 317432 208084 317484
rect 209136 317432 209188 317484
rect 209688 317432 209740 317484
rect 210332 317432 210384 317484
rect 211068 317432 211120 317484
rect 211160 317432 211212 317484
rect 212080 317432 212132 317484
rect 212816 317432 212868 317484
rect 213736 317432 213788 317484
rect 276664 317432 276716 317484
rect 236184 317407 236236 317416
rect 236184 317373 236193 317407
rect 236193 317373 236227 317407
rect 236227 317373 236236 317407
rect 236184 317364 236236 317373
rect 237656 317364 237708 317416
rect 238576 317364 238628 317416
rect 238944 317407 238996 317416
rect 238944 317373 238953 317407
rect 238953 317373 238987 317407
rect 238987 317373 238996 317407
rect 238944 317364 238996 317373
rect 240508 317364 240560 317416
rect 241244 317364 241296 317416
rect 248144 317364 248196 317416
rect 248328 317364 248380 317416
rect 266912 317364 266964 317416
rect 267648 317364 267700 317416
rect 267740 317364 267792 317416
rect 268936 317364 268988 317416
rect 238852 316140 238904 316192
rect 239956 316140 240008 316192
rect 251364 316140 251416 316192
rect 252468 316140 252520 316192
rect 95240 316072 95292 316124
rect 95884 316072 95936 316124
rect 244096 316072 244148 316124
rect 256976 316072 257028 316124
rect 257804 316072 257856 316124
rect 75920 316004 75972 316056
rect 76472 316004 76524 316056
rect 93952 316004 94004 316056
rect 94596 316004 94648 316056
rect 234896 316004 234948 316056
rect 235632 316004 235684 316056
rect 238852 316004 238904 316056
rect 239772 316004 239824 316056
rect 70400 315936 70452 315988
rect 71044 315936 71096 315988
rect 71872 315936 71924 315988
rect 72700 315936 72752 315988
rect 73160 315936 73212 315988
rect 73988 315936 74040 315988
rect 76012 315936 76064 315988
rect 76932 315936 76984 315988
rect 81532 315936 81584 315988
rect 82268 315936 82320 315988
rect 88432 315936 88484 315988
rect 88892 315936 88944 315988
rect 92572 315936 92624 315988
rect 93308 315936 93360 315988
rect 93860 315936 93912 315988
rect 94228 315936 94280 315988
rect 96620 315936 96672 315988
rect 97540 315936 97592 315988
rect 228732 315936 228784 315988
rect 229008 315936 229060 315988
rect 234620 315936 234672 315988
rect 235448 315936 235500 315988
rect 236000 315936 236052 315988
rect 236460 315936 236512 315988
rect 237472 315936 237524 315988
rect 238116 315936 238168 315988
rect 238760 315936 238812 315988
rect 239312 315936 239364 315988
rect 240140 315936 240192 315988
rect 240968 315936 241020 315988
rect 241520 315936 241572 315988
rect 242164 315936 242216 315988
rect 242900 315936 242952 315988
rect 243084 315936 243136 315988
rect 270500 316004 270552 316056
rect 271696 316004 271748 316056
rect 252560 315936 252612 315988
rect 253388 315936 253440 315988
rect 258816 315936 258868 315988
rect 259368 315936 259420 315988
rect 259460 315936 259512 315988
rect 260012 315936 260064 315988
rect 261300 315936 261352 315988
rect 262128 315936 262180 315988
rect 262312 315936 262364 315988
rect 157800 315868 157852 315920
rect 158444 315868 158496 315920
rect 244096 315868 244148 315920
rect 265256 315936 265308 315988
rect 266084 315936 266136 315988
rect 271236 315936 271288 315988
rect 271788 315936 271840 315988
rect 266452 315868 266504 315920
rect 267556 315868 267608 315920
rect 262404 315732 262456 315784
rect 230572 315324 230624 315376
rect 231492 315324 231544 315376
rect 73252 315256 73304 315308
rect 73620 315256 73672 315308
rect 246488 315188 246540 315240
rect 246948 315188 247000 315240
rect 255320 314984 255372 315036
rect 256424 314984 256476 315036
rect 257436 314984 257488 315036
rect 257896 314984 257948 315036
rect 267832 314644 267884 314696
rect 268108 314644 268160 314696
rect 241612 314100 241664 314152
rect 242624 314100 242676 314152
rect 250536 313896 250588 313948
rect 250996 313896 251048 313948
rect 264152 313896 264204 313948
rect 264704 313896 264756 313948
rect 262312 312740 262364 312792
rect 262772 312740 262824 312792
rect 262220 312672 262272 312724
rect 262496 312672 262548 312724
rect 150900 312604 150952 312656
rect 151176 312604 151228 312656
rect 105084 311924 105136 311976
rect 233332 311788 233384 311840
rect 234344 311788 234396 311840
rect 105176 311720 105228 311772
rect 248512 311584 248564 311636
rect 249432 311584 249484 311636
rect 249892 311584 249944 311636
rect 250628 311584 250680 311636
rect 223672 311176 223724 311228
rect 224868 311176 224920 311228
rect 247224 309748 247276 309800
rect 248328 309748 248380 309800
rect 251732 309544 251784 309596
rect 77576 309272 77628 309324
rect 193956 309204 194008 309256
rect 70860 309179 70912 309188
rect 70860 309145 70869 309179
rect 70869 309145 70903 309179
rect 70903 309145 70912 309179
rect 70860 309136 70912 309145
rect 77576 309136 77628 309188
rect 78956 309136 79008 309188
rect 79416 309136 79468 309188
rect 84660 309136 84712 309188
rect 85120 309136 85172 309188
rect 151084 309136 151136 309188
rect 162124 309179 162176 309188
rect 162124 309145 162133 309179
rect 162133 309145 162167 309179
rect 162167 309145 162176 309179
rect 162124 309136 162176 309145
rect 198004 309179 198056 309188
rect 198004 309145 198013 309179
rect 198013 309145 198047 309179
rect 198047 309145 198056 309179
rect 198004 309136 198056 309145
rect 204904 309179 204956 309188
rect 204904 309145 204913 309179
rect 204913 309145 204947 309179
rect 204947 309145 204956 309179
rect 204904 309136 204956 309145
rect 251272 309136 251324 309188
rect 251456 309136 251508 309188
rect 259184 309136 259236 309188
rect 259276 309136 259328 309188
rect 270776 309136 270828 309188
rect 271512 309136 271564 309188
rect 245568 309111 245620 309120
rect 245568 309077 245577 309111
rect 245577 309077 245611 309111
rect 245611 309077 245620 309111
rect 245568 309068 245620 309077
rect 254032 309111 254084 309120
rect 254032 309077 254041 309111
rect 254041 309077 254075 309111
rect 254075 309077 254084 309111
rect 254032 309068 254084 309077
rect 264704 309068 264756 309120
rect 325056 309068 325108 309120
rect 264796 309000 264848 309052
rect 94044 307887 94096 307896
rect 94044 307853 94053 307887
rect 94053 307853 94087 307887
rect 94087 307853 94096 307887
rect 94044 307844 94096 307853
rect 70860 307819 70912 307828
rect 70860 307785 70869 307819
rect 70869 307785 70903 307819
rect 70903 307785 70912 307819
rect 70860 307776 70912 307785
rect 73528 307776 73580 307828
rect 73620 307776 73672 307828
rect 92848 307819 92900 307828
rect 92848 307785 92857 307819
rect 92857 307785 92891 307819
rect 92891 307785 92900 307819
rect 92848 307776 92900 307785
rect 193864 307819 193916 307828
rect 193864 307785 193873 307819
rect 193873 307785 193907 307819
rect 193907 307785 193916 307819
rect 193864 307776 193916 307785
rect 236184 307819 236236 307828
rect 236184 307785 236193 307819
rect 236193 307785 236227 307819
rect 236227 307785 236236 307819
rect 236184 307776 236236 307785
rect 238944 307819 238996 307828
rect 238944 307785 238953 307819
rect 238953 307785 238987 307819
rect 238987 307785 238996 307819
rect 238944 307776 238996 307785
rect 94044 307751 94096 307760
rect 94044 307717 94053 307751
rect 94053 307717 94087 307751
rect 94087 307717 94096 307751
rect 94044 307708 94096 307717
rect 247040 307300 247092 307352
rect 248144 307300 248196 307352
rect 255320 307096 255372 307148
rect 256516 307096 256568 307148
rect 224960 307028 225012 307080
rect 226156 307028 226208 307080
rect 230572 307028 230624 307080
rect 231584 307028 231636 307080
rect 231860 307028 231912 307080
rect 233056 307028 233108 307080
rect 233240 307028 233292 307080
rect 234528 307028 234580 307080
rect 234620 307028 234672 307080
rect 235816 307028 235868 307080
rect 236000 307028 236052 307080
rect 237288 307028 237340 307080
rect 237380 307028 237432 307080
rect 238668 307028 238720 307080
rect 238852 307028 238904 307080
rect 239864 307028 239916 307080
rect 240140 307028 240192 307080
rect 241428 307028 241480 307080
rect 241520 307028 241572 307080
rect 242808 307028 242860 307080
rect 244280 307028 244332 307080
rect 245476 307028 245528 307080
rect 245660 307028 245712 307080
rect 246856 307028 246908 307080
rect 248420 307028 248472 307080
rect 249708 307028 249760 307080
rect 249800 307028 249852 307080
rect 251088 307028 251140 307080
rect 252560 307028 252612 307080
rect 253848 307028 253900 307080
rect 253940 307028 253992 307080
rect 255136 307028 255188 307080
rect 255412 307028 255464 307080
rect 256424 307028 256476 307080
rect 256700 307028 256752 307080
rect 257988 307028 258040 307080
rect 259644 307028 259696 307080
rect 260748 307028 260800 307080
rect 262220 307028 262272 307080
rect 263324 307028 263376 307080
rect 267740 307028 267792 307080
rect 268936 307028 268988 307080
rect 270500 307028 270552 307080
rect 271604 307028 271656 307080
rect 230756 306960 230808 307012
rect 231768 306960 231820 307012
rect 238760 306960 238812 307012
rect 240048 306960 240100 307012
rect 255504 306960 255556 307012
rect 256608 306960 256660 307012
rect 259460 306960 259512 307012
rect 260656 306960 260708 307012
rect 262404 306960 262456 307012
rect 263508 306960 263560 307012
rect 266452 306960 266504 307012
rect 267556 306960 267608 307012
rect 251272 306935 251324 306944
rect 251272 306901 251281 306935
rect 251281 306901 251315 306935
rect 251315 306901 251324 306935
rect 251272 306892 251324 306901
rect 242900 306824 242952 306876
rect 243912 306824 243964 306876
rect 236184 306688 236236 306740
rect 237104 306688 237156 306740
rect 266544 306348 266596 306400
rect 267096 306348 267148 306400
rect 262312 306008 262364 306060
rect 263232 306008 263284 306060
rect 269120 305736 269172 305788
rect 270224 305736 270276 305788
rect 267096 303603 267148 303612
rect 267096 303569 267105 303603
rect 267105 303569 267139 303603
rect 267139 303569 267148 303603
rect 267096 303560 267148 303569
rect 70584 302268 70636 302320
rect 233424 302268 233476 302320
rect 259184 302268 259236 302320
rect 105176 302200 105228 302252
rect 106556 302200 106608 302252
rect 106740 302200 106792 302252
rect 211804 302200 211856 302252
rect 211988 302200 212040 302252
rect 232044 302200 232096 302252
rect 233148 302200 233200 302252
rect 234436 302200 234488 302252
rect 238944 302200 238996 302252
rect 70492 302132 70544 302184
rect 237472 302132 237524 302184
rect 238392 302132 238444 302184
rect 239772 302132 239824 302184
rect 259184 302132 259236 302184
rect 265808 302175 265860 302184
rect 265808 302141 265817 302175
rect 265817 302141 265851 302175
rect 265851 302141 265860 302175
rect 265808 302132 265860 302141
rect 259552 302064 259604 302116
rect 260472 302064 260524 302116
rect 92848 299548 92900 299600
rect 70676 299480 70728 299532
rect 70860 299480 70912 299532
rect 234252 299480 234304 299532
rect 234344 299480 234396 299532
rect 245568 299523 245620 299532
rect 245568 299489 245577 299523
rect 245577 299489 245611 299523
rect 245611 299489 245620 299523
rect 245568 299480 245620 299489
rect 250812 299480 250864 299532
rect 250996 299480 251048 299532
rect 255044 299480 255096 299532
rect 255228 299523 255280 299532
rect 255228 299489 255237 299523
rect 255237 299489 255271 299523
rect 255271 299489 255280 299523
rect 255228 299480 255280 299489
rect 266084 299480 266136 299532
rect 266176 299480 266228 299532
rect 267832 299480 267884 299532
rect 268752 299480 268804 299532
rect 324964 299523 325016 299532
rect 324964 299489 324973 299523
rect 324973 299489 325007 299523
rect 325007 299489 325016 299523
rect 324964 299480 325016 299489
rect 70492 299455 70544 299464
rect 70492 299421 70501 299455
rect 70501 299421 70535 299455
rect 70535 299421 70544 299455
rect 70492 299412 70544 299421
rect 73436 299412 73488 299464
rect 73528 299412 73580 299464
rect 92848 299412 92900 299464
rect 151084 299455 151136 299464
rect 151084 299421 151093 299455
rect 151093 299421 151127 299455
rect 151127 299421 151136 299455
rect 151084 299412 151136 299421
rect 227352 299455 227404 299464
rect 227352 299421 227361 299455
rect 227361 299421 227395 299455
rect 227395 299421 227404 299455
rect 227352 299412 227404 299421
rect 251272 299455 251324 299464
rect 251272 299421 251281 299455
rect 251281 299421 251315 299455
rect 251315 299421 251324 299455
rect 251272 299412 251324 299421
rect 267096 299455 267148 299464
rect 267096 299421 267105 299455
rect 267105 299421 267139 299455
rect 267139 299421 267148 299455
rect 267096 299412 267148 299421
rect 271512 299455 271564 299464
rect 271512 299421 271521 299455
rect 271521 299421 271555 299455
rect 271555 299421 271564 299455
rect 271512 299412 271564 299421
rect 89996 298188 90048 298240
rect 90180 298188 90232 298240
rect 94044 298163 94096 298172
rect 94044 298129 94053 298163
rect 94053 298129 94087 298163
rect 94087 298129 94096 298163
rect 94044 298120 94096 298129
rect 105084 298163 105136 298172
rect 105084 298129 105093 298163
rect 105093 298129 105127 298163
rect 105127 298129 105136 298163
rect 105084 298120 105136 298129
rect 255228 298163 255280 298172
rect 255228 298129 255237 298163
rect 255237 298129 255271 298163
rect 255271 298129 255280 298163
rect 255228 298120 255280 298129
rect 70768 298095 70820 298104
rect 70768 298061 70777 298095
rect 70777 298061 70811 298095
rect 70811 298061 70820 298095
rect 70768 298052 70820 298061
rect 73436 298052 73488 298104
rect 73528 298052 73580 298104
rect 193864 298095 193916 298104
rect 193864 298061 193873 298095
rect 193873 298061 193907 298095
rect 193907 298061 193916 298095
rect 193864 298052 193916 298061
rect 242624 298095 242676 298104
rect 242624 298061 242633 298095
rect 242633 298061 242667 298095
rect 242667 298061 242676 298095
rect 242624 298052 242676 298061
rect 243912 298095 243964 298104
rect 243912 298061 243921 298095
rect 243921 298061 243955 298095
rect 243955 298061 243964 298095
rect 243912 298052 243964 298061
rect 246948 298095 247000 298104
rect 246948 298061 246957 298095
rect 246957 298061 246991 298095
rect 246991 298061 247000 298095
rect 246948 298052 247000 298061
rect 248236 298095 248288 298104
rect 248236 298061 248245 298095
rect 248245 298061 248279 298095
rect 248279 298061 248288 298095
rect 248236 298052 248288 298061
rect 255228 298027 255280 298036
rect 255228 297993 255237 298027
rect 255237 297993 255271 298027
rect 255271 297993 255280 298027
rect 255228 297984 255280 297993
rect 259184 297440 259236 297492
rect 268844 297372 268896 297424
rect 269028 297372 269080 297424
rect 252192 297236 252244 297288
rect 234896 296760 234948 296812
rect 235724 296760 235776 296812
rect 72148 296667 72200 296676
rect 72148 296633 72157 296667
rect 72157 296633 72191 296667
rect 72191 296633 72200 296667
rect 72148 296624 72200 296633
rect 235724 296667 235776 296676
rect 235724 296633 235733 296667
rect 235733 296633 235767 296667
rect 235767 296633 235776 296667
rect 235724 296624 235776 296633
rect 244372 296284 244424 296336
rect 245384 296284 245436 296336
rect 249892 296284 249944 296336
rect 250904 296284 250956 296336
rect 245752 294584 245804 294636
rect 246764 294584 246816 294636
rect 247224 294584 247276 294636
rect 248052 294584 248104 294636
rect 248512 294584 248564 294636
rect 249524 294584 249576 294636
rect 252744 294584 252796 294636
rect 253664 294584 253716 294636
rect 271512 293539 271564 293548
rect 271512 293505 271521 293539
rect 271521 293505 271555 293539
rect 271555 293505 271564 293539
rect 271512 293496 271564 293505
rect 265900 292612 265952 292664
rect 265900 292476 265952 292528
rect 105176 292408 105228 292460
rect 105360 292408 105412 292460
rect 265992 292408 266044 292460
rect 78956 289892 79008 289944
rect 70584 289824 70636 289876
rect 77576 289824 77628 289876
rect 77668 289824 77720 289876
rect 78864 289824 78916 289876
rect 81716 289824 81768 289876
rect 81808 289824 81860 289876
rect 151084 289867 151136 289876
rect 151084 289833 151093 289867
rect 151093 289833 151127 289867
rect 151127 289833 151136 289867
rect 151084 289824 151136 289833
rect 227444 289824 227496 289876
rect 249432 289824 249484 289876
rect 249616 289824 249668 289876
rect 250812 289824 250864 289876
rect 250996 289824 251048 289876
rect 259276 289867 259328 289876
rect 259276 289833 259285 289867
rect 259285 289833 259319 289867
rect 259319 289833 259328 289867
rect 259276 289824 259328 289833
rect 325056 289756 325108 289808
rect 70768 288439 70820 288448
rect 70768 288405 70777 288439
rect 70777 288405 70811 288439
rect 70811 288405 70820 288439
rect 70768 288396 70820 288405
rect 94044 288396 94096 288448
rect 94136 288396 94188 288448
rect 193864 288439 193916 288448
rect 193864 288405 193873 288439
rect 193873 288405 193907 288439
rect 193907 288405 193916 288439
rect 193864 288396 193916 288405
rect 242624 288439 242676 288448
rect 242624 288405 242633 288439
rect 242633 288405 242667 288439
rect 242667 288405 242676 288439
rect 242624 288396 242676 288405
rect 243820 288396 243872 288448
rect 246948 288439 247000 288448
rect 246948 288405 246957 288439
rect 246957 288405 246991 288439
rect 246991 288405 247000 288439
rect 246948 288396 247000 288405
rect 248236 288439 248288 288448
rect 248236 288405 248245 288439
rect 248245 288405 248279 288439
rect 248279 288405 248288 288439
rect 248236 288396 248288 288405
rect 255228 288439 255280 288448
rect 255228 288405 255237 288439
rect 255237 288405 255271 288439
rect 255271 288405 255280 288439
rect 255228 288396 255280 288405
rect 72332 288328 72384 288380
rect 267188 287759 267240 287768
rect 267188 287725 267197 287759
rect 267197 287725 267231 287759
rect 267231 287725 267240 287759
rect 267188 287716 267240 287725
rect 268844 287716 268896 287768
rect 269028 287716 269080 287768
rect 235724 287147 235776 287156
rect 235724 287113 235733 287147
rect 235733 287113 235767 287147
rect 235767 287113 235776 287147
rect 235724 287104 235776 287113
rect 90088 287036 90140 287088
rect 90272 287036 90324 287088
rect 233976 287036 234028 287088
rect 234068 287036 234120 287088
rect 264520 284248 264572 284300
rect 264704 284248 264756 284300
rect 70768 282888 70820 282940
rect 77576 282956 77628 283008
rect 105176 282956 105228 283008
rect 78772 282888 78824 282940
rect 70860 282820 70912 282872
rect 77484 282820 77536 282872
rect 106556 282888 106608 282940
rect 106740 282888 106792 282940
rect 211804 282888 211856 282940
rect 211988 282888 212040 282940
rect 227260 282888 227312 282940
rect 227444 282888 227496 282940
rect 267280 282888 267332 282940
rect 105176 282752 105228 282804
rect 324964 280211 325016 280220
rect 324964 280177 324973 280211
rect 324973 280177 325007 280211
rect 325007 280177 325016 280211
rect 324964 280168 325016 280177
rect 105176 280143 105228 280152
rect 105176 280109 105185 280143
rect 105185 280109 105219 280143
rect 105219 280109 105228 280143
rect 105176 280100 105228 280109
rect 106648 280143 106700 280152
rect 106648 280109 106657 280143
rect 106657 280109 106691 280143
rect 106691 280109 106700 280143
rect 106648 280100 106700 280109
rect 151084 280143 151136 280152
rect 151084 280109 151093 280143
rect 151093 280109 151127 280143
rect 151127 280109 151136 280143
rect 151084 280100 151136 280109
rect 73436 278808 73488 278860
rect 73528 278808 73580 278860
rect 243820 278851 243872 278860
rect 243820 278817 243829 278851
rect 243829 278817 243863 278851
rect 243863 278817 243872 278851
rect 243820 278808 243872 278817
rect 78864 278783 78916 278792
rect 78864 278749 78873 278783
rect 78873 278749 78907 278783
rect 78907 278749 78916 278783
rect 78864 278740 78916 278749
rect 81624 278740 81676 278792
rect 81716 278672 81768 278724
rect 268844 278060 268896 278112
rect 269028 278060 269080 278112
rect 72332 277380 72384 277432
rect 72516 277380 72568 277432
rect 94136 277380 94188 277432
rect 94320 277380 94372 277432
rect 243820 277423 243872 277432
rect 243820 277389 243829 277423
rect 243829 277389 243863 277423
rect 243863 277389 243872 277423
rect 243820 277380 243872 277389
rect 81716 275952 81768 276004
rect 81900 275952 81952 276004
rect 264704 274592 264756 274644
rect 90088 273300 90140 273352
rect 106832 273232 106884 273284
rect 268660 273275 268712 273284
rect 268660 273241 268669 273275
rect 268669 273241 268703 273275
rect 268703 273241 268712 273275
rect 268660 273232 268712 273241
rect 105176 273139 105228 273148
rect 105176 273105 105185 273139
rect 105185 273105 105219 273139
rect 105219 273105 105228 273139
rect 105176 273096 105228 273105
rect 70768 270512 70820 270564
rect 70860 270512 70912 270564
rect 151084 270555 151136 270564
rect 151084 270521 151093 270555
rect 151093 270521 151127 270555
rect 151127 270521 151136 270555
rect 151084 270512 151136 270521
rect 77484 270444 77536 270496
rect 77576 270444 77628 270496
rect 78680 270444 78732 270496
rect 78864 270444 78916 270496
rect 105176 270487 105228 270496
rect 105176 270453 105185 270487
rect 105185 270453 105219 270487
rect 105219 270453 105228 270487
rect 105176 270444 105228 270453
rect 106832 270487 106884 270496
rect 106832 270453 106841 270487
rect 106841 270453 106875 270487
rect 106875 270453 106884 270487
rect 106832 270444 106884 270453
rect 242532 270444 242584 270496
rect 242624 270444 242676 270496
rect 249616 270487 249668 270496
rect 249616 270453 249625 270487
rect 249625 270453 249659 270487
rect 249659 270453 249668 270487
rect 249616 270444 249668 270453
rect 250996 270487 251048 270496
rect 250996 270453 251005 270487
rect 251005 270453 251039 270487
rect 251039 270453 251048 270487
rect 250996 270444 251048 270453
rect 252284 270487 252336 270496
rect 252284 270453 252293 270487
rect 252293 270453 252327 270487
rect 252327 270453 252336 270487
rect 252284 270444 252336 270453
rect 259276 270487 259328 270496
rect 259276 270453 259285 270487
rect 259285 270453 259319 270487
rect 259319 270453 259328 270487
rect 259276 270444 259328 270453
rect 325056 270444 325108 270496
rect 234160 270376 234212 270428
rect 92756 269084 92808 269136
rect 92848 269084 92900 269136
rect 193680 269084 193732 269136
rect 193864 269084 193916 269136
rect 243820 269152 243872 269204
rect 255228 269084 255280 269136
rect 255320 269084 255372 269136
rect 243728 269016 243780 269068
rect 268752 268200 268804 268252
rect 269028 268200 269080 268252
rect 72424 267724 72476 267776
rect 72608 267724 72660 267776
rect 73436 267724 73488 267776
rect 73620 267724 73672 267776
rect 89996 267767 90048 267776
rect 89996 267733 90005 267767
rect 90005 267733 90039 267767
rect 90039 267733 90048 267767
rect 89996 267724 90048 267733
rect 268660 267767 268712 267776
rect 268660 267733 268669 267767
rect 268669 267733 268703 267767
rect 268703 267733 268712 267767
rect 268660 267724 268712 267733
rect 264612 264979 264664 264988
rect 264612 264945 264621 264979
rect 264621 264945 264655 264979
rect 264655 264945 264664 264979
rect 264612 264936 264664 264945
rect 70492 264052 70544 264104
rect 70676 264052 70728 264104
rect 70768 263576 70820 263628
rect 73436 263576 73488 263628
rect 84476 263576 84528 263628
rect 84660 263576 84712 263628
rect 211804 263576 211856 263628
rect 211988 263576 212040 263628
rect 227260 263576 227312 263628
rect 227444 263576 227496 263628
rect 70676 263508 70728 263560
rect 73528 263440 73580 263492
rect 105176 263483 105228 263492
rect 105176 263449 105185 263483
rect 105185 263449 105219 263483
rect 105219 263449 105228 263483
rect 105176 263440 105228 263449
rect 92756 260856 92808 260908
rect 106924 260856 106976 260908
rect 234068 260899 234120 260908
rect 234068 260865 234077 260899
rect 234077 260865 234111 260899
rect 234111 260865 234120 260899
rect 234068 260856 234120 260865
rect 249616 260899 249668 260908
rect 249616 260865 249625 260899
rect 249625 260865 249659 260899
rect 249659 260865 249668 260899
rect 249616 260856 249668 260865
rect 250996 260899 251048 260908
rect 250996 260865 251005 260899
rect 251005 260865 251039 260899
rect 251039 260865 251048 260899
rect 250996 260856 251048 260865
rect 252284 260899 252336 260908
rect 252284 260865 252293 260899
rect 252293 260865 252327 260899
rect 252327 260865 252336 260899
rect 252284 260856 252336 260865
rect 259276 260899 259328 260908
rect 259276 260865 259285 260899
rect 259285 260865 259319 260899
rect 259319 260865 259328 260899
rect 259276 260856 259328 260865
rect 324964 260899 325016 260908
rect 324964 260865 324973 260899
rect 324973 260865 325007 260899
rect 325007 260865 325016 260899
rect 324964 260856 325016 260865
rect 89996 260788 90048 260840
rect 90088 260788 90140 260840
rect 105176 260831 105228 260840
rect 105176 260797 105185 260831
rect 105185 260797 105219 260831
rect 105219 260797 105228 260831
rect 105176 260788 105228 260797
rect 151084 260831 151136 260840
rect 151084 260797 151093 260831
rect 151093 260797 151127 260831
rect 151127 260797 151136 260831
rect 151084 260788 151136 260797
rect 92848 260720 92900 260772
rect 70676 259360 70728 259412
rect 268752 258748 268804 258800
rect 269028 258748 269080 258800
rect 89996 253920 90048 253972
rect 70492 253852 70544 253904
rect 70676 253852 70728 253904
rect 106924 253988 106976 254040
rect 106832 253852 106884 253904
rect 90088 253784 90140 253836
rect 105176 253827 105228 253836
rect 105176 253793 105185 253827
rect 105185 253793 105219 253827
rect 105219 253793 105228 253827
rect 105176 253784 105228 253793
rect 73528 252560 73580 252612
rect 94044 251200 94096 251252
rect 94136 251200 94188 251252
rect 151084 251243 151136 251252
rect 151084 251209 151093 251243
rect 151093 251209 151127 251243
rect 151127 251209 151136 251243
rect 151084 251200 151136 251209
rect 234068 251200 234120 251252
rect 234160 251200 234212 251252
rect 324780 251200 324832 251252
rect 324964 251200 325016 251252
rect 105176 251132 105228 251184
rect 252284 251175 252336 251184
rect 252284 251141 252293 251175
rect 252293 251141 252327 251175
rect 252327 251141 252336 251175
rect 252284 251132 252336 251141
rect 324780 251107 324832 251116
rect 324780 251073 324789 251107
rect 324789 251073 324823 251107
rect 324823 251073 324832 251107
rect 324780 251064 324832 251073
rect 81716 250996 81768 251048
rect 81716 250860 81768 250912
rect 72148 249772 72200 249824
rect 72424 249772 72476 249824
rect 92664 249772 92716 249824
rect 92848 249772 92900 249824
rect 193680 249772 193732 249824
rect 193864 249772 193916 249824
rect 243636 249772 243688 249824
rect 243820 249772 243872 249824
rect 246948 249772 247000 249824
rect 247132 249772 247184 249824
rect 78772 248412 78824 248464
rect 78956 248412 79008 248464
rect 77668 244944 77720 244996
rect 77852 244944 77904 244996
rect 94136 244944 94188 244996
rect 268752 244672 268804 244724
rect 269028 244672 269080 244724
rect 70676 244332 70728 244384
rect 70492 244264 70544 244316
rect 84476 244264 84528 244316
rect 84660 244264 84712 244316
rect 211804 244264 211856 244316
rect 211988 244264 212040 244316
rect 227260 244264 227312 244316
rect 227444 244264 227496 244316
rect 268660 244264 268712 244316
rect 268844 244264 268896 244316
rect 324872 241544 324924 241596
rect 70768 241519 70820 241528
rect 70768 241485 70777 241519
rect 70777 241485 70811 241519
rect 70811 241485 70820 241519
rect 70768 241476 70820 241485
rect 73712 241476 73764 241528
rect 81716 241476 81768 241528
rect 105084 241519 105136 241528
rect 105084 241485 105093 241519
rect 105093 241485 105127 241519
rect 105127 241485 105136 241519
rect 105084 241476 105136 241485
rect 252284 241519 252336 241528
rect 252284 241485 252293 241519
rect 252293 241485 252327 241519
rect 252327 241485 252336 241519
rect 252284 241476 252336 241485
rect 81808 241408 81860 241460
rect 324872 241451 324924 241460
rect 324872 241417 324881 241451
rect 324881 241417 324915 241451
rect 324915 241417 324924 241451
rect 324872 241408 324924 241417
rect 72240 240116 72292 240168
rect 72424 240116 72476 240168
rect 78772 240116 78824 240168
rect 234068 240116 234120 240168
rect 234160 240116 234212 240168
rect 242348 240116 242400 240168
rect 242532 240116 242584 240168
rect 255228 240116 255280 240168
rect 255320 240116 255372 240168
rect 78864 240048 78916 240100
rect 268752 239436 268804 239488
rect 269028 239436 269080 239488
rect 81808 234608 81860 234660
rect 70492 234540 70544 234592
rect 70676 234540 70728 234592
rect 70768 234583 70820 234592
rect 70768 234549 70777 234583
rect 70777 234549 70811 234583
rect 70811 234549 70820 234583
rect 70768 234540 70820 234549
rect 95700 234608 95752 234660
rect 105084 234608 105136 234660
rect 234068 234608 234120 234660
rect 325056 234608 325108 234660
rect 95608 234540 95660 234592
rect 81808 234472 81860 234524
rect 105176 234472 105228 234524
rect 234160 234472 234212 234524
rect 70768 231863 70820 231872
rect 70768 231829 70777 231863
rect 70777 231829 70811 231863
rect 70811 231829 70820 231863
rect 70768 231820 70820 231829
rect 72148 231820 72200 231872
rect 72424 231820 72476 231872
rect 73436 231820 73488 231872
rect 73712 231820 73764 231872
rect 94136 231820 94188 231872
rect 150992 231820 151044 231872
rect 151084 231820 151136 231872
rect 89996 230460 90048 230512
rect 90180 230460 90232 230512
rect 90824 230460 90876 230512
rect 90916 230460 90968 230512
rect 193680 230460 193732 230512
rect 193864 230460 193916 230512
rect 243636 230460 243688 230512
rect 243820 230460 243872 230512
rect 246948 230460 247000 230512
rect 247132 230460 247184 230512
rect 250812 230460 250864 230512
rect 250996 230460 251048 230512
rect 252100 230460 252152 230512
rect 252284 230460 252336 230512
rect 255228 230460 255280 230512
rect 255320 230460 255372 230512
rect 259092 230460 259144 230512
rect 259276 230460 259328 230512
rect 265992 230503 266044 230512
rect 265992 230469 266001 230503
rect 266001 230469 266035 230503
rect 266035 230469 266044 230503
rect 265992 230460 266044 230469
rect 106556 230392 106608 230444
rect 268752 229712 268804 229764
rect 269028 229712 269080 229764
rect 78956 229032 79008 229084
rect 255228 229032 255280 229084
rect 255504 229032 255556 229084
rect 77760 225632 77812 225684
rect 70676 225020 70728 225072
rect 70492 224952 70544 225004
rect 84476 224952 84528 225004
rect 84660 224952 84712 225004
rect 94136 225020 94188 225072
rect 105084 224995 105136 225004
rect 105084 224961 105093 224995
rect 105093 224961 105127 224995
rect 105127 224961 105136 224995
rect 105084 224952 105136 224961
rect 211804 224952 211856 225004
rect 211988 224952 212040 225004
rect 227260 224952 227312 225004
rect 227444 224952 227496 225004
rect 234160 225020 234212 225072
rect 268660 224952 268712 225004
rect 268844 224952 268896 225004
rect 94044 224884 94096 224936
rect 234068 224884 234120 224936
rect 268752 224476 268804 224528
rect 269028 224476 269080 224528
rect 72148 222164 72200 222216
rect 72424 222164 72476 222216
rect 81716 222164 81768 222216
rect 81808 222164 81860 222216
rect 105084 222207 105136 222216
rect 105084 222173 105093 222207
rect 105093 222173 105127 222207
rect 105127 222173 105136 222207
rect 105084 222164 105136 222173
rect 324872 222164 324924 222216
rect 325148 222164 325200 222216
rect 106464 220915 106516 220924
rect 106464 220881 106473 220915
rect 106473 220881 106507 220915
rect 106507 220881 106516 220915
rect 106464 220872 106516 220881
rect 90640 220804 90692 220856
rect 91008 220804 91060 220856
rect 242348 220804 242400 220856
rect 242532 220804 242584 220856
rect 106464 220736 106516 220788
rect 106648 220736 106700 220788
rect 91008 220711 91060 220720
rect 91008 220677 91017 220711
rect 91017 220677 91051 220711
rect 91051 220677 91060 220711
rect 91008 220668 91060 220677
rect 78772 219487 78824 219496
rect 78772 219453 78781 219487
rect 78781 219453 78815 219487
rect 78815 219453 78824 219487
rect 78772 219444 78824 219453
rect 265992 218059 266044 218068
rect 265992 218025 266001 218059
rect 266001 218025 266035 218059
rect 266035 218025 266044 218059
rect 265992 218016 266044 218025
rect 77576 217336 77628 217388
rect 233792 216631 233844 216640
rect 233792 216597 233801 216631
rect 233801 216597 233835 216631
rect 233835 216597 233844 216631
rect 233792 216588 233844 216597
rect 95700 215296 95752 215348
rect 105084 215296 105136 215348
rect 70492 215228 70544 215280
rect 70676 215228 70728 215280
rect 70768 215271 70820 215280
rect 70768 215237 70777 215271
rect 70777 215237 70811 215271
rect 70811 215237 70820 215271
rect 70768 215228 70820 215237
rect 95608 215228 95660 215280
rect 325148 215364 325200 215416
rect 325056 215228 325108 215280
rect 105176 215160 105228 215212
rect 70768 212551 70820 212560
rect 70768 212517 70777 212551
rect 70777 212517 70811 212551
rect 70811 212517 70820 212551
rect 70768 212508 70820 212517
rect 72148 212508 72200 212560
rect 72424 212508 72476 212560
rect 73436 212508 73488 212560
rect 73712 212508 73764 212560
rect 94136 212508 94188 212560
rect 94320 212508 94372 212560
rect 150992 212508 151044 212560
rect 151084 212508 151136 212560
rect 91100 212440 91152 212492
rect 78680 211148 78732 211200
rect 78772 211148 78824 211200
rect 243728 211148 243780 211200
rect 243820 211148 243872 211200
rect 255320 211148 255372 211200
rect 91192 211080 91244 211132
rect 242348 211080 242400 211132
rect 242532 211080 242584 211132
rect 255596 211012 255648 211064
rect 268752 210400 268804 210452
rect 269028 210400 269080 210452
rect 235724 209720 235776 209772
rect 233792 208403 233844 208412
rect 233792 208369 233801 208403
rect 233801 208369 233835 208403
rect 233835 208369 233844 208403
rect 233792 208360 233844 208369
rect 255412 206184 255464 206236
rect 255596 206184 255648 206236
rect 70676 205708 70728 205760
rect 70492 205640 70544 205692
rect 77484 205683 77536 205692
rect 77484 205649 77493 205683
rect 77493 205649 77527 205683
rect 77527 205649 77536 205683
rect 77484 205640 77536 205649
rect 84476 205640 84528 205692
rect 84660 205640 84712 205692
rect 89996 205640 90048 205692
rect 94136 205708 94188 205760
rect 105084 205683 105136 205692
rect 105084 205649 105093 205683
rect 105093 205649 105127 205683
rect 105127 205649 105136 205683
rect 105084 205640 105136 205649
rect 211804 205640 211856 205692
rect 211988 205640 212040 205692
rect 227260 205640 227312 205692
rect 227444 205640 227496 205692
rect 268660 205640 268712 205692
rect 268844 205640 268896 205692
rect 94044 205572 94096 205624
rect 90088 205504 90140 205556
rect 233792 203532 233844 203584
rect 234344 203532 234396 203584
rect 72148 202852 72200 202904
rect 72424 202852 72476 202904
rect 77484 202895 77536 202904
rect 77484 202861 77493 202895
rect 77493 202861 77527 202895
rect 77527 202861 77536 202895
rect 77484 202852 77536 202861
rect 105084 202895 105136 202904
rect 105084 202861 105093 202895
rect 105093 202861 105127 202895
rect 105127 202861 105136 202895
rect 105084 202852 105136 202861
rect 106556 202852 106608 202904
rect 106740 202852 106792 202904
rect 324872 202852 324924 202904
rect 325148 202852 325200 202904
rect 91008 202827 91060 202836
rect 91008 202793 91017 202827
rect 91017 202793 91051 202827
rect 91051 202793 91060 202827
rect 91008 202784 91060 202793
rect 94044 202827 94096 202836
rect 94044 202793 94053 202827
rect 94053 202793 94087 202827
rect 94087 202793 94096 202827
rect 94044 202784 94096 202793
rect 193680 201424 193732 201476
rect 193864 201424 193916 201476
rect 246948 201424 247000 201476
rect 247132 201424 247184 201476
rect 252284 201467 252336 201476
rect 252284 201433 252293 201467
rect 252293 201433 252327 201467
rect 252327 201433 252336 201467
rect 252284 201424 252336 201433
rect 268752 200948 268804 201000
rect 269028 200948 269080 201000
rect 235540 200175 235592 200184
rect 235540 200141 235549 200175
rect 235549 200141 235583 200175
rect 235583 200141 235592 200175
rect 235540 200132 235592 200141
rect 81716 195984 81768 196036
rect 70492 195916 70544 195968
rect 70676 195916 70728 195968
rect 70768 195959 70820 195968
rect 70768 195925 70777 195959
rect 70777 195925 70811 195959
rect 70811 195925 70820 195959
rect 95700 195984 95752 196036
rect 105084 195984 105136 196036
rect 106740 195984 106792 196036
rect 70768 195916 70820 195925
rect 81808 195916 81860 195968
rect 95608 195916 95660 195968
rect 325148 196052 325200 196104
rect 106832 195916 106884 195968
rect 325056 195916 325108 195968
rect 105176 195848 105228 195900
rect 92756 193264 92808 193316
rect 92940 193264 92992 193316
rect 70768 193239 70820 193248
rect 70768 193205 70777 193239
rect 70777 193205 70811 193239
rect 70811 193205 70820 193239
rect 70768 193196 70820 193205
rect 72148 193196 72200 193248
rect 72424 193196 72476 193248
rect 73436 193196 73488 193248
rect 73712 193196 73764 193248
rect 94136 193196 94188 193248
rect 150992 193196 151044 193248
rect 151084 193196 151136 193248
rect 264612 192559 264664 192568
rect 264612 192525 264621 192559
rect 264621 192525 264655 192559
rect 264655 192525 264664 192559
rect 264612 192516 264664 192525
rect 243728 191836 243780 191888
rect 243820 191836 243872 191888
rect 252284 191879 252336 191888
rect 252284 191845 252293 191879
rect 252293 191845 252327 191879
rect 252327 191845 252336 191879
rect 252284 191836 252336 191845
rect 72056 191768 72108 191820
rect 72148 191768 72200 191820
rect 73344 191768 73396 191820
rect 73436 191768 73488 191820
rect 242348 191768 242400 191820
rect 242532 191768 242584 191820
rect 268752 191088 268804 191140
rect 269028 191088 269080 191140
rect 255320 190476 255372 190528
rect 255412 190476 255464 190528
rect 260288 190408 260340 190460
rect 260472 190408 260524 190460
rect 70676 186396 70728 186448
rect 70492 186328 70544 186380
rect 77576 186396 77628 186448
rect 267280 186396 267332 186448
rect 78772 186371 78824 186380
rect 78772 186337 78781 186371
rect 78781 186337 78815 186371
rect 78815 186337 78824 186371
rect 78772 186328 78824 186337
rect 84476 186328 84528 186380
rect 84660 186328 84712 186380
rect 105084 186371 105136 186380
rect 105084 186337 105093 186371
rect 105093 186337 105127 186371
rect 105127 186337 105136 186371
rect 105084 186328 105136 186337
rect 211804 186328 211856 186380
rect 211988 186328 212040 186380
rect 227260 186328 227312 186380
rect 227444 186328 227496 186380
rect 267096 186328 267148 186380
rect 268660 186328 268712 186380
rect 268844 186328 268896 186380
rect 77484 186260 77536 186312
rect 264612 185691 264664 185700
rect 264612 185657 264621 185691
rect 264621 185657 264655 185691
rect 264655 185657 264664 185691
rect 264612 185648 264664 185657
rect 204904 183608 204956 183660
rect 78772 183583 78824 183592
rect 78772 183549 78781 183583
rect 78781 183549 78815 183583
rect 78815 183549 78824 183583
rect 78772 183540 78824 183549
rect 91008 183583 91060 183592
rect 91008 183549 91017 183583
rect 91017 183549 91051 183583
rect 91051 183549 91060 183583
rect 91008 183540 91060 183549
rect 105084 183583 105136 183592
rect 105084 183549 105093 183583
rect 105093 183549 105127 183583
rect 105127 183549 105136 183583
rect 105084 183540 105136 183549
rect 106648 183540 106700 183592
rect 106924 183540 106976 183592
rect 204720 183540 204772 183592
rect 324872 183540 324924 183592
rect 325148 183540 325200 183592
rect 77484 183515 77536 183524
rect 77484 183481 77493 183515
rect 77493 183481 77527 183515
rect 77527 183481 77536 183515
rect 77484 183472 77536 183481
rect 193680 182112 193732 182164
rect 193864 182112 193916 182164
rect 246948 182112 247000 182164
rect 247132 182112 247184 182164
rect 250812 182112 250864 182164
rect 250996 182112 251048 182164
rect 252100 182112 252152 182164
rect 252284 182112 252336 182164
rect 259092 182112 259144 182164
rect 259276 182112 259328 182164
rect 268752 181432 268804 181484
rect 269028 181432 269080 181484
rect 265992 180956 266044 181008
rect 91008 180863 91060 180872
rect 91008 180829 91017 180863
rect 91017 180829 91051 180863
rect 91051 180829 91060 180863
rect 91008 180820 91060 180829
rect 265992 180820 266044 180872
rect 235724 180752 235776 180804
rect 265992 179367 266044 179376
rect 265992 179333 266001 179367
rect 266001 179333 266035 179367
rect 266035 179333 266044 179367
rect 265992 179324 266044 179333
rect 267280 179367 267332 179376
rect 267280 179333 267289 179367
rect 267289 179333 267323 179367
rect 267323 179333 267332 179367
rect 267280 179324 267332 179333
rect 91008 178687 91060 178696
rect 91008 178653 91017 178687
rect 91017 178653 91051 178687
rect 91051 178653 91060 178687
rect 91008 178644 91060 178653
rect 95516 176672 95568 176724
rect 105084 176672 105136 176724
rect 70492 176604 70544 176656
rect 70676 176604 70728 176656
rect 70768 176647 70820 176656
rect 70768 176613 70777 176647
rect 70777 176613 70811 176647
rect 70811 176613 70820 176647
rect 70768 176604 70820 176613
rect 95608 176604 95660 176656
rect 325148 176740 325200 176792
rect 325056 176604 325108 176656
rect 105176 176536 105228 176588
rect 72332 174063 72384 174072
rect 72332 174029 72341 174063
rect 72341 174029 72375 174063
rect 72375 174029 72384 174063
rect 72332 174020 72384 174029
rect 89996 173952 90048 174004
rect 90180 173952 90232 174004
rect 70768 173927 70820 173936
rect 70768 173893 70777 173927
rect 70777 173893 70811 173927
rect 70811 173893 70820 173927
rect 70768 173884 70820 173893
rect 73436 173884 73488 173936
rect 73620 173884 73672 173936
rect 77576 173884 77628 173936
rect 78772 173884 78824 173936
rect 78864 173884 78916 173936
rect 81808 173884 81860 173936
rect 81900 173884 81952 173936
rect 94136 173884 94188 173936
rect 94228 173884 94280 173936
rect 106740 173884 106792 173936
rect 106924 173884 106976 173936
rect 150992 173884 151044 173936
rect 151084 173884 151136 173936
rect 204720 173884 204772 173936
rect 204904 173884 204956 173936
rect 211712 173884 211764 173936
rect 211988 173884 212040 173936
rect 227168 173884 227220 173936
rect 227444 173884 227496 173936
rect 243728 172524 243780 172576
rect 243820 172524 243872 172576
rect 73344 172456 73396 172508
rect 73436 172456 73488 172508
rect 94136 172456 94188 172508
rect 94320 172456 94372 172508
rect 242532 172499 242584 172508
rect 242532 172465 242541 172499
rect 242541 172465 242575 172499
rect 242575 172465 242584 172499
rect 242532 172456 242584 172465
rect 243820 172388 243872 172440
rect 243912 172388 243964 172440
rect 268752 171572 268804 171624
rect 269028 171572 269080 171624
rect 72332 171139 72384 171148
rect 72332 171105 72341 171139
rect 72341 171105 72375 171139
rect 72375 171105 72384 171139
rect 72332 171096 72384 171105
rect 91192 171096 91244 171148
rect 235632 171139 235684 171148
rect 235632 171105 235641 171139
rect 235641 171105 235675 171139
rect 235675 171105 235684 171139
rect 235632 171096 235684 171105
rect 255320 171096 255372 171148
rect 255412 171096 255464 171148
rect 265992 169779 266044 169788
rect 265992 169745 266001 169779
rect 266001 169745 266035 169779
rect 266035 169745 266044 169779
rect 265992 169736 266044 169745
rect 267280 169779 267332 169788
rect 267280 169745 267289 169779
rect 267289 169745 267323 169779
rect 267323 169745 267332 169779
rect 267280 169736 267332 169745
rect 264612 169711 264664 169720
rect 264612 169677 264621 169711
rect 264621 169677 264655 169711
rect 264655 169677 264664 169711
rect 264612 169668 264664 169677
rect 104900 169056 104952 169108
rect 105084 169056 105136 169108
rect 77392 167628 77444 167680
rect 77576 167628 77628 167680
rect 78680 167628 78732 167680
rect 78864 167628 78916 167680
rect 81808 167628 81860 167680
rect 81992 167628 82044 167680
rect 70676 167084 70728 167136
rect 70492 167016 70544 167068
rect 84476 167016 84528 167068
rect 84660 167016 84712 167068
rect 211804 167016 211856 167068
rect 211988 167016 212040 167068
rect 227260 167016 227312 167068
rect 227444 167016 227496 167068
rect 324872 166948 324924 167000
rect 325056 166948 325108 167000
rect 106648 164203 106700 164212
rect 106648 164169 106657 164203
rect 106657 164169 106691 164203
rect 106691 164169 106700 164203
rect 106648 164160 106700 164169
rect 151084 164203 151136 164212
rect 151084 164169 151093 164203
rect 151093 164169 151127 164203
rect 151127 164169 151136 164203
rect 151084 164160 151136 164169
rect 211896 164203 211948 164212
rect 211896 164169 211905 164203
rect 211905 164169 211939 164203
rect 211939 164169 211948 164203
rect 211896 164160 211948 164169
rect 227352 164203 227404 164212
rect 227352 164169 227361 164203
rect 227361 164169 227395 164203
rect 227395 164169 227404 164203
rect 227352 164160 227404 164169
rect 204812 164092 204864 164144
rect 204904 164092 204956 164144
rect 242532 162911 242584 162920
rect 242532 162877 242541 162911
rect 242541 162877 242575 162911
rect 242575 162877 242584 162911
rect 242532 162868 242584 162877
rect 193864 162843 193916 162852
rect 193864 162809 193873 162843
rect 193873 162809 193907 162843
rect 193907 162809 193916 162843
rect 193864 162800 193916 162809
rect 234160 162800 234212 162852
rect 234344 162800 234396 162852
rect 250812 162800 250864 162852
rect 250996 162800 251048 162852
rect 252100 162800 252152 162852
rect 252284 162800 252336 162852
rect 259092 162800 259144 162852
rect 259276 162800 259328 162852
rect 268752 162324 268804 162376
rect 269028 162324 269080 162376
rect 81900 161415 81952 161424
rect 81900 161381 81909 161415
rect 81909 161381 81943 161415
rect 81943 161381 81952 161415
rect 81900 161372 81952 161381
rect 234160 161415 234212 161424
rect 234160 161381 234169 161415
rect 234169 161381 234203 161415
rect 234203 161381 234212 161415
rect 234160 161372 234212 161381
rect 243820 161415 243872 161424
rect 243820 161381 243829 161415
rect 243829 161381 243863 161415
rect 243863 161381 243872 161415
rect 243820 161372 243872 161381
rect 264612 160123 264664 160132
rect 264612 160089 264621 160123
rect 264621 160089 264655 160123
rect 264655 160089 264664 160123
rect 264612 160080 264664 160089
rect 265992 160055 266044 160064
rect 265992 160021 266001 160055
rect 266001 160021 266035 160055
rect 266035 160021 266044 160055
rect 265992 160012 266044 160021
rect 267280 160055 267332 160064
rect 267280 160021 267289 160055
rect 267289 160021 267323 160055
rect 267323 160021 267332 160055
rect 267280 160012 267332 160021
rect 70768 157428 70820 157480
rect 89996 157428 90048 157480
rect 105084 157360 105136 157412
rect 70492 157292 70544 157344
rect 70768 157292 70820 157344
rect 89996 157292 90048 157344
rect 106648 157335 106700 157344
rect 106648 157301 106657 157335
rect 106657 157301 106691 157335
rect 106691 157301 106700 157335
rect 106648 157292 106700 157301
rect 211896 157335 211948 157344
rect 211896 157301 211905 157335
rect 211905 157301 211939 157335
rect 211939 157301 211948 157335
rect 211896 157292 211948 157301
rect 227352 157335 227404 157344
rect 227352 157301 227361 157335
rect 227361 157301 227395 157335
rect 227395 157301 227404 157335
rect 227352 157292 227404 157301
rect 325148 157428 325200 157480
rect 105176 157224 105228 157276
rect 325056 157224 325108 157276
rect 94136 156612 94188 156664
rect 70676 154615 70728 154624
rect 70676 154581 70685 154615
rect 70685 154581 70719 154615
rect 70719 154581 70728 154615
rect 70676 154572 70728 154581
rect 73528 154572 73580 154624
rect 73620 154572 73672 154624
rect 151084 154615 151136 154624
rect 151084 154581 151093 154615
rect 151093 154581 151127 154615
rect 151127 154581 151136 154615
rect 151084 154572 151136 154581
rect 325056 154504 325108 154556
rect 325240 154504 325292 154556
rect 193864 153255 193916 153264
rect 193864 153221 193873 153255
rect 193873 153221 193907 153255
rect 193907 153221 193916 153255
rect 193864 153212 193916 153221
rect 73436 153187 73488 153196
rect 73436 153153 73445 153187
rect 73445 153153 73479 153187
rect 73479 153153 73488 153187
rect 73436 153144 73488 153153
rect 77484 153144 77536 153196
rect 78772 153144 78824 153196
rect 242532 153187 242584 153196
rect 242532 153153 242541 153187
rect 242541 153153 242575 153187
rect 242575 153153 242584 153187
rect 242532 153144 242584 153153
rect 77668 153008 77720 153060
rect 78956 153008 79008 153060
rect 268752 152464 268804 152516
rect 269028 152464 269080 152516
rect 72148 151784 72200 151836
rect 72332 151784 72384 151836
rect 234160 151827 234212 151836
rect 234160 151793 234169 151827
rect 234169 151793 234203 151827
rect 234203 151793 234212 151827
rect 234160 151784 234212 151793
rect 243820 151827 243872 151836
rect 243820 151793 243829 151827
rect 243829 151793 243863 151827
rect 243863 151793 243872 151827
rect 243820 151784 243872 151793
rect 264520 150424 264572 150476
rect 264612 150424 264664 150476
rect 265992 150467 266044 150476
rect 265992 150433 266001 150467
rect 266001 150433 266035 150467
rect 266035 150433 266044 150467
rect 265992 150424 266044 150433
rect 267280 150467 267332 150476
rect 267280 150433 267289 150467
rect 267289 150433 267323 150467
rect 267323 150433 267332 150467
rect 267280 150424 267332 150433
rect 70492 147636 70544 147688
rect 70768 147636 70820 147688
rect 84476 147636 84528 147688
rect 84660 147636 84712 147688
rect 105176 147704 105228 147756
rect 106556 147636 106608 147688
rect 106740 147636 106792 147688
rect 211804 147636 211856 147688
rect 211988 147636 212040 147688
rect 227260 147636 227312 147688
rect 227444 147636 227496 147688
rect 268660 147636 268712 147688
rect 268844 147636 268896 147688
rect 105084 147568 105136 147620
rect 94320 146956 94372 147008
rect 234160 144916 234212 144968
rect 73436 144891 73488 144900
rect 73436 144857 73445 144891
rect 73445 144857 73479 144891
rect 73479 144857 73488 144891
rect 73436 144848 73488 144857
rect 106648 144891 106700 144900
rect 106648 144857 106657 144891
rect 106657 144857 106691 144891
rect 106691 144857 106700 144891
rect 106648 144848 106700 144857
rect 151084 144891 151136 144900
rect 151084 144857 151093 144891
rect 151093 144857 151127 144891
rect 151127 144857 151136 144891
rect 151084 144848 151136 144857
rect 211896 144891 211948 144900
rect 211896 144857 211905 144891
rect 211905 144857 211939 144891
rect 211939 144857 211948 144891
rect 211896 144848 211948 144857
rect 227352 144891 227404 144900
rect 227352 144857 227361 144891
rect 227361 144857 227395 144891
rect 227395 144857 227404 144891
rect 227352 144848 227404 144857
rect 81900 144823 81952 144832
rect 81900 144789 81909 144823
rect 81909 144789 81943 144823
rect 81943 144789 81952 144823
rect 81900 144780 81952 144789
rect 204812 144780 204864 144832
rect 204904 144780 204956 144832
rect 234252 144780 234304 144832
rect 242532 143599 242584 143608
rect 242532 143565 242541 143599
rect 242541 143565 242575 143599
rect 242575 143565 242584 143599
rect 242532 143556 242584 143565
rect 243636 143556 243688 143608
rect 243820 143556 243872 143608
rect 72148 143488 72200 143540
rect 72332 143488 72384 143540
rect 81900 143488 81952 143540
rect 82084 143488 82136 143540
rect 105084 143531 105136 143540
rect 105084 143497 105093 143531
rect 105093 143497 105127 143531
rect 105127 143497 105136 143531
rect 105084 143488 105136 143497
rect 193864 143531 193916 143540
rect 193864 143497 193873 143531
rect 193873 143497 193907 143531
rect 193907 143497 193916 143531
rect 193864 143488 193916 143497
rect 246948 143488 247000 143540
rect 247132 143488 247184 143540
rect 248236 143488 248288 143540
rect 248420 143488 248472 143540
rect 249432 143488 249484 143540
rect 249616 143488 249668 143540
rect 250996 143488 251048 143540
rect 251180 143488 251232 143540
rect 252100 143488 252152 143540
rect 252284 143488 252336 143540
rect 259092 143488 259144 143540
rect 259276 143488 259328 143540
rect 264796 143488 264848 143540
rect 264980 143488 265032 143540
rect 73528 143463 73580 143472
rect 73528 143429 73537 143463
rect 73537 143429 73571 143463
rect 73571 143429 73580 143463
rect 73528 143420 73580 143429
rect 268752 142808 268804 142860
rect 269028 142808 269080 142860
rect 234252 142060 234304 142112
rect 264520 140768 264572 140820
rect 264612 140768 264664 140820
rect 265992 140743 266044 140752
rect 265992 140709 266001 140743
rect 266001 140709 266035 140743
rect 266035 140709 266044 140743
rect 265992 140700 266044 140709
rect 267280 140743 267332 140752
rect 267280 140709 267289 140743
rect 267289 140709 267323 140743
rect 267323 140709 267332 140743
rect 267280 140700 267332 140709
rect 324964 137980 325016 138032
rect 105084 137955 105136 137964
rect 105084 137921 105093 137955
rect 105093 137921 105127 137955
rect 105127 137921 105136 137955
rect 105084 137912 105136 137921
rect 106648 137955 106700 137964
rect 106648 137921 106657 137955
rect 106657 137921 106691 137955
rect 106691 137921 106700 137955
rect 106648 137912 106700 137921
rect 211896 137955 211948 137964
rect 211896 137921 211905 137955
rect 211905 137921 211939 137955
rect 211939 137921 211948 137955
rect 211896 137912 211948 137921
rect 227352 137955 227404 137964
rect 227352 137921 227361 137955
rect 227361 137921 227395 137955
rect 227395 137921 227404 137955
rect 227352 137912 227404 137921
rect 325056 137912 325108 137964
rect 151084 135303 151136 135312
rect 151084 135269 151093 135303
rect 151093 135269 151127 135303
rect 151127 135269 151136 135303
rect 151084 135260 151136 135269
rect 325056 135192 325108 135244
rect 325240 135192 325292 135244
rect 91008 133900 91060 133952
rect 91192 133900 91244 133952
rect 193864 133943 193916 133952
rect 193864 133909 193873 133943
rect 193873 133909 193907 133943
rect 193907 133909 193916 133943
rect 193864 133900 193916 133909
rect 243636 133900 243688 133952
rect 243820 133900 243872 133952
rect 72332 133875 72384 133884
rect 72332 133841 72341 133875
rect 72341 133841 72375 133875
rect 72375 133841 72384 133875
rect 72332 133832 72384 133841
rect 242532 133875 242584 133884
rect 242532 133841 242541 133875
rect 242541 133841 242575 133875
rect 242575 133841 242584 133875
rect 242532 133832 242584 133841
rect 243820 133807 243872 133816
rect 243820 133773 243829 133807
rect 243829 133773 243863 133807
rect 243863 133773 243872 133807
rect 243820 133764 243872 133773
rect 268752 133152 268804 133204
rect 269028 133152 269080 133204
rect 73620 131520 73672 131572
rect 264520 131112 264572 131164
rect 264612 131112 264664 131164
rect 265992 131155 266044 131164
rect 265992 131121 266001 131155
rect 266001 131121 266035 131155
rect 266035 131121 266044 131155
rect 265992 131112 266044 131121
rect 267280 131155 267332 131164
rect 267280 131121 267289 131155
rect 267289 131121 267323 131155
rect 267323 131121 267332 131155
rect 267280 131112 267332 131121
rect 70676 128392 70728 128444
rect 70768 128392 70820 128444
rect 70492 128324 70544 128376
rect 70584 128256 70636 128308
rect 84476 128324 84528 128376
rect 84660 128324 84712 128376
rect 105176 128392 105228 128444
rect 211804 128324 211856 128376
rect 211988 128324 212040 128376
rect 227260 128324 227312 128376
rect 227444 128324 227496 128376
rect 268660 128324 268712 128376
rect 268844 128324 268896 128376
rect 105084 128256 105136 128308
rect 70492 125536 70544 125588
rect 70676 125536 70728 125588
rect 90088 125536 90140 125588
rect 90180 125536 90232 125588
rect 92848 125536 92900 125588
rect 92940 125536 92992 125588
rect 151084 125579 151136 125588
rect 151084 125545 151093 125579
rect 151093 125545 151127 125579
rect 151127 125545 151136 125579
rect 151084 125536 151136 125545
rect 211896 125579 211948 125588
rect 211896 125545 211905 125579
rect 211905 125545 211939 125579
rect 211939 125545 211948 125579
rect 211896 125536 211948 125545
rect 227352 125579 227404 125588
rect 227352 125545 227361 125579
rect 227361 125545 227395 125579
rect 227395 125545 227404 125579
rect 227352 125536 227404 125545
rect 70584 125468 70636 125520
rect 70768 125468 70820 125520
rect 72332 124219 72384 124228
rect 72332 124185 72341 124219
rect 72341 124185 72375 124219
rect 72375 124185 72384 124219
rect 72332 124176 72384 124185
rect 106464 124176 106516 124228
rect 106740 124176 106792 124228
rect 234252 124176 234304 124228
rect 242532 124219 242584 124228
rect 242532 124185 242541 124219
rect 242541 124185 242575 124219
rect 242575 124185 242584 124219
rect 242532 124176 242584 124185
rect 243820 124219 243872 124228
rect 243820 124185 243829 124219
rect 243829 124185 243863 124219
rect 243863 124185 243872 124219
rect 243820 124176 243872 124185
rect 70768 124108 70820 124160
rect 70860 124108 70912 124160
rect 91008 124108 91060 124160
rect 91192 124108 91244 124160
rect 105084 124151 105136 124160
rect 105084 124117 105093 124151
rect 105093 124117 105127 124151
rect 105127 124117 105136 124151
rect 105084 124108 105136 124117
rect 193864 124151 193916 124160
rect 193864 124117 193873 124151
rect 193873 124117 193907 124151
rect 193907 124117 193916 124151
rect 193864 124108 193916 124117
rect 252284 124151 252336 124160
rect 252284 124117 252293 124151
rect 252293 124117 252327 124151
rect 252327 124117 252336 124151
rect 252284 124108 252336 124117
rect 255228 124151 255280 124160
rect 255228 124117 255237 124151
rect 255237 124117 255271 124151
rect 255271 124117 255280 124151
rect 255228 124108 255280 124117
rect 106464 124083 106516 124092
rect 106464 124049 106473 124083
rect 106473 124049 106507 124083
rect 106507 124049 106516 124083
rect 106464 124040 106516 124049
rect 268752 123496 268804 123548
rect 269028 123496 269080 123548
rect 243820 122791 243872 122800
rect 243820 122757 243829 122791
rect 243829 122757 243863 122791
rect 243863 122757 243872 122791
rect 243820 122748 243872 122757
rect 268660 122791 268712 122800
rect 268660 122757 268669 122791
rect 268669 122757 268703 122791
rect 268703 122757 268712 122791
rect 268660 122748 268712 122757
rect 264520 121456 264572 121508
rect 264612 121456 264664 121508
rect 265992 121431 266044 121440
rect 265992 121397 266001 121431
rect 266001 121397 266035 121431
rect 266035 121397 266044 121431
rect 265992 121388 266044 121397
rect 267280 121388 267332 121440
rect 234252 119391 234304 119400
rect 234252 119357 234261 119391
rect 234261 119357 234295 119391
rect 234295 119357 234304 119391
rect 234252 119348 234304 119357
rect 95608 118736 95660 118788
rect 324964 118668 325016 118720
rect 95608 118600 95660 118652
rect 211896 118643 211948 118652
rect 211896 118609 211905 118643
rect 211905 118609 211939 118643
rect 211939 118609 211948 118643
rect 211896 118600 211948 118609
rect 227352 118643 227404 118652
rect 227352 118609 227361 118643
rect 227361 118609 227395 118643
rect 227395 118609 227404 118643
rect 227352 118600 227404 118609
rect 325056 118600 325108 118652
rect 94044 118396 94096 118448
rect 94136 118328 94188 118380
rect 151084 115991 151136 116000
rect 151084 115957 151093 115991
rect 151093 115957 151127 115991
rect 151127 115957 151136 115991
rect 151084 115948 151136 115957
rect 204904 115948 204956 116000
rect 205088 115948 205140 116000
rect 78864 115880 78916 115932
rect 89996 115880 90048 115932
rect 90180 115880 90232 115932
rect 92756 115880 92808 115932
rect 92940 115880 92992 115932
rect 325056 115880 325108 115932
rect 325240 115880 325292 115932
rect 106556 114588 106608 114640
rect 234068 114588 234120 114640
rect 72148 114520 72200 114572
rect 72240 114520 72292 114572
rect 73436 114520 73488 114572
rect 73528 114520 73580 114572
rect 105176 114520 105228 114572
rect 193864 114563 193916 114572
rect 193864 114529 193873 114563
rect 193873 114529 193907 114563
rect 193907 114529 193916 114563
rect 193864 114520 193916 114529
rect 252284 114563 252336 114572
rect 252284 114529 252293 114563
rect 252293 114529 252327 114563
rect 252327 114529 252336 114563
rect 252284 114520 252336 114529
rect 259092 114520 259144 114572
rect 259276 114520 259328 114572
rect 90916 114495 90968 114504
rect 90916 114461 90925 114495
rect 90925 114461 90959 114495
rect 90959 114461 90968 114495
rect 90916 114452 90968 114461
rect 234160 114495 234212 114504
rect 234160 114461 234169 114495
rect 234169 114461 234203 114495
rect 234203 114461 234212 114495
rect 234160 114452 234212 114461
rect 242532 114495 242584 114504
rect 242532 114461 242541 114495
rect 242541 114461 242575 114495
rect 242575 114461 242584 114495
rect 242532 114452 242584 114461
rect 268752 113840 268804 113892
rect 269028 113840 269080 113892
rect 243820 113203 243872 113212
rect 243820 113169 243829 113203
rect 243829 113169 243863 113203
rect 243863 113169 243872 113203
rect 243820 113160 243872 113169
rect 268844 113160 268896 113212
rect 264520 111800 264572 111852
rect 264612 111800 264664 111852
rect 265992 111843 266044 111852
rect 265992 111809 266001 111843
rect 266001 111809 266035 111843
rect 266035 111809 266044 111843
rect 265992 111800 266044 111809
rect 267280 111800 267332 111852
rect 264612 111707 264664 111716
rect 264612 111673 264621 111707
rect 264621 111673 264655 111707
rect 264655 111673 264664 111707
rect 264612 111664 264664 111673
rect 70676 109080 70728 109132
rect 70492 109012 70544 109064
rect 77576 109080 77628 109132
rect 81808 109080 81860 109132
rect 84476 109012 84528 109064
rect 84660 109012 84712 109064
rect 105176 109080 105228 109132
rect 106556 109080 106608 109132
rect 211804 109012 211856 109064
rect 211988 109012 212040 109064
rect 227260 109012 227312 109064
rect 227444 109012 227496 109064
rect 268660 109012 268712 109064
rect 268844 109012 268896 109064
rect 77484 108944 77536 108996
rect 81716 108944 81768 108996
rect 105084 108944 105136 108996
rect 106556 108944 106608 108996
rect 268752 108536 268804 108588
rect 269028 108536 269080 108588
rect 78772 106335 78824 106344
rect 78772 106301 78781 106335
rect 78781 106301 78815 106335
rect 78815 106301 78824 106335
rect 78772 106292 78824 106301
rect 204720 106292 204772 106344
rect 204904 106292 204956 106344
rect 255228 106335 255280 106344
rect 255228 106301 255237 106335
rect 255237 106301 255271 106335
rect 255271 106301 255280 106335
rect 255228 106292 255280 106301
rect 72240 106267 72292 106276
rect 72240 106233 72249 106267
rect 72249 106233 72283 106267
rect 72283 106233 72292 106267
rect 72240 106224 72292 106233
rect 73528 106267 73580 106276
rect 73528 106233 73537 106267
rect 73537 106233 73571 106267
rect 73571 106233 73580 106267
rect 73528 106224 73580 106233
rect 151084 106267 151136 106276
rect 151084 106233 151093 106267
rect 151093 106233 151127 106267
rect 151127 106233 151136 106267
rect 151084 106224 151136 106233
rect 211896 106267 211948 106276
rect 211896 106233 211905 106267
rect 211905 106233 211939 106267
rect 211939 106233 211948 106267
rect 211896 106224 211948 106233
rect 227352 106267 227404 106276
rect 227352 106233 227361 106267
rect 227361 106233 227395 106267
rect 227395 106233 227404 106267
rect 227352 106224 227404 106233
rect 243820 104932 243872 104984
rect 91008 104864 91060 104916
rect 234252 104864 234304 104916
rect 242532 104907 242584 104916
rect 242532 104873 242541 104907
rect 242541 104873 242575 104907
rect 242575 104873 242584 104907
rect 242532 104864 242584 104873
rect 243636 104864 243688 104916
rect 70860 104796 70912 104848
rect 94044 104839 94096 104848
rect 94044 104805 94053 104839
rect 94053 104805 94087 104839
rect 94087 104805 94096 104839
rect 94044 104796 94096 104805
rect 105084 104839 105136 104848
rect 105084 104805 105093 104839
rect 105093 104805 105127 104839
rect 105127 104805 105136 104839
rect 105084 104796 105136 104805
rect 193864 104839 193916 104848
rect 193864 104805 193873 104839
rect 193873 104805 193907 104839
rect 193907 104805 193916 104839
rect 193864 104796 193916 104805
rect 246948 104839 247000 104848
rect 246948 104805 246957 104839
rect 246957 104805 246991 104839
rect 246991 104805 247000 104839
rect 246948 104796 247000 104805
rect 252284 104796 252336 104848
rect 255228 104839 255280 104848
rect 255228 104805 255237 104839
rect 255237 104805 255271 104839
rect 255271 104805 255280 104839
rect 255228 104796 255280 104805
rect 259276 104839 259328 104848
rect 259276 104805 259285 104839
rect 259285 104805 259319 104839
rect 259319 104805 259328 104839
rect 259276 104796 259328 104805
rect 106648 103479 106700 103488
rect 106648 103445 106657 103479
rect 106657 103445 106691 103479
rect 106691 103445 106700 103479
rect 106648 103436 106700 103445
rect 268660 103436 268712 103488
rect 264612 102187 264664 102196
rect 264612 102153 264621 102187
rect 264621 102153 264655 102187
rect 264655 102153 264664 102187
rect 264612 102144 264664 102153
rect 265992 102119 266044 102128
rect 265992 102085 266001 102119
rect 266001 102085 266035 102119
rect 266035 102085 266044 102119
rect 265992 102076 266044 102085
rect 267280 102119 267332 102128
rect 267280 102085 267289 102119
rect 267289 102085 267323 102119
rect 267323 102085 267332 102119
rect 267280 102076 267332 102085
rect 324780 101396 324832 101448
rect 324964 101396 325016 101448
rect 234252 100036 234304 100088
rect 211896 99331 211948 99340
rect 211896 99297 211905 99331
rect 211905 99297 211939 99331
rect 211939 99297 211948 99331
rect 211896 99288 211948 99297
rect 227352 99331 227404 99340
rect 227352 99297 227361 99331
rect 227361 99297 227395 99331
rect 227395 99297 227404 99331
rect 227352 99288 227404 99297
rect 72240 96747 72292 96756
rect 72240 96713 72249 96747
rect 72249 96713 72283 96747
rect 72283 96713 72292 96747
rect 72240 96704 72292 96713
rect 151084 96679 151136 96688
rect 151084 96645 151093 96679
rect 151093 96645 151127 96679
rect 151127 96645 151136 96679
rect 151084 96636 151136 96645
rect 204720 96636 204772 96688
rect 204904 96636 204956 96688
rect 235724 96611 235776 96620
rect 235724 96577 235733 96611
rect 235733 96577 235767 96611
rect 235767 96577 235776 96611
rect 235724 96568 235776 96577
rect 70768 95319 70820 95328
rect 70768 95285 70777 95319
rect 70777 95285 70811 95319
rect 70811 95285 70820 95319
rect 70768 95276 70820 95285
rect 70492 95208 70544 95260
rect 70676 95208 70728 95260
rect 73620 95208 73672 95260
rect 91008 95208 91060 95260
rect 91100 95208 91152 95260
rect 94044 95251 94096 95260
rect 94044 95217 94053 95251
rect 94053 95217 94087 95251
rect 94087 95217 94096 95251
rect 94044 95208 94096 95217
rect 105176 95208 105228 95260
rect 193864 95251 193916 95260
rect 193864 95217 193873 95251
rect 193873 95217 193907 95251
rect 193907 95217 193916 95251
rect 193864 95208 193916 95217
rect 234160 95251 234212 95260
rect 234160 95217 234169 95251
rect 234169 95217 234203 95251
rect 234203 95217 234212 95251
rect 234160 95208 234212 95217
rect 243636 95208 243688 95260
rect 243820 95208 243872 95260
rect 246948 95251 247000 95260
rect 246948 95217 246957 95251
rect 246957 95217 246991 95251
rect 246991 95217 247000 95251
rect 246948 95208 247000 95217
rect 252100 95251 252152 95260
rect 252100 95217 252109 95251
rect 252109 95217 252143 95251
rect 252143 95217 252152 95251
rect 252100 95208 252152 95217
rect 259276 95251 259328 95260
rect 259276 95217 259285 95251
rect 259285 95217 259319 95251
rect 259319 95217 259328 95251
rect 259276 95208 259328 95217
rect 70768 95140 70820 95192
rect 70952 95140 71004 95192
rect 242532 95183 242584 95192
rect 242532 95149 242541 95183
rect 242541 95149 242575 95183
rect 242575 95149 242584 95183
rect 242532 95140 242584 95149
rect 268752 94324 268804 94376
rect 269028 94324 269080 94376
rect 106556 93848 106608 93900
rect 268568 93891 268620 93900
rect 268568 93857 268577 93891
rect 268577 93857 268611 93891
rect 268611 93857 268620 93891
rect 268568 93848 268620 93857
rect 78864 93780 78916 93832
rect 264520 92488 264572 92540
rect 264612 92488 264664 92540
rect 265992 92531 266044 92540
rect 265992 92497 266001 92531
rect 266001 92497 266035 92531
rect 266035 92497 266044 92531
rect 265992 92488 266044 92497
rect 267280 92531 267332 92540
rect 267280 92497 267289 92531
rect 267289 92497 267323 92531
rect 267323 92497 267332 92531
rect 267280 92488 267332 92497
rect 264612 92395 264664 92404
rect 264612 92361 264621 92395
rect 264621 92361 264655 92395
rect 264655 92361 264664 92395
rect 264612 92352 264664 92361
rect 234160 91783 234212 91792
rect 234160 91749 234169 91783
rect 234169 91749 234203 91783
rect 234203 91749 234212 91783
rect 234160 91740 234212 91749
rect 70676 89768 70728 89820
rect 70492 89700 70544 89752
rect 84476 89700 84528 89752
rect 84660 89700 84712 89752
rect 105176 89768 105228 89820
rect 106556 89768 106608 89820
rect 211804 89700 211856 89752
rect 211988 89700 212040 89752
rect 227260 89700 227312 89752
rect 227444 89700 227496 89752
rect 105084 89632 105136 89684
rect 234344 87048 234396 87100
rect 204720 86980 204772 87032
rect 204904 86980 204956 87032
rect 235724 87023 235776 87032
rect 235724 86989 235733 87023
rect 235733 86989 235767 87023
rect 235767 86989 235776 87023
rect 235724 86980 235776 86989
rect 255228 87023 255280 87032
rect 255228 86989 255237 87023
rect 255237 86989 255271 87023
rect 255271 86989 255280 87023
rect 255228 86980 255280 86989
rect 151084 86955 151136 86964
rect 151084 86921 151093 86955
rect 151093 86921 151127 86955
rect 151127 86921 151136 86955
rect 151084 86912 151136 86921
rect 211896 86955 211948 86964
rect 211896 86921 211905 86955
rect 211905 86921 211939 86955
rect 211939 86921 211948 86955
rect 211896 86912 211948 86921
rect 227352 86955 227404 86964
rect 227352 86921 227361 86955
rect 227361 86921 227395 86955
rect 227395 86921 227404 86955
rect 227352 86912 227404 86921
rect 89996 86887 90048 86896
rect 89996 86853 90005 86887
rect 90005 86853 90039 86887
rect 90039 86853 90048 86887
rect 89996 86844 90048 86853
rect 92756 86887 92808 86896
rect 92756 86853 92765 86887
rect 92765 86853 92799 86887
rect 92799 86853 92808 86887
rect 92756 86844 92808 86853
rect 106648 85595 106700 85604
rect 106648 85561 106657 85595
rect 106657 85561 106691 85595
rect 106691 85561 106700 85595
rect 106648 85552 106700 85561
rect 242532 85595 242584 85604
rect 242532 85561 242541 85595
rect 242541 85561 242575 85595
rect 242575 85561 242584 85595
rect 242532 85552 242584 85561
rect 72148 85527 72200 85536
rect 72148 85493 72157 85527
rect 72157 85493 72191 85527
rect 72191 85493 72200 85527
rect 72148 85484 72200 85493
rect 73436 85527 73488 85536
rect 73436 85493 73445 85527
rect 73445 85493 73479 85527
rect 73479 85493 73488 85527
rect 73436 85484 73488 85493
rect 77484 85527 77536 85536
rect 77484 85493 77493 85527
rect 77493 85493 77527 85527
rect 77527 85493 77536 85527
rect 77484 85484 77536 85493
rect 81716 85527 81768 85536
rect 81716 85493 81725 85527
rect 81725 85493 81759 85527
rect 81759 85493 81768 85527
rect 81716 85484 81768 85493
rect 94044 85527 94096 85536
rect 94044 85493 94053 85527
rect 94053 85493 94087 85527
rect 94087 85493 94096 85527
rect 94044 85484 94096 85493
rect 105084 85527 105136 85536
rect 105084 85493 105093 85527
rect 105093 85493 105127 85527
rect 105127 85493 105136 85527
rect 105084 85484 105136 85493
rect 193864 85527 193916 85536
rect 193864 85493 193873 85527
rect 193873 85493 193907 85527
rect 193907 85493 193916 85527
rect 193864 85484 193916 85493
rect 204720 85527 204772 85536
rect 204720 85493 204729 85527
rect 204729 85493 204763 85527
rect 204763 85493 204772 85527
rect 204720 85484 204772 85493
rect 234252 85484 234304 85536
rect 246948 85527 247000 85536
rect 246948 85493 246957 85527
rect 246957 85493 246991 85527
rect 246991 85493 247000 85527
rect 246948 85484 247000 85493
rect 252284 85527 252336 85536
rect 252284 85493 252293 85527
rect 252293 85493 252327 85527
rect 252327 85493 252336 85527
rect 252284 85484 252336 85493
rect 255228 85527 255280 85536
rect 255228 85493 255237 85527
rect 255237 85493 255271 85527
rect 255271 85493 255280 85527
rect 255228 85484 255280 85493
rect 259276 85527 259328 85536
rect 259276 85493 259285 85527
rect 259285 85493 259319 85527
rect 259319 85493 259328 85527
rect 259276 85484 259328 85493
rect 268752 84872 268804 84924
rect 269028 84872 269080 84924
rect 78680 84303 78732 84312
rect 78680 84269 78689 84303
rect 78689 84269 78723 84303
rect 78723 84269 78732 84303
rect 78680 84260 78732 84269
rect 78680 84124 78732 84176
rect 78864 84056 78916 84108
rect 104992 84056 105044 84108
rect 264612 82875 264664 82884
rect 264612 82841 264621 82875
rect 264621 82841 264655 82875
rect 264655 82841 264664 82875
rect 264612 82832 264664 82841
rect 78864 82764 78916 82816
rect 265992 82807 266044 82816
rect 265992 82773 266001 82807
rect 266001 82773 266035 82807
rect 266035 82773 266044 82807
rect 265992 82764 266044 82773
rect 267280 82807 267332 82816
rect 267280 82773 267289 82807
rect 267289 82773 267323 82807
rect 267323 82773 267332 82807
rect 267280 82764 267332 82773
rect 94320 80928 94372 80980
rect 324964 80044 325016 80096
rect 325056 79908 325108 79960
rect 89996 77299 90048 77308
rect 89996 77265 90005 77299
rect 90005 77265 90039 77299
rect 90039 77265 90048 77299
rect 89996 77256 90048 77265
rect 92756 77299 92808 77308
rect 92756 77265 92765 77299
rect 92765 77265 92799 77299
rect 92799 77265 92808 77299
rect 92756 77256 92808 77265
rect 151084 77299 151136 77308
rect 151084 77265 151093 77299
rect 151093 77265 151127 77299
rect 151127 77265 151136 77299
rect 151084 77256 151136 77265
rect 211988 77256 212040 77308
rect 227444 77256 227496 77308
rect 93860 77188 93912 77240
rect 93952 77188 94004 77240
rect 235724 77231 235776 77240
rect 235724 77197 235733 77231
rect 235733 77197 235767 77231
rect 235767 77197 235776 77231
rect 235724 77188 235776 77197
rect 325056 77188 325108 77240
rect 93952 77052 94004 77104
rect 93860 76984 93912 77036
rect 72148 75939 72200 75948
rect 72148 75905 72157 75939
rect 72157 75905 72191 75939
rect 72191 75905 72200 75939
rect 72148 75896 72200 75905
rect 73528 75896 73580 75948
rect 77576 75896 77628 75948
rect 81808 75896 81860 75948
rect 193864 75939 193916 75948
rect 193864 75905 193873 75939
rect 193873 75905 193907 75939
rect 193907 75905 193916 75939
rect 193864 75896 193916 75905
rect 204904 75896 204956 75948
rect 234160 75939 234212 75948
rect 234160 75905 234169 75939
rect 234169 75905 234203 75939
rect 234203 75905 234212 75939
rect 234160 75896 234212 75905
rect 243636 75896 243688 75948
rect 243820 75896 243872 75948
rect 246948 75939 247000 75948
rect 246948 75905 246957 75939
rect 246957 75905 246991 75939
rect 246991 75905 247000 75939
rect 246948 75896 247000 75905
rect 252284 75939 252336 75948
rect 252284 75905 252293 75939
rect 252293 75905 252327 75939
rect 252327 75905 252336 75939
rect 252284 75896 252336 75905
rect 255228 75939 255280 75948
rect 255228 75905 255237 75939
rect 255237 75905 255271 75939
rect 255271 75905 255280 75939
rect 255228 75896 255280 75905
rect 259276 75939 259328 75948
rect 259276 75905 259285 75939
rect 259285 75905 259319 75939
rect 259319 75905 259328 75939
rect 259276 75896 259328 75905
rect 106556 75828 106608 75880
rect 211988 75828 212040 75880
rect 242532 75871 242584 75880
rect 242532 75837 242541 75871
rect 242541 75837 242575 75871
rect 242575 75837 242584 75871
rect 242532 75828 242584 75837
rect 268752 75080 268804 75132
rect 269028 75080 269080 75132
rect 104992 74579 105044 74588
rect 104992 74545 105001 74579
rect 105001 74545 105035 74579
rect 105035 74545 105044 74579
rect 104992 74536 105044 74545
rect 94320 74468 94372 74520
rect 264520 73176 264572 73228
rect 264612 73176 264664 73228
rect 265992 73219 266044 73228
rect 265992 73185 266001 73219
rect 266001 73185 266035 73219
rect 266035 73185 266044 73219
rect 265992 73176 266044 73185
rect 267280 73219 267332 73228
rect 267280 73185 267289 73219
rect 267289 73185 267323 73219
rect 267323 73185 267332 73219
rect 267280 73176 267332 73185
rect 72148 72471 72200 72480
rect 72148 72437 72157 72471
rect 72157 72437 72191 72471
rect 72191 72437 72200 72471
rect 72148 72428 72200 72437
rect 70492 71408 70544 71460
rect 70676 71408 70728 71460
rect 70768 70456 70820 70508
rect 77576 70456 77628 70508
rect 81808 70456 81860 70508
rect 268660 70388 268712 70440
rect 268844 70388 268896 70440
rect 70676 70320 70728 70372
rect 77484 70320 77536 70372
rect 81808 70320 81860 70372
rect 211896 70363 211948 70372
rect 211896 70329 211905 70363
rect 211905 70329 211939 70363
rect 211939 70329 211948 70363
rect 211896 70320 211948 70329
rect 72148 67711 72200 67720
rect 72148 67677 72157 67711
rect 72157 67677 72191 67711
rect 72191 67677 72200 67711
rect 72148 67668 72200 67677
rect 234068 67600 234120 67652
rect 234252 67600 234304 67652
rect 235724 67643 235776 67652
rect 235724 67609 235733 67643
rect 235733 67609 235767 67643
rect 235767 67609 235776 67643
rect 235724 67600 235776 67609
rect 324964 67643 325016 67652
rect 324964 67609 324973 67643
rect 324973 67609 325007 67643
rect 325007 67609 325016 67643
rect 324964 67600 325016 67609
rect 70676 67575 70728 67584
rect 70676 67541 70685 67575
rect 70685 67541 70719 67575
rect 70719 67541 70728 67575
rect 70676 67532 70728 67541
rect 89996 67575 90048 67584
rect 89996 67541 90005 67575
rect 90005 67541 90039 67575
rect 90039 67541 90048 67575
rect 89996 67532 90048 67541
rect 92756 67575 92808 67584
rect 92756 67541 92765 67575
rect 92765 67541 92799 67575
rect 92799 67541 92808 67575
rect 92756 67532 92808 67541
rect 151084 67575 151136 67584
rect 151084 67541 151093 67575
rect 151093 67541 151127 67575
rect 151127 67541 151136 67575
rect 151084 67532 151136 67541
rect 70492 67124 70544 67176
rect 70676 67124 70728 67176
rect 91100 66308 91152 66360
rect 106464 66351 106516 66360
rect 106464 66317 106473 66351
rect 106473 66317 106507 66351
rect 106507 66317 106516 66351
rect 106464 66308 106516 66317
rect 84568 66240 84620 66292
rect 84660 66240 84712 66292
rect 91008 66240 91060 66292
rect 104992 66283 105044 66292
rect 104992 66249 105001 66283
rect 105001 66249 105035 66283
rect 105035 66249 105044 66283
rect 104992 66240 105044 66249
rect 242532 66283 242584 66292
rect 242532 66249 242541 66283
rect 242541 66249 242575 66283
rect 242575 66249 242584 66283
rect 242532 66240 242584 66249
rect 72148 66172 72200 66224
rect 77392 66172 77444 66224
rect 77484 66172 77536 66224
rect 106464 66172 106516 66224
rect 106556 66172 106608 66224
rect 193864 66215 193916 66224
rect 193864 66181 193873 66215
rect 193873 66181 193907 66215
rect 193907 66181 193916 66215
rect 193864 66172 193916 66181
rect 204904 66215 204956 66224
rect 204904 66181 204913 66215
rect 204913 66181 204947 66215
rect 204947 66181 204956 66215
rect 204904 66172 204956 66181
rect 234068 66215 234120 66224
rect 234068 66181 234077 66215
rect 234077 66181 234111 66215
rect 234111 66181 234120 66215
rect 234068 66172 234120 66181
rect 246948 66215 247000 66224
rect 246948 66181 246957 66215
rect 246957 66181 246991 66215
rect 246991 66181 247000 66215
rect 246948 66172 247000 66181
rect 252284 66215 252336 66224
rect 252284 66181 252293 66215
rect 252293 66181 252327 66215
rect 252327 66181 252336 66215
rect 252284 66172 252336 66181
rect 255228 66215 255280 66224
rect 255228 66181 255237 66215
rect 255237 66181 255271 66215
rect 255271 66181 255280 66215
rect 255228 66172 255280 66181
rect 259276 66215 259328 66224
rect 259276 66181 259285 66215
rect 259285 66181 259319 66215
rect 259319 66181 259328 66215
rect 259276 66172 259328 66181
rect 262036 66172 262088 66224
rect 262220 66172 262272 66224
rect 268752 65492 268804 65544
rect 269028 65492 269080 65544
rect 78680 64923 78732 64932
rect 78680 64889 78689 64923
rect 78689 64889 78723 64923
rect 78723 64889 78732 64923
rect 78680 64880 78732 64889
rect 94136 64923 94188 64932
rect 94136 64889 94145 64923
rect 94145 64889 94179 64923
rect 94179 64889 94188 64923
rect 94136 64880 94188 64889
rect 104992 64812 105044 64864
rect 105268 64812 105320 64864
rect 267280 63495 267332 63504
rect 267280 63461 267289 63495
rect 267289 63461 267323 63495
rect 267323 63461 267332 63495
rect 267280 63452 267332 63461
rect 78680 61412 78732 61464
rect 78956 61412 79008 61464
rect 94136 60027 94188 60036
rect 94136 59993 94145 60027
rect 94145 59993 94179 60027
rect 94179 59993 94188 60027
rect 94136 59984 94188 59993
rect 89996 58055 90048 58064
rect 89996 58021 90005 58055
rect 90005 58021 90039 58055
rect 90039 58021 90048 58055
rect 89996 58012 90048 58021
rect 92756 58055 92808 58064
rect 92756 58021 92765 58055
rect 92765 58021 92799 58055
rect 92799 58021 92808 58055
rect 92756 58012 92808 58021
rect 70768 57944 70820 57996
rect 151084 57987 151136 57996
rect 151084 57953 151093 57987
rect 151093 57953 151127 57987
rect 151127 57953 151136 57987
rect 151084 57944 151136 57953
rect 211988 57876 212040 57928
rect 227444 57876 227496 57928
rect 235724 57919 235776 57928
rect 235724 57885 235733 57919
rect 235733 57885 235767 57919
rect 235767 57885 235776 57919
rect 235724 57876 235776 57885
rect 234252 57808 234304 57860
rect 91008 56652 91060 56704
rect 72056 56627 72108 56636
rect 72056 56593 72065 56627
rect 72065 56593 72099 56627
rect 72099 56593 72108 56627
rect 72056 56584 72108 56593
rect 193864 56627 193916 56636
rect 193864 56593 193873 56627
rect 193873 56593 193907 56627
rect 193907 56593 193916 56627
rect 193864 56584 193916 56593
rect 204904 56627 204956 56636
rect 204904 56593 204913 56627
rect 204913 56593 204947 56627
rect 204947 56593 204956 56627
rect 204904 56584 204956 56593
rect 243636 56584 243688 56636
rect 243820 56584 243872 56636
rect 246948 56627 247000 56636
rect 246948 56593 246957 56627
rect 246957 56593 246991 56627
rect 246991 56593 247000 56627
rect 246948 56584 247000 56593
rect 252284 56627 252336 56636
rect 252284 56593 252293 56627
rect 252293 56593 252327 56627
rect 252327 56593 252336 56627
rect 252284 56584 252336 56593
rect 255228 56627 255280 56636
rect 255228 56593 255237 56627
rect 255237 56593 255271 56627
rect 255271 56593 255280 56627
rect 255228 56584 255280 56593
rect 259276 56627 259328 56636
rect 259276 56593 259285 56627
rect 259285 56593 259319 56627
rect 259319 56593 259328 56627
rect 259276 56584 259328 56593
rect 96988 56559 97040 56568
rect 96988 56525 96997 56559
rect 96997 56525 97031 56559
rect 97031 56525 97040 56559
rect 96988 56516 97040 56525
rect 242532 56559 242584 56568
rect 242532 56525 242541 56559
rect 242541 56525 242575 56559
rect 242575 56525 242584 56559
rect 242532 56516 242584 56525
rect 268752 55836 268804 55888
rect 269028 55836 269080 55888
rect 90916 55267 90968 55276
rect 90916 55233 90925 55267
rect 90925 55233 90959 55267
rect 90959 55233 90968 55267
rect 90916 55224 90968 55233
rect 267280 53839 267332 53848
rect 267280 53805 267289 53839
rect 267289 53805 267323 53839
rect 267323 53805 267332 53839
rect 267280 53796 267332 53805
rect 264612 53771 264664 53780
rect 264612 53737 264621 53771
rect 264621 53737 264655 53771
rect 264655 53737 264664 53771
rect 264612 53728 264664 53737
rect 70492 53116 70544 53168
rect 70676 53116 70728 53168
rect 81808 51756 81860 51808
rect 70768 51076 70820 51128
rect 70676 51008 70728 51060
rect 106556 51008 106608 51060
rect 106740 51008 106792 51060
rect 227352 51051 227404 51060
rect 227352 51017 227361 51051
rect 227361 51017 227395 51051
rect 227395 51017 227404 51051
rect 227352 51008 227404 51017
rect 211896 50711 211948 50720
rect 211896 50677 211905 50711
rect 211905 50677 211939 50711
rect 211939 50677 211948 50711
rect 211896 50668 211948 50677
rect 94136 50643 94188 50652
rect 94136 50609 94145 50643
rect 94145 50609 94179 50643
rect 94179 50609 94188 50643
rect 94136 50600 94188 50609
rect 262036 49376 262088 49428
rect 262220 49376 262272 49428
rect 73436 48356 73488 48408
rect 72056 48288 72108 48340
rect 72240 48288 72292 48340
rect 73528 48288 73580 48340
rect 78772 48288 78824 48340
rect 78956 48288 79008 48340
rect 84568 48288 84620 48340
rect 84660 48288 84712 48340
rect 92756 48288 92808 48340
rect 234068 48288 234120 48340
rect 234252 48288 234304 48340
rect 235724 48331 235776 48340
rect 235724 48297 235733 48331
rect 235733 48297 235767 48331
rect 235767 48297 235776 48331
rect 235724 48288 235776 48297
rect 151084 48263 151136 48272
rect 151084 48229 151093 48263
rect 151093 48229 151127 48263
rect 151127 48229 151136 48263
rect 151084 48220 151136 48229
rect 324596 48220 324648 48272
rect 324780 48220 324832 48272
rect 92848 48152 92900 48204
rect 96988 47039 97040 47048
rect 96988 47005 96997 47039
rect 96997 47005 97031 47039
rect 97031 47005 97040 47039
rect 96988 46996 97040 47005
rect 90916 46928 90968 46980
rect 91008 46928 91060 46980
rect 104900 46928 104952 46980
rect 105268 46928 105320 46980
rect 242532 46971 242584 46980
rect 242532 46937 242541 46971
rect 242541 46937 242575 46971
rect 242575 46937 242584 46971
rect 242532 46928 242584 46937
rect 72240 46860 72292 46912
rect 73528 46860 73580 46912
rect 96988 46903 97040 46912
rect 96988 46869 96997 46903
rect 96997 46869 97031 46903
rect 97031 46869 97040 46903
rect 96988 46860 97040 46869
rect 193864 46903 193916 46912
rect 193864 46869 193873 46903
rect 193873 46869 193907 46903
rect 193907 46869 193916 46903
rect 193864 46860 193916 46869
rect 204904 46903 204956 46912
rect 204904 46869 204913 46903
rect 204913 46869 204947 46903
rect 204947 46869 204956 46903
rect 204904 46860 204956 46869
rect 234068 46903 234120 46912
rect 234068 46869 234077 46903
rect 234077 46869 234111 46903
rect 234111 46869 234120 46903
rect 234068 46860 234120 46869
rect 246948 46903 247000 46912
rect 246948 46869 246957 46903
rect 246957 46869 246991 46903
rect 246991 46869 247000 46903
rect 246948 46860 247000 46869
rect 250996 46903 251048 46912
rect 250996 46869 251005 46903
rect 251005 46869 251039 46903
rect 251039 46869 251048 46903
rect 250996 46860 251048 46869
rect 252284 46903 252336 46912
rect 252284 46869 252293 46903
rect 252293 46869 252327 46903
rect 252327 46869 252336 46903
rect 252284 46860 252336 46869
rect 255228 46903 255280 46912
rect 255228 46869 255237 46903
rect 255237 46869 255271 46903
rect 255271 46869 255280 46903
rect 255228 46860 255280 46869
rect 259276 46903 259328 46912
rect 259276 46869 259285 46903
rect 259285 46869 259319 46903
rect 259319 46869 259328 46903
rect 259276 46860 259328 46869
rect 324596 46860 324648 46912
rect 91008 46792 91060 46844
rect 91192 46792 91244 46844
rect 268752 46180 268804 46232
rect 269028 46180 269080 46232
rect 264612 44319 264664 44328
rect 264612 44285 264621 44319
rect 264621 44285 264655 44319
rect 264655 44285 264664 44319
rect 264612 44276 264664 44285
rect 267280 44115 267332 44124
rect 267280 44081 267289 44115
rect 267289 44081 267323 44115
rect 267323 44081 267332 44115
rect 267280 44072 267332 44081
rect 70492 41352 70544 41404
rect 70676 41352 70728 41404
rect 70584 41284 70636 41336
rect 70768 41284 70820 41336
rect 89996 41284 90048 41336
rect 104900 41284 104952 41336
rect 105176 41284 105228 41336
rect 89996 41148 90048 41200
rect 77392 38700 77444 38752
rect 78772 38675 78824 38684
rect 78772 38641 78781 38675
rect 78781 38641 78815 38675
rect 78815 38641 78824 38675
rect 78772 38632 78824 38641
rect 81808 38632 81860 38684
rect 151084 38675 151136 38684
rect 151084 38641 151093 38675
rect 151093 38641 151127 38675
rect 151127 38641 151136 38675
rect 151084 38632 151136 38641
rect 234068 38675 234120 38684
rect 234068 38641 234077 38675
rect 234077 38641 234111 38675
rect 234111 38641 234120 38675
rect 234068 38632 234120 38641
rect 77392 38564 77444 38616
rect 106832 38607 106884 38616
rect 106832 38573 106841 38607
rect 106841 38573 106875 38607
rect 106875 38573 106884 38607
rect 106832 38564 106884 38573
rect 211988 38564 212040 38616
rect 235724 38607 235776 38616
rect 235724 38573 235733 38607
rect 235733 38573 235767 38607
rect 235767 38573 235776 38607
rect 235724 38564 235776 38573
rect 324872 38539 324924 38548
rect 324872 38505 324881 38539
rect 324881 38505 324915 38539
rect 324915 38505 324924 38539
rect 324872 38496 324924 38505
rect 72056 37315 72108 37324
rect 72056 37281 72065 37315
rect 72065 37281 72099 37315
rect 72099 37281 72108 37315
rect 72056 37272 72108 37281
rect 73436 37315 73488 37324
rect 73436 37281 73445 37315
rect 73445 37281 73479 37315
rect 73479 37281 73488 37315
rect 73436 37272 73488 37281
rect 78772 37315 78824 37324
rect 78772 37281 78781 37315
rect 78781 37281 78815 37315
rect 78815 37281 78824 37315
rect 78772 37272 78824 37281
rect 96988 37315 97040 37324
rect 96988 37281 96997 37315
rect 96997 37281 97031 37315
rect 97031 37281 97040 37315
rect 96988 37272 97040 37281
rect 204904 37315 204956 37324
rect 204904 37281 204913 37315
rect 204913 37281 204947 37315
rect 204947 37281 204956 37315
rect 204904 37272 204956 37281
rect 243636 37272 243688 37324
rect 243820 37272 243872 37324
rect 246948 37315 247000 37324
rect 246948 37281 246957 37315
rect 246957 37281 246991 37315
rect 246991 37281 247000 37315
rect 246948 37272 247000 37281
rect 250996 37315 251048 37324
rect 250996 37281 251005 37315
rect 251005 37281 251039 37315
rect 251039 37281 251048 37315
rect 250996 37272 251048 37281
rect 252284 37315 252336 37324
rect 252284 37281 252293 37315
rect 252293 37281 252327 37315
rect 252327 37281 252336 37315
rect 252284 37272 252336 37281
rect 255228 37315 255280 37324
rect 255228 37281 255237 37315
rect 255237 37281 255271 37315
rect 255271 37281 255280 37315
rect 255228 37272 255280 37281
rect 259276 37315 259328 37324
rect 259276 37281 259285 37315
rect 259285 37281 259319 37315
rect 259319 37281 259328 37315
rect 259276 37272 259328 37281
rect 242532 37247 242584 37256
rect 242532 37213 242541 37247
rect 242541 37213 242575 37247
rect 242575 37213 242584 37247
rect 242532 37204 242584 37213
rect 73436 36295 73488 36304
rect 73436 36261 73445 36295
rect 73445 36261 73479 36295
rect 73479 36261 73488 36295
rect 73436 36252 73488 36261
rect 267372 35776 267424 35828
rect 70492 33804 70544 33856
rect 70676 33804 70728 33856
rect 262036 33192 262088 33244
rect 264428 33192 264480 33244
rect 264612 33192 264664 33244
rect 268752 32172 268804 32224
rect 269028 32172 269080 32224
rect 70768 31764 70820 31816
rect 94136 31764 94188 31816
rect 70676 31696 70728 31748
rect 105176 31764 105228 31816
rect 324872 31764 324924 31816
rect 105084 31696 105136 31748
rect 227260 31696 227312 31748
rect 227444 31696 227496 31748
rect 324872 31628 324924 31680
rect 94136 31560 94188 31612
rect 106832 31603 106884 31612
rect 106832 31569 106841 31603
rect 106841 31569 106875 31603
rect 106875 31569 106884 31603
rect 106832 31560 106884 31569
rect 262036 29656 262088 29708
rect 84660 29044 84712 29096
rect 72056 28976 72108 29028
rect 72240 28976 72292 29028
rect 73528 28976 73580 29028
rect 84568 28976 84620 29028
rect 91008 28976 91060 29028
rect 91192 28976 91244 29028
rect 193956 28976 194008 29028
rect 211896 29019 211948 29028
rect 211896 28985 211905 29019
rect 211905 28985 211939 29019
rect 211939 28985 211948 29019
rect 211896 28976 211948 28985
rect 235724 29019 235776 29028
rect 235724 28985 235733 29019
rect 235733 28985 235767 29019
rect 235767 28985 235776 29019
rect 235724 28976 235776 28985
rect 89996 28951 90048 28960
rect 89996 28917 90005 28951
rect 90005 28917 90039 28951
rect 90039 28917 90048 28951
rect 89996 28908 90048 28917
rect 96988 28951 97040 28960
rect 96988 28917 96997 28951
rect 96997 28917 97031 28951
rect 97031 28917 97040 28951
rect 96988 28908 97040 28917
rect 151084 28951 151136 28960
rect 151084 28917 151093 28951
rect 151093 28917 151127 28951
rect 151127 28917 151136 28951
rect 151084 28908 151136 28917
rect 92848 27684 92900 27736
rect 92756 27616 92808 27668
rect 242532 27659 242584 27668
rect 242532 27625 242541 27659
rect 242541 27625 242575 27659
rect 242575 27625 242584 27659
rect 242532 27616 242584 27625
rect 77484 27591 77536 27600
rect 77484 27557 77493 27591
rect 77493 27557 77527 27591
rect 77527 27557 77536 27591
rect 77484 27548 77536 27557
rect 78956 27548 79008 27600
rect 91008 27548 91060 27600
rect 204904 27591 204956 27600
rect 204904 27557 204913 27591
rect 204913 27557 204947 27591
rect 204947 27557 204956 27591
rect 204904 27548 204956 27557
rect 248236 27591 248288 27600
rect 248236 27557 248245 27591
rect 248245 27557 248279 27591
rect 248279 27557 248288 27591
rect 248236 27548 248288 27557
rect 249616 27591 249668 27600
rect 249616 27557 249625 27591
rect 249625 27557 249659 27591
rect 249659 27557 249668 27591
rect 249616 27548 249668 27557
rect 255228 27591 255280 27600
rect 255228 27557 255237 27591
rect 255237 27557 255271 27591
rect 255271 27557 255280 27591
rect 255228 27548 255280 27557
rect 268752 26868 268804 26920
rect 269028 26868 269080 26920
rect 260472 26188 260524 26240
rect 264428 24828 264480 24880
rect 264704 24828 264756 24880
rect 262036 23332 262088 23384
rect 262220 23332 262272 23384
rect 259184 22763 259236 22772
rect 259184 22729 259193 22763
rect 259193 22729 259227 22763
rect 259227 22729 259236 22763
rect 259184 22720 259236 22729
rect 70492 22652 70544 22704
rect 70676 22652 70728 22704
rect 72240 22108 72292 22160
rect 72148 22040 72200 22092
rect 96988 21947 97040 21956
rect 96988 21913 96997 21947
rect 96997 21913 97031 21947
rect 97031 21913 97040 21947
rect 96988 21904 97040 21913
rect 250812 19864 250864 19916
rect 250996 19864 251048 19916
rect 89996 19363 90048 19372
rect 89996 19329 90005 19363
rect 90005 19329 90039 19363
rect 90039 19329 90048 19363
rect 89996 19320 90048 19329
rect 151084 19363 151136 19372
rect 151084 19329 151093 19363
rect 151093 19329 151127 19363
rect 151127 19329 151136 19363
rect 151084 19320 151136 19329
rect 193772 19295 193824 19304
rect 193772 19261 193781 19295
rect 193781 19261 193815 19295
rect 193815 19261 193824 19295
rect 193772 19252 193824 19261
rect 227352 19295 227404 19304
rect 227352 19261 227361 19295
rect 227361 19261 227395 19295
rect 227395 19261 227404 19295
rect 227352 19252 227404 19261
rect 234344 19252 234396 19304
rect 234620 19252 234672 19304
rect 235724 19295 235776 19304
rect 235724 19261 235733 19295
rect 235733 19261 235767 19295
rect 235767 19261 235776 19295
rect 235724 19252 235776 19261
rect 245292 19252 245344 19304
rect 245568 19252 245620 19304
rect 77484 18003 77536 18012
rect 77484 17969 77493 18003
rect 77493 17969 77527 18003
rect 77527 17969 77536 18003
rect 77484 17960 77536 17969
rect 78864 18003 78916 18012
rect 78864 17969 78873 18003
rect 78873 17969 78907 18003
rect 78907 17969 78916 18003
rect 78864 17960 78916 17969
rect 91008 17960 91060 18012
rect 204904 18003 204956 18012
rect 204904 17969 204913 18003
rect 204913 17969 204947 18003
rect 204947 17969 204956 18003
rect 204904 17960 204956 17969
rect 243728 17960 243780 18012
rect 243820 17960 243872 18012
rect 248236 18003 248288 18012
rect 248236 17969 248245 18003
rect 248245 17969 248279 18003
rect 248279 17969 248288 18003
rect 248236 17960 248288 17969
rect 249616 18003 249668 18012
rect 249616 17969 249625 18003
rect 249625 17969 249659 18003
rect 249659 17969 249668 18003
rect 249616 17960 249668 17969
rect 255228 18003 255280 18012
rect 255228 17969 255237 18003
rect 255237 17969 255271 18003
rect 255271 17969 255280 18003
rect 255228 17960 255280 17969
rect 73436 17892 73488 17944
rect 268752 17212 268804 17264
rect 269028 17212 269080 17264
rect 248236 17076 248288 17128
rect 248420 17076 248472 17128
rect 219072 16532 219124 16584
rect 219348 16532 219400 16584
rect 169484 16396 169536 16448
rect 285680 16396 285732 16448
rect 170864 16328 170916 16380
rect 288440 16328 288492 16380
rect 172152 16260 172204 16312
rect 292580 16260 292632 16312
rect 173624 16192 173676 16244
rect 296720 16192 296772 16244
rect 176292 16124 176344 16176
rect 303620 16124 303672 16176
rect 206744 16056 206796 16108
rect 391940 16056 391992 16108
rect 212264 15988 212316 16040
rect 407120 15988 407172 16040
rect 216312 15920 216364 15972
rect 420920 15920 420972 15972
rect 477500 15852 477552 15904
rect 202788 15104 202840 15156
rect 379520 15104 379572 15156
rect 204076 15036 204128 15088
rect 382372 15036 382424 15088
rect 202696 14968 202748 15020
rect 380900 14968 380952 15020
rect 203892 14900 203944 14952
rect 383660 14900 383712 14952
rect 205456 14832 205508 14884
rect 387800 14832 387852 14884
rect 203984 14764 204036 14816
rect 386420 14764 386472 14816
rect 206836 14696 206888 14748
rect 390560 14696 390612 14748
rect 237104 14628 237156 14680
rect 478880 14628 478932 14680
rect 238576 14560 238628 14612
rect 484400 14560 484452 14612
rect 238392 14492 238444 14544
rect 485780 14492 485832 14544
rect 239680 14424 239732 14476
rect 487160 14424 487212 14476
rect 201224 14356 201276 14408
rect 375380 14356 375432 14408
rect 170956 14288 171008 14340
rect 287060 14288 287112 14340
rect 169576 14220 169628 14272
rect 284300 14220 284352 14272
rect 168196 14152 168248 14204
rect 282920 14152 282972 14204
rect 168012 14084 168064 14136
rect 281540 14084 281592 14136
rect 166724 14016 166776 14068
rect 278872 14016 278924 14068
rect 168288 13948 168340 14000
rect 280160 13948 280212 14000
rect 168104 13880 168156 13932
rect 278780 13880 278832 13932
rect 166816 13812 166868 13864
rect 277400 13812 277452 13864
rect 248144 13744 248196 13796
rect 510620 13744 510672 13796
rect 248052 13676 248104 13728
rect 513380 13676 513432 13728
rect 249524 13608 249576 13660
rect 517520 13608 517572 13660
rect 250904 13540 250956 13592
rect 520280 13540 520332 13592
rect 252192 13472 252244 13524
rect 524420 13472 524472 13524
rect 253664 13404 253716 13456
rect 528560 13404 528612 13456
rect 255044 13336 255096 13388
rect 531320 13336 531372 13388
rect 256332 13268 256384 13320
rect 535460 13268 535512 13320
rect 257804 13200 257856 13252
rect 538220 13200 538272 13252
rect 542360 13132 542412 13184
rect 255136 13107 255188 13116
rect 255136 13073 255145 13107
rect 255145 13073 255179 13107
rect 255179 13073 255188 13107
rect 255136 13064 255188 13073
rect 546500 13064 546552 13116
rect 246764 12996 246816 13048
rect 506480 12996 506532 13048
rect 245384 12928 245436 12980
rect 502340 12928 502392 12980
rect 243820 12860 243872 12912
rect 499580 12860 499632 12912
rect 242440 12792 242492 12844
rect 495440 12792 495492 12844
rect 241152 12724 241204 12776
rect 492680 12724 492732 12776
rect 240048 12656 240100 12708
rect 488540 12656 488592 12708
rect 239956 12588 240008 12640
rect 485872 12588 485924 12640
rect 70676 12520 70728 12572
rect 238668 12520 238720 12572
rect 483020 12520 483072 12572
rect 70492 12452 70544 12504
rect 91008 12452 91060 12504
rect 94136 12452 94188 12504
rect 165344 12452 165396 12504
rect 271880 12452 271932 12504
rect 90916 12384 90968 12436
rect 193772 12427 193824 12436
rect 193772 12393 193781 12427
rect 193781 12393 193815 12427
rect 193815 12393 193824 12427
rect 193772 12384 193824 12393
rect 217876 12384 217928 12436
rect 423680 12384 423732 12436
rect 94228 12316 94280 12368
rect 219164 12316 219216 12368
rect 426440 12316 426492 12368
rect 220544 12248 220596 12300
rect 430580 12248 430632 12300
rect 220636 12180 220688 12232
rect 433340 12180 433392 12232
rect 221924 12112 221976 12164
rect 437480 12112 437532 12164
rect 223396 12044 223448 12096
rect 441620 12044 441672 12096
rect 224684 11976 224736 12028
rect 444380 11976 444432 12028
rect 226064 11908 226116 11960
rect 448520 11908 448572 11960
rect 451280 11840 451332 11892
rect 228824 11772 228876 11824
rect 455420 11772 455472 11824
rect 230296 11704 230348 11756
rect 459652 11704 459704 11756
rect 216404 11636 216456 11688
rect 419540 11636 419592 11688
rect 215116 11568 215168 11620
rect 416872 11568 416924 11620
rect 213644 11500 213696 11552
rect 412640 11500 412692 11552
rect 212356 11432 212408 11484
rect 408500 11432 408552 11484
rect 210976 11364 211028 11416
rect 405740 11364 405792 11416
rect 209596 11296 209648 11348
rect 401600 11296 401652 11348
rect 208032 11228 208084 11280
rect 398840 11228 398892 11280
rect 208124 11160 208176 11212
rect 394700 11160 394752 11212
rect 165436 11092 165488 11144
rect 274640 11092 274692 11144
rect 253664 11024 253716 11076
rect 253848 11024 253900 11076
rect 255136 11067 255188 11076
rect 255136 11033 255145 11067
rect 255145 11033 255179 11067
rect 255179 11033 255188 11067
rect 255136 11024 255188 11033
rect 183376 10956 183428 11008
rect 322940 10956 322992 11008
rect 184664 10888 184716 10940
rect 327080 10888 327132 10940
rect 184572 10820 184624 10872
rect 331312 10820 331364 10872
rect 186136 10752 186188 10804
rect 333980 10752 334032 10804
rect 187424 10684 187476 10736
rect 338120 10684 338172 10736
rect 188804 10616 188856 10668
rect 340880 10616 340932 10668
rect 190276 10548 190328 10600
rect 345020 10548 345072 10600
rect 191564 10480 191616 10532
rect 347780 10480 347832 10532
rect 192944 10412 192996 10464
rect 351920 10412 351972 10464
rect 194324 10344 194376 10396
rect 356152 10344 356204 10396
rect 195796 10276 195848 10328
rect 358820 10276 358872 10328
rect 181904 10208 181956 10260
rect 320180 10208 320232 10260
rect 180524 10140 180576 10192
rect 316040 10140 316092 10192
rect 179144 10072 179196 10124
rect 313372 10072 313424 10124
rect 177856 10004 177908 10056
rect 309140 10004 309192 10056
rect 176384 9936 176436 9988
rect 305000 9936 305052 9988
rect 175004 9868 175056 9920
rect 302240 9868 302292 9920
rect 173716 9800 173768 9852
rect 298100 9800 298152 9852
rect 162124 9732 162176 9784
rect 172336 9732 172388 9784
rect 295340 9732 295392 9784
rect 161940 9664 161992 9716
rect 172244 9664 172296 9716
rect 291200 9664 291252 9716
rect 90916 9596 90968 9648
rect 94228 9639 94280 9648
rect 94228 9605 94237 9639
rect 94237 9605 94271 9639
rect 94271 9605 94280 9639
rect 94228 9596 94280 9605
rect 154396 9596 154448 9648
rect 250352 9596 250404 9648
rect 250904 9596 250956 9648
rect 520372 9596 520424 9648
rect 155776 9528 155828 9580
rect 90916 9460 90968 9512
rect 155684 9460 155736 9512
rect 246764 9528 246816 9580
rect 157064 9392 157116 9444
rect 245568 9460 245620 9512
rect 245476 9392 245528 9444
rect 252192 9528 252244 9580
rect 523868 9528 523920 9580
rect 253756 9460 253808 9512
rect 527456 9460 527508 9512
rect 253848 9392 253900 9444
rect 256424 9392 256476 9444
rect 156972 9324 157024 9376
rect 244004 9324 244056 9376
rect 158536 9256 158588 9308
rect 246856 9256 246908 9308
rect 249524 9324 249576 9376
rect 531044 9392 531096 9444
rect 534540 9324 534592 9376
rect 252652 9256 252704 9308
rect 158444 9188 158496 9240
rect 159916 9120 159968 9172
rect 256240 9188 256292 9240
rect 256516 9256 256568 9308
rect 538128 9256 538180 9308
rect 257804 9188 257856 9240
rect 257896 9188 257948 9240
rect 541716 9188 541768 9240
rect 159824 9052 159876 9104
rect 255136 9120 255188 9172
rect 259828 9120 259880 9172
rect 260656 9120 260708 9172
rect 548892 9120 548944 9172
rect 267372 9052 267424 9104
rect 267464 9052 267516 9104
rect 566740 9052 566792 9104
rect 162676 8984 162728 9036
rect 267004 8984 267056 9036
rect 267556 8984 267608 9036
rect 570236 8984 570288 9036
rect 153016 8916 153068 8968
rect 164056 8916 164108 8968
rect 270500 8916 270552 8968
rect 271696 8916 271748 8968
rect 581092 8916 581144 8968
rect 154304 8848 154356 8900
rect 205640 8780 205692 8832
rect 215116 8780 215168 8832
rect 224960 8780 225012 8832
rect 152924 8712 152976 8764
rect 238392 8712 238444 8764
rect 248788 8848 248840 8900
rect 516784 8848 516836 8900
rect 242716 8780 242768 8832
rect 241980 8712 242032 8764
rect 248144 8712 248196 8764
rect 248420 8712 248472 8764
rect 513196 8780 513248 8832
rect 509608 8712 509660 8764
rect 152832 8644 152884 8696
rect 236000 8644 236052 8696
rect 243176 8644 243228 8696
rect 176476 8440 176528 8492
rect 197176 8576 197228 8628
rect 506020 8644 506072 8696
rect 249340 8576 249392 8628
rect 502432 8576 502484 8628
rect 181996 8508 182048 8560
rect 191656 8372 191708 8424
rect 234436 8372 234488 8424
rect 242900 8508 242952 8560
rect 498936 8508 498988 8560
rect 239772 8440 239824 8492
rect 495348 8440 495400 8492
rect 241336 8372 241388 8424
rect 491760 8372 491812 8424
rect 73344 8347 73396 8356
rect 73344 8313 73353 8347
rect 73353 8313 73387 8347
rect 73387 8313 73396 8347
rect 73344 8304 73396 8313
rect 165528 8304 165580 8356
rect 274088 8304 274140 8356
rect 216496 8236 216548 8288
rect 419172 8236 419224 8288
rect 216588 8168 216640 8220
rect 422760 8168 422812 8220
rect 217968 8100 218020 8152
rect 426348 8100 426400 8152
rect 219256 8032 219308 8084
rect 429936 8032 429988 8084
rect 140504 7964 140556 8016
rect 202696 7964 202748 8016
rect 220728 7964 220780 8016
rect 433524 7964 433576 8016
rect 141976 7896 142028 7948
rect 206284 7896 206336 7948
rect 218704 7896 218756 7948
rect 219256 7896 219308 7948
rect 222016 7896 222068 7948
rect 437020 7896 437072 7948
rect 143356 7828 143408 7880
rect 209872 7828 209924 7880
rect 223488 7828 223540 7880
rect 440608 7828 440660 7880
rect 144552 7760 144604 7812
rect 213460 7760 213512 7812
rect 224776 7760 224828 7812
rect 444196 7760 444248 7812
rect 146116 7692 146168 7744
rect 217048 7692 217100 7744
rect 226156 7692 226208 7744
rect 447784 7692 447836 7744
rect 147496 7624 147548 7676
rect 220544 7624 220596 7676
rect 227628 7624 227680 7676
rect 451372 7624 451424 7676
rect 148784 7556 148836 7608
rect 224132 7556 224184 7608
rect 227536 7556 227588 7608
rect 454868 7556 454920 7608
rect 215208 7488 215260 7540
rect 415676 7488 415728 7540
rect 156604 7420 156656 7472
rect 213736 7420 213788 7472
rect 412088 7420 412140 7472
rect 212448 7352 212500 7404
rect 408592 7352 408644 7404
rect 211068 7284 211120 7336
rect 404912 7284 404964 7336
rect 209688 7216 209740 7268
rect 401324 7216 401376 7268
rect 208216 7148 208268 7200
rect 397828 7148 397880 7200
rect 206928 7080 206980 7132
rect 394240 7080 394292 7132
rect 198004 7012 198056 7064
rect 204812 7012 204864 7064
rect 205548 7012 205600 7064
rect 390652 7012 390704 7064
rect 161296 6944 161348 6996
rect 263416 6944 263468 6996
rect 241428 6919 241480 6928
rect 241428 6885 241437 6919
rect 241437 6885 241471 6919
rect 241471 6885 241480 6919
rect 241428 6876 241480 6885
rect 248328 6876 248380 6928
rect 180616 6808 180668 6860
rect 319260 6808 319312 6860
rect 182088 6740 182140 6792
rect 322848 6740 322900 6792
rect 183468 6672 183520 6724
rect 326436 6672 326488 6724
rect 161940 6604 161992 6656
rect 184756 6604 184808 6656
rect 330024 6604 330076 6656
rect 129464 6536 129516 6588
rect 170588 6536 170640 6588
rect 186228 6536 186280 6588
rect 333612 6536 333664 6588
rect 130844 6468 130896 6520
rect 174176 6468 174228 6520
rect 187516 6468 187568 6520
rect 337108 6468 337160 6520
rect 132224 6400 132276 6452
rect 177764 6400 177816 6452
rect 188896 6400 188948 6452
rect 340696 6400 340748 6452
rect 133788 6332 133840 6384
rect 181352 6332 181404 6384
rect 190368 6332 190420 6384
rect 344284 6332 344336 6384
rect 135168 6264 135220 6316
rect 184848 6264 184900 6316
rect 191748 6264 191800 6316
rect 347872 6264 347924 6316
rect 136548 6196 136600 6248
rect 188436 6196 188488 6248
rect 193036 6196 193088 6248
rect 351368 6196 351420 6248
rect 136456 6128 136508 6180
rect 192024 6128 192076 6180
rect 193128 6128 193180 6180
rect 354956 6128 355008 6180
rect 180708 6060 180760 6112
rect 315764 6060 315816 6112
rect 179236 5992 179288 6044
rect 312176 5992 312228 6044
rect 177948 5924 178000 5976
rect 308588 5924 308640 5976
rect 176568 5856 176620 5908
rect 305092 5856 305144 5908
rect 175096 5788 175148 5840
rect 301412 5788 301464 5840
rect 173808 5720 173860 5772
rect 297916 5720 297968 5772
rect 172428 5652 172480 5704
rect 294328 5652 294380 5704
rect 171048 5584 171100 5636
rect 290740 5584 290792 5636
rect 157156 5516 157208 5568
rect 169668 5516 169720 5568
rect 286968 5516 287020 5568
rect 287060 5516 287112 5568
rect 288348 5516 288400 5568
rect 367744 5516 367796 5568
rect 368204 5516 368256 5568
rect 148968 5448 149020 5500
rect 226524 5448 226576 5500
rect 245384 5448 245436 5500
rect 252376 5448 252428 5500
rect 526260 5448 526312 5500
rect 148876 5380 148928 5432
rect 227720 5380 227772 5432
rect 253664 5380 253716 5432
rect 529848 5380 529900 5432
rect 150256 5312 150308 5364
rect 230112 5312 230164 5364
rect 249708 5312 249760 5364
rect 533436 5312 533488 5364
rect 58808 5244 58860 5296
rect 89812 5244 89864 5296
rect 150348 5244 150400 5296
rect 231308 5244 231360 5296
rect 256608 5244 256660 5296
rect 536932 5244 536984 5296
rect 55220 5176 55272 5228
rect 88432 5176 88484 5228
rect 151636 5176 151688 5228
rect 233700 5176 233752 5228
rect 257988 5176 258040 5228
rect 540520 5176 540572 5228
rect 51632 5108 51684 5160
rect 87052 5108 87104 5160
rect 151728 5108 151780 5160
rect 234804 5108 234856 5160
rect 251456 5108 251508 5160
rect 255136 5108 255188 5160
rect 260748 5108 260800 5160
rect 48228 5040 48280 5092
rect 85672 5040 85724 5092
rect 116952 5040 117004 5092
rect 117228 5040 117280 5092
rect 153108 5040 153160 5092
rect 237196 5040 237248 5092
rect 242808 5040 242860 5092
rect 264612 5040 264664 5092
rect 264888 5040 264940 5092
rect 544108 5108 544160 5160
rect 7656 4972 7708 5024
rect 72148 4972 72200 5024
rect 154488 4972 154540 5024
rect 240784 4972 240836 5024
rect 244188 4972 244240 5024
rect 252468 4972 252520 5024
rect 261024 4972 261076 5024
rect 262128 4972 262180 5024
rect 2872 4904 2924 4956
rect 70768 4904 70820 4956
rect 155868 4904 155920 4956
rect 244372 4904 244424 4956
rect 572 4836 624 4888
rect 69020 4836 69072 4888
rect 157248 4836 157300 4888
rect 247960 4836 248012 4888
rect 1676 4768 1728 4820
rect 70492 4768 70544 4820
rect 215116 4768 215168 4820
rect 215576 4768 215628 4820
rect 147588 4700 147640 4752
rect 146208 4632 146260 4684
rect 218980 4632 219032 4684
rect 219256 4632 219308 4684
rect 144736 4564 144788 4616
rect 215852 4564 215904 4616
rect 144644 4496 144696 4548
rect 212264 4496 212316 4548
rect 215116 4496 215168 4548
rect 222936 4564 222988 4616
rect 216036 4496 216088 4548
rect 268108 4904 268160 4956
rect 547696 5040 547748 5092
rect 551192 4972 551244 5024
rect 561956 4904 562008 4956
rect 259276 4836 259328 4888
rect 268752 4836 268804 4888
rect 572628 4836 572680 4888
rect 143448 4428 143500 4480
rect 208676 4428 208728 4480
rect 209044 4428 209096 4480
rect 211804 4428 211856 4480
rect 215300 4428 215352 4480
rect 249064 4700 249116 4752
rect 271696 4768 271748 4820
rect 271788 4768 271840 4820
rect 579804 4768 579856 4820
rect 522672 4700 522724 4752
rect 251088 4632 251140 4684
rect 519084 4632 519136 4684
rect 142068 4360 142120 4412
rect 205088 4360 205140 4412
rect 231860 4360 231912 4412
rect 244188 4428 244240 4480
rect 140596 4292 140648 4344
rect 201500 4292 201552 4344
rect 36176 4088 36228 4140
rect 81532 4088 81584 4140
rect 34980 4020 35032 4072
rect 81808 4020 81860 4072
rect 82636 4088 82688 4140
rect 84844 4088 84896 4140
rect 87328 4088 87380 4140
rect 88248 4088 88300 4140
rect 89720 4088 89772 4140
rect 91744 4088 91796 4140
rect 93308 4088 93360 4140
rect 93768 4088 93820 4140
rect 94504 4088 94556 4140
rect 95884 4088 95936 4140
rect 96896 4088 96948 4140
rect 97908 4088 97960 4140
rect 102784 4088 102836 4140
rect 103428 4088 103480 4140
rect 105176 4088 105228 4140
rect 106280 4088 106332 4140
rect 106832 4088 106884 4140
rect 107568 4088 107620 4140
rect 107844 4088 107896 4140
rect 108764 4088 108816 4140
rect 125324 4088 125376 4140
rect 134524 4156 134576 4208
rect 139308 4224 139360 4276
rect 198004 4224 198056 4276
rect 202144 4224 202196 4276
rect 232504 4292 232556 4344
rect 84384 4020 84436 4072
rect 86132 4020 86184 4072
rect 89076 4020 89128 4072
rect 96712 4020 96764 4072
rect 101588 4020 101640 4072
rect 104992 4020 105044 4072
rect 114284 4020 114336 4072
rect 127532 4020 127584 4072
rect 30288 3952 30340 4004
rect 80336 3952 80388 4004
rect 81440 3952 81492 4004
rect 88984 3952 89036 4004
rect 96620 3952 96672 4004
rect 110328 3952 110380 4004
rect 114744 3952 114796 4004
rect 115664 3952 115716 4004
rect 27896 3884 27948 3936
rect 71872 3884 71924 3936
rect 80060 3884 80112 3936
rect 20720 3816 20772 3868
rect 76012 3816 76064 3868
rect 21916 3748 21968 3800
rect 12440 3680 12492 3732
rect 73160 3748 73212 3800
rect 78864 3816 78916 3868
rect 79048 3816 79100 3868
rect 96988 3884 97040 3936
rect 100484 3884 100536 3936
rect 103704 3884 103756 3936
rect 121368 3884 121420 3936
rect 145564 4088 145616 4140
rect 193864 4156 193916 4208
rect 225328 4156 225380 4208
rect 231952 4224 232004 4276
rect 257436 4564 257488 4616
rect 515588 4564 515640 4616
rect 512000 4496 512052 4548
rect 249248 4428 249300 4480
rect 508412 4428 508464 4480
rect 504824 4360 504876 4412
rect 501236 4292 501288 4344
rect 497740 4224 497792 4276
rect 228916 4156 228968 4208
rect 494152 4156 494204 4208
rect 183744 4088 183796 4140
rect 184756 4088 184808 4140
rect 328828 4088 328880 4140
rect 345020 4088 345072 4140
rect 354588 4088 354640 4140
rect 368020 4088 368072 4140
rect 368204 4088 368256 4140
rect 369124 4088 369176 4140
rect 446588 4088 446640 4140
rect 128176 4020 128228 4072
rect 148324 4020 148376 4072
rect 153844 4020 153896 4072
rect 156328 4020 156380 4072
rect 164700 4020 164752 4072
rect 186044 4020 186096 4072
rect 187608 4020 187660 4072
rect 335912 4020 335964 4072
rect 336004 4020 336056 4072
rect 364892 4020 364944 4072
rect 364984 4020 365036 4072
rect 453672 4020 453724 4072
rect 129004 3952 129056 4004
rect 129648 3952 129700 4004
rect 169392 3952 169444 4004
rect 331864 3952 331916 4004
rect 340236 3952 340288 4004
rect 382280 3952 382332 4004
rect 149244 3884 149296 3936
rect 151176 3884 151228 3936
rect 155132 3884 155184 3936
rect 190828 3884 190880 3936
rect 194508 3884 194560 3936
rect 357348 3884 357400 3936
rect 360936 3884 360988 3936
rect 361028 3884 361080 3936
rect 369124 3884 369176 3936
rect 95700 3816 95752 3868
rect 111616 3816 111668 3868
rect 119436 3816 119488 3868
rect 122656 3816 122708 3868
rect 151544 3816 151596 3868
rect 152464 3816 152516 3868
rect 194416 3816 194468 3868
rect 200028 3816 200080 3868
rect 371608 3816 371660 3868
rect 371884 3884 371936 3936
rect 467932 3884 467984 3936
rect 482284 3816 482336 3868
rect 77484 3748 77536 3800
rect 77852 3748 77904 3800
rect 93952 3748 94004 3800
rect 115848 3748 115900 3800
rect 130200 3748 130252 3800
rect 131028 3748 131080 3800
rect 172980 3748 173032 3800
rect 201408 3748 201460 3800
rect 378784 3748 378836 3800
rect 382372 3748 382424 3800
rect 383568 3748 383620 3800
rect 92112 3680 92164 3732
rect 100116 3680 100168 3732
rect 115756 3680 115808 3732
rect 131396 3680 131448 3732
rect 132408 3680 132460 3732
rect 176568 3680 176620 3732
rect 179328 3680 179380 3732
rect 204168 3680 204220 3732
rect 385868 3680 385920 3732
rect 390560 3680 390612 3732
rect 391848 3680 391900 3732
rect 11244 3612 11296 3664
rect 73252 3612 73304 3664
rect 75460 3612 75512 3664
rect 95240 3612 95292 3664
rect 98092 3612 98144 3664
rect 102600 3612 102652 3664
rect 111156 3612 111208 3664
rect 8852 3544 8904 3596
rect 71780 3544 71832 3596
rect 74264 3544 74316 3596
rect 95424 3544 95476 3596
rect 6460 3476 6512 3528
rect 71964 3476 72016 3528
rect 73068 3476 73120 3528
rect 95332 3476 95384 3528
rect 99288 3476 99340 3528
rect 100024 3476 100076 3528
rect 103980 3476 104032 3528
rect 104808 3476 104860 3528
rect 111064 3476 111116 3528
rect 112352 3476 112404 3528
rect 113088 3612 113140 3664
rect 123024 3612 123076 3664
rect 113824 3544 113876 3596
rect 117136 3544 117188 3596
rect 115940 3476 115992 3528
rect 4068 3408 4120 3460
rect 70400 3408 70452 3460
rect 16028 3340 16080 3392
rect 16488 3340 16540 3392
rect 17224 3340 17276 3392
rect 17868 3340 17920 3392
rect 24308 3340 24360 3392
rect 24768 3340 24820 3392
rect 25504 3340 25556 3392
rect 26148 3340 26200 3392
rect 26700 3340 26752 3392
rect 27528 3340 27580 3392
rect 33876 3340 33928 3392
rect 34428 3340 34480 3392
rect 76656 3408 76708 3460
rect 79784 3340 79836 3392
rect 93860 3408 93912 3460
rect 95700 3408 95752 3460
rect 96528 3408 96580 3460
rect 110236 3408 110288 3460
rect 82544 3340 82596 3392
rect 88432 3340 88484 3392
rect 88524 3340 88576 3392
rect 98276 3340 98328 3392
rect 108948 3340 109000 3392
rect 111156 3340 111208 3392
rect 111708 3408 111760 3460
rect 118240 3408 118292 3460
rect 113548 3340 113600 3392
rect 114376 3340 114428 3392
rect 122564 3476 122616 3528
rect 153936 3612 153988 3664
rect 155224 3612 155276 3664
rect 199200 3612 199252 3664
rect 208308 3612 208360 3664
rect 396632 3612 396684 3664
rect 408500 3612 408552 3664
rect 409696 3612 409748 3664
rect 126612 3544 126664 3596
rect 126888 3544 126940 3596
rect 162308 3544 162360 3596
rect 164792 3544 164844 3596
rect 164884 3544 164936 3596
rect 167092 3544 167144 3596
rect 167644 3544 167696 3596
rect 168288 3544 168340 3596
rect 211068 3544 211120 3596
rect 213828 3544 213880 3596
rect 414480 3544 414532 3596
rect 477500 3544 477552 3596
rect 478696 3544 478748 3596
rect 123484 3476 123536 3528
rect 124220 3476 124272 3528
rect 124312 3476 124364 3528
rect 133236 3476 133288 3528
rect 136088 3476 136140 3528
rect 141424 3476 141476 3528
rect 144460 3476 144512 3528
rect 145656 3476 145708 3528
rect 148048 3476 148100 3528
rect 193220 3476 193272 3528
rect 219164 3476 219216 3528
rect 428740 3476 428792 3528
rect 433340 3476 433392 3528
rect 434628 3476 434680 3528
rect 451280 3476 451332 3528
rect 452476 3476 452528 3528
rect 502340 3476 502392 3528
rect 503628 3476 503680 3528
rect 520280 3476 520332 3528
rect 521476 3476 521528 3528
rect 563060 3476 563112 3528
rect 564348 3476 564400 3528
rect 581000 3476 581052 3528
rect 582196 3476 582248 3528
rect 118608 3408 118660 3460
rect 133144 3408 133196 3460
rect 139676 3408 139728 3460
rect 140688 3408 140740 3460
rect 200396 3408 200448 3460
rect 222108 3408 222160 3460
rect 435824 3408 435876 3460
rect 118516 3340 118568 3392
rect 45744 3204 45796 3256
rect 46848 3204 46900 3256
rect 46940 3204 46992 3256
rect 48136 3204 48188 3256
rect 50528 3204 50580 3256
rect 50988 3204 51040 3256
rect 84476 3272 84528 3324
rect 84936 3272 84988 3324
rect 93124 3272 93176 3324
rect 116584 3272 116636 3324
rect 121828 3272 121880 3324
rect 125416 3340 125468 3392
rect 125508 3340 125560 3392
rect 151268 3340 151320 3392
rect 159364 3340 159416 3392
rect 164884 3340 164936 3392
rect 182548 3340 182600 3392
rect 278780 3340 278832 3392
rect 280068 3340 280120 3392
rect 300124 3340 300176 3392
rect 157524 3272 157576 3324
rect 157984 3272 158036 3324
rect 83004 3204 83056 3256
rect 83832 3204 83884 3256
rect 97264 3204 97316 3256
rect 108856 3204 108908 3256
rect 109960 3204 110012 3256
rect 124036 3204 124088 3256
rect 158720 3204 158772 3256
rect 159456 3272 159508 3324
rect 163504 3204 163556 3256
rect 44548 3136 44600 3188
rect 43352 3068 43404 3120
rect 54024 3136 54076 3188
rect 80152 3136 80204 3188
rect 80244 3136 80296 3188
rect 114468 3136 114520 3188
rect 122748 3136 122800 3188
rect 150440 3136 150492 3188
rect 161112 3136 161164 3188
rect 168196 3136 168248 3188
rect 168288 3136 168340 3188
rect 175188 3272 175240 3324
rect 300308 3272 300360 3324
rect 305000 3340 305052 3392
rect 306196 3340 306248 3392
rect 307024 3340 307076 3392
rect 329104 3340 329156 3392
rect 310980 3272 311032 3324
rect 311164 3272 311216 3324
rect 325240 3272 325292 3324
rect 325332 3272 325384 3324
rect 347780 3272 347832 3324
rect 349068 3272 349120 3324
rect 359648 3340 359700 3392
rect 439412 3340 439464 3392
rect 432328 3272 432380 3324
rect 221740 3204 221792 3256
rect 276664 3204 276716 3256
rect 400220 3204 400272 3256
rect 203892 3136 203944 3188
rect 267372 3136 267424 3188
rect 364524 3136 364576 3188
rect 365720 3136 365772 3188
rect 366916 3136 366968 3188
rect 367008 3136 367060 3188
rect 375196 3136 375248 3188
rect 375288 3136 375340 3188
rect 460848 3136 460900 3188
rect 62396 3068 62448 3120
rect 63408 3068 63460 3120
rect 37372 3000 37424 3052
rect 61200 3000 61252 3052
rect 91284 3068 91336 3120
rect 119896 3068 119948 3120
rect 142068 3068 142120 3120
rect 145472 3068 145524 3120
rect 153844 3068 153896 3120
rect 195612 3068 195664 3120
rect 257804 3068 257856 3120
rect 350264 3068 350316 3120
rect 353944 3068 353996 3120
rect 63592 3000 63644 3052
rect 64696 3000 64748 3052
rect 60004 2932 60056 2984
rect 89996 3000 90048 3052
rect 117044 3000 117096 3052
rect 134892 3000 134944 3052
rect 135904 3000 135956 3052
rect 137928 3000 137980 3052
rect 67180 2932 67232 2984
rect 92756 2932 92808 2984
rect 117228 2932 117280 2984
rect 132592 2932 132644 2984
rect 138480 2932 138532 2984
rect 143264 3000 143316 3052
rect 152740 3000 152792 3052
rect 153200 3000 153252 3052
rect 187240 3000 187292 3052
rect 188988 3000 189040 3052
rect 249800 3000 249852 3052
rect 321652 3000 321704 3052
rect 322204 3000 322256 3052
rect 346676 3000 346728 3052
rect 353760 3000 353812 3052
rect 425152 3068 425204 3120
rect 157248 2932 157300 2984
rect 163504 2932 163556 2984
rect 163596 2932 163648 2984
rect 196808 2932 196860 2984
rect 242900 2932 242952 2984
rect 307392 2932 307444 2984
rect 313924 2932 313976 2984
rect 52828 2864 52880 2916
rect 69388 2864 69440 2916
rect 69480 2864 69532 2916
rect 119988 2864 120040 2916
rect 140872 2864 140924 2916
rect 65984 2796 66036 2848
rect 68192 2796 68244 2848
rect 68284 2796 68336 2848
rect 92572 2796 92624 2848
rect 116952 2796 117004 2848
rect 133788 2796 133840 2848
rect 137284 2796 137336 2848
rect 151728 2864 151780 2916
rect 180156 2864 180208 2916
rect 314568 2864 314620 2916
rect 318064 2932 318116 2984
rect 318156 2932 318208 2984
rect 339500 2932 339552 2984
rect 345664 2932 345716 2984
rect 348424 2932 348476 2984
rect 349804 2932 349856 2984
rect 417976 3000 418028 3052
rect 332416 2864 332468 2916
rect 342904 2864 342956 2916
rect 149704 2796 149756 2848
rect 160744 2796 160796 2848
rect 163596 2796 163648 2848
rect 189632 2796 189684 2848
rect 343088 2796 343140 2848
rect 347044 2864 347096 2916
rect 410892 2932 410944 2984
rect 403716 2864 403768 2916
rect 389456 2796 389508 2848
rect 70676 960 70728 1012
rect 146576 552 146628 604
rect 146852 552 146904 604
rect 271880 552 271932 604
rect 272892 552 272944 604
rect 274640 552 274692 604
rect 275284 552 275336 604
rect 277400 552 277452 604
rect 277676 552 277728 604
rect 280160 552 280212 604
rect 281264 552 281316 604
rect 281540 552 281592 604
rect 282460 552 282512 604
rect 282920 552 282972 604
rect 283656 552 283708 604
rect 285680 552 285732 604
rect 285956 552 286008 604
rect 288440 552 288492 604
rect 289544 552 289596 604
rect 291200 552 291252 604
rect 291936 552 291988 604
rect 292580 552 292632 604
rect 293132 552 293184 604
rect 295340 552 295392 604
rect 295524 552 295576 604
rect 298100 552 298152 604
rect 299112 552 299164 604
rect 303620 552 303672 604
rect 303804 552 303856 604
rect 309140 552 309192 604
rect 309784 552 309836 604
rect 316040 552 316092 604
rect 316960 552 317012 604
rect 322940 552 322992 604
rect 324044 552 324096 604
rect 327080 552 327132 604
rect 327632 552 327684 604
rect 333980 552 334032 604
rect 334716 552 334768 604
rect 340880 552 340932 604
rect 341892 552 341944 604
rect 351920 552 351972 604
rect 352564 552 352616 604
rect 358820 552 358872 604
rect 359740 552 359792 604
rect 369860 552 369912 604
rect 370412 552 370464 604
rect 375380 552 375432 604
rect 376392 552 376444 604
rect 376760 552 376812 604
rect 377588 552 377640 604
rect 379520 552 379572 604
rect 379980 552 380032 604
rect 394700 552 394752 604
rect 395436 552 395488 604
rect 401600 552 401652 604
rect 402520 552 402572 604
rect 405740 552 405792 604
rect 406108 552 406160 604
rect 412640 552 412692 604
rect 413284 552 413336 604
rect 419540 552 419592 604
rect 420368 552 420420 604
rect 420920 552 420972 604
rect 421564 552 421616 604
rect 423680 552 423732 604
rect 423956 552 424008 604
rect 426440 552 426492 604
rect 427544 552 427596 604
rect 430580 552 430632 604
rect 431132 552 431184 604
rect 437480 552 437532 604
rect 438216 552 438268 604
rect 455420 552 455472 604
rect 456064 552 456116 604
rect 462320 552 462372 604
rect 463240 552 463292 604
rect 466460 552 466512 604
rect 466828 552 466880 604
rect 469220 552 469272 604
rect 470324 552 470376 604
rect 478880 552 478932 604
rect 479892 552 479944 604
rect 489920 552 489972 604
rect 490564 552 490616 604
rect 495440 552 495492 604
rect 496544 552 496596 604
rect 499580 552 499632 604
rect 500132 552 500184 604
rect 506480 552 506532 604
rect 507216 552 507268 604
rect 510620 552 510672 604
rect 510804 552 510856 604
rect 513380 552 513432 604
rect 514392 552 514444 604
rect 524420 552 524472 604
rect 525064 552 525116 604
rect 531320 552 531372 604
rect 532240 552 532292 604
rect 538220 552 538272 604
rect 539324 552 539376 604
rect 542360 552 542412 604
rect 542912 552 542964 604
rect 549260 552 549312 604
rect 550088 552 550140 604
rect 556160 552 556212 604
rect 557172 552 557224 604
rect 576860 552 576912 604
rect 577412 552 577464 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 78586 656024 78642 656033
rect 78586 655959 78642 655968
rect 187698 656024 187754 656033
rect 187698 655959 187754 655968
rect 78494 654936 78550 654945
rect 78494 654871 78550 654880
rect 78402 653168 78458 653177
rect 78402 653103 78458 653112
rect 78310 652080 78366 652089
rect 78310 652015 78366 652024
rect 78218 647592 78274 647601
rect 78218 647527 78274 647536
rect 75826 568168 75882 568177
rect 75826 568103 75882 568112
rect 73066 567896 73122 567905
rect 73066 567831 73122 567840
rect 70950 523696 71006 523705
rect 70950 523631 71006 523640
rect 70964 521900 70992 523631
rect 73080 521914 73108 567831
rect 75840 524414 75868 568103
rect 77206 568032 77262 568041
rect 77206 567967 77262 567976
rect 74724 524408 74776 524414
rect 74724 524350 74776 524356
rect 75828 524408 75880 524414
rect 75828 524350 75880 524356
rect 72818 521886 73108 521914
rect 74736 521900 74764 524350
rect 77220 522050 77248 567967
rect 78128 567248 78180 567254
rect 78128 567190 78180 567196
rect 77128 522022 77248 522050
rect 77128 521914 77156 522022
rect 76682 521886 77156 521914
rect 78140 521914 78168 567190
rect 78232 523666 78260 647527
rect 78324 523938 78352 652015
rect 78312 523932 78364 523938
rect 78312 523874 78364 523880
rect 78416 523870 78444 653103
rect 78404 523864 78456 523870
rect 78404 523806 78456 523812
rect 78508 523802 78536 654871
rect 78496 523796 78548 523802
rect 78496 523738 78548 523744
rect 78600 523734 78628 655959
rect 187712 655586 187740 655959
rect 156604 655580 156656 655586
rect 156604 655522 156656 655528
rect 187700 655580 187752 655586
rect 187700 655522 187752 655528
rect 78678 650448 78734 650457
rect 78678 650383 78734 650392
rect 78692 524006 78720 650383
rect 78770 649224 78826 649233
rect 78770 649159 78826 649168
rect 78784 524074 78812 649159
rect 78862 589656 78918 589665
rect 78862 589591 78918 589600
rect 78876 524142 78904 589591
rect 103334 570344 103390 570353
rect 103334 570279 103390 570288
rect 94870 570208 94926 570217
rect 94870 570143 94926 570152
rect 98366 570208 98422 570217
rect 98366 570143 98422 570152
rect 101770 570208 101826 570217
rect 101770 570143 101826 570152
rect 86774 568576 86830 568585
rect 86774 568511 86830 568520
rect 85488 567724 85540 567730
rect 85488 567666 85540 567672
rect 81348 567384 81400 567390
rect 81348 567326 81400 567332
rect 81360 524414 81388 567326
rect 82728 567316 82780 567322
rect 82728 567258 82780 567264
rect 80428 524408 80480 524414
rect 80428 524350 80480 524356
rect 81348 524408 81400 524414
rect 81348 524350 81400 524356
rect 78864 524136 78916 524142
rect 78864 524078 78916 524084
rect 78772 524068 78824 524074
rect 78772 524010 78824 524016
rect 78680 524000 78732 524006
rect 78680 523942 78732 523948
rect 78588 523728 78640 523734
rect 78588 523670 78640 523676
rect 78220 523660 78272 523666
rect 78220 523602 78272 523608
rect 78140 521886 78522 521914
rect 80440 521900 80468 524350
rect 82740 521914 82768 567258
rect 85500 524414 85528 567666
rect 86132 525156 86184 525162
rect 86132 525098 86184 525104
rect 84292 524408 84344 524414
rect 84292 524350 84344 524356
rect 85488 524408 85540 524414
rect 85488 524350 85540 524356
rect 82386 521886 82768 521914
rect 84304 521900 84332 524350
rect 86144 521900 86172 525098
rect 86788 523530 86816 568511
rect 93766 568304 93822 568313
rect 93766 568239 93822 568248
rect 93780 568138 93808 568239
rect 93768 568132 93820 568138
rect 93768 568074 93820 568080
rect 94884 567866 94912 570143
rect 95146 568576 95202 568585
rect 95146 568511 95148 568520
rect 95200 568511 95202 568520
rect 95148 568482 95200 568488
rect 95146 568440 95202 568449
rect 95146 568375 95202 568384
rect 94872 567860 94924 567866
rect 94872 567802 94924 567808
rect 91098 567760 91154 567769
rect 91098 567695 91100 567704
rect 91152 567695 91154 567704
rect 91100 567666 91152 567672
rect 95160 567594 95188 568375
rect 98380 568342 98408 570143
rect 98368 568336 98420 568342
rect 96526 568304 96582 568313
rect 96526 568239 96582 568248
rect 97906 568304 97962 568313
rect 98368 568278 98420 568284
rect 100666 568304 100722 568313
rect 97906 568239 97962 568248
rect 100666 568239 100668 568248
rect 96540 568002 96568 568239
rect 97920 568206 97948 568239
rect 100720 568239 100722 568248
rect 100668 568210 100720 568216
rect 97908 568200 97960 568206
rect 97908 568142 97960 568148
rect 101784 568138 101812 570143
rect 101954 568576 102010 568585
rect 101954 568511 102010 568520
rect 102966 568576 103022 568585
rect 102966 568511 103022 568520
rect 103150 568576 103206 568585
rect 103150 568511 103152 568520
rect 101772 568132 101824 568138
rect 101772 568074 101824 568080
rect 96528 567996 96580 568002
rect 96528 567938 96580 567944
rect 97906 567760 97962 567769
rect 97906 567695 97962 567704
rect 100666 567760 100722 567769
rect 100666 567695 100668 567704
rect 97920 567662 97948 567695
rect 100720 567695 100722 567704
rect 100668 567666 100720 567672
rect 97908 567656 97960 567662
rect 97908 567598 97960 567604
rect 95148 567588 95200 567594
rect 95148 567530 95200 567536
rect 88338 567488 88394 567497
rect 88338 567423 88394 567432
rect 88352 567390 88380 567423
rect 88340 567384 88392 567390
rect 86958 567352 87014 567361
rect 88340 567326 88392 567332
rect 89994 567352 90050 567361
rect 86958 567287 87014 567296
rect 89994 567287 89996 567296
rect 86972 567254 87000 567287
rect 90048 567287 90050 567296
rect 89996 567258 90048 567264
rect 86960 567248 87012 567254
rect 86960 567190 87012 567196
rect 93674 567216 93730 567225
rect 93674 567151 93730 567160
rect 95054 567216 95110 567225
rect 95054 567151 95110 567160
rect 96434 567216 96490 567225
rect 96434 567151 96490 567160
rect 99194 567216 99250 567225
rect 99194 567151 99250 567160
rect 91836 525224 91888 525230
rect 91836 525166 91888 525172
rect 89996 525088 90048 525094
rect 89996 525030 90048 525036
rect 88064 524136 88116 524142
rect 88064 524078 88116 524084
rect 86776 523524 86828 523530
rect 86776 523466 86828 523472
rect 88076 521900 88104 524078
rect 90008 521900 90036 525030
rect 91848 521900 91876 525166
rect 93688 524754 93716 567151
rect 93768 525292 93820 525298
rect 93768 525234 93820 525240
rect 93676 524748 93728 524754
rect 93676 524690 93728 524696
rect 93780 521900 93808 525234
rect 95068 524414 95096 567151
rect 95700 525360 95752 525366
rect 95700 525302 95752 525308
rect 95056 524408 95108 524414
rect 95056 524350 95108 524356
rect 95712 521900 95740 525302
rect 96448 524278 96476 567151
rect 97632 525428 97684 525434
rect 97632 525370 97684 525376
rect 96436 524272 96488 524278
rect 96436 524214 96488 524220
rect 97644 521900 97672 525370
rect 99208 524346 99236 567151
rect 101404 525564 101456 525570
rect 101404 525506 101456 525512
rect 99472 525496 99524 525502
rect 99472 525438 99524 525444
rect 99196 524340 99248 524346
rect 99196 524282 99248 524288
rect 99484 521900 99512 525438
rect 101416 521900 101444 525506
rect 101968 524210 101996 568511
rect 102046 568304 102102 568313
rect 102046 568239 102102 568248
rect 102060 567934 102088 568239
rect 102048 567928 102100 567934
rect 102048 567870 102100 567876
rect 102980 567798 103008 568511
rect 103204 568511 103206 568520
rect 103152 568482 103204 568488
rect 103164 568070 103192 568482
rect 103152 568064 103204 568070
rect 103152 568006 103204 568012
rect 102968 567792 103020 567798
rect 102968 567734 103020 567740
rect 101956 524204 102008 524210
rect 101956 524146 102008 524152
rect 103348 524142 103376 570279
rect 109038 570208 109094 570217
rect 109038 570143 109094 570152
rect 112258 570208 112314 570217
rect 112258 570143 112314 570152
rect 117962 570208 118018 570217
rect 117962 570143 118018 570152
rect 119986 570208 120042 570217
rect 119986 570143 120042 570152
rect 104070 568576 104126 568585
rect 104070 568511 104126 568520
rect 104806 568576 104862 568585
rect 104806 568511 104862 568520
rect 105266 568576 105322 568585
rect 105266 568511 105322 568520
rect 106186 568576 106242 568585
rect 106186 568511 106242 568520
rect 106646 568576 106702 568585
rect 106646 568511 106702 568520
rect 107566 568576 107622 568585
rect 107566 568511 107622 568520
rect 107750 568576 107806 568585
rect 107750 568511 107806 568520
rect 108946 568576 109002 568585
rect 108946 568511 109002 568520
rect 104084 567866 104112 568511
rect 104072 567860 104124 567866
rect 104072 567802 104124 567808
rect 104820 524890 104848 568511
rect 105280 568002 105308 568511
rect 105268 567996 105320 568002
rect 105268 567938 105320 567944
rect 104808 524884 104860 524890
rect 104808 524826 104860 524832
rect 106200 524822 106228 568511
rect 106660 568206 106688 568511
rect 106648 568200 106700 568206
rect 106648 568142 106700 568148
rect 107580 524958 107608 568511
rect 107764 568342 107792 568511
rect 107752 568336 107804 568342
rect 107752 568278 107804 568284
rect 108960 525026 108988 568511
rect 109052 568274 109080 570143
rect 110326 568576 110382 568585
rect 110326 568511 110382 568520
rect 110694 568576 110750 568585
rect 110694 568511 110750 568520
rect 111706 568576 111762 568585
rect 111706 568511 111762 568520
rect 110340 568478 110368 568511
rect 110328 568472 110380 568478
rect 109866 568440 109922 568449
rect 110328 568414 110380 568420
rect 109866 568375 109922 568384
rect 109040 568268 109092 568274
rect 109040 568210 109092 568216
rect 109880 567934 109908 568375
rect 110708 568138 110736 568511
rect 110696 568132 110748 568138
rect 110696 568074 110748 568080
rect 109868 567928 109920 567934
rect 109868 567870 109920 567876
rect 110326 567760 110382 567769
rect 110326 567695 110382 567704
rect 110340 567526 110368 567695
rect 110328 567520 110380 567526
rect 110328 567462 110380 567468
rect 110708 567254 110736 568074
rect 110696 567248 110748 567254
rect 110696 567190 110748 567196
rect 111720 525774 111748 568511
rect 112272 568070 112300 570143
rect 113638 569800 113694 569809
rect 113638 569735 113694 569744
rect 112260 568064 112312 568070
rect 112260 568006 112312 568012
rect 113652 567866 113680 569735
rect 114466 569664 114522 569673
rect 114466 569599 114522 569608
rect 117134 569664 117190 569673
rect 117134 569599 117190 569608
rect 113640 567860 113692 567866
rect 113640 567802 113692 567808
rect 111708 525768 111760 525774
rect 111708 525710 111760 525716
rect 108948 525020 109000 525026
rect 108948 524962 109000 524968
rect 107568 524952 107620 524958
rect 107568 524894 107620 524900
rect 106188 524816 106240 524822
rect 106188 524758 106240 524764
rect 103336 524136 103388 524142
rect 103336 524078 103388 524084
rect 109040 524000 109092 524006
rect 109040 523942 109092 523948
rect 107108 523660 107160 523666
rect 107108 523602 107160 523608
rect 103336 523592 103388 523598
rect 103336 523534 103388 523540
rect 103348 521900 103376 523534
rect 105176 523524 105228 523530
rect 105176 523466 105228 523472
rect 105188 521900 105216 523466
rect 107120 521900 107148 523602
rect 109052 521900 109080 523942
rect 114480 523938 114508 569599
rect 114742 568712 114798 568721
rect 114742 568647 114798 568656
rect 114756 568002 114784 568647
rect 115846 568576 115902 568585
rect 115846 568511 115902 568520
rect 115860 568206 115888 568511
rect 117148 568342 117176 569599
rect 117976 568410 118004 570143
rect 118330 569800 118386 569809
rect 118330 569735 118386 569744
rect 118054 568712 118110 568721
rect 118054 568647 118110 568656
rect 117964 568404 118016 568410
rect 117964 568346 118016 568352
rect 117136 568336 117188 568342
rect 117136 568278 117188 568284
rect 117148 568206 117176 568278
rect 115848 568200 115900 568206
rect 115848 568142 115900 568148
rect 117136 568200 117188 568206
rect 117136 568142 117188 568148
rect 114744 567996 114796 568002
rect 114744 567938 114796 567944
rect 118068 567866 118096 568647
rect 118056 567860 118108 567866
rect 118056 567802 118108 567808
rect 118344 567322 118372 569735
rect 119434 569120 119490 569129
rect 119434 569055 119490 569064
rect 119250 568984 119306 568993
rect 119250 568919 119306 568928
rect 119264 568002 119292 568919
rect 119448 568546 119476 569055
rect 119436 568540 119488 568546
rect 119436 568482 119488 568488
rect 119252 567996 119304 568002
rect 119252 567938 119304 567944
rect 118332 567316 118384 567322
rect 118332 567258 118384 567264
rect 118514 566536 118570 566545
rect 118514 566471 118570 566480
rect 118528 524006 118556 566471
rect 120000 525706 120028 570143
rect 120722 569800 120778 569809
rect 120722 569735 120778 569744
rect 120078 569664 120134 569673
rect 120078 569599 120134 569608
rect 120092 568070 120120 569599
rect 120080 568064 120132 568070
rect 120080 568006 120132 568012
rect 120632 567384 120684 567390
rect 120630 567352 120632 567361
rect 120684 567352 120686 567361
rect 120630 567287 120686 567296
rect 120736 567254 120764 569735
rect 120998 569120 121054 569129
rect 120998 569055 121054 569064
rect 121012 568342 121040 569055
rect 122746 568848 122802 568857
rect 122746 568783 122802 568792
rect 121000 568336 121052 568342
rect 121000 568278 121052 568284
rect 121276 567316 121328 567322
rect 121276 567258 121328 567264
rect 120724 567248 120776 567254
rect 120724 567190 120776 567196
rect 119988 525700 120040 525706
rect 119988 525642 120040 525648
rect 120448 524068 120500 524074
rect 120448 524010 120500 524016
rect 118516 524000 118568 524006
rect 118516 523942 118568 523948
rect 110972 523932 111024 523938
rect 110972 523874 111024 523880
rect 114468 523932 114520 523938
rect 114468 523874 114520 523880
rect 110984 521900 111012 523874
rect 114744 523864 114796 523870
rect 114744 523806 114796 523812
rect 112812 523524 112864 523530
rect 112812 523466 112864 523472
rect 112824 521900 112852 523466
rect 114756 521900 114784 523806
rect 116676 523796 116728 523802
rect 116676 523738 116728 523744
rect 116688 521900 116716 523738
rect 118516 523728 118568 523734
rect 118516 523670 118568 523676
rect 118528 521900 118556 523670
rect 120460 521900 120488 524010
rect 120736 523326 120764 567190
rect 121288 524074 121316 567258
rect 122656 567248 122708 567254
rect 122656 567190 122708 567196
rect 122102 566128 122158 566137
rect 122102 566063 122158 566072
rect 121276 524068 121328 524074
rect 121276 524010 121328 524016
rect 120724 523320 120776 523326
rect 120724 523262 120776 523268
rect 122116 523258 122144 566063
rect 122104 523252 122156 523258
rect 122104 523194 122156 523200
rect 122668 521914 122696 567190
rect 122760 523938 122788 568783
rect 126610 568576 126666 568585
rect 126610 568511 126666 568520
rect 128450 568576 128506 568585
rect 128450 568511 128452 568520
rect 124126 568304 124182 568313
rect 124126 568239 124182 568248
rect 124310 568304 124366 568313
rect 124310 568239 124312 568248
rect 124140 568138 124168 568239
rect 124364 568239 124366 568248
rect 125506 568304 125562 568313
rect 126624 568274 126652 568511
rect 128504 568511 128506 568520
rect 132408 568540 132460 568546
rect 128452 568482 128504 568488
rect 132408 568482 132460 568488
rect 125506 568239 125562 568248
rect 126612 568268 126664 568274
rect 124312 568210 124364 568216
rect 123484 568132 123536 568138
rect 123484 568074 123536 568080
rect 124128 568132 124180 568138
rect 124128 568074 124180 568080
rect 123496 567225 123524 568074
rect 125520 567934 125548 568239
rect 126612 568210 126664 568216
rect 128464 568206 128492 568482
rect 128452 568200 128504 568206
rect 128452 568142 128504 568148
rect 125508 567928 125560 567934
rect 125508 567870 125560 567876
rect 124862 567760 124918 567769
rect 124862 567695 124918 567704
rect 124876 567458 124904 567695
rect 124864 567452 124916 567458
rect 124864 567394 124916 567400
rect 127624 567452 127676 567458
rect 127624 567394 127676 567400
rect 128268 567452 128320 567458
rect 128268 567394 128320 567400
rect 123482 567216 123538 567225
rect 123482 567151 123538 567160
rect 122748 523932 122800 523938
rect 122748 523874 122800 523880
rect 123496 523666 123524 567151
rect 124312 523864 124364 523870
rect 124312 523806 124364 523812
rect 123484 523660 123536 523666
rect 123484 523602 123536 523608
rect 122406 521886 122696 521914
rect 124324 521900 124352 523806
rect 124876 523462 124904 567394
rect 125416 567384 125468 567390
rect 125046 567352 125102 567361
rect 125416 567326 125468 567332
rect 125046 567287 125102 567296
rect 124864 523456 124916 523462
rect 124864 523398 124916 523404
rect 125060 523394 125088 567287
rect 125322 567216 125378 567225
rect 125322 567151 125378 567160
rect 125336 523977 125364 567151
rect 125322 523968 125378 523977
rect 125322 523903 125378 523912
rect 125428 523870 125456 567326
rect 127636 567225 127664 567394
rect 126886 567216 126942 567225
rect 126886 567151 126942 567160
rect 127622 567216 127678 567225
rect 127622 567151 127678 567160
rect 128174 567216 128230 567225
rect 128174 567151 128230 567160
rect 125416 523864 125468 523870
rect 126900 523841 126928 567151
rect 125416 523806 125468 523812
rect 126886 523832 126942 523841
rect 126886 523767 126942 523776
rect 126152 523728 126204 523734
rect 126152 523670 126204 523676
rect 125048 523388 125100 523394
rect 125048 523330 125100 523336
rect 126164 521900 126192 523670
rect 127636 523530 127664 567151
rect 128188 525638 128216 567151
rect 128176 525632 128228 525638
rect 128176 525574 128228 525580
rect 127624 523524 127676 523530
rect 127624 523466 127676 523472
rect 128280 521914 128308 567394
rect 130016 523796 130068 523802
rect 130016 523738 130068 523744
rect 128110 521886 128308 521914
rect 130028 521900 130056 523738
rect 132420 521914 132448 568482
rect 135904 568472 135956 568478
rect 135904 568414 135956 568420
rect 133788 523864 133840 523870
rect 133788 523806 133840 523812
rect 131882 521886 132448 521914
rect 133800 521900 133828 523806
rect 135720 523320 135772 523326
rect 135720 523262 135772 523268
rect 135732 521900 135760 523262
rect 135916 523190 135944 568414
rect 137284 568404 137336 568410
rect 137284 568346 137336 568352
rect 137296 523326 137324 568346
rect 140044 568336 140096 568342
rect 140044 568278 140096 568284
rect 145562 568304 145618 568313
rect 138664 567520 138716 567526
rect 138664 567462 138716 567468
rect 137284 523320 137336 523326
rect 137284 523262 137336 523268
rect 137652 523252 137704 523258
rect 137652 523194 137704 523200
rect 135904 523184 135956 523190
rect 135904 523126 135956 523132
rect 137664 521900 137692 523194
rect 138676 523122 138704 567462
rect 140056 523666 140084 568278
rect 144920 568268 144972 568274
rect 145562 568239 145618 568248
rect 144920 568210 144972 568216
rect 144184 568064 144236 568070
rect 144184 568006 144236 568012
rect 142896 567996 142948 568002
rect 142896 567938 142948 567944
rect 142804 567860 142856 567866
rect 142804 567802 142856 567808
rect 139492 523660 139544 523666
rect 139492 523602 139544 523608
rect 140044 523660 140096 523666
rect 140044 523602 140096 523608
rect 138664 523116 138716 523122
rect 138664 523058 138716 523064
rect 139504 521900 139532 523602
rect 141424 523388 141476 523394
rect 141424 523330 141476 523336
rect 141436 521900 141464 523330
rect 142816 523054 142844 567802
rect 142908 523258 142936 567938
rect 143356 523456 143408 523462
rect 143356 523398 143408 523404
rect 142896 523252 142948 523258
rect 142896 523194 142948 523200
rect 142804 523048 142856 523054
rect 142804 522990 142856 522996
rect 143368 521900 143396 523398
rect 144196 523394 144224 568006
rect 144184 523388 144236 523394
rect 144184 523330 144236 523336
rect 144932 521914 144960 568210
rect 145576 524113 145604 568239
rect 149060 568200 149112 568206
rect 149060 568142 149112 568148
rect 146944 568132 146996 568138
rect 146944 568074 146996 568080
rect 145562 524104 145618 524113
rect 145562 524039 145618 524048
rect 146956 523462 146984 568074
rect 147128 523524 147180 523530
rect 147128 523466 147180 523472
rect 146944 523456 146996 523462
rect 146944 523398 146996 523404
rect 144932 521886 145222 521914
rect 147140 521900 147168 523466
rect 149072 521900 149100 568142
rect 152464 567928 152516 567934
rect 152464 567870 152516 567876
rect 150992 524748 151044 524754
rect 150992 524690 151044 524696
rect 151004 521900 151032 524690
rect 152476 524249 152504 567870
rect 155224 567656 155276 567662
rect 155224 567598 155276 567604
rect 153844 567588 153896 567594
rect 153844 567530 153896 567536
rect 153856 524414 153884 567530
rect 155236 524414 155264 567598
rect 156616 524498 156644 655522
rect 188342 654936 188398 654945
rect 188342 654871 188398 654880
rect 156696 567792 156748 567798
rect 156696 567734 156748 567740
rect 156156 524470 156644 524498
rect 152832 524408 152884 524414
rect 152832 524350 152884 524356
rect 153844 524408 153896 524414
rect 153844 524350 153896 524356
rect 154764 524408 154816 524414
rect 154764 524350 154816 524356
rect 155224 524408 155276 524414
rect 155224 524350 155276 524356
rect 152462 524240 152518 524249
rect 152462 524175 152518 524184
rect 152844 521900 152872 524350
rect 154776 521900 154804 524350
rect 155960 523592 156012 523598
rect 156156 523546 156184 524470
rect 156708 524346 156736 567734
rect 156788 567724 156840 567730
rect 156788 567666 156840 567672
rect 156420 524340 156472 524346
rect 156420 524282 156472 524288
rect 156696 524340 156748 524346
rect 156696 524282 156748 524288
rect 156012 523540 156184 523546
rect 155960 523534 156184 523540
rect 155972 523518 156184 523534
rect 156432 521914 156460 524282
rect 156800 524278 156828 567666
rect 181444 525768 181496 525774
rect 181444 525710 181496 525716
rect 175740 525020 175792 525026
rect 175740 524962 175792 524968
rect 173808 524952 173860 524958
rect 173808 524894 173860 524900
rect 170036 524884 170088 524890
rect 170036 524826 170088 524832
rect 158536 524408 158588 524414
rect 158536 524350 158588 524356
rect 162400 524408 162452 524414
rect 162400 524350 162452 524356
rect 156788 524272 156840 524278
rect 156788 524214 156840 524220
rect 156432 521886 156722 521914
rect 158548 521900 158576 524350
rect 160468 523592 160520 523598
rect 160468 523534 160520 523540
rect 160480 521900 160508 523534
rect 162412 521900 162440 524350
rect 166172 524340 166224 524346
rect 166172 524282 166224 524288
rect 164332 524204 164384 524210
rect 164332 524146 164384 524152
rect 164344 521900 164372 524146
rect 166184 521900 166212 524282
rect 168104 524136 168156 524142
rect 168104 524078 168156 524084
rect 168116 521900 168144 524078
rect 170048 521900 170076 524826
rect 171968 524816 172020 524822
rect 171968 524758 172020 524764
rect 171980 521900 172008 524758
rect 173820 521900 173848 524894
rect 175752 521900 175780 524962
rect 177672 523184 177724 523190
rect 177672 523126 177724 523132
rect 177684 521900 177712 523126
rect 179512 523116 179564 523122
rect 179512 523058 179564 523064
rect 179524 521900 179552 523058
rect 181456 521900 181484 525710
rect 188356 525570 188384 654871
rect 188434 653168 188490 653177
rect 188434 653103 188490 653112
rect 188344 525564 188396 525570
rect 188344 525506 188396 525512
rect 188448 525502 188476 653103
rect 188526 652080 188582 652089
rect 188526 652015 188582 652024
rect 188436 525496 188488 525502
rect 188436 525438 188488 525444
rect 188540 525434 188568 652015
rect 188618 650448 188674 650457
rect 188618 650383 188674 650392
rect 188528 525428 188580 525434
rect 188528 525370 188580 525376
rect 188632 525366 188660 650383
rect 188710 649224 188766 649233
rect 188710 649159 188766 649168
rect 188620 525360 188672 525366
rect 188620 525302 188672 525308
rect 188724 525298 188752 649159
rect 188802 647592 188858 647601
rect 188802 647527 188858 647536
rect 188712 525292 188764 525298
rect 188712 525234 188764 525240
rect 188816 525230 188844 647527
rect 188894 589656 188950 589665
rect 188894 589591 188950 589600
rect 188804 525224 188856 525230
rect 188804 525166 188856 525172
rect 188908 525162 188936 589591
rect 202786 570208 202842 570217
rect 202786 570143 202842 570152
rect 220726 570208 220782 570217
rect 220726 570143 220782 570152
rect 238758 570208 238814 570217
rect 238758 570143 238814 570152
rect 195978 568576 196034 568585
rect 195978 568511 196034 568520
rect 197450 568576 197506 568585
rect 197450 568511 197506 568520
rect 202234 568576 202290 568585
rect 202234 568511 202290 568520
rect 194414 568440 194470 568449
rect 194414 568375 194470 568384
rect 194428 567633 194456 568375
rect 194414 567624 194470 567633
rect 194414 567559 194416 567568
rect 194468 567559 194470 567568
rect 194416 567530 194468 567536
rect 194428 567499 194456 567530
rect 194784 525700 194836 525706
rect 194784 525642 194836 525648
rect 188896 525156 188948 525162
rect 188896 525098 188948 525104
rect 185308 524068 185360 524074
rect 185308 524010 185360 524016
rect 183376 523320 183428 523326
rect 183376 523262 183428 523268
rect 183388 521900 183416 523262
rect 185320 521900 185348 524010
rect 191012 524000 191064 524006
rect 191012 523942 191064 523948
rect 189080 523388 189132 523394
rect 189080 523330 189132 523336
rect 187148 523252 187200 523258
rect 187148 523194 187200 523200
rect 187160 521900 187188 523194
rect 189092 521900 189120 523330
rect 191024 521900 191052 523942
rect 192852 523456 192904 523462
rect 192852 523398 192904 523404
rect 192864 521900 192892 523398
rect 194796 521900 194824 525642
rect 195992 525094 196020 568511
rect 195980 525088 196032 525094
rect 195980 525030 196032 525036
rect 197464 523705 197492 568511
rect 202248 568070 202276 568511
rect 202236 568064 202288 568070
rect 202236 568006 202288 568012
rect 202248 567322 202276 568006
rect 202236 567316 202288 567322
rect 202236 567258 202288 567264
rect 202418 523968 202474 523977
rect 198648 523932 198700 523938
rect 202800 523938 202828 570143
rect 217874 569664 217930 569673
rect 217874 569599 217930 569608
rect 204166 568576 204222 568585
rect 204166 568511 204222 568520
rect 204810 568576 204866 568585
rect 204810 568511 204866 568520
rect 205546 568576 205602 568585
rect 205546 568511 205602 568520
rect 207018 568576 207074 568585
rect 207018 568511 207074 568520
rect 209594 568576 209650 568585
rect 209594 568511 209596 568520
rect 203706 568440 203762 568449
rect 203706 568375 203762 568384
rect 203720 568002 203748 568375
rect 203708 567996 203760 568002
rect 203708 567938 203760 567944
rect 203720 567254 203748 567938
rect 203708 567248 203760 567254
rect 203708 567190 203760 567196
rect 204180 524074 204208 568511
rect 204824 567934 204852 568511
rect 204812 567928 204864 567934
rect 204812 567870 204864 567876
rect 204824 567390 204852 567870
rect 204812 567384 204864 567390
rect 204812 567326 204864 567332
rect 204350 524240 204406 524249
rect 204350 524175 204406 524184
rect 204168 524068 204220 524074
rect 204168 524010 204220 524016
rect 202418 523903 202474 523912
rect 202788 523932 202840 523938
rect 198648 523874 198700 523880
rect 197450 523696 197506 523705
rect 196716 523660 196768 523666
rect 197450 523631 197506 523640
rect 196716 523602 196768 523608
rect 196728 521900 196756 523602
rect 198660 521900 198688 523874
rect 200488 523524 200540 523530
rect 200488 523466 200540 523472
rect 200500 521900 200528 523466
rect 202432 521900 202460 523903
rect 202788 523874 202840 523880
rect 204364 521900 204392 524175
rect 205560 524006 205588 568511
rect 207032 567458 207060 568511
rect 209648 568511 209650 568520
rect 211894 568576 211950 568585
rect 211894 568511 211950 568520
rect 213090 568576 213146 568585
rect 213090 568511 213146 568520
rect 214102 568576 214158 568585
rect 214102 568511 214158 568520
rect 215574 568576 215630 568585
rect 215574 568511 215630 568520
rect 217138 568576 217194 568585
rect 217138 568511 217194 568520
rect 209596 568482 209648 568488
rect 209608 568206 209636 568482
rect 209596 568200 209648 568206
rect 209596 568142 209648 568148
rect 211908 568070 211936 568511
rect 211896 568064 211948 568070
rect 211896 568006 211948 568012
rect 213104 568002 213132 568511
rect 213092 567996 213144 568002
rect 213092 567938 213144 567944
rect 214116 567934 214144 568511
rect 215588 568274 215616 568511
rect 217152 568342 217180 568511
rect 217140 568336 217192 568342
rect 217140 568278 217192 568284
rect 215576 568268 215628 568274
rect 215576 568210 215628 568216
rect 214104 567928 214156 567934
rect 214104 567870 214156 567876
rect 208308 567860 208360 567866
rect 208308 567802 208360 567808
rect 208320 567458 208348 567802
rect 207020 567452 207072 567458
rect 207020 567394 207072 567400
rect 208308 567452 208360 567458
rect 208308 567394 208360 567400
rect 209056 567390 209084 567421
rect 209044 567384 209096 567390
rect 209042 567352 209044 567361
rect 209096 567352 209098 567361
rect 211066 567352 211122 567361
rect 209042 567287 209098 567296
rect 210424 567316 210476 567322
rect 206296 567254 206324 567285
rect 206284 567248 206336 567254
rect 206282 567216 206284 567225
rect 206336 567216 206338 567225
rect 206282 567151 206338 567160
rect 206926 567216 206982 567225
rect 206926 567151 206982 567160
rect 208306 567216 208362 567225
rect 208306 567151 208362 567160
rect 205548 524000 205600 524006
rect 205548 523942 205600 523948
rect 206190 523832 206246 523841
rect 206190 523767 206246 523776
rect 206204 521900 206232 523767
rect 206296 523734 206324 567151
rect 206940 523734 206968 567151
rect 208124 525632 208176 525638
rect 208124 525574 208176 525580
rect 206284 523728 206336 523734
rect 206284 523670 206336 523676
rect 206928 523728 206980 523734
rect 206928 523670 206980 523676
rect 208136 521900 208164 525574
rect 208320 524414 208348 567151
rect 208308 524408 208360 524414
rect 208308 524350 208360 524356
rect 209056 523802 209084 567287
rect 211066 567287 211122 567296
rect 210424 567258 210476 567264
rect 210436 567225 210464 567258
rect 209686 567216 209742 567225
rect 209686 567151 209742 567160
rect 210422 567216 210478 567225
rect 210422 567151 210478 567160
rect 210974 567216 211030 567225
rect 210974 567151 211030 567160
rect 209700 524278 209728 567151
rect 209688 524272 209740 524278
rect 209688 524214 209740 524220
rect 210054 524104 210110 524113
rect 210054 524039 210110 524048
rect 209044 523796 209096 523802
rect 209044 523738 209096 523744
rect 210068 521900 210096 524039
rect 210436 523870 210464 567151
rect 210988 523870 211016 567151
rect 211080 524346 211108 567287
rect 215588 567254 215616 568210
rect 217152 567866 217180 568278
rect 217888 568138 217916 569599
rect 218978 568576 219034 568585
rect 218978 568511 219034 568520
rect 218992 568206 219020 568511
rect 220082 568440 220138 568449
rect 220082 568375 220138 568384
rect 218980 568200 219032 568206
rect 218980 568142 219032 568148
rect 217876 568132 217928 568138
rect 217876 568074 217928 568080
rect 217140 567860 217192 567866
rect 217140 567802 217192 567808
rect 217888 567390 217916 568074
rect 220096 567866 220124 568375
rect 220084 567860 220136 567866
rect 220084 567802 220136 567808
rect 217876 567384 217928 567390
rect 217876 567326 217928 567332
rect 217966 567352 218022 567361
rect 220096 567322 220124 567802
rect 217966 567287 218022 567296
rect 220084 567316 220136 567322
rect 215576 567248 215628 567254
rect 212446 567216 212502 567225
rect 212446 567151 212502 567160
rect 213826 567216 213882 567225
rect 213826 567151 213882 567160
rect 215206 567216 215262 567225
rect 215576 567190 215628 567196
rect 216586 567216 216642 567225
rect 215206 567151 215262 567160
rect 216586 567151 216642 567160
rect 217874 567216 217930 567225
rect 217874 567151 217930 567160
rect 211068 524340 211120 524346
rect 211068 524282 211120 524288
rect 212460 524210 212488 567151
rect 213840 524226 213868 567151
rect 212448 524204 212500 524210
rect 213840 524198 213960 524226
rect 212448 524146 212500 524152
rect 213932 524074 213960 524198
rect 213828 524068 213880 524074
rect 213828 524010 213880 524016
rect 213920 524068 213972 524074
rect 213920 524010 213972 524016
rect 211988 523932 212040 523938
rect 211988 523874 212040 523880
rect 210424 523864 210476 523870
rect 210424 523806 210476 523812
rect 210976 523864 211028 523870
rect 210976 523806 211028 523812
rect 212000 521900 212028 523874
rect 213840 521900 213868 524010
rect 215220 523938 215248 567151
rect 216600 524006 216628 567151
rect 215760 524000 215812 524006
rect 215760 523942 215812 523948
rect 216588 524000 216640 524006
rect 216588 523942 216640 523948
rect 215208 523932 215260 523938
rect 215208 523874 215260 523880
rect 215772 521900 215800 523942
rect 217888 523734 217916 567151
rect 217980 523870 218008 567287
rect 220084 567258 220136 567264
rect 219346 567216 219402 567225
rect 219346 567151 219402 567160
rect 217968 523864 218020 523870
rect 217968 523806 218020 523812
rect 219360 523802 219388 567151
rect 219532 524408 219584 524414
rect 219532 524350 219584 524356
rect 219348 523796 219400 523802
rect 219348 523738 219400 523744
rect 217692 523728 217744 523734
rect 217692 523670 217744 523676
rect 217876 523728 217928 523734
rect 217876 523670 217928 523676
rect 217704 521900 217732 523670
rect 219544 521900 219572 524350
rect 220740 523326 220768 570143
rect 221462 568576 221518 568585
rect 221462 568511 221518 568520
rect 222382 568576 222438 568585
rect 222382 568511 222438 568520
rect 223670 568576 223726 568585
rect 223670 568511 223726 568520
rect 225878 568576 225934 568585
rect 225878 568511 225934 568520
rect 226246 568576 226302 568585
rect 226246 568511 226302 568520
rect 227166 568576 227222 568585
rect 227166 568511 227222 568520
rect 227626 568576 227682 568585
rect 227626 568511 227682 568520
rect 228362 568576 228418 568585
rect 228362 568511 228418 568520
rect 229006 568576 229062 568585
rect 229006 568511 229062 568520
rect 229374 568576 229430 568585
rect 229374 568511 229430 568520
rect 230386 568576 230442 568585
rect 230386 568511 230442 568520
rect 231766 568576 231822 568585
rect 231766 568511 231822 568520
rect 233054 568576 233110 568585
rect 233054 568511 233110 568520
rect 234526 568576 234582 568585
rect 234526 568511 234582 568520
rect 235906 568576 235962 568585
rect 235906 568511 235962 568520
rect 237286 568576 237342 568585
rect 237286 568511 237342 568520
rect 238666 568576 238722 568585
rect 238666 568511 238722 568520
rect 221476 568070 221504 568511
rect 221464 568064 221516 568070
rect 221464 568006 221516 568012
rect 222396 568002 222424 568511
rect 222384 567996 222436 568002
rect 222384 567938 222436 567944
rect 223684 567934 223712 568511
rect 225892 568342 225920 568511
rect 226154 568440 226210 568449
rect 226154 568375 226210 568384
rect 225880 568336 225932 568342
rect 224774 568304 224830 568313
rect 225880 568278 225932 568284
rect 224774 568239 224776 568248
rect 224828 568239 224830 568248
rect 224776 568210 224828 568216
rect 223672 567928 223724 567934
rect 223672 567870 223724 567876
rect 222106 567216 222162 567225
rect 222106 567151 222162 567160
rect 223486 567216 223542 567225
rect 223486 567151 223542 567160
rect 224866 567216 224922 567225
rect 224866 567151 224922 567160
rect 221464 524272 221516 524278
rect 221464 524214 221516 524220
rect 220728 523320 220780 523326
rect 220728 523262 220780 523268
rect 221476 521900 221504 524214
rect 222120 523394 222148 567151
rect 223396 524340 223448 524346
rect 223396 524282 223448 524288
rect 222108 523388 222160 523394
rect 222108 523330 222160 523336
rect 223408 521900 223436 524282
rect 223500 523530 223528 567151
rect 223488 523524 223540 523530
rect 223488 523466 223540 523472
rect 224880 523462 224908 567151
rect 225328 524136 225380 524142
rect 225328 524078 225380 524084
rect 224868 523456 224920 523462
rect 224868 523398 224920 523404
rect 225340 521900 225368 524078
rect 226168 523598 226196 568375
rect 226260 523666 226288 568511
rect 227180 568138 227208 568511
rect 227168 568132 227220 568138
rect 227168 568074 227220 568080
rect 227640 524346 227668 568511
rect 228376 568206 228404 568511
rect 228364 568200 228416 568206
rect 228364 568142 228416 568148
rect 229020 524414 229048 568511
rect 229388 567866 229416 568511
rect 229376 567860 229428 567866
rect 229376 567802 229428 567808
rect 229008 524408 229060 524414
rect 229008 524350 229060 524356
rect 227628 524340 227680 524346
rect 227628 524282 227680 524288
rect 230400 524210 230428 568511
rect 230478 568168 230534 568177
rect 230478 568103 230534 568112
rect 230492 568070 230520 568103
rect 230480 568064 230532 568070
rect 230480 568006 230532 568012
rect 231780 524278 231808 568511
rect 231950 568168 232006 568177
rect 231950 568103 232006 568112
rect 231858 568032 231914 568041
rect 231858 567967 231860 567976
rect 231912 567967 231914 567976
rect 231860 567938 231912 567944
rect 231964 567934 231992 568103
rect 231952 567928 232004 567934
rect 231952 567870 232004 567876
rect 231768 524272 231820 524278
rect 231768 524214 231820 524220
rect 227168 524204 227220 524210
rect 227168 524146 227220 524152
rect 230388 524204 230440 524210
rect 230388 524146 230440 524152
rect 226248 523660 226300 523666
rect 226248 523602 226300 523608
rect 226156 523592 226208 523598
rect 226156 523534 226208 523540
rect 227180 521900 227208 524146
rect 229100 524068 229152 524074
rect 229100 524010 229152 524016
rect 229112 521900 229140 524010
rect 232872 524000 232924 524006
rect 232872 523942 232924 523948
rect 231032 523932 231084 523938
rect 231032 523874 231084 523880
rect 231044 521900 231072 523874
rect 232884 521900 232912 523942
rect 233068 523938 233096 568511
rect 233146 568440 233202 568449
rect 233146 568375 233202 568384
rect 233160 524142 233188 568375
rect 233238 568304 233294 568313
rect 233238 568239 233240 568248
rect 233292 568239 233294 568248
rect 233240 568210 233292 568216
rect 233148 524136 233200 524142
rect 233148 524078 233200 524084
rect 234540 524074 234568 568511
rect 234618 568440 234674 568449
rect 234618 568375 234674 568384
rect 234632 568342 234660 568375
rect 234620 568336 234672 568342
rect 234620 568278 234672 568284
rect 234528 524068 234580 524074
rect 234528 524010 234580 524016
rect 235920 524006 235948 568511
rect 235998 568168 236054 568177
rect 235998 568103 236000 568112
rect 236052 568103 236054 568112
rect 236000 568074 236052 568080
rect 235908 524000 235960 524006
rect 235908 523942 235960 523948
rect 237300 523938 237328 568511
rect 237378 568304 237434 568313
rect 237378 568239 237434 568248
rect 237392 568206 237420 568239
rect 237380 568200 237432 568206
rect 237380 568142 237432 568148
rect 233056 523932 233108 523938
rect 233056 523874 233108 523880
rect 237288 523932 237340 523938
rect 237288 523874 237340 523880
rect 238680 523870 238708 568511
rect 238772 567866 238800 570143
rect 240046 568576 240102 568585
rect 240046 568511 240102 568520
rect 238760 567860 238812 567866
rect 238760 567802 238812 567808
rect 240060 523870 240088 568511
rect 252192 567588 252244 567594
rect 252192 567530 252244 567536
rect 252204 561626 252232 567530
rect 252204 561598 252600 561626
rect 252572 557598 252600 561598
rect 252560 557592 252612 557598
rect 252560 557534 252612 557540
rect 257988 557524 258040 557530
rect 257988 557466 258040 557472
rect 258000 555506 258028 557466
rect 258000 555478 258120 555506
rect 258092 551682 258120 555478
rect 258080 551676 258132 551682
rect 258080 551618 258132 551624
rect 259736 551676 259788 551682
rect 259736 551618 259788 551624
rect 259748 549234 259776 551618
rect 259736 549228 259788 549234
rect 259736 549170 259788 549176
rect 261484 549228 261536 549234
rect 261484 549170 261536 549176
rect 261496 541006 261524 549170
rect 261484 541000 261536 541006
rect 261484 540942 261536 540948
rect 263600 540932 263652 540938
rect 263600 540874 263652 540880
rect 263612 538898 263640 540874
rect 263600 538892 263652 538898
rect 263600 538834 263652 538840
rect 272064 538892 272116 538898
rect 272064 538834 272116 538840
rect 272076 534614 272104 538834
rect 272064 534608 272116 534614
rect 272064 534550 272116 534556
rect 273904 534608 273956 534614
rect 273904 534550 273956 534556
rect 253848 524408 253900 524414
rect 253848 524350 253900 524356
rect 252008 524340 252060 524346
rect 252008 524282 252060 524288
rect 234804 523864 234856 523870
rect 234804 523806 234856 523812
rect 238668 523864 238720 523870
rect 238668 523806 238720 523812
rect 240048 523864 240100 523870
rect 240048 523806 240100 523812
rect 234816 521900 234844 523806
rect 238300 523796 238352 523802
rect 238300 523738 238352 523744
rect 236736 523728 236788 523734
rect 236736 523670 236788 523676
rect 236748 521900 236776 523670
rect 238312 521914 238340 523738
rect 250076 523660 250128 523666
rect 250076 523602 250128 523608
rect 248144 523592 248196 523598
rect 248144 523534 248196 523540
rect 244372 523524 244424 523530
rect 244372 523466 244424 523472
rect 242440 523388 242492 523394
rect 242440 523330 242492 523336
rect 240508 523320 240560 523326
rect 240508 523262 240560 523268
rect 238312 521886 238694 521914
rect 240520 521900 240548 523262
rect 242452 521900 242480 523330
rect 244384 521900 244412 523466
rect 246212 523456 246264 523462
rect 246212 523398 246264 523404
rect 246224 521900 246252 523398
rect 248156 521900 248184 523534
rect 250088 521900 250116 523602
rect 252020 521900 252048 524282
rect 253860 521900 253888 524350
rect 257712 524272 257764 524278
rect 257712 524214 257764 524220
rect 255780 524204 255832 524210
rect 255780 524146 255832 524152
rect 255792 521900 255820 524146
rect 257724 521900 257752 524214
rect 259552 524136 259604 524142
rect 259552 524078 259604 524084
rect 259564 521900 259592 524078
rect 263416 524068 263468 524074
rect 263416 524010 263468 524016
rect 261484 524000 261536 524006
rect 261484 523942 261536 523948
rect 261496 521900 261524 523942
rect 263428 521900 263456 524010
rect 267188 523932 267240 523938
rect 267188 523874 267240 523880
rect 265348 523864 265400 523870
rect 265348 523806 265400 523812
rect 265360 521900 265388 523806
rect 267200 521900 267228 523874
rect 273916 523802 273944 534550
rect 269120 523796 269172 523802
rect 269120 523738 269172 523744
rect 273904 523796 273956 523802
rect 273904 523738 273956 523744
rect 275376 523796 275428 523802
rect 275376 523738 275428 523744
rect 269132 521900 269160 523738
rect 271052 523728 271104 523734
rect 271052 523670 271104 523676
rect 271064 521900 271092 523670
rect 273994 520976 274050 520985
rect 273994 520911 274050 520920
rect 273904 516792 273956 516798
rect 273904 516734 273956 516740
rect 273812 516384 273864 516390
rect 273812 516326 273864 516332
rect 273626 515264 273682 515273
rect 273626 515199 273682 515208
rect 273640 514826 273668 515199
rect 273628 514820 273680 514826
rect 273628 514762 273680 514768
rect 273534 511456 273590 511465
rect 273534 511391 273590 511400
rect 273548 510678 273576 511391
rect 273536 510672 273588 510678
rect 273536 510614 273588 510620
rect 273718 507648 273774 507657
rect 273718 507583 273774 507592
rect 273732 506598 273760 507583
rect 273720 506592 273772 506598
rect 273720 506534 273772 506540
rect 273534 505744 273590 505753
rect 273534 505679 273590 505688
rect 273548 505238 273576 505679
rect 273536 505232 273588 505238
rect 273536 505174 273588 505180
rect 273534 503840 273590 503849
rect 273534 503775 273590 503784
rect 273548 495530 273576 503775
rect 273626 501936 273682 501945
rect 273626 501871 273682 501880
rect 273640 501090 273668 501871
rect 273628 501084 273680 501090
rect 273628 501026 273680 501032
rect 273718 500032 273774 500041
rect 273718 499967 273774 499976
rect 273732 499662 273760 499967
rect 273720 499656 273772 499662
rect 273720 499598 273772 499604
rect 273718 498128 273774 498137
rect 273718 498063 273774 498072
rect 273732 496942 273760 498063
rect 273720 496936 273772 496942
rect 273720 496878 273772 496884
rect 273718 496224 273774 496233
rect 273718 496159 273774 496168
rect 273732 495650 273760 496159
rect 273720 495644 273772 495650
rect 273720 495586 273772 495592
rect 273548 495502 273760 495530
rect 273626 494320 273682 494329
rect 273626 494255 273682 494264
rect 273640 494154 273668 494255
rect 273628 494148 273680 494154
rect 273628 494090 273680 494096
rect 273626 492416 273682 492425
rect 273626 492351 273682 492360
rect 273640 491434 273668 492351
rect 273628 491428 273680 491434
rect 273628 491370 273680 491376
rect 273442 490512 273498 490521
rect 273442 490447 273498 490456
rect 273456 490006 273484 490447
rect 273444 490000 273496 490006
rect 273444 489942 273496 489948
rect 273628 488708 273680 488714
rect 273628 488650 273680 488656
rect 273640 488617 273668 488650
rect 273626 488608 273682 488617
rect 273626 488543 273682 488552
rect 273534 486704 273590 486713
rect 273534 486639 273590 486648
rect 273548 485926 273576 486639
rect 273536 485920 273588 485926
rect 273536 485862 273588 485868
rect 273626 484800 273682 484809
rect 273626 484735 273682 484744
rect 273640 484498 273668 484735
rect 273628 484492 273680 484498
rect 273628 484434 273680 484440
rect 273626 482896 273682 482905
rect 273626 482831 273682 482840
rect 273640 481778 273668 482831
rect 273628 481772 273680 481778
rect 273628 481714 273680 481720
rect 273626 480992 273682 481001
rect 273626 480927 273682 480936
rect 273640 480350 273668 480927
rect 273628 480344 273680 480350
rect 273628 480286 273680 480292
rect 273626 479088 273682 479097
rect 273626 479023 273682 479032
rect 273640 478922 273668 479023
rect 273628 478916 273680 478922
rect 273628 478858 273680 478864
rect 273626 477184 273682 477193
rect 273626 477119 273682 477128
rect 273640 476134 273668 477119
rect 273628 476128 273680 476134
rect 273628 476070 273680 476076
rect 273626 475280 273682 475289
rect 273626 475215 273682 475224
rect 273640 474842 273668 475215
rect 273628 474836 273680 474842
rect 273628 474778 273680 474784
rect 273536 474020 273588 474026
rect 273536 473962 273588 473968
rect 273548 472274 273576 473962
rect 273628 473408 273680 473414
rect 273626 473376 273628 473385
rect 273680 473376 273682 473385
rect 273626 473311 273682 473320
rect 273548 472246 273668 472274
rect 273444 472048 273496 472054
rect 273444 471990 273496 471996
rect 273352 470620 273404 470626
rect 273352 470562 273404 470568
rect 273258 463856 273314 463865
rect 273258 463791 273314 463800
rect 273272 463758 273300 463791
rect 273260 463752 273312 463758
rect 273260 463694 273312 463700
rect 273258 461952 273314 461961
rect 273258 461887 273314 461896
rect 273272 460970 273300 461887
rect 273260 460964 273312 460970
rect 273260 460906 273312 460912
rect 273260 460080 273312 460086
rect 273258 460048 273260 460057
rect 273312 460048 273314 460057
rect 273258 459983 273314 459992
rect 273260 458176 273312 458182
rect 273258 458144 273260 458153
rect 273312 458144 273314 458153
rect 273258 458079 273314 458088
rect 273260 456272 273312 456278
rect 273258 456240 273260 456249
rect 273312 456240 273314 456249
rect 273258 456175 273314 456184
rect 273260 454368 273312 454374
rect 273258 454336 273260 454345
rect 273312 454336 273314 454345
rect 273258 454271 273314 454280
rect 273260 452464 273312 452470
rect 273258 452432 273260 452441
rect 273312 452432 273314 452441
rect 273258 452367 273314 452376
rect 273364 450537 273392 470562
rect 273350 450528 273406 450537
rect 273350 450463 273406 450472
rect 273456 448633 273484 471990
rect 273534 471472 273590 471481
rect 273534 471407 273590 471416
rect 273548 470694 273576 471407
rect 273536 470688 273588 470694
rect 273536 470630 273588 470636
rect 273534 469568 273590 469577
rect 273534 469503 273590 469512
rect 273548 469334 273576 469503
rect 273536 469328 273588 469334
rect 273536 469270 273588 469276
rect 273534 467664 273590 467673
rect 273534 467599 273590 467608
rect 273548 466546 273576 467599
rect 273536 466540 273588 466546
rect 273536 466482 273588 466488
rect 273534 465760 273590 465769
rect 273534 465695 273590 465704
rect 273442 448624 273498 448633
rect 273442 448559 273498 448568
rect 273444 447092 273496 447098
rect 273444 447034 273496 447040
rect 273456 446729 273484 447034
rect 273442 446720 273498 446729
rect 273442 446655 273498 446664
rect 273444 444848 273496 444854
rect 273442 444816 273444 444825
rect 273496 444816 273498 444825
rect 273442 444751 273498 444760
rect 273444 442944 273496 442950
rect 273442 442912 273444 442921
rect 273496 442912 273498 442921
rect 273442 442847 273498 442856
rect 273444 441312 273496 441318
rect 273444 441254 273496 441260
rect 273456 441017 273484 441254
rect 273442 441008 273498 441017
rect 273442 440943 273498 440952
rect 273444 439748 273496 439754
rect 273444 439690 273496 439696
rect 273456 439113 273484 439690
rect 273442 439104 273498 439113
rect 273442 439039 273498 439048
rect 273260 433424 273312 433430
rect 273258 433392 273260 433401
rect 273312 433392 273314 433401
rect 273258 433327 273314 433336
rect 273260 431520 273312 431526
rect 273258 431488 273260 431497
rect 273312 431488 273314 431497
rect 273258 431423 273314 431432
rect 273260 429616 273312 429622
rect 273258 429584 273260 429593
rect 273312 429584 273314 429593
rect 273258 429519 273314 429528
rect 273260 427712 273312 427718
rect 273258 427680 273260 427689
rect 273312 427680 273314 427689
rect 273258 427615 273314 427624
rect 273260 425808 273312 425814
rect 273258 425776 273260 425785
rect 273312 425776 273314 425785
rect 273258 425711 273314 425720
rect 273444 424040 273496 424046
rect 273444 423982 273496 423988
rect 273456 423881 273484 423982
rect 273442 423872 273498 423881
rect 273442 423807 273498 423816
rect 273444 422068 273496 422074
rect 273444 422010 273496 422016
rect 273456 421977 273484 422010
rect 273442 421968 273498 421977
rect 273442 421903 273498 421912
rect 273444 420096 273496 420102
rect 273442 420064 273444 420073
rect 273496 420064 273498 420073
rect 273442 419999 273498 420008
rect 273442 418160 273498 418169
rect 273442 418095 273444 418104
rect 273496 418095 273498 418104
rect 273444 418066 273496 418072
rect 273444 416288 273496 416294
rect 273442 416256 273444 416265
rect 273496 416256 273498 416265
rect 273442 416191 273498 416200
rect 273444 414384 273496 414390
rect 273442 414352 273444 414361
rect 273496 414352 273498 414361
rect 273442 414287 273498 414296
rect 273444 412480 273496 412486
rect 273442 412448 273444 412457
rect 273496 412448 273498 412457
rect 273442 412383 273498 412392
rect 273444 410576 273496 410582
rect 273442 410544 273444 410553
rect 273496 410544 273498 410553
rect 273442 410479 273498 410488
rect 273444 408672 273496 408678
rect 273442 408640 273444 408649
rect 273496 408640 273498 408649
rect 273442 408575 273498 408584
rect 273444 406768 273496 406774
rect 273442 406736 273444 406745
rect 273496 406736 273498 406745
rect 273442 406671 273498 406680
rect 273444 402960 273496 402966
rect 273442 402928 273444 402937
rect 273496 402928 273498 402937
rect 273442 402863 273498 402872
rect 273444 401056 273496 401062
rect 273442 401024 273444 401033
rect 273496 401024 273498 401033
rect 273442 400959 273498 400968
rect 273444 400172 273496 400178
rect 273444 400114 273496 400120
rect 273456 399129 273484 400114
rect 273442 399120 273498 399129
rect 273442 399055 273498 399064
rect 273444 397452 273496 397458
rect 273444 397394 273496 397400
rect 273456 397225 273484 397394
rect 273442 397216 273498 397225
rect 273442 397151 273498 397160
rect 273260 396840 273312 396846
rect 273260 396782 273312 396788
rect 273272 336297 273300 396782
rect 273444 396024 273496 396030
rect 273444 395966 273496 395972
rect 273456 395321 273484 395966
rect 273442 395312 273498 395321
rect 273442 395247 273498 395256
rect 273444 394664 273496 394670
rect 273444 394606 273496 394612
rect 273456 393417 273484 394606
rect 273442 393408 273498 393417
rect 273442 393343 273498 393352
rect 273444 391944 273496 391950
rect 273444 391886 273496 391892
rect 273456 391513 273484 391886
rect 273442 391504 273498 391513
rect 273442 391439 273498 391448
rect 273548 390674 273576 465695
rect 273456 390646 273576 390674
rect 273456 389450 273484 390646
rect 273536 390516 273588 390522
rect 273536 390458 273588 390464
rect 273548 389609 273576 390458
rect 273534 389600 273590 389609
rect 273534 389535 273590 389544
rect 273456 389422 273576 389450
rect 273444 389224 273496 389230
rect 273444 389166 273496 389172
rect 273352 388068 273404 388074
rect 273352 388010 273404 388016
rect 273364 385014 273392 388010
rect 273352 385008 273404 385014
rect 273352 384950 273404 384956
rect 273456 383874 273484 389166
rect 273548 388074 273576 389422
rect 273536 388068 273588 388074
rect 273536 388010 273588 388016
rect 273640 387954 273668 472246
rect 273548 387926 273668 387954
rect 273548 385801 273576 387926
rect 273628 387796 273680 387802
rect 273628 387738 273680 387744
rect 273640 387705 273668 387738
rect 273626 387696 273682 387705
rect 273626 387631 273682 387640
rect 273628 387592 273680 387598
rect 273628 387534 273680 387540
rect 273534 385792 273590 385801
rect 273534 385727 273590 385736
rect 273364 383846 273484 383874
rect 273364 383586 273392 383846
rect 273352 383580 273404 383586
rect 273352 383522 273404 383528
rect 273640 383466 273668 387534
rect 273364 383438 273668 383466
rect 273258 336288 273314 336297
rect 273258 336223 273314 336232
rect 273364 331362 273392 383438
rect 273444 383376 273496 383382
rect 273444 383318 273496 383324
rect 273352 331356 273404 331362
rect 273352 331298 273404 331304
rect 273352 331220 273404 331226
rect 273352 331162 273404 331168
rect 273364 330585 273392 331162
rect 273350 330576 273406 330585
rect 273350 330511 273406 330520
rect 273456 324873 273484 383318
rect 273534 381984 273590 381993
rect 273534 381919 273590 381928
rect 273548 380254 273576 381919
rect 273626 380352 273682 380361
rect 273626 380287 273682 380296
rect 273536 380248 273588 380254
rect 273536 380190 273588 380196
rect 273640 380186 273668 380287
rect 273628 380180 273680 380186
rect 273628 380122 273680 380128
rect 273536 378956 273588 378962
rect 273536 378898 273588 378904
rect 273548 374542 273576 378898
rect 273628 374672 273680 374678
rect 273628 374614 273680 374620
rect 273536 374536 273588 374542
rect 273536 374478 273588 374484
rect 273640 368665 273668 374614
rect 273626 368656 273682 368665
rect 273626 368591 273682 368600
rect 273732 362914 273760 495502
rect 273824 374678 273852 516326
rect 273812 374672 273864 374678
rect 273812 374614 273864 374620
rect 273812 374536 273864 374542
rect 273812 374478 273864 374484
rect 273824 364857 273852 374478
rect 273810 364848 273866 364857
rect 273810 364783 273866 364792
rect 273720 362908 273772 362914
rect 273720 362850 273772 362856
rect 273536 361072 273588 361078
rect 273534 361040 273536 361049
rect 273588 361040 273590 361049
rect 273534 360975 273590 360984
rect 273812 359712 273864 359718
rect 273812 359654 273864 359660
rect 273824 359145 273852 359654
rect 273810 359136 273866 359145
rect 273810 359071 273866 359080
rect 273812 353456 273864 353462
rect 273810 353424 273812 353433
rect 273864 353424 273866 353433
rect 273810 353359 273866 353368
rect 273536 349648 273588 349654
rect 273534 349616 273536 349625
rect 273588 349616 273590 349625
rect 273534 349551 273590 349560
rect 273536 347744 273588 347750
rect 273534 347712 273536 347721
rect 273588 347712 273590 347721
rect 273534 347647 273590 347656
rect 273536 345908 273588 345914
rect 273536 345850 273588 345856
rect 273548 345817 273576 345850
rect 273534 345808 273590 345817
rect 273534 345743 273590 345752
rect 273628 344004 273680 344010
rect 273628 343946 273680 343952
rect 273640 343913 273668 343946
rect 273626 343904 273682 343913
rect 273626 343839 273682 343848
rect 273536 342168 273588 342174
rect 273536 342110 273588 342116
rect 273548 342009 273576 342110
rect 273534 342000 273590 342009
rect 273534 341935 273590 341944
rect 273536 340128 273588 340134
rect 273534 340096 273536 340105
rect 273588 340096 273590 340105
rect 273534 340031 273590 340040
rect 273916 338201 273944 516734
rect 274008 346390 274036 520911
rect 274270 519072 274326 519081
rect 275388 519042 275416 523738
rect 274270 519007 274326 519016
rect 275376 519036 275428 519042
rect 274284 518974 274312 519007
rect 275376 518978 275428 518984
rect 278780 519036 278832 519042
rect 278780 518978 278832 518984
rect 274272 518968 274324 518974
rect 274272 518910 274324 518916
rect 274086 517168 274142 517177
rect 274086 517103 274142 517112
rect 274100 349110 274128 517103
rect 278792 517070 278820 518978
rect 301504 518968 301556 518974
rect 301504 518910 301556 518916
rect 278780 517064 278832 517070
rect 278780 517006 278832 517012
rect 280068 517064 280120 517070
rect 280068 517006 280120 517012
rect 280080 516866 280108 517006
rect 280068 516860 280120 516866
rect 280068 516802 280120 516808
rect 275376 516724 275428 516730
rect 275376 516666 275428 516672
rect 274364 516588 274416 516594
rect 274364 516530 274416 516536
rect 274178 513360 274234 513369
rect 274178 513295 274234 513304
rect 274192 350470 274220 513295
rect 274270 509552 274326 509561
rect 274270 509487 274326 509496
rect 274284 353258 274312 509487
rect 274376 362953 274404 516530
rect 274456 516520 274508 516526
rect 274456 516462 274508 516468
rect 274468 378962 274496 516462
rect 274548 516452 274600 516458
rect 274548 516394 274600 516400
rect 274456 378956 274508 378962
rect 274456 378898 274508 378904
rect 274456 378820 274508 378826
rect 274456 378762 274508 378768
rect 274468 378185 274496 378762
rect 274454 378176 274510 378185
rect 274454 378111 274510 378120
rect 274454 376272 274510 376281
rect 274454 376207 274510 376216
rect 274468 376038 274496 376207
rect 274456 376032 274508 376038
rect 274456 375974 274508 375980
rect 274456 374672 274508 374678
rect 274456 374614 274508 374620
rect 274468 374377 274496 374614
rect 274454 374368 274510 374377
rect 274454 374303 274510 374312
rect 274454 372464 274510 372473
rect 274454 372399 274510 372408
rect 274468 371890 274496 372399
rect 274456 371884 274508 371890
rect 274456 371826 274508 371832
rect 274454 370560 274510 370569
rect 274454 370495 274456 370504
rect 274508 370495 274510 370504
rect 274456 370466 274508 370472
rect 274560 366761 274588 516394
rect 275284 512032 275336 512038
rect 275284 511974 275336 511980
rect 275192 491360 275244 491366
rect 275192 491302 275244 491308
rect 275100 489932 275152 489938
rect 275100 489874 275152 489880
rect 275008 488640 275060 488646
rect 275008 488582 275060 488588
rect 274916 488572 274968 488578
rect 274916 488514 274968 488520
rect 274824 487212 274876 487218
rect 274824 487154 274876 487160
rect 274732 485852 274784 485858
rect 274732 485794 274784 485800
rect 274640 484424 274692 484430
rect 274640 484366 274692 484372
rect 274652 437209 274680 484366
rect 274638 437200 274694 437209
rect 274638 437135 274694 437144
rect 274744 435305 274772 485794
rect 274730 435296 274786 435305
rect 274730 435231 274786 435240
rect 274836 433430 274864 487154
rect 274824 433424 274876 433430
rect 274824 433366 274876 433372
rect 274928 431526 274956 488514
rect 274916 431520 274968 431526
rect 274916 431462 274968 431468
rect 275020 429622 275048 488582
rect 275008 429616 275060 429622
rect 275008 429558 275060 429564
rect 275112 427718 275140 489874
rect 275100 427712 275152 427718
rect 275100 427654 275152 427660
rect 275204 425814 275232 491302
rect 275192 425808 275244 425814
rect 275192 425750 275244 425756
rect 275192 396636 275244 396642
rect 275192 396578 275244 396584
rect 275100 396568 275152 396574
rect 275100 396510 275152 396516
rect 275008 396500 275060 396506
rect 275008 396442 275060 396448
rect 274916 396432 274968 396438
rect 274916 396374 274968 396380
rect 274824 396364 274876 396370
rect 274824 396306 274876 396312
rect 274638 383888 274694 383897
rect 274638 383823 274694 383832
rect 274652 378894 274680 383823
rect 274640 378888 274692 378894
rect 274640 378830 274692 378836
rect 274546 366752 274602 366761
rect 274546 366687 274602 366696
rect 274362 362944 274418 362953
rect 274362 362879 274418 362888
rect 274364 355972 274416 355978
rect 274364 355914 274416 355920
rect 274376 355337 274404 355914
rect 274362 355328 274418 355337
rect 274362 355263 274418 355272
rect 274836 353462 274864 396306
rect 274824 353456 274876 353462
rect 274824 353398 274876 353404
rect 274272 353252 274324 353258
rect 274272 353194 274324 353200
rect 274928 351642 274956 396374
rect 274560 351614 274956 351642
rect 274560 351529 274588 351614
rect 274546 351520 274602 351529
rect 274546 351455 274602 351464
rect 274180 350464 274232 350470
rect 274180 350406 274232 350412
rect 275020 349654 275048 396442
rect 275008 349648 275060 349654
rect 275008 349590 275060 349596
rect 274088 349104 274140 349110
rect 274088 349046 274140 349052
rect 275112 347750 275140 396510
rect 275100 347744 275152 347750
rect 275100 347686 275152 347692
rect 273996 346384 274048 346390
rect 273996 346326 274048 346332
rect 275204 345914 275232 396578
rect 275296 355978 275324 511974
rect 275388 359718 275416 516666
rect 275468 516656 275520 516662
rect 275468 516598 275520 516604
rect 275480 361078 275508 516598
rect 279424 509312 279476 509318
rect 279424 509254 279476 509260
rect 275560 506524 275612 506530
rect 275560 506466 275612 506472
rect 275572 401062 275600 506466
rect 275652 505164 275704 505170
rect 275652 505106 275704 505112
rect 275664 402966 275692 505106
rect 276664 503736 276716 503742
rect 276664 503678 276716 503684
rect 275744 495508 275796 495514
rect 275744 495450 275796 495456
rect 275756 420102 275784 495450
rect 275836 494080 275888 494086
rect 275836 494022 275888 494028
rect 275848 422074 275876 494022
rect 275928 492720 275980 492726
rect 275928 492662 275980 492668
rect 275940 424046 275968 492662
rect 276572 480276 276624 480282
rect 276572 480218 276624 480224
rect 276480 474768 276532 474774
rect 276480 474710 276532 474716
rect 276388 469260 276440 469266
rect 276388 469202 276440 469208
rect 276296 467968 276348 467974
rect 276296 467910 276348 467916
rect 276204 467900 276256 467906
rect 276204 467842 276256 467848
rect 276112 466472 276164 466478
rect 276112 466414 276164 466420
rect 276020 465112 276072 465118
rect 276020 465054 276072 465060
rect 276032 460086 276060 465054
rect 276020 460080 276072 460086
rect 276020 460022 276072 460028
rect 276124 458182 276152 466414
rect 276112 458176 276164 458182
rect 276112 458118 276164 458124
rect 276216 456278 276244 467842
rect 276204 456272 276256 456278
rect 276204 456214 276256 456220
rect 276308 454374 276336 467910
rect 276296 454368 276348 454374
rect 276296 454310 276348 454316
rect 276400 452470 276428 469202
rect 276388 452464 276440 452470
rect 276388 452406 276440 452412
rect 276492 444854 276520 474710
rect 276480 444848 276532 444854
rect 276480 444790 276532 444796
rect 276584 442950 276612 480218
rect 276572 442944 276624 442950
rect 276572 442886 276624 442892
rect 275928 424040 275980 424046
rect 275928 423982 275980 423988
rect 275836 422068 275888 422074
rect 275836 422010 275888 422016
rect 275744 420096 275796 420102
rect 275744 420038 275796 420044
rect 276676 406774 276704 503678
rect 276756 502512 276808 502518
rect 276756 502454 276808 502460
rect 276768 408678 276796 502454
rect 276848 501016 276900 501022
rect 276848 500958 276900 500964
rect 276860 410582 276888 500958
rect 276940 499588 276992 499594
rect 276940 499530 276992 499536
rect 276952 412486 276980 499530
rect 277032 498228 277084 498234
rect 277032 498170 277084 498176
rect 277044 414390 277072 498170
rect 278596 496868 278648 496874
rect 278596 496810 278648 496816
rect 278044 494148 278096 494154
rect 278044 494090 278096 494096
rect 277216 483064 277268 483070
rect 277216 483006 277268 483012
rect 277124 463752 277176 463758
rect 277124 463694 277176 463700
rect 277032 414384 277084 414390
rect 277032 414326 277084 414332
rect 276940 412480 276992 412486
rect 276940 412422 276992 412428
rect 276848 410576 276900 410582
rect 276848 410518 276900 410524
rect 276756 408672 276808 408678
rect 276756 408614 276808 408620
rect 276664 406768 276716 406774
rect 276664 406710 276716 406716
rect 275652 402960 275704 402966
rect 275652 402902 275704 402908
rect 275560 401056 275612 401062
rect 275560 400998 275612 401004
rect 275744 396772 275796 396778
rect 275744 396714 275796 396720
rect 275560 392012 275612 392018
rect 275560 391954 275612 391960
rect 275468 361072 275520 361078
rect 275468 361014 275520 361020
rect 275376 359712 275428 359718
rect 275376 359654 275428 359660
rect 275284 355972 275336 355978
rect 275284 355914 275336 355920
rect 275192 345908 275244 345914
rect 275192 345850 275244 345856
rect 273902 338192 273958 338201
rect 273902 338127 273958 338136
rect 273812 335300 273864 335306
rect 273812 335242 273864 335248
rect 273824 334393 273852 335242
rect 273810 334384 273866 334393
rect 273810 334319 273866 334328
rect 274272 332512 274324 332518
rect 274270 332480 274272 332489
rect 274324 332480 274326 332489
rect 274270 332415 274326 332424
rect 273536 331356 273588 331362
rect 273536 331298 273588 331304
rect 273548 326777 273576 331298
rect 273996 329792 274048 329798
rect 273996 329734 274048 329740
rect 274008 328681 274036 329734
rect 273994 328672 274050 328681
rect 273994 328607 274050 328616
rect 273534 326768 273590 326777
rect 273534 326703 273590 326712
rect 273442 324864 273498 324873
rect 273442 324799 273498 324808
rect 273536 323332 273588 323338
rect 273536 323274 273588 323280
rect 273548 322969 273576 323274
rect 273534 322960 273590 322969
rect 273534 322895 273590 322904
rect 275572 321298 275600 391954
rect 275652 390584 275704 390590
rect 275652 390526 275704 390532
rect 275664 323338 275692 390526
rect 275756 342174 275784 396714
rect 275928 396704 275980 396710
rect 275928 396646 275980 396652
rect 275836 392080 275888 392086
rect 275836 392022 275888 392028
rect 275744 342168 275796 342174
rect 275744 342110 275796 342116
rect 275848 340134 275876 392022
rect 275940 344010 275968 396646
rect 277136 386374 277164 463694
rect 277228 439754 277256 483006
rect 277308 481704 277360 481710
rect 277308 481646 277360 481652
rect 277320 441318 277348 481646
rect 277308 441312 277360 441318
rect 277308 441254 277360 441260
rect 277216 439748 277268 439754
rect 277216 439690 277268 439696
rect 277124 386368 277176 386374
rect 277124 386310 277176 386316
rect 278056 368490 278084 494090
rect 278136 488708 278188 488714
rect 278136 488650 278188 488656
rect 278148 371210 278176 488650
rect 278228 485920 278280 485926
rect 278228 485862 278280 485868
rect 278240 372570 278268 485862
rect 278320 484492 278372 484498
rect 278320 484434 278372 484440
rect 278332 373998 278360 484434
rect 278412 481772 278464 481778
rect 278412 481714 278464 481720
rect 278424 375358 278452 481714
rect 278504 480344 278556 480350
rect 278504 480286 278556 480292
rect 278516 381154 278544 480286
rect 278608 416294 278636 496810
rect 278688 460964 278740 460970
rect 278688 460906 278740 460912
rect 278596 416288 278648 416294
rect 278596 416230 278648 416236
rect 278700 387734 278728 460906
rect 278688 387728 278740 387734
rect 278688 387670 278740 387676
rect 278516 381126 278636 381154
rect 278608 376718 278636 381126
rect 278596 376712 278648 376718
rect 278596 376654 278648 376660
rect 278412 375352 278464 375358
rect 278412 375294 278464 375300
rect 278320 373992 278372 373998
rect 278320 373934 278372 373940
rect 278228 372564 278280 372570
rect 278228 372506 278280 372512
rect 278136 371204 278188 371210
rect 278136 371146 278188 371152
rect 278044 368484 278096 368490
rect 278044 368426 278096 368432
rect 275928 344004 275980 344010
rect 275928 343946 275980 343952
rect 275836 340128 275888 340134
rect 275836 340070 275888 340076
rect 279436 332518 279464 509254
rect 279516 495576 279568 495582
rect 279516 495518 279568 495524
rect 279528 418130 279556 495518
rect 279516 418124 279568 418130
rect 279516 418066 279568 418072
rect 280080 396137 280108 516802
rect 298744 514820 298796 514826
rect 298744 514762 298796 514768
rect 297364 510672 297416 510678
rect 297364 510614 297416 510620
rect 294604 506592 294656 506598
rect 294604 506534 294656 506540
rect 291844 505232 291896 505238
rect 291844 505174 291896 505180
rect 290464 501084 290516 501090
rect 290464 501026 290516 501032
rect 287704 499656 287756 499662
rect 287704 499598 287756 499604
rect 286324 496936 286376 496942
rect 286324 496878 286376 496884
rect 284944 495644 284996 495650
rect 284944 495586 284996 495592
rect 283564 491428 283616 491434
rect 283564 491370 283616 491376
rect 280804 490000 280856 490006
rect 280804 489942 280856 489948
rect 280066 396128 280122 396137
rect 280066 396063 280122 396072
rect 280816 369850 280844 489942
rect 280804 369844 280856 369850
rect 280804 369786 280856 369792
rect 283576 369782 283604 491370
rect 283564 369776 283616 369782
rect 283564 369718 283616 369724
rect 284956 366926 284984 495586
rect 284944 366920 284996 366926
rect 284944 366862 284996 366868
rect 286336 365702 286364 496878
rect 286324 365696 286376 365702
rect 286324 365638 286376 365644
rect 287716 364342 287744 499598
rect 287704 364336 287756 364342
rect 287704 364278 287756 364284
rect 290476 362846 290504 501026
rect 290464 362840 290516 362846
rect 290464 362782 290516 362788
rect 291856 356046 291884 505174
rect 291844 356040 291896 356046
rect 291844 355982 291896 355988
rect 294616 354686 294644 506534
rect 294604 354680 294656 354686
rect 294604 354622 294656 354628
rect 297376 351898 297404 510614
rect 297364 351892 297416 351898
rect 297364 351834 297416 351840
rect 298756 349042 298784 514762
rect 298744 349036 298796 349042
rect 298744 348978 298796 348984
rect 301516 347750 301544 518910
rect 337750 517440 337806 517449
rect 337750 517375 337806 517384
rect 320180 516860 320232 516866
rect 320180 516802 320232 516808
rect 320192 516769 320220 516802
rect 337764 516798 337792 517375
rect 337752 516792 337804 516798
rect 320178 516760 320234 516769
rect 337752 516734 337804 516740
rect 338396 516792 338448 516798
rect 338396 516734 338448 516740
rect 340880 516792 340932 516798
rect 340880 516734 340932 516740
rect 398838 516760 398894 516769
rect 320178 516695 320234 516704
rect 338408 516497 338436 516734
rect 340892 516497 340920 516734
rect 398838 516695 398840 516704
rect 398892 516695 398894 516704
rect 398840 516666 398892 516672
rect 400220 516656 400272 516662
rect 400218 516624 400220 516633
rect 400272 516624 400274 516633
rect 400218 516559 400274 516568
rect 401598 516624 401654 516633
rect 401598 516559 401600 516568
rect 401652 516559 401654 516568
rect 401600 516530 401652 516536
rect 403348 516520 403400 516526
rect 338394 516488 338450 516497
rect 338394 516423 338450 516432
rect 340878 516488 340934 516497
rect 340878 516423 340934 516432
rect 403346 516488 403348 516497
rect 403400 516488 403402 516497
rect 403346 516423 403402 516432
rect 404358 516488 404414 516497
rect 404358 516423 404360 516432
rect 404412 516423 404414 516432
rect 406014 516488 406070 516497
rect 406014 516423 406016 516432
rect 404360 516394 404412 516400
rect 406068 516423 406070 516432
rect 406016 516394 406068 516400
rect 320178 512136 320234 512145
rect 320178 512071 320234 512080
rect 320192 512038 320220 512071
rect 320180 512032 320232 512038
rect 320180 511974 320232 511980
rect 320364 509312 320416 509318
rect 320364 509254 320416 509260
rect 316682 509144 316738 509153
rect 316682 509079 316738 509088
rect 302884 507884 302936 507890
rect 302884 507826 302936 507832
rect 301504 347744 301556 347750
rect 301504 347686 301556 347692
rect 302896 335306 302924 507826
rect 315304 478916 315356 478922
rect 315304 478858 315356 478864
rect 312544 476128 312596 476134
rect 312544 476070 312596 476076
rect 309784 474836 309836 474842
rect 309784 474778 309836 474784
rect 308404 473408 308456 473414
rect 308404 473350 308456 473356
rect 305644 470688 305696 470694
rect 305644 470630 305696 470636
rect 304264 469328 304316 469334
rect 304264 469270 304316 469276
rect 302976 466540 303028 466546
rect 302976 466482 303028 466488
rect 302988 384946 303016 466482
rect 302976 384940 303028 384946
rect 302976 384882 303028 384888
rect 304276 383654 304304 469270
rect 304264 383648 304316 383654
rect 304264 383590 304316 383596
rect 305656 382226 305684 470630
rect 305644 382220 305696 382226
rect 305644 382162 305696 382168
rect 308416 380866 308444 473350
rect 308404 380860 308456 380866
rect 308404 380802 308456 380808
rect 309796 379506 309824 474778
rect 309784 379500 309836 379506
rect 309784 379442 309836 379448
rect 312556 376786 312584 476070
rect 315316 376854 315344 478858
rect 315304 376848 315356 376854
rect 315304 376790 315356 376796
rect 312544 376780 312596 376786
rect 312544 376722 312596 376728
rect 302884 335300 302936 335306
rect 302884 335242 302936 335248
rect 279424 332512 279476 332518
rect 279424 332454 279476 332460
rect 316696 329798 316724 509079
rect 319442 507920 319498 507929
rect 319442 507855 319498 507864
rect 320180 507884 320232 507890
rect 318800 366308 318852 366314
rect 318800 366250 318852 366256
rect 318812 363497 318840 366250
rect 318798 363488 318854 363497
rect 318798 363423 318854 363432
rect 319456 331226 319484 507855
rect 320180 507826 320232 507832
rect 319812 506524 319864 506530
rect 319812 506466 319864 506472
rect 319824 506297 319852 506466
rect 320192 506297 320220 507826
rect 320376 507521 320404 509254
rect 320362 507512 320418 507521
rect 320362 507447 320418 507456
rect 319810 506288 319866 506297
rect 319810 506223 319866 506232
rect 320178 506288 320234 506297
rect 320178 506223 320234 506232
rect 320180 505164 320232 505170
rect 320180 505106 320232 505112
rect 319996 503736 320048 503742
rect 319996 503678 320048 503684
rect 319812 501016 319864 501022
rect 319810 500984 319812 500993
rect 319864 500984 319866 500993
rect 319810 500919 319866 500928
rect 320008 500857 320036 503678
rect 320192 503169 320220 505106
rect 320730 504792 320786 504801
rect 320730 504727 320786 504736
rect 320546 503704 320602 503713
rect 320546 503639 320602 503648
rect 320178 503160 320234 503169
rect 320178 503095 320234 503104
rect 320272 502580 320324 502586
rect 320272 502522 320324 502528
rect 319994 500848 320050 500857
rect 319994 500783 320050 500792
rect 320284 499633 320312 502522
rect 320362 502480 320418 502489
rect 320362 502415 320418 502424
rect 320270 499624 320326 499633
rect 320180 499588 320232 499594
rect 320270 499559 320326 499568
rect 320180 499530 320232 499536
rect 319812 498228 319864 498234
rect 319812 498170 319864 498176
rect 319824 498001 319852 498170
rect 319810 497992 319866 498001
rect 319810 497927 319866 497936
rect 320192 497321 320220 499530
rect 320270 497856 320326 497865
rect 320270 497791 320326 497800
rect 320178 497312 320234 497321
rect 320178 497247 320234 497256
rect 320180 496868 320232 496874
rect 320180 496810 320232 496816
rect 319812 495576 319864 495582
rect 319812 495518 319864 495524
rect 319824 495281 319852 495518
rect 319996 495508 320048 495514
rect 319996 495450 320048 495456
rect 319810 495272 319866 495281
rect 319810 495207 319866 495216
rect 319812 494080 319864 494086
rect 319812 494022 319864 494028
rect 319824 493785 319852 494022
rect 319810 493776 319866 493785
rect 319810 493711 319866 493720
rect 320008 492697 320036 495450
rect 320192 495009 320220 496810
rect 320178 495000 320234 495009
rect 320178 494935 320234 494944
rect 320180 492720 320232 492726
rect 319994 492688 320050 492697
rect 320180 492662 320232 492668
rect 319994 492623 320050 492632
rect 319812 491360 319864 491366
rect 319812 491302 319864 491308
rect 319824 491201 319852 491302
rect 319810 491192 319866 491201
rect 319810 491127 319866 491136
rect 320192 490385 320220 492662
rect 320178 490376 320234 490385
rect 320178 490311 320234 490320
rect 320180 489932 320232 489938
rect 320180 489874 320232 489880
rect 320088 489864 320140 489870
rect 320086 489832 320088 489841
rect 320140 489832 320142 489841
rect 320086 489767 320142 489776
rect 319812 488640 319864 488646
rect 319812 488582 319864 488588
rect 319720 488572 319772 488578
rect 319720 488514 319772 488520
rect 319732 486713 319760 488514
rect 319824 487937 319852 488582
rect 320192 487937 320220 489874
rect 320284 488481 320312 497791
rect 320376 493513 320404 502415
rect 320454 496632 320510 496641
rect 320454 496567 320510 496576
rect 320362 493504 320418 493513
rect 320362 493439 320418 493448
rect 320270 488472 320326 488481
rect 320270 488407 320326 488416
rect 319810 487928 319866 487937
rect 319810 487863 319866 487872
rect 320178 487928 320234 487937
rect 320178 487863 320234 487872
rect 320270 487384 320326 487393
rect 320270 487319 320326 487328
rect 320180 487212 320232 487218
rect 320180 487154 320232 487160
rect 319718 486704 319774 486713
rect 319718 486639 319774 486648
rect 319812 485852 319864 485858
rect 319812 485794 319864 485800
rect 319824 485625 319852 485794
rect 319810 485616 319866 485625
rect 319810 485551 319866 485560
rect 320192 484537 320220 487154
rect 320178 484528 320234 484537
rect 320178 484463 320234 484472
rect 320180 484424 320232 484430
rect 320180 484366 320232 484372
rect 319812 483064 319864 483070
rect 319810 483032 319812 483041
rect 319864 483032 319866 483041
rect 319810 482967 319866 482976
rect 320192 482089 320220 484366
rect 320178 482080 320234 482089
rect 320178 482015 320234 482024
rect 320180 481704 320232 481710
rect 320180 481646 320232 481652
rect 319812 480276 319864 480282
rect 319812 480218 319864 480224
rect 319824 479777 319852 480218
rect 320192 479777 320220 481646
rect 320284 480486 320312 487319
rect 320376 484129 320404 493439
rect 320468 487393 320496 496567
rect 320560 494601 320588 503639
rect 320638 500168 320694 500177
rect 320638 500103 320694 500112
rect 320652 495514 320680 500103
rect 320744 499066 320772 504727
rect 320822 501392 320878 501401
rect 320878 501350 320956 501378
rect 320822 501327 320878 501336
rect 320744 499038 320864 499066
rect 320730 498944 320786 498953
rect 320730 498879 320786 498888
rect 320640 495508 320692 495514
rect 320640 495450 320692 495456
rect 320546 494592 320602 494601
rect 320546 494527 320602 494536
rect 320454 487384 320510 487393
rect 320454 487319 320510 487328
rect 320456 487280 320508 487286
rect 320456 487222 320508 487228
rect 320468 486169 320496 487222
rect 320560 486266 320588 494527
rect 320744 492386 320772 498879
rect 320836 495553 320864 499038
rect 320822 495544 320878 495553
rect 320822 495479 320878 495488
rect 320836 492386 320864 495479
rect 320732 492380 320784 492386
rect 320732 492322 320784 492328
rect 320824 492380 320876 492386
rect 320824 492322 320876 492328
rect 320638 492280 320694 492289
rect 320928 492266 320956 501350
rect 320694 492238 320956 492266
rect 320638 492215 320694 492224
rect 320732 492176 320784 492182
rect 320732 492118 320784 492124
rect 320824 492176 320876 492182
rect 320824 492118 320876 492124
rect 320640 490952 320692 490958
rect 320638 490920 320640 490929
rect 320692 490920 320694 490929
rect 320638 490855 320694 490864
rect 320640 489932 320692 489938
rect 320640 489874 320692 489880
rect 320652 486266 320680 489874
rect 320744 489870 320772 492118
rect 320836 489870 320864 492118
rect 320732 489864 320784 489870
rect 320732 489806 320784 489812
rect 320824 489864 320876 489870
rect 320824 489806 320876 489812
rect 320824 489456 320876 489462
rect 320824 489398 320876 489404
rect 320730 488472 320786 488481
rect 320730 488407 320786 488416
rect 320548 486260 320600 486266
rect 320548 486202 320600 486208
rect 320640 486260 320692 486266
rect 320640 486202 320692 486208
rect 320454 486160 320510 486169
rect 320454 486095 320510 486104
rect 320362 484120 320418 484129
rect 320362 484055 320418 484064
rect 320272 480480 320324 480486
rect 320272 480422 320324 480428
rect 320272 480344 320324 480350
rect 320272 480286 320324 480292
rect 319810 479768 319866 479777
rect 319810 479703 319866 479712
rect 320178 479768 320234 479777
rect 320178 479703 320234 479712
rect 320180 479324 320232 479330
rect 320180 479266 320232 479272
rect 320192 476882 320220 479266
rect 320180 476876 320232 476882
rect 320180 476818 320232 476824
rect 320178 476776 320234 476785
rect 320284 476762 320312 480286
rect 320376 476898 320404 484055
rect 320468 482866 320496 486095
rect 320548 486056 320600 486062
rect 320548 485998 320600 486004
rect 320640 486056 320692 486062
rect 320640 485998 320692 486004
rect 320560 484945 320588 485998
rect 320546 484936 320602 484945
rect 320546 484871 320602 484880
rect 320456 482860 320508 482866
rect 320456 482802 320508 482808
rect 320456 482724 320508 482730
rect 320456 482666 320508 482672
rect 320468 481545 320496 482666
rect 320560 482474 320588 484871
rect 320652 482730 320680 485998
rect 320744 482769 320772 488407
rect 320730 482760 320786 482769
rect 320640 482724 320692 482730
rect 320836 482730 320864 489398
rect 320730 482695 320786 482704
rect 320824 482724 320876 482730
rect 320640 482666 320692 482672
rect 320824 482666 320876 482672
rect 320638 482624 320694 482633
rect 320928 482610 320956 492238
rect 320694 482582 320956 482610
rect 320638 482559 320694 482568
rect 320560 482446 320772 482474
rect 320548 482384 320600 482390
rect 320548 482326 320600 482332
rect 320638 482352 320694 482361
rect 320454 481536 320510 481545
rect 320454 481471 320510 481480
rect 320468 477018 320496 481471
rect 320560 480321 320588 482326
rect 320638 482287 320694 482296
rect 320546 480312 320602 480321
rect 320546 480247 320602 480256
rect 320456 477012 320508 477018
rect 320456 476954 320508 476960
rect 320376 476870 320496 476898
rect 320362 476776 320418 476785
rect 320284 476734 320362 476762
rect 320178 476711 320234 476720
rect 320362 476711 320418 476720
rect 320192 474774 320220 476711
rect 320272 476672 320324 476678
rect 320272 476614 320324 476620
rect 320180 474768 320232 474774
rect 320180 474710 320232 474716
rect 320178 474464 320234 474473
rect 320178 474399 320234 474408
rect 320192 472054 320220 474399
rect 320284 473385 320312 476614
rect 320376 474026 320404 476711
rect 320468 475969 320496 476870
rect 320454 475960 320510 475969
rect 320454 475895 320510 475904
rect 320456 475856 320508 475862
rect 320456 475798 320508 475804
rect 320364 474020 320416 474026
rect 320364 473962 320416 473968
rect 320468 473906 320496 475798
rect 320376 473878 320496 473906
rect 320270 473376 320326 473385
rect 320270 473311 320326 473320
rect 320270 473240 320326 473249
rect 320270 473175 320326 473184
rect 320180 472048 320232 472054
rect 320180 471990 320232 471996
rect 320178 471064 320234 471073
rect 320178 470999 320234 471008
rect 320192 468738 320220 470999
rect 320284 470626 320312 473175
rect 320376 472297 320404 473878
rect 320560 473362 320588 480247
rect 320652 479097 320680 482287
rect 320744 479210 320772 482446
rect 320824 480480 320876 480486
rect 320824 480422 320876 480428
rect 320836 479466 320864 480422
rect 320824 479460 320876 479466
rect 320824 479402 320876 479408
rect 320928 479346 320956 482582
rect 320836 479330 320956 479346
rect 320824 479324 320956 479330
rect 320876 479318 320956 479324
rect 320824 479266 320876 479272
rect 320744 479182 320864 479210
rect 320638 479088 320694 479097
rect 320694 479046 320772 479074
rect 320638 479023 320694 479032
rect 320640 478984 320692 478990
rect 320640 478926 320692 478932
rect 320652 478009 320680 478926
rect 320638 478000 320694 478009
rect 320638 477935 320694 477944
rect 320640 477012 320692 477018
rect 320640 476954 320692 476960
rect 320652 475930 320680 476954
rect 320744 476066 320772 479046
rect 320732 476060 320784 476066
rect 320732 476002 320784 476008
rect 320730 475960 320786 475969
rect 320640 475924 320692 475930
rect 320730 475895 320786 475904
rect 320640 475866 320692 475872
rect 320638 475824 320694 475833
rect 320638 475759 320694 475768
rect 320468 473334 320588 473362
rect 320362 472288 320418 472297
rect 320362 472223 320418 472232
rect 320362 472152 320418 472161
rect 320362 472087 320418 472096
rect 320272 470620 320324 470626
rect 320272 470562 320324 470568
rect 320272 470484 320324 470490
rect 320272 470426 320324 470432
rect 320284 470121 320312 470426
rect 320270 470112 320326 470121
rect 320270 470047 320326 470056
rect 320270 469840 320326 469849
rect 320270 469775 320326 469784
rect 320100 468710 320220 468738
rect 320100 467702 320128 468710
rect 320178 468616 320234 468625
rect 320178 468551 320234 468560
rect 320088 467696 320140 467702
rect 320088 467638 320140 467644
rect 320192 466478 320220 468551
rect 320284 467906 320312 469775
rect 320376 469266 320404 472087
rect 320468 471073 320496 473334
rect 320546 473240 320602 473249
rect 320546 473175 320602 473184
rect 320454 471064 320510 471073
rect 320454 470999 320510 471008
rect 320454 470928 320510 470937
rect 320454 470863 320510 470872
rect 320364 469260 320416 469266
rect 320364 469202 320416 469208
rect 320362 469160 320418 469169
rect 320362 469095 320418 469104
rect 320272 467900 320324 467906
rect 320272 467842 320324 467848
rect 320376 467786 320404 469095
rect 320468 467974 320496 470863
rect 320456 467968 320508 467974
rect 320456 467910 320508 467916
rect 320560 467838 320588 473175
rect 320652 468897 320680 475759
rect 320744 474473 320772 475895
rect 320836 475833 320864 479182
rect 320822 475824 320878 475833
rect 320822 475759 320824 475768
rect 320876 475759 320878 475768
rect 320824 475730 320876 475736
rect 320836 475699 320864 475730
rect 320822 475552 320878 475561
rect 320822 475487 320878 475496
rect 320730 474464 320786 474473
rect 320730 474399 320786 474408
rect 320638 468888 320694 468897
rect 320638 468823 320694 468832
rect 320548 467832 320600 467838
rect 320272 467764 320324 467770
rect 320376 467758 320496 467786
rect 320548 467774 320600 467780
rect 320272 467706 320324 467712
rect 320180 466472 320232 466478
rect 320180 466414 320232 466420
rect 320178 465216 320234 465225
rect 320178 465151 320234 465160
rect 320192 465118 320220 465151
rect 320180 465112 320232 465118
rect 320180 465054 320232 465060
rect 320178 464944 320234 464953
rect 320178 464879 320234 464888
rect 320192 457162 320220 464879
rect 320180 457156 320232 457162
rect 320180 457098 320232 457104
rect 320284 457042 320312 467706
rect 320364 467628 320416 467634
rect 320364 467570 320416 467576
rect 320192 457014 320312 457042
rect 320192 452334 320220 457014
rect 320376 456958 320404 467570
rect 320468 457502 320496 467758
rect 320548 467696 320600 467702
rect 320652 467673 320680 468823
rect 320744 467770 320772 474399
rect 320732 467764 320784 467770
rect 320732 467706 320784 467712
rect 320548 467638 320600 467644
rect 320638 467664 320694 467673
rect 320456 457496 320508 457502
rect 320456 457438 320508 457444
rect 320364 456952 320416 456958
rect 320364 456894 320416 456900
rect 320364 456680 320416 456686
rect 320364 456622 320416 456628
rect 320456 456680 320508 456686
rect 320456 456622 320508 456628
rect 320180 452328 320232 452334
rect 320180 452270 320232 452276
rect 320376 447370 320404 456622
rect 320468 447370 320496 456622
rect 320560 447370 320588 467638
rect 320638 467599 320694 467608
rect 320640 467560 320692 467566
rect 320640 467502 320692 467508
rect 320652 457502 320680 467502
rect 320732 467424 320784 467430
rect 320732 467366 320784 467372
rect 320640 457496 320692 457502
rect 320640 457438 320692 457444
rect 320744 456958 320772 467366
rect 320836 457366 320864 475487
rect 320824 457360 320876 457366
rect 320824 457302 320876 457308
rect 320732 456952 320784 456958
rect 320732 456894 320784 456900
rect 320640 456544 320692 456550
rect 320640 456486 320692 456492
rect 320652 449886 320680 456486
rect 320640 449880 320692 449886
rect 320640 449822 320692 449828
rect 320364 447364 320416 447370
rect 320364 447306 320416 447312
rect 320456 447364 320508 447370
rect 320456 447306 320508 447312
rect 320548 447364 320600 447370
rect 320548 447306 320600 447312
rect 320456 447228 320508 447234
rect 320456 447170 320508 447176
rect 320548 447228 320600 447234
rect 320548 447170 320600 447176
rect 320364 447024 320416 447030
rect 320364 446966 320416 446972
rect 320272 431996 320324 432002
rect 320272 431938 320324 431944
rect 320284 427786 320312 431938
rect 320272 427780 320324 427786
rect 320272 427722 320324 427728
rect 320180 398880 320232 398886
rect 320180 398822 320232 398828
rect 320192 392170 320220 398822
rect 320100 392142 320220 392170
rect 320100 391898 320128 392142
rect 320180 392080 320232 392086
rect 320178 392048 320180 392057
rect 320232 392048 320234 392057
rect 320178 391983 320234 391992
rect 320272 392012 320324 392018
rect 320272 391954 320324 391960
rect 320100 391870 320220 391898
rect 320088 390584 320140 390590
rect 320088 390526 320140 390532
rect 320100 389065 320128 390526
rect 320192 390522 320220 391870
rect 320180 390516 320232 390522
rect 320180 390458 320232 390464
rect 320284 389881 320312 391954
rect 320376 391950 320404 446966
rect 320468 442377 320496 447170
rect 320560 442474 320588 447170
rect 320640 447160 320692 447166
rect 320640 447102 320692 447108
rect 320548 442468 320600 442474
rect 320548 442410 320600 442416
rect 320454 442368 320510 442377
rect 320454 442303 320510 442312
rect 320548 442196 320600 442202
rect 320548 442138 320600 442144
rect 320456 442060 320508 442066
rect 320456 442002 320508 442008
rect 320468 394670 320496 442002
rect 320560 396030 320588 442138
rect 320652 397458 320680 447102
rect 320836 446962 320956 446978
rect 320824 446956 320956 446962
rect 320876 446950 320956 446956
rect 320824 446898 320876 446904
rect 320732 446888 320784 446894
rect 320732 446830 320784 446836
rect 320744 442474 320772 446830
rect 320824 446820 320876 446826
rect 320824 446762 320876 446768
rect 320732 442468 320784 442474
rect 320732 442410 320784 442416
rect 320730 442368 320786 442377
rect 320730 442303 320786 442312
rect 320744 400178 320772 442303
rect 320836 432002 320864 446762
rect 320824 431996 320876 432002
rect 320824 431938 320876 431944
rect 320824 427780 320876 427786
rect 320824 427722 320876 427728
rect 320732 400172 320784 400178
rect 320732 400114 320784 400120
rect 320836 398886 320864 427722
rect 320824 398880 320876 398886
rect 320824 398822 320876 398828
rect 320640 397452 320692 397458
rect 320640 397394 320692 397400
rect 320548 396024 320600 396030
rect 320548 395966 320600 395972
rect 320456 394664 320508 394670
rect 320456 394606 320508 394612
rect 320364 391944 320416 391950
rect 320364 391886 320416 391892
rect 320270 389872 320326 389881
rect 320270 389807 320326 389816
rect 320272 389224 320324 389230
rect 320272 389166 320324 389172
rect 320086 389056 320142 389065
rect 320086 388991 320142 389000
rect 320180 387864 320232 387870
rect 320180 387806 320232 387812
rect 320192 386345 320220 387806
rect 320284 387569 320312 389166
rect 320928 387818 320956 446950
rect 338672 396840 338724 396846
rect 338670 396808 338672 396817
rect 338724 396808 338726 396817
rect 338670 396743 338726 396752
rect 397458 396808 397514 396817
rect 397458 396743 397460 396752
rect 397512 396743 397514 396752
rect 397460 396714 397512 396720
rect 398840 396704 398892 396710
rect 398838 396672 398840 396681
rect 398892 396672 398894 396681
rect 398838 396607 398894 396616
rect 400218 396672 400274 396681
rect 400218 396607 400220 396616
rect 400272 396607 400274 396616
rect 400220 396578 400272 396584
rect 401600 396568 401652 396574
rect 401598 396536 401600 396545
rect 401652 396536 401654 396545
rect 401598 396471 401654 396480
rect 403346 396536 403402 396545
rect 403346 396471 403348 396480
rect 403400 396471 403402 396480
rect 404358 396536 404414 396545
rect 404358 396471 404414 396480
rect 406014 396536 406070 396545
rect 406014 396471 406070 396480
rect 403348 396442 403400 396448
rect 404372 396438 404400 396471
rect 406028 396438 406056 396471
rect 404360 396432 404412 396438
rect 404360 396374 404412 396380
rect 406016 396432 406068 396438
rect 406016 396374 406068 396380
rect 320836 387802 320956 387818
rect 320824 387796 320956 387802
rect 320876 387790 320956 387796
rect 320824 387738 320876 387744
rect 320364 387728 320416 387734
rect 320364 387670 320416 387676
rect 320270 387560 320326 387569
rect 320270 387495 320326 387504
rect 320376 386481 320404 387670
rect 320362 386472 320418 386481
rect 320362 386407 320418 386416
rect 320272 386368 320324 386374
rect 320178 386336 320234 386345
rect 320272 386310 320324 386316
rect 320178 386271 320234 386280
rect 320180 385008 320232 385014
rect 320180 384950 320232 384956
rect 320192 383761 320220 384950
rect 320178 383752 320234 383761
rect 320178 383687 320234 383696
rect 320180 383648 320232 383654
rect 320180 383590 320232 383596
rect 320192 383058 320220 383590
rect 320284 383217 320312 386310
rect 320364 384940 320416 384946
rect 320364 384882 320416 384888
rect 320270 383208 320326 383217
rect 320270 383143 320326 383152
rect 320192 383030 320312 383058
rect 320180 380860 320232 380866
rect 320180 380802 320232 380808
rect 320088 380248 320140 380254
rect 320088 380190 320140 380196
rect 320100 379386 320128 380190
rect 320192 379545 320220 380802
rect 320284 379681 320312 383030
rect 320376 380905 320404 384882
rect 320638 384840 320694 384849
rect 320638 384775 320694 384784
rect 320548 382220 320600 382226
rect 320548 382162 320600 382168
rect 320362 380896 320418 380905
rect 320362 380831 320418 380840
rect 320456 380180 320508 380186
rect 320456 380122 320508 380128
rect 320270 379672 320326 379681
rect 320270 379607 320326 379616
rect 320178 379536 320234 379545
rect 320178 379471 320234 379480
rect 320272 379500 320324 379506
rect 320272 379442 320324 379448
rect 320100 379358 320220 379386
rect 320192 377777 320220 379358
rect 320178 377768 320234 377777
rect 320178 377703 320234 377712
rect 319996 376848 320048 376854
rect 319996 376790 320048 376796
rect 320178 376816 320234 376825
rect 319812 376780 319864 376786
rect 319812 376722 319864 376728
rect 319824 375193 319852 376722
rect 319810 375184 319866 375193
rect 319810 375119 319866 375128
rect 320008 373833 320036 376790
rect 320178 376751 320234 376760
rect 320192 375465 320220 376751
rect 320284 376145 320312 379442
rect 320468 379001 320496 380122
rect 320454 378992 320510 379001
rect 320454 378927 320510 378936
rect 320364 378888 320416 378894
rect 320364 378830 320416 378836
rect 320376 376689 320404 378830
rect 320362 376680 320418 376689
rect 320362 376615 320418 376624
rect 320364 376576 320416 376582
rect 320364 376518 320416 376524
rect 320270 376136 320326 376145
rect 320270 376071 320326 376080
rect 320178 375456 320234 375465
rect 320178 375391 320234 375400
rect 320192 374082 320220 375391
rect 320272 375352 320324 375358
rect 320272 375294 320324 375300
rect 320100 374054 320220 374082
rect 319994 373824 320050 373833
rect 319994 373759 320050 373768
rect 320100 373538 320128 374054
rect 320180 373992 320232 373998
rect 320180 373934 320232 373940
rect 320008 373510 320128 373538
rect 319904 371884 319956 371890
rect 319904 371826 319956 371832
rect 319812 369776 319864 369782
rect 319812 369718 319864 369724
rect 319824 365673 319852 369718
rect 319916 369102 319944 371826
rect 320008 370530 320036 373510
rect 320086 373144 320142 373153
rect 320086 373079 320142 373088
rect 320100 372978 320128 373079
rect 320088 372972 320140 372978
rect 320088 372914 320140 372920
rect 320192 372745 320220 373934
rect 320178 372736 320234 372745
rect 320178 372671 320234 372680
rect 320284 371521 320312 375294
rect 320376 372609 320404 376518
rect 320362 372600 320418 372609
rect 320362 372535 320418 372544
rect 320364 372496 320416 372502
rect 320364 372438 320416 372444
rect 320270 371512 320326 371521
rect 320270 371447 320326 371456
rect 320272 371204 320324 371210
rect 320272 371146 320324 371152
rect 319996 370524 320048 370530
rect 319996 370466 320048 370472
rect 320008 369510 320036 370466
rect 320180 369844 320232 369850
rect 320180 369786 320232 369792
rect 319996 369504 320048 369510
rect 319996 369446 320048 369452
rect 319904 369096 319956 369102
rect 319904 369038 319956 369044
rect 320192 368529 320220 369786
rect 320178 368520 320234 368529
rect 320178 368455 320234 368464
rect 320284 367985 320312 371146
rect 320376 369209 320404 372438
rect 320468 369753 320496 378927
rect 320560 378457 320588 382162
rect 320652 381410 320680 384775
rect 320730 383616 320786 383625
rect 320730 383551 320786 383560
rect 320640 381404 320692 381410
rect 320640 381346 320692 381352
rect 320638 381304 320694 381313
rect 320638 381239 320694 381248
rect 320652 379778 320680 381239
rect 320640 379772 320692 379778
rect 320640 379714 320692 379720
rect 320744 379658 320772 383551
rect 320822 382528 320878 382537
rect 320822 382463 320878 382472
rect 320836 380322 320864 382463
rect 320824 380316 320876 380322
rect 320824 380258 320876 380264
rect 320822 380216 320878 380225
rect 320822 380151 320878 380160
rect 320652 379630 320772 379658
rect 320546 378448 320602 378457
rect 320546 378383 320602 378392
rect 320548 378344 320600 378350
rect 320548 378286 320600 378292
rect 320560 376038 320588 378286
rect 320548 376032 320600 376038
rect 320548 375974 320600 375980
rect 320560 374474 320588 375974
rect 320548 374468 320600 374474
rect 320548 374410 320600 374416
rect 320546 374368 320602 374377
rect 320652 374354 320680 379630
rect 320732 379568 320784 379574
rect 320732 379510 320784 379516
rect 320744 376825 320772 379510
rect 320836 378826 320864 380151
rect 320824 378820 320876 378826
rect 320824 378762 320876 378768
rect 320836 377890 320864 378762
rect 320836 377862 320956 377890
rect 320822 377768 320878 377777
rect 320822 377703 320878 377712
rect 320730 376816 320786 376825
rect 320730 376751 320786 376760
rect 320602 374326 320680 374354
rect 320546 374303 320602 374312
rect 320560 371890 320588 374303
rect 320640 374264 320692 374270
rect 320640 374206 320692 374212
rect 320652 372337 320680 374206
rect 320638 372328 320694 372337
rect 320638 372263 320694 372272
rect 320548 371884 320600 371890
rect 320548 371826 320600 371832
rect 320652 370530 320680 372263
rect 320836 371618 320864 377703
rect 320824 371612 320876 371618
rect 320824 371554 320876 371560
rect 320822 371240 320878 371249
rect 320928 371226 320956 377862
rect 320878 371198 320956 371226
rect 320822 371175 320878 371184
rect 320836 371074 320864 371175
rect 320824 371068 320876 371074
rect 320824 371010 320876 371016
rect 320640 370524 320692 370530
rect 320640 370466 320692 370472
rect 320824 370524 320876 370530
rect 320876 370484 320956 370512
rect 320824 370466 320876 370472
rect 320640 370320 320692 370326
rect 320640 370262 320692 370268
rect 320454 369744 320510 369753
rect 320454 369679 320510 369688
rect 320652 369594 320680 370262
rect 320468 369566 320680 369594
rect 320362 369200 320418 369209
rect 320362 369135 320418 369144
rect 320364 369096 320416 369102
rect 320364 369038 320416 369044
rect 320270 367976 320326 367985
rect 320270 367911 320326 367920
rect 320272 367872 320324 367878
rect 320272 367814 320324 367820
rect 320180 365764 320232 365770
rect 320180 365706 320232 365712
rect 319810 365664 319866 365673
rect 319810 365599 319866 365608
rect 320192 364993 320220 365706
rect 320178 364984 320234 364993
rect 320178 364919 320234 364928
rect 320284 364426 320312 367814
rect 320376 365838 320404 369038
rect 320468 368626 320496 369566
rect 320640 369504 320692 369510
rect 320640 369446 320692 369452
rect 320730 369472 320786 369481
rect 320456 368620 320508 368626
rect 320456 368562 320508 368568
rect 320456 368484 320508 368490
rect 320456 368426 320508 368432
rect 320364 365832 320416 365838
rect 320364 365774 320416 365780
rect 320364 365696 320416 365702
rect 320364 365638 320416 365644
rect 320192 364398 320312 364426
rect 320008 363798 320036 363829
rect 319996 363792 320048 363798
rect 319994 363760 319996 363769
rect 320048 363760 320050 363769
rect 319994 363695 320050 363704
rect 319812 362840 319864 362846
rect 319812 362782 319864 362788
rect 319824 361457 319852 362782
rect 319810 361448 319866 361457
rect 319810 361383 319866 361392
rect 320008 359854 320036 363695
rect 320088 362704 320140 362710
rect 320086 362672 320088 362681
rect 320140 362672 320142 362681
rect 320086 362607 320142 362616
rect 320192 361457 320220 364398
rect 320272 364336 320324 364342
rect 320272 364278 320324 364284
rect 320178 361448 320234 361457
rect 320178 361383 320234 361392
rect 320192 360346 320220 361383
rect 320284 361049 320312 364278
rect 320376 362137 320404 365638
rect 320468 364449 320496 368426
rect 320652 366217 320680 369446
rect 320730 369407 320786 369416
rect 320638 366208 320694 366217
rect 320638 366143 320694 366152
rect 320652 365378 320680 366143
rect 320560 365350 320680 365378
rect 320454 364440 320510 364449
rect 320454 364375 320510 364384
rect 320456 362908 320508 362914
rect 320456 362850 320508 362856
rect 320362 362128 320418 362137
rect 320362 362063 320418 362072
rect 320468 361978 320496 362850
rect 320376 361950 320496 361978
rect 320270 361040 320326 361049
rect 320270 360975 320326 360984
rect 320272 360936 320324 360942
rect 320272 360878 320324 360884
rect 320284 360369 320312 360878
rect 320100 360318 320220 360346
rect 320270 360360 320326 360369
rect 320100 360074 320128 360318
rect 320270 360295 320326 360304
rect 320284 360194 320312 360295
rect 320272 360188 320324 360194
rect 320272 360130 320324 360136
rect 320100 360046 320220 360074
rect 319996 359848 320048 359854
rect 319996 359790 320048 359796
rect 320192 356930 320220 360046
rect 320272 360052 320324 360058
rect 320272 359994 320324 360000
rect 320284 357921 320312 359994
rect 320376 358601 320404 361950
rect 320456 360256 320508 360262
rect 320456 360198 320508 360204
rect 320468 359825 320496 360198
rect 320454 359816 320510 359825
rect 320454 359751 320510 359760
rect 320362 358592 320418 358601
rect 320362 358527 320418 358536
rect 320270 357912 320326 357921
rect 320270 357847 320326 357856
rect 320180 356924 320232 356930
rect 320180 356866 320232 356872
rect 320178 356824 320234 356833
rect 320178 356759 320234 356768
rect 320192 356046 320220 356759
rect 320180 356040 320232 356046
rect 320180 355982 320232 355988
rect 320178 355600 320234 355609
rect 320178 355535 320234 355544
rect 320192 354686 320220 355535
rect 320180 354680 320232 354686
rect 320180 354622 320232 354628
rect 320178 354512 320234 354521
rect 320178 354447 320234 354456
rect 320192 353258 320220 354447
rect 320284 353433 320312 357847
rect 320560 357105 320588 365350
rect 320638 364984 320694 364993
rect 320638 364919 320694 364928
rect 320546 357096 320602 357105
rect 320546 357031 320602 357040
rect 320364 356924 320416 356930
rect 320364 356866 320416 356872
rect 320270 353424 320326 353433
rect 320270 353359 320326 353368
rect 320270 353288 320326 353297
rect 320180 353252 320232 353258
rect 320270 353223 320326 353232
rect 320180 353194 320232 353200
rect 320178 352608 320234 352617
rect 320178 352543 320234 352552
rect 320192 351234 320220 352543
rect 320284 351898 320312 353223
rect 320376 352481 320404 356866
rect 320652 356017 320680 364919
rect 320744 360942 320772 369407
rect 320822 368520 320878 368529
rect 320928 368506 320956 370484
rect 320878 368478 320956 368506
rect 320822 368455 320878 368464
rect 320822 367296 320878 367305
rect 320822 367231 320878 367240
rect 320732 360936 320784 360942
rect 320732 360878 320784 360884
rect 320836 360754 320864 367231
rect 320744 360726 320864 360754
rect 320744 360058 320772 360726
rect 320928 360618 320956 368478
rect 320836 360590 320956 360618
rect 320836 360330 320864 360590
rect 320824 360324 320876 360330
rect 320824 360266 320876 360272
rect 320732 360052 320784 360058
rect 320732 359994 320784 360000
rect 320744 359922 320956 359938
rect 320732 359916 320956 359922
rect 320784 359910 320956 359916
rect 320732 359858 320784 359864
rect 320824 359848 320876 359854
rect 320730 359816 320786 359825
rect 320824 359790 320876 359796
rect 320730 359751 320786 359760
rect 320638 356008 320694 356017
rect 320638 355943 320694 355952
rect 320640 355904 320692 355910
rect 320640 355846 320692 355852
rect 320362 352472 320418 352481
rect 320362 352407 320418 352416
rect 320272 351892 320324 351898
rect 320272 351834 320324 351840
rect 320652 351257 320680 355846
rect 320638 351248 320694 351257
rect 320192 351206 320312 351234
rect 320284 350470 320312 351206
rect 320638 351183 320694 351192
rect 320362 350976 320418 350985
rect 320362 350911 320418 350920
rect 320272 350464 320324 350470
rect 320272 350406 320324 350412
rect 320178 349752 320234 349761
rect 320178 349687 320234 349696
rect 320192 349110 320220 349687
rect 320180 349104 320232 349110
rect 320180 349046 320232 349052
rect 320376 349042 320404 350911
rect 320744 350169 320772 359751
rect 320836 354657 320864 359790
rect 320822 354648 320878 354657
rect 320822 354583 320878 354592
rect 320822 353288 320878 353297
rect 320928 353274 320956 359910
rect 320878 353246 320956 353274
rect 320822 353223 320878 353232
rect 320730 350160 320786 350169
rect 320730 350095 320786 350104
rect 320364 349036 320416 349042
rect 320364 348978 320416 348984
rect 320178 348664 320234 348673
rect 320178 348599 320234 348608
rect 320192 347750 320220 348599
rect 320180 347744 320232 347750
rect 320180 347686 320232 347692
rect 320180 346384 320232 346390
rect 320178 346352 320180 346361
rect 320232 346352 320234 346361
rect 320178 346287 320234 346296
rect 319444 331220 319496 331226
rect 319444 331162 319496 331168
rect 316684 329792 316736 329798
rect 316684 329734 316736 329740
rect 275652 323332 275704 323338
rect 275652 323274 275704 323280
rect 273444 321292 273496 321298
rect 273444 321234 273496 321240
rect 275560 321292 275612 321298
rect 275560 321234 275612 321240
rect 273456 321065 273484 321234
rect 273442 321056 273498 321065
rect 273442 320991 273498 321000
rect 70306 320648 70362 320657
rect 70242 320620 70306 320634
rect 70228 320606 70306 320620
rect 49608 318776 49660 318782
rect 70228 318753 70256 320606
rect 70306 320583 70362 320592
rect 267384 320334 267674 320362
rect 70412 320198 70610 320226
rect 70780 320198 70978 320226
rect 77404 320198 77602 320226
rect 81912 320198 82110 320226
rect 90468 320198 90850 320226
rect 104452 320198 104834 320226
rect 105004 320198 105202 320226
rect 163976 320198 164174 320226
rect 231504 320210 231794 320226
rect 230664 320204 230716 320210
rect 70412 319410 70440 320198
rect 70780 319410 70808 320198
rect 71056 320062 71438 320090
rect 70412 319382 70532 319410
rect 70780 319382 70900 319410
rect 49608 318718 49660 318724
rect 69018 318744 69074 318753
rect 46848 318708 46900 318714
rect 46848 318650 46900 318656
rect 39948 318640 40000 318646
rect 23386 318608 23442 318617
rect 39948 318582 40000 318588
rect 23386 318543 23442 318552
rect 17866 318472 17922 318481
rect 17866 318407 17922 318416
rect 16486 318336 16542 318345
rect 16486 318271 16542 318280
rect 15106 318200 15162 318209
rect 15106 318135 15162 318144
rect 13726 318064 13782 318073
rect 13726 317999 13782 318008
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2884 480 2912 4898
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 480 4108 3402
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 6472 480 6500 3470
rect 7668 480 7696 4966
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8864 480 8892 3538
rect 10046 3496 10102 3505
rect 10046 3431 10102 3440
rect 10060 480 10088 3431
rect 11256 480 11284 3606
rect 12452 480 12480 3674
rect 13740 3482 13768 317999
rect 15120 3482 15148 318135
rect 13648 3454 13768 3482
rect 14844 3454 15148 3482
rect 13648 480 13676 3454
rect 14844 480 14872 3454
rect 16500 3398 16528 318271
rect 17880 3398 17908 318407
rect 20720 3868 20772 3874
rect 20720 3810 20772 3816
rect 19522 3768 19578 3777
rect 19522 3703 19578 3712
rect 18326 3632 18382 3641
rect 18326 3567 18382 3576
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 16040 480 16068 3334
rect 17236 480 17264 3334
rect 18340 480 18368 3567
rect 19536 480 19564 3703
rect 20732 480 20760 3810
rect 21916 3800 21968 3806
rect 21916 3742 21968 3748
rect 21928 480 21956 3742
rect 23400 3482 23428 318543
rect 38568 318504 38620 318510
rect 38568 318446 38620 318452
rect 34428 318436 34480 318442
rect 34428 318378 34480 318384
rect 33048 318368 33100 318374
rect 33048 318310 33100 318316
rect 27528 318300 27580 318306
rect 27528 318242 27580 318248
rect 26148 318164 26200 318170
rect 26148 318106 26200 318112
rect 24768 318096 24820 318102
rect 24768 318038 24820 318044
rect 23124 3454 23428 3482
rect 23124 480 23152 3454
rect 24780 3398 24808 318038
rect 26160 3398 26188 318106
rect 27540 3398 27568 318242
rect 31668 318232 31720 318238
rect 31668 318174 31720 318180
rect 30288 4004 30340 4010
rect 30288 3946 30340 3952
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 29090 3904 29146 3913
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 25504 3392 25556 3398
rect 25504 3334 25556 3340
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 26700 3392 26752 3398
rect 26700 3334 26752 3340
rect 27528 3392 27580 3398
rect 27528 3334 27580 3340
rect 24320 480 24348 3334
rect 25516 480 25544 3334
rect 26712 480 26740 3334
rect 27908 480 27936 3878
rect 29090 3839 29146 3848
rect 29104 480 29132 3839
rect 30300 480 30328 3946
rect 31680 3482 31708 318174
rect 33060 3482 33088 318310
rect 31496 3454 31708 3482
rect 32692 3454 33088 3482
rect 31496 480 31524 3454
rect 32692 480 32720 3454
rect 34440 3398 34468 318378
rect 36176 4140 36228 4146
rect 36176 4082 36228 4088
rect 34980 4072 35032 4078
rect 34980 4014 35032 4020
rect 33876 3392 33928 3398
rect 33876 3334 33928 3340
rect 34428 3392 34480 3398
rect 34428 3334 34480 3340
rect 33888 480 33916 3334
rect 34992 480 35020 4014
rect 36188 480 36216 4082
rect 37372 3052 37424 3058
rect 37372 2994 37424 3000
rect 37384 480 37412 2994
rect 38580 480 38608 318446
rect 39960 3482 39988 318582
rect 41328 318572 41380 318578
rect 41328 318514 41380 318520
rect 41340 3482 41368 318514
rect 42154 4040 42210 4049
rect 42154 3975 42210 3984
rect 39776 3454 39988 3482
rect 40972 3454 41368 3482
rect 39776 480 39804 3454
rect 40972 480 41000 3454
rect 42168 480 42196 3975
rect 46860 3262 46888 318650
rect 48136 318028 48188 318034
rect 48136 317970 48188 317976
rect 48148 3262 48176 317970
rect 48228 5092 48280 5098
rect 48228 5034 48280 5040
rect 45744 3256 45796 3262
rect 45744 3198 45796 3204
rect 46848 3256 46900 3262
rect 46848 3198 46900 3204
rect 46940 3256 46992 3262
rect 46940 3198 46992 3204
rect 48136 3256 48188 3262
rect 48136 3198 48188 3204
rect 44548 3188 44600 3194
rect 44548 3130 44600 3136
rect 43352 3120 43404 3126
rect 43352 3062 43404 3068
rect 43364 480 43392 3062
rect 44560 480 44588 3130
rect 45756 480 45784 3198
rect 46952 480 46980 3198
rect 48240 2530 48268 5034
rect 49620 3482 49648 318718
rect 69018 318679 69074 318688
rect 70214 318744 70270 318753
rect 70214 318679 70270 318688
rect 50988 317960 51040 317966
rect 50988 317902 51040 317908
rect 48148 2502 48268 2530
rect 49344 3454 49648 3482
rect 48148 480 48176 2502
rect 49344 480 49372 3454
rect 51000 3262 51028 317902
rect 56416 317892 56468 317898
rect 56416 317834 56468 317840
rect 55220 5228 55272 5234
rect 55220 5170 55272 5176
rect 51632 5160 51684 5166
rect 51632 5102 51684 5108
rect 50528 3256 50580 3262
rect 50528 3198 50580 3204
rect 50988 3256 51040 3262
rect 50988 3198 51040 3204
rect 50540 480 50568 3198
rect 51644 480 51672 5102
rect 54024 3188 54076 3194
rect 54024 3130 54076 3136
rect 52828 2916 52880 2922
rect 52828 2858 52880 2864
rect 52840 480 52868 2858
rect 54036 480 54064 3130
rect 55232 480 55260 5170
rect 56428 480 56456 317834
rect 57888 317824 57940 317830
rect 57888 317766 57940 317772
rect 57900 3482 57928 317766
rect 64788 317756 64840 317762
rect 64788 317698 64840 317704
rect 63408 317688 63460 317694
rect 63408 317630 63460 317636
rect 58808 5296 58860 5302
rect 58808 5238 58860 5244
rect 57624 3454 57928 3482
rect 57624 480 57652 3454
rect 58820 480 58848 5238
rect 63420 3126 63448 317630
rect 64696 317552 64748 317558
rect 64696 317494 64748 317500
rect 62396 3120 62448 3126
rect 62396 3062 62448 3068
rect 63408 3120 63460 3126
rect 63408 3062 63460 3068
rect 61200 3052 61252 3058
rect 61200 2994 61252 3000
rect 60004 2984 60056 2990
rect 60004 2926 60056 2932
rect 60016 480 60044 2926
rect 61212 480 61240 2994
rect 62408 480 62436 3062
rect 64708 3058 64736 317494
rect 63592 3052 63644 3058
rect 63592 2994 63644 3000
rect 64696 3052 64748 3058
rect 64696 2994 64748 3000
rect 63604 480 63632 2994
rect 64800 480 64828 317698
rect 68284 317484 68336 317490
rect 68284 317426 68336 317432
rect 67180 2984 67232 2990
rect 68296 2938 68324 317426
rect 69032 4894 69060 318679
rect 69664 317484 69716 317490
rect 69664 317426 69716 317432
rect 69020 4888 69072 4894
rect 69020 4830 69072 4836
rect 69676 3074 69704 317426
rect 70400 315988 70452 315994
rect 70400 315930 70452 315936
rect 70412 3466 70440 315930
rect 70504 313970 70532 319382
rect 70504 313942 70624 313970
rect 70596 302326 70624 313942
rect 70872 309194 70900 319382
rect 71056 315994 71084 320062
rect 71044 315988 71096 315994
rect 71044 315930 71096 315936
rect 70860 309188 70912 309194
rect 70860 309130 70912 309136
rect 70860 307828 70912 307834
rect 70860 307770 70912 307776
rect 70584 302320 70636 302326
rect 70584 302262 70636 302268
rect 70492 302184 70544 302190
rect 70492 302126 70544 302132
rect 70504 299470 70532 302126
rect 70872 299538 70900 307770
rect 70676 299532 70728 299538
rect 70676 299474 70728 299480
rect 70860 299532 70912 299538
rect 70860 299474 70912 299480
rect 70492 299464 70544 299470
rect 70492 299406 70544 299412
rect 70688 299418 70716 299474
rect 70688 299390 70808 299418
rect 70780 298110 70808 299390
rect 70768 298104 70820 298110
rect 70768 298046 70820 298052
rect 70584 289876 70636 289882
rect 70584 289818 70636 289824
rect 70596 280106 70624 289818
rect 70768 288448 70820 288454
rect 70768 288390 70820 288396
rect 70780 282946 70808 288390
rect 70768 282940 70820 282946
rect 70768 282882 70820 282888
rect 70860 282872 70912 282878
rect 70860 282814 70912 282820
rect 70596 280078 70716 280106
rect 70688 264110 70716 280078
rect 70872 270570 70900 282814
rect 70768 270564 70820 270570
rect 70768 270506 70820 270512
rect 70860 270564 70912 270570
rect 70860 270506 70912 270512
rect 70492 264104 70544 264110
rect 70492 264046 70544 264052
rect 70676 264104 70728 264110
rect 70676 264046 70728 264052
rect 70504 253910 70532 264046
rect 70780 263634 70808 270506
rect 70768 263628 70820 263634
rect 70768 263570 70820 263576
rect 70676 263560 70728 263566
rect 70676 263502 70728 263508
rect 70688 259418 70716 263502
rect 70676 259412 70728 259418
rect 70676 259354 70728 259360
rect 70492 253904 70544 253910
rect 70492 253846 70544 253852
rect 70676 253904 70728 253910
rect 70676 253846 70728 253852
rect 70688 244390 70716 253846
rect 70676 244384 70728 244390
rect 70676 244326 70728 244332
rect 70492 244316 70544 244322
rect 70492 244258 70544 244264
rect 70504 234598 70532 244258
rect 70768 241528 70820 241534
rect 70768 241470 70820 241476
rect 70780 234598 70808 241470
rect 70492 234592 70544 234598
rect 70492 234534 70544 234540
rect 70676 234592 70728 234598
rect 70676 234534 70728 234540
rect 70768 234592 70820 234598
rect 70768 234534 70820 234540
rect 70688 225078 70716 234534
rect 70768 231872 70820 231878
rect 70768 231814 70820 231820
rect 70676 225072 70728 225078
rect 70676 225014 70728 225020
rect 70492 225004 70544 225010
rect 70492 224946 70544 224952
rect 70504 215286 70532 224946
rect 70780 215286 70808 231814
rect 70492 215280 70544 215286
rect 70492 215222 70544 215228
rect 70676 215280 70728 215286
rect 70676 215222 70728 215228
rect 70768 215280 70820 215286
rect 70768 215222 70820 215228
rect 70688 205766 70716 215222
rect 70768 212560 70820 212566
rect 70768 212502 70820 212508
rect 70676 205760 70728 205766
rect 70676 205702 70728 205708
rect 70492 205692 70544 205698
rect 70492 205634 70544 205640
rect 70504 195974 70532 205634
rect 70780 195974 70808 212502
rect 70492 195968 70544 195974
rect 70492 195910 70544 195916
rect 70676 195968 70728 195974
rect 70676 195910 70728 195916
rect 70768 195968 70820 195974
rect 70768 195910 70820 195916
rect 70688 186454 70716 195910
rect 70768 193248 70820 193254
rect 70768 193190 70820 193196
rect 70676 186448 70728 186454
rect 70676 186390 70728 186396
rect 70492 186380 70544 186386
rect 70492 186322 70544 186328
rect 70504 176662 70532 186322
rect 70780 176662 70808 193190
rect 70492 176656 70544 176662
rect 70492 176598 70544 176604
rect 70676 176656 70728 176662
rect 70676 176598 70728 176604
rect 70768 176656 70820 176662
rect 70768 176598 70820 176604
rect 70688 167142 70716 176598
rect 70768 173936 70820 173942
rect 70768 173878 70820 173884
rect 70676 167136 70728 167142
rect 70676 167078 70728 167084
rect 70492 167068 70544 167074
rect 70492 167010 70544 167016
rect 70504 157350 70532 167010
rect 70780 157486 70808 173878
rect 70768 157480 70820 157486
rect 70768 157422 70820 157428
rect 70492 157344 70544 157350
rect 70492 157286 70544 157292
rect 70768 157344 70820 157350
rect 70768 157286 70820 157292
rect 70676 154624 70728 154630
rect 70676 154566 70728 154572
rect 70492 147688 70544 147694
rect 70492 147630 70544 147636
rect 70504 140026 70532 147630
rect 70688 140434 70716 154566
rect 70780 147694 70808 157286
rect 70768 147688 70820 147694
rect 70768 147630 70820 147636
rect 70688 140406 70992 140434
rect 70504 139998 70716 140026
rect 70688 128450 70716 139998
rect 70964 135289 70992 140406
rect 70766 135280 70822 135289
rect 70766 135215 70822 135224
rect 70950 135280 71006 135289
rect 70950 135215 71006 135224
rect 70780 128450 70808 135215
rect 70676 128444 70728 128450
rect 70676 128386 70728 128392
rect 70768 128444 70820 128450
rect 70768 128386 70820 128392
rect 70492 128376 70544 128382
rect 70492 128318 70544 128324
rect 70504 125594 70532 128318
rect 70584 128308 70636 128314
rect 70584 128250 70636 128256
rect 70492 125588 70544 125594
rect 70492 125530 70544 125536
rect 70596 125526 70624 128250
rect 70676 125588 70728 125594
rect 70676 125530 70728 125536
rect 70584 125520 70636 125526
rect 70584 125462 70636 125468
rect 70688 109138 70716 125530
rect 70768 125520 70820 125526
rect 70768 125462 70820 125468
rect 70780 124166 70808 125462
rect 70768 124160 70820 124166
rect 70768 124102 70820 124108
rect 70860 124160 70912 124166
rect 70860 124102 70912 124108
rect 70676 109132 70728 109138
rect 70676 109074 70728 109080
rect 70492 109064 70544 109070
rect 70492 109006 70544 109012
rect 70504 95266 70532 109006
rect 70872 104854 70900 124102
rect 70860 104848 70912 104854
rect 70860 104790 70912 104796
rect 70768 95328 70820 95334
rect 70768 95270 70820 95276
rect 70492 95260 70544 95266
rect 70492 95202 70544 95208
rect 70676 95260 70728 95266
rect 70676 95202 70728 95208
rect 70688 89826 70716 95202
rect 70780 95198 70808 95270
rect 70768 95192 70820 95198
rect 70768 95134 70820 95140
rect 70952 95192 71004 95198
rect 70952 95134 71004 95140
rect 70676 89820 70728 89826
rect 70676 89762 70728 89768
rect 70492 89752 70544 89758
rect 70492 89694 70544 89700
rect 70504 83858 70532 89694
rect 70504 83830 70716 83858
rect 70688 71466 70716 83830
rect 70964 77353 70992 95134
rect 70766 77344 70822 77353
rect 70766 77279 70822 77288
rect 70950 77344 71006 77353
rect 70950 77279 71006 77288
rect 70492 71460 70544 71466
rect 70492 71402 70544 71408
rect 70676 71460 70728 71466
rect 70676 71402 70728 71408
rect 70504 67182 70532 71402
rect 70780 70514 70808 77279
rect 70768 70508 70820 70514
rect 70768 70450 70820 70456
rect 70676 70372 70728 70378
rect 70676 70314 70728 70320
rect 70688 67590 70716 70314
rect 70676 67584 70728 67590
rect 70676 67526 70728 67532
rect 70492 67176 70544 67182
rect 70492 67118 70544 67124
rect 70676 67176 70728 67182
rect 70676 67118 70728 67124
rect 70688 53174 70716 67118
rect 70768 57996 70820 58002
rect 70768 57938 70820 57944
rect 70492 53168 70544 53174
rect 70492 53110 70544 53116
rect 70676 53168 70728 53174
rect 70676 53110 70728 53116
rect 70504 41410 70532 53110
rect 70780 51134 70808 57938
rect 70768 51128 70820 51134
rect 70768 51070 70820 51076
rect 70676 51060 70728 51066
rect 70676 51002 70728 51008
rect 70688 46186 70716 51002
rect 70596 46158 70716 46186
rect 70492 41404 70544 41410
rect 70492 41346 70544 41352
rect 70596 41342 70624 46158
rect 70676 41404 70728 41410
rect 70676 41346 70728 41352
rect 70584 41336 70636 41342
rect 70584 41278 70636 41284
rect 70688 33862 70716 41346
rect 70768 41336 70820 41342
rect 70768 41278 70820 41284
rect 70492 33856 70544 33862
rect 70492 33798 70544 33804
rect 70676 33856 70728 33862
rect 70676 33798 70728 33804
rect 70504 22710 70532 33798
rect 70780 31822 70808 41278
rect 70768 31816 70820 31822
rect 70768 31758 70820 31764
rect 70676 31748 70728 31754
rect 70676 31690 70728 31696
rect 70688 22930 70716 31690
rect 70688 22902 70808 22930
rect 70492 22704 70544 22710
rect 70492 22646 70544 22652
rect 70676 22704 70728 22710
rect 70676 22646 70728 22652
rect 70688 12578 70716 22646
rect 70676 12572 70728 12578
rect 70676 12514 70728 12520
rect 70492 12504 70544 12510
rect 70492 12446 70544 12452
rect 70504 4826 70532 12446
rect 70780 4962 70808 22902
rect 70768 4956 70820 4962
rect 70768 4898 70820 4904
rect 70492 4820 70544 4826
rect 70492 4762 70544 4768
rect 71792 4162 71820 320076
rect 71976 320062 72266 320090
rect 72436 320062 72634 320090
rect 72712 320062 73094 320090
rect 73462 320062 73568 320090
rect 71872 315988 71924 315994
rect 71872 315930 71924 315936
rect 71700 4134 71820 4162
rect 70400 3460 70452 3466
rect 70400 3402 70452 3408
rect 71700 3369 71728 4134
rect 71884 4026 71912 315930
rect 71792 3998 71912 4026
rect 71792 3602 71820 3998
rect 71872 3936 71924 3942
rect 71872 3878 71924 3884
rect 71780 3596 71832 3602
rect 71780 3538 71832 3544
rect 71686 3360 71742 3369
rect 71686 3295 71742 3304
rect 67180 2926 67232 2932
rect 65984 2848 66036 2854
rect 65984 2790 66036 2796
rect 65996 480 66024 2790
rect 67192 480 67220 2926
rect 68204 2910 68324 2938
rect 69400 3046 69704 3074
rect 69400 2922 69428 3046
rect 69388 2916 69440 2922
rect 68204 2854 68232 2910
rect 69388 2858 69440 2864
rect 69480 2916 69532 2922
rect 69480 2858 69532 2864
rect 68192 2848 68244 2854
rect 68192 2790 68244 2796
rect 68284 2848 68336 2854
rect 68284 2790 68336 2796
rect 68296 480 68324 2790
rect 69492 480 69520 2858
rect 70676 1012 70728 1018
rect 70676 954 70728 960
rect 70688 480 70716 954
rect 71884 480 71912 3878
rect 71976 3534 72004 320062
rect 72436 309312 72464 320062
rect 72712 315994 72740 320062
rect 72700 315988 72752 315994
rect 72700 315930 72752 315936
rect 73160 315988 73212 315994
rect 73160 315930 73212 315936
rect 72344 309284 72464 309312
rect 72344 309210 72372 309284
rect 72252 309182 72372 309210
rect 72252 302410 72280 309182
rect 72252 302382 72372 302410
rect 72344 302138 72372 302382
rect 72160 302110 72372 302138
rect 72160 296682 72188 302110
rect 72148 296676 72200 296682
rect 72148 296618 72200 296624
rect 72332 288380 72384 288386
rect 72332 288322 72384 288328
rect 72344 287065 72372 288322
rect 72330 287056 72386 287065
rect 72330 286991 72386 287000
rect 72514 287056 72570 287065
rect 72514 286991 72570 287000
rect 72528 277438 72556 286991
rect 72332 277432 72384 277438
rect 72330 277400 72332 277409
rect 72516 277432 72568 277438
rect 72384 277400 72386 277409
rect 72516 277374 72568 277380
rect 72606 277400 72662 277409
rect 72330 277335 72386 277344
rect 72606 277335 72662 277344
rect 72620 267782 72648 277335
rect 72424 267776 72476 267782
rect 72424 267718 72476 267724
rect 72608 267776 72660 267782
rect 72608 267718 72660 267724
rect 72436 249830 72464 267718
rect 72148 249824 72200 249830
rect 72424 249824 72476 249830
rect 72200 249772 72280 249778
rect 72148 249766 72280 249772
rect 72424 249766 72476 249772
rect 72160 249750 72280 249766
rect 72252 240174 72280 249750
rect 72240 240168 72292 240174
rect 72240 240110 72292 240116
rect 72424 240168 72476 240174
rect 72424 240110 72476 240116
rect 72436 231878 72464 240110
rect 72148 231872 72200 231878
rect 72148 231814 72200 231820
rect 72424 231872 72476 231878
rect 72424 231814 72476 231820
rect 72160 222222 72188 231814
rect 72148 222216 72200 222222
rect 72148 222158 72200 222164
rect 72424 222216 72476 222222
rect 72424 222158 72476 222164
rect 72436 212566 72464 222158
rect 72148 212560 72200 212566
rect 72148 212502 72200 212508
rect 72424 212560 72476 212566
rect 72424 212502 72476 212508
rect 72160 202910 72188 212502
rect 72148 202904 72200 202910
rect 72148 202846 72200 202852
rect 72424 202904 72476 202910
rect 72424 202846 72476 202852
rect 72436 193254 72464 202846
rect 72148 193248 72200 193254
rect 72148 193190 72200 193196
rect 72424 193248 72476 193254
rect 72424 193190 72476 193196
rect 72160 191826 72188 193190
rect 72056 191820 72108 191826
rect 72056 191762 72108 191768
rect 72148 191820 72200 191826
rect 72148 191762 72200 191768
rect 72068 182209 72096 191762
rect 72054 182200 72110 182209
rect 72054 182135 72110 182144
rect 72330 182200 72386 182209
rect 72330 182135 72386 182144
rect 72344 174078 72372 182135
rect 72332 174072 72384 174078
rect 72332 174014 72384 174020
rect 72332 171148 72384 171154
rect 72332 171090 72384 171096
rect 72344 151842 72372 171090
rect 72148 151836 72200 151842
rect 72148 151778 72200 151784
rect 72332 151836 72384 151842
rect 72332 151778 72384 151784
rect 72160 143546 72188 151778
rect 72148 143540 72200 143546
rect 72148 143482 72200 143488
rect 72332 143540 72384 143546
rect 72332 143482 72384 143488
rect 72344 133890 72372 143482
rect 72332 133884 72384 133890
rect 72332 133826 72384 133832
rect 72332 124228 72384 124234
rect 72332 124170 72384 124176
rect 72344 116090 72372 124170
rect 72252 116062 72372 116090
rect 72252 114578 72280 116062
rect 72148 114572 72200 114578
rect 72148 114514 72200 114520
rect 72240 114572 72292 114578
rect 72240 114514 72292 114520
rect 72160 108984 72188 114514
rect 72160 108956 72280 108984
rect 72252 106282 72280 108956
rect 72240 106276 72292 106282
rect 72240 106218 72292 106224
rect 72240 96756 72292 96762
rect 72240 96698 72292 96704
rect 72252 87145 72280 96698
rect 72238 87136 72294 87145
rect 72238 87071 72294 87080
rect 72146 87000 72202 87009
rect 72146 86935 72202 86944
rect 72160 85542 72188 86935
rect 72148 85536 72200 85542
rect 72148 85478 72200 85484
rect 72148 75948 72200 75954
rect 72148 75890 72200 75896
rect 72160 72486 72188 75890
rect 72148 72480 72200 72486
rect 72148 72422 72200 72428
rect 72148 67720 72200 67726
rect 72148 67662 72200 67668
rect 72160 66230 72188 67662
rect 72148 66224 72200 66230
rect 72148 66166 72200 66172
rect 72056 56636 72108 56642
rect 72056 56578 72108 56584
rect 72068 48346 72096 56578
rect 72056 48340 72108 48346
rect 72056 48282 72108 48288
rect 72240 48340 72292 48346
rect 72240 48282 72292 48288
rect 72252 46918 72280 48282
rect 72240 46912 72292 46918
rect 72240 46854 72292 46860
rect 72056 37324 72108 37330
rect 72056 37266 72108 37272
rect 72068 29034 72096 37266
rect 72056 29028 72108 29034
rect 72056 28970 72108 28976
rect 72240 29028 72292 29034
rect 72240 28970 72292 28976
rect 72252 22166 72280 28970
rect 72240 22160 72292 22166
rect 72240 22102 72292 22108
rect 72148 22092 72200 22098
rect 72148 22034 72200 22040
rect 72160 5030 72188 22034
rect 72148 5024 72200 5030
rect 72148 4966 72200 4972
rect 73172 3806 73200 315930
rect 73252 315308 73304 315314
rect 73252 315250 73304 315256
rect 73160 3800 73212 3806
rect 73160 3742 73212 3748
rect 73264 3670 73292 315250
rect 73540 310570 73568 320062
rect 73632 320062 73922 320090
rect 74000 320062 74290 320090
rect 73632 315314 73660 320062
rect 74000 315994 74028 320062
rect 74736 318073 74764 320076
rect 75104 318209 75132 320076
rect 75564 318345 75592 320076
rect 75932 318481 75960 320076
rect 76116 320062 76406 320090
rect 76484 320062 76774 320090
rect 76944 320062 77234 320090
rect 75918 318472 75974 318481
rect 75918 318407 75974 318416
rect 75550 318336 75606 318345
rect 75550 318271 75606 318280
rect 75090 318200 75146 318209
rect 75090 318135 75146 318144
rect 74722 318064 74778 318073
rect 74722 317999 74778 318008
rect 75920 316056 75972 316062
rect 75920 315998 75972 316004
rect 73988 315988 74040 315994
rect 73988 315930 74040 315936
rect 73620 315308 73672 315314
rect 73620 315250 73672 315256
rect 73540 310542 73660 310570
rect 73632 307834 73660 310542
rect 73528 307828 73580 307834
rect 73528 307770 73580 307776
rect 73620 307828 73672 307834
rect 73620 307770 73672 307776
rect 73540 299470 73568 307770
rect 73436 299464 73488 299470
rect 73436 299406 73488 299412
rect 73528 299464 73580 299470
rect 73528 299406 73580 299412
rect 73448 298110 73476 299406
rect 73436 298104 73488 298110
rect 73436 298046 73488 298052
rect 73528 298104 73580 298110
rect 73528 298046 73580 298052
rect 73540 278866 73568 298046
rect 73436 278860 73488 278866
rect 73436 278802 73488 278808
rect 73528 278860 73580 278866
rect 73528 278802 73580 278808
rect 73448 277409 73476 278802
rect 73434 277400 73490 277409
rect 73434 277335 73490 277344
rect 73618 277400 73674 277409
rect 73618 277335 73674 277344
rect 73632 267782 73660 277335
rect 73436 267776 73488 267782
rect 73436 267718 73488 267724
rect 73620 267776 73672 267782
rect 73620 267718 73672 267724
rect 73448 263634 73476 267718
rect 73436 263628 73488 263634
rect 73436 263570 73488 263576
rect 73528 263492 73580 263498
rect 73528 263434 73580 263440
rect 73540 252618 73568 263434
rect 73528 252612 73580 252618
rect 73528 252554 73580 252560
rect 73712 241528 73764 241534
rect 73712 241470 73764 241476
rect 73724 231878 73752 241470
rect 73436 231872 73488 231878
rect 73434 231840 73436 231849
rect 73712 231872 73764 231878
rect 73488 231840 73490 231849
rect 73434 231775 73490 231784
rect 73710 231840 73712 231849
rect 73764 231840 73766 231849
rect 73710 231775 73766 231784
rect 73724 212566 73752 231775
rect 73436 212560 73488 212566
rect 73434 212528 73436 212537
rect 73712 212560 73764 212566
rect 73488 212528 73490 212537
rect 73434 212463 73490 212472
rect 73710 212528 73712 212537
rect 73764 212528 73766 212537
rect 73710 212463 73766 212472
rect 73724 193254 73752 212463
rect 73436 193248 73488 193254
rect 73436 193190 73488 193196
rect 73712 193248 73764 193254
rect 73712 193190 73764 193196
rect 73448 191826 73476 193190
rect 73344 191820 73396 191826
rect 73344 191762 73396 191768
rect 73436 191820 73488 191826
rect 73436 191762 73488 191768
rect 73356 182209 73384 191762
rect 73342 182200 73398 182209
rect 73342 182135 73398 182144
rect 73618 182200 73674 182209
rect 73618 182135 73674 182144
rect 73632 173942 73660 182135
rect 73436 173936 73488 173942
rect 73436 173878 73488 173884
rect 73620 173936 73672 173942
rect 73620 173878 73672 173884
rect 73448 172514 73476 173878
rect 73344 172508 73396 172514
rect 73344 172450 73396 172456
rect 73436 172508 73488 172514
rect 73436 172450 73488 172456
rect 73356 162897 73384 172450
rect 73342 162888 73398 162897
rect 73342 162823 73398 162832
rect 73618 162888 73674 162897
rect 73618 162823 73674 162832
rect 73632 154630 73660 162823
rect 73528 154624 73580 154630
rect 73448 154572 73528 154578
rect 73448 154566 73580 154572
rect 73620 154624 73672 154630
rect 73620 154566 73672 154572
rect 73448 154550 73568 154566
rect 73448 153202 73476 154550
rect 73436 153196 73488 153202
rect 73436 153138 73488 153144
rect 73436 144900 73488 144906
rect 73436 144842 73488 144848
rect 73448 143562 73476 144842
rect 73448 143534 73568 143562
rect 73540 143478 73568 143534
rect 73528 143472 73580 143478
rect 73528 143414 73580 143420
rect 73620 131572 73672 131578
rect 73620 131514 73672 131520
rect 73632 116090 73660 131514
rect 73540 116062 73660 116090
rect 73540 114578 73568 116062
rect 73436 114572 73488 114578
rect 73436 114514 73488 114520
rect 73528 114572 73580 114578
rect 73528 114514 73580 114520
rect 73448 108882 73476 114514
rect 73448 108854 73568 108882
rect 73540 106282 73568 108854
rect 73528 106276 73580 106282
rect 73528 106218 73580 106224
rect 73620 95260 73672 95266
rect 73620 95202 73672 95208
rect 73632 87009 73660 95202
rect 73434 87000 73490 87009
rect 73434 86935 73490 86944
rect 73618 87000 73674 87009
rect 73618 86935 73674 86944
rect 73448 85542 73476 86935
rect 73436 85536 73488 85542
rect 73436 85478 73488 85484
rect 73528 75948 73580 75954
rect 73528 75890 73580 75896
rect 73540 62778 73568 75890
rect 73448 62750 73568 62778
rect 73448 48414 73476 62750
rect 73436 48408 73488 48414
rect 73436 48350 73488 48356
rect 73528 48340 73580 48346
rect 73528 48282 73580 48288
rect 73540 46918 73568 48282
rect 73528 46912 73580 46918
rect 73528 46854 73580 46860
rect 73436 37324 73488 37330
rect 73436 37266 73488 37272
rect 73448 36310 73476 37266
rect 73436 36304 73488 36310
rect 73436 36246 73488 36252
rect 73528 29028 73580 29034
rect 73528 28970 73580 28976
rect 73540 22658 73568 28970
rect 73448 22630 73568 22658
rect 73448 17950 73476 22630
rect 73436 17944 73488 17950
rect 73436 17886 73488 17892
rect 73344 8356 73396 8362
rect 73344 8298 73396 8304
rect 73252 3664 73304 3670
rect 73252 3606 73304 3612
rect 71964 3528 72016 3534
rect 71964 3470 72016 3476
rect 73068 3528 73120 3534
rect 73356 3505 73384 8298
rect 75932 3777 75960 315998
rect 76012 315988 76064 315994
rect 76012 315930 76064 315936
rect 76024 3874 76052 315930
rect 76012 3868 76064 3874
rect 76012 3810 76064 3816
rect 75918 3768 75974 3777
rect 75918 3703 75974 3712
rect 75460 3664 75512 3670
rect 76116 3641 76144 320062
rect 76484 316062 76512 320062
rect 76472 316056 76524 316062
rect 76472 315998 76524 316004
rect 76944 315994 76972 320062
rect 77404 319410 77432 320198
rect 77404 319382 77524 319410
rect 77496 318764 77524 319382
rect 77496 318736 77616 318764
rect 76932 315988 76984 315994
rect 76932 315930 76984 315936
rect 77588 309330 77616 318736
rect 78048 318617 78076 320076
rect 78034 318608 78090 318617
rect 78034 318543 78090 318552
rect 78416 318170 78444 320076
rect 78876 318442 78904 320076
rect 78864 318436 78916 318442
rect 78864 318378 78916 318384
rect 79244 318306 79272 320076
rect 79428 320062 79718 320090
rect 80086 320062 80192 320090
rect 79232 318300 79284 318306
rect 79232 318242 79284 318248
rect 78404 318164 78456 318170
rect 78404 318106 78456 318112
rect 77576 309324 77628 309330
rect 77576 309266 77628 309272
rect 79428 309194 79456 320062
rect 77576 309188 77628 309194
rect 77576 309130 77628 309136
rect 78956 309188 79008 309194
rect 78956 309130 79008 309136
rect 79416 309188 79468 309194
rect 79416 309130 79468 309136
rect 77588 309074 77616 309130
rect 77588 309046 77708 309074
rect 77680 289882 77708 309046
rect 78968 289950 78996 309130
rect 78956 289944 79008 289950
rect 78956 289886 79008 289892
rect 77576 289876 77628 289882
rect 77576 289818 77628 289824
rect 77668 289876 77720 289882
rect 77668 289818 77720 289824
rect 78864 289876 78916 289882
rect 78864 289818 78916 289824
rect 77588 283014 77616 289818
rect 78876 288402 78904 289818
rect 78784 288374 78904 288402
rect 77576 283008 77628 283014
rect 77576 282950 77628 282956
rect 78784 282946 78812 288374
rect 78772 282940 78824 282946
rect 78772 282882 78824 282888
rect 77484 282872 77536 282878
rect 77484 282814 77536 282820
rect 77496 270502 77524 282814
rect 78864 278792 78916 278798
rect 78864 278734 78916 278740
rect 78876 270502 78904 278734
rect 77484 270496 77536 270502
rect 77484 270438 77536 270444
rect 77576 270496 77628 270502
rect 77576 270438 77628 270444
rect 78680 270496 78732 270502
rect 78680 270438 78732 270444
rect 78864 270496 78916 270502
rect 78864 270438 78916 270444
rect 77588 253178 77616 270438
rect 78692 267753 78720 270438
rect 78678 267744 78734 267753
rect 78678 267679 78734 267688
rect 78954 267744 79010 267753
rect 78954 267679 79010 267688
rect 77496 253150 77616 253178
rect 77496 248441 77524 253150
rect 78968 248470 78996 267679
rect 78772 248464 78824 248470
rect 77482 248432 77538 248441
rect 77482 248367 77538 248376
rect 77850 248432 77906 248441
rect 78772 248406 78824 248412
rect 78956 248464 79008 248470
rect 78956 248406 79008 248412
rect 77850 248367 77906 248376
rect 77864 245002 77892 248367
rect 77668 244996 77720 245002
rect 77668 244938 77720 244944
rect 77852 244996 77904 245002
rect 77852 244938 77904 244944
rect 77680 230466 77708 244938
rect 78784 240174 78812 248406
rect 78772 240168 78824 240174
rect 78772 240110 78824 240116
rect 78864 240100 78916 240106
rect 78864 240042 78916 240048
rect 77680 230438 77800 230466
rect 77772 225690 77800 230438
rect 78876 229106 78904 240042
rect 78876 229090 78996 229106
rect 78876 229084 79008 229090
rect 78876 229078 78956 229084
rect 78956 229026 79008 229032
rect 78968 228995 78996 229026
rect 77760 225684 77812 225690
rect 77760 225626 77812 225632
rect 78772 219496 78824 219502
rect 78772 219438 78824 219444
rect 77576 217388 77628 217394
rect 77576 217330 77628 217336
rect 77588 212514 77616 217330
rect 77496 212486 77616 212514
rect 77496 205698 77524 212486
rect 78784 211206 78812 219438
rect 78680 211200 78732 211206
rect 78680 211142 78732 211148
rect 78772 211200 78824 211206
rect 78772 211142 78824 211148
rect 77484 205692 77536 205698
rect 77484 205634 77536 205640
rect 78692 203538 78720 211142
rect 78692 203510 78812 203538
rect 77484 202904 77536 202910
rect 77482 202872 77484 202881
rect 78784 202881 78812 203510
rect 77536 202872 77538 202881
rect 77482 202807 77538 202816
rect 78770 202872 78826 202881
rect 78770 202807 78826 202816
rect 78862 202736 78918 202745
rect 78862 202671 78918 202680
rect 77574 195800 77630 195809
rect 77574 195735 77630 195744
rect 77588 186454 77616 195735
rect 78876 193202 78904 202671
rect 78784 193174 78904 193202
rect 77576 186448 77628 186454
rect 77576 186390 77628 186396
rect 78784 186386 78812 193174
rect 78772 186380 78824 186386
rect 78772 186322 78824 186328
rect 77484 186312 77536 186318
rect 77484 186254 77536 186260
rect 77496 183530 77524 186254
rect 78784 183598 78812 183629
rect 78772 183592 78824 183598
rect 78824 183540 78904 183546
rect 78772 183534 78904 183540
rect 77484 183524 77536 183530
rect 78784 183518 78904 183534
rect 77484 183466 77536 183472
rect 78876 183410 78904 183518
rect 78784 183382 78904 183410
rect 78784 173942 78812 183382
rect 77576 173936 77628 173942
rect 77576 173878 77628 173884
rect 78772 173936 78824 173942
rect 78772 173878 78824 173884
rect 78864 173936 78916 173942
rect 78864 173878 78916 173884
rect 77588 167686 77616 173878
rect 78876 167686 78904 173878
rect 77392 167680 77444 167686
rect 77392 167622 77444 167628
rect 77576 167680 77628 167686
rect 77576 167622 77628 167628
rect 78680 167680 78732 167686
rect 78680 167622 78732 167628
rect 78864 167680 78916 167686
rect 78864 167622 78916 167628
rect 77404 162874 77432 167622
rect 78692 162874 78720 167622
rect 77404 162846 77524 162874
rect 78692 162846 78812 162874
rect 77496 153202 77524 162846
rect 78784 153202 78812 162846
rect 77484 153196 77536 153202
rect 77484 153138 77536 153144
rect 78772 153196 78824 153202
rect 78772 153138 78824 153144
rect 77668 153060 77720 153066
rect 77668 153002 77720 153008
rect 78956 153060 79008 153066
rect 78956 153002 79008 153008
rect 77680 125633 77708 153002
rect 78968 125633 78996 153002
rect 77482 125624 77538 125633
rect 77482 125559 77538 125568
rect 77666 125624 77722 125633
rect 77666 125559 77722 125568
rect 78770 125624 78826 125633
rect 78770 125559 78826 125568
rect 78954 125624 79010 125633
rect 78954 125559 79010 125568
rect 77496 120714 77524 125559
rect 78784 120714 78812 125559
rect 77496 120686 77616 120714
rect 78784 120686 78904 120714
rect 77588 109138 77616 120686
rect 78876 115938 78904 120686
rect 78864 115932 78916 115938
rect 78864 115874 78916 115880
rect 77576 109132 77628 109138
rect 77576 109074 77628 109080
rect 77484 108996 77536 109002
rect 77484 108938 77536 108944
rect 77496 96642 77524 108938
rect 78772 106344 78824 106350
rect 78772 106286 78824 106292
rect 78784 101402 78812 106286
rect 78784 101374 78904 101402
rect 77496 96614 77616 96642
rect 77588 87145 77616 96614
rect 78876 93838 78904 101374
rect 78864 93832 78916 93838
rect 78864 93774 78916 93780
rect 77574 87136 77630 87145
rect 77574 87071 77630 87080
rect 77482 87000 77538 87009
rect 77482 86935 77538 86944
rect 77496 85542 77524 86935
rect 77484 85536 77536 85542
rect 77484 85478 77536 85484
rect 78680 84312 78732 84318
rect 78680 84254 78732 84260
rect 78692 84182 78720 84254
rect 78680 84176 78732 84182
rect 78680 84118 78732 84124
rect 78864 84108 78916 84114
rect 78864 84050 78916 84056
rect 78876 82822 78904 84050
rect 78864 82816 78916 82822
rect 78864 82758 78916 82764
rect 77576 75948 77628 75954
rect 77576 75890 77628 75896
rect 77588 70514 77616 75890
rect 77576 70508 77628 70514
rect 77576 70450 77628 70456
rect 77484 70372 77536 70378
rect 77484 70314 77536 70320
rect 77496 66230 77524 70314
rect 77392 66224 77444 66230
rect 77392 66166 77444 66172
rect 77484 66224 77536 66230
rect 77484 66166 77536 66172
rect 77404 38758 77432 66166
rect 78680 64932 78732 64938
rect 78680 64874 78732 64880
rect 78692 61470 78720 64874
rect 78680 61464 78732 61470
rect 78680 61406 78732 61412
rect 78956 61464 79008 61470
rect 78956 61406 79008 61412
rect 78968 48346 78996 61406
rect 78772 48340 78824 48346
rect 78772 48282 78824 48288
rect 78956 48340 79008 48346
rect 78956 48282 79008 48288
rect 77392 38752 77444 38758
rect 77392 38694 77444 38700
rect 78784 38690 78812 48282
rect 78772 38684 78824 38690
rect 78772 38626 78824 38632
rect 77392 38616 77444 38622
rect 77392 38558 77444 38564
rect 77404 29050 77432 38558
rect 78772 37324 78824 37330
rect 78772 37266 78824 37272
rect 78784 29050 78812 37266
rect 77404 29022 77524 29050
rect 78784 29022 78996 29050
rect 77496 27606 77524 29022
rect 78968 27606 78996 29022
rect 77484 27600 77536 27606
rect 77484 27542 77536 27548
rect 78956 27600 79008 27606
rect 78956 27542 79008 27548
rect 77484 18012 77536 18018
rect 77484 17954 77536 17960
rect 78864 18012 78916 18018
rect 78864 17954 78916 17960
rect 77496 3806 77524 17954
rect 78876 3874 78904 17954
rect 80060 3936 80112 3942
rect 80164 3913 80192 320062
rect 80348 320062 80546 320090
rect 80348 4010 80376 320062
rect 80900 318170 80928 320076
rect 81360 318442 81388 320076
rect 81728 318510 81756 320076
rect 81912 319410 81940 320198
rect 82280 320062 82570 320090
rect 82938 320062 83044 320090
rect 81912 319382 82032 319410
rect 81716 318504 81768 318510
rect 81716 318446 81768 318452
rect 81348 318436 81400 318442
rect 81348 318378 81400 318384
rect 80888 318164 80940 318170
rect 80888 318106 80940 318112
rect 82004 316010 82032 319382
rect 81532 315988 81584 315994
rect 81532 315930 81584 315936
rect 81636 315982 82032 316010
rect 82280 315994 82308 320062
rect 82268 315988 82320 315994
rect 81544 4146 81572 315930
rect 81636 302138 81664 315982
rect 82268 315930 82320 315936
rect 81636 302110 81756 302138
rect 81728 289882 81756 302110
rect 81716 289876 81768 289882
rect 81716 289818 81768 289824
rect 81808 289876 81860 289882
rect 81808 289818 81860 289824
rect 81820 287065 81848 289818
rect 81622 287056 81678 287065
rect 81622 286991 81678 287000
rect 81806 287056 81862 287065
rect 81806 286991 81862 287000
rect 81636 278798 81664 286991
rect 81624 278792 81676 278798
rect 81624 278734 81676 278740
rect 81716 278724 81768 278730
rect 81716 278666 81768 278672
rect 81728 276010 81756 278666
rect 81716 276004 81768 276010
rect 81716 275946 81768 275952
rect 81900 276004 81952 276010
rect 81900 275946 81952 275952
rect 81912 258097 81940 275946
rect 81714 258088 81770 258097
rect 81714 258023 81770 258032
rect 81898 258088 81954 258097
rect 81898 258023 81954 258032
rect 81728 251054 81756 258023
rect 81716 251048 81768 251054
rect 81716 250990 81768 250996
rect 81716 250912 81768 250918
rect 81716 250854 81768 250860
rect 81728 241534 81756 250854
rect 81716 241528 81768 241534
rect 81716 241470 81768 241476
rect 81808 241460 81860 241466
rect 81808 241402 81860 241408
rect 81820 234666 81848 241402
rect 81808 234660 81860 234666
rect 81808 234602 81860 234608
rect 81808 234524 81860 234530
rect 81808 234466 81860 234472
rect 81820 222222 81848 234466
rect 81716 222216 81768 222222
rect 81714 222184 81716 222193
rect 81808 222216 81860 222222
rect 81768 222184 81770 222193
rect 81808 222158 81860 222164
rect 81714 222119 81770 222128
rect 81806 222048 81862 222057
rect 81806 221983 81862 221992
rect 81820 205578 81848 221983
rect 81728 205550 81848 205578
rect 81728 196042 81756 205550
rect 81716 196036 81768 196042
rect 81716 195978 81768 195984
rect 81808 195968 81860 195974
rect 81808 195910 81860 195916
rect 81820 186266 81848 195910
rect 81728 186238 81848 186266
rect 81728 183569 81756 186238
rect 81714 183560 81770 183569
rect 81714 183495 81770 183504
rect 81898 183560 81954 183569
rect 81898 183495 81954 183504
rect 81912 173942 81940 183495
rect 81808 173936 81860 173942
rect 81808 173878 81860 173884
rect 81900 173936 81952 173942
rect 81900 173878 81952 173884
rect 81820 167686 81848 173878
rect 81808 167680 81860 167686
rect 81808 167622 81860 167628
rect 81992 167680 82044 167686
rect 81992 167622 82044 167628
rect 82004 162874 82032 167622
rect 81912 162846 82032 162874
rect 81912 161430 81940 162846
rect 81900 161424 81952 161430
rect 81900 161366 81952 161372
rect 81900 144832 81952 144838
rect 81900 144774 81952 144780
rect 81912 143546 81940 144774
rect 81900 143540 81952 143546
rect 81900 143482 81952 143488
rect 82084 143540 82136 143546
rect 82084 143482 82136 143488
rect 82096 133929 82124 143482
rect 81898 133920 81954 133929
rect 81898 133855 81954 133864
rect 82082 133920 82138 133929
rect 82082 133855 82138 133864
rect 81912 125633 81940 133855
rect 81714 125624 81770 125633
rect 81714 125559 81770 125568
rect 81898 125624 81954 125633
rect 81898 125559 81954 125568
rect 81728 120714 81756 125559
rect 81728 120686 81848 120714
rect 81820 109138 81848 120686
rect 81808 109132 81860 109138
rect 81808 109074 81860 109080
rect 81716 108996 81768 109002
rect 81716 108938 81768 108944
rect 81728 96642 81756 108938
rect 81728 96614 81848 96642
rect 81820 87145 81848 96614
rect 81806 87136 81862 87145
rect 81806 87071 81862 87080
rect 81714 87000 81770 87009
rect 81714 86935 81770 86944
rect 81728 85542 81756 86935
rect 81716 85536 81768 85542
rect 81716 85478 81768 85484
rect 81808 75948 81860 75954
rect 81808 75890 81860 75896
rect 81820 70514 81848 75890
rect 81808 70508 81860 70514
rect 81808 70450 81860 70456
rect 81808 70372 81860 70378
rect 81808 70314 81860 70320
rect 81820 66337 81848 70314
rect 81806 66328 81862 66337
rect 81806 66263 81862 66272
rect 81806 66056 81862 66065
rect 81806 65991 81862 66000
rect 81820 51814 81848 65991
rect 81808 51808 81860 51814
rect 81808 51750 81860 51756
rect 81808 38684 81860 38690
rect 81808 38626 81860 38632
rect 81820 35306 81848 38626
rect 81728 35278 81848 35306
rect 81728 31634 81756 35278
rect 81728 31606 81940 31634
rect 81912 22114 81940 31606
rect 81728 22086 81940 22114
rect 81728 12458 81756 22086
rect 81728 12430 81848 12458
rect 81532 4140 81584 4146
rect 81532 4082 81584 4088
rect 81820 4078 81848 12430
rect 82636 4140 82688 4146
rect 82636 4082 82688 4088
rect 81808 4072 81860 4078
rect 81808 4014 81860 4020
rect 80336 4004 80388 4010
rect 80336 3946 80388 3952
rect 81440 4004 81492 4010
rect 81440 3946 81492 3952
rect 80060 3878 80112 3884
rect 80150 3904 80206 3913
rect 78864 3868 78916 3874
rect 78864 3810 78916 3816
rect 79048 3868 79100 3874
rect 79048 3810 79100 3816
rect 77484 3800 77536 3806
rect 77484 3742 77536 3748
rect 77852 3800 77904 3806
rect 77852 3742 77904 3748
rect 75460 3606 75512 3612
rect 76102 3632 76158 3641
rect 74264 3596 74316 3602
rect 74264 3538 74316 3544
rect 73068 3470 73120 3476
rect 73342 3496 73398 3505
rect 73080 480 73108 3470
rect 73342 3431 73398 3440
rect 74276 480 74304 3538
rect 75472 480 75500 3606
rect 76102 3567 76158 3576
rect 76656 3460 76708 3466
rect 76656 3402 76708 3408
rect 76668 480 76696 3402
rect 77864 480 77892 3742
rect 79060 480 79088 3810
rect 79784 3392 79836 3398
rect 79784 3334 79836 3340
rect 79796 3233 79824 3334
rect 80072 3233 80100 3878
rect 80150 3839 80206 3848
rect 80150 3360 80206 3369
rect 80150 3295 80206 3304
rect 79782 3224 79838 3233
rect 79782 3159 79838 3168
rect 80058 3224 80114 3233
rect 80164 3194 80192 3295
rect 80058 3159 80114 3168
rect 80152 3188 80204 3194
rect 80152 3130 80204 3136
rect 80244 3188 80296 3194
rect 80244 3130 80296 3136
rect 80256 480 80284 3130
rect 81452 480 81480 3946
rect 82544 3392 82596 3398
rect 82542 3360 82544 3369
rect 82596 3360 82598 3369
rect 82542 3295 82598 3304
rect 82648 480 82676 4082
rect 83016 3262 83044 320062
rect 83384 318102 83412 320076
rect 83752 318646 83780 320076
rect 83740 318640 83792 318646
rect 83740 318582 83792 318588
rect 84212 318578 84240 320076
rect 84304 320062 84594 320090
rect 84672 320062 85054 320090
rect 85132 320062 85422 320090
rect 84200 318572 84252 318578
rect 84200 318514 84252 318520
rect 83372 318096 83424 318102
rect 83372 318038 83424 318044
rect 84304 4049 84332 320062
rect 84672 316010 84700 320062
rect 84936 317824 84988 317830
rect 84396 315982 84700 316010
rect 84856 317784 84936 317812
rect 84396 4078 84424 315982
rect 84660 309188 84712 309194
rect 84660 309130 84712 309136
rect 84672 304314 84700 309130
rect 84580 304286 84700 304314
rect 84580 299418 84608 304286
rect 84580 299390 84700 299418
rect 84672 263634 84700 299390
rect 84476 263628 84528 263634
rect 84476 263570 84528 263576
rect 84660 263628 84712 263634
rect 84660 263570 84712 263576
rect 84488 263514 84516 263570
rect 84488 263486 84608 263514
rect 84580 253994 84608 263486
rect 84580 253966 84700 253994
rect 84672 244322 84700 253966
rect 84476 244316 84528 244322
rect 84476 244258 84528 244264
rect 84660 244316 84712 244322
rect 84660 244258 84712 244264
rect 84488 244202 84516 244258
rect 84488 244174 84608 244202
rect 84580 234682 84608 244174
rect 84580 234654 84700 234682
rect 84672 225010 84700 234654
rect 84476 225004 84528 225010
rect 84476 224946 84528 224952
rect 84660 225004 84712 225010
rect 84660 224946 84712 224952
rect 84488 224890 84516 224946
rect 84488 224862 84608 224890
rect 84580 215370 84608 224862
rect 84580 215342 84700 215370
rect 84672 205698 84700 215342
rect 84476 205692 84528 205698
rect 84476 205634 84528 205640
rect 84660 205692 84712 205698
rect 84660 205634 84712 205640
rect 84488 205578 84516 205634
rect 84488 205550 84608 205578
rect 84580 196058 84608 205550
rect 84580 196030 84700 196058
rect 84672 186386 84700 196030
rect 84476 186380 84528 186386
rect 84476 186322 84528 186328
rect 84660 186380 84712 186386
rect 84660 186322 84712 186328
rect 84488 186266 84516 186322
rect 84488 186238 84608 186266
rect 84580 179194 84608 186238
rect 84580 179166 84700 179194
rect 84672 167074 84700 179166
rect 84476 167068 84528 167074
rect 84476 167010 84528 167016
rect 84660 167068 84712 167074
rect 84660 167010 84712 167016
rect 84488 166954 84516 167010
rect 84488 166926 84608 166954
rect 84580 159338 84608 166926
rect 84580 159310 84700 159338
rect 84672 147694 84700 159310
rect 84476 147688 84528 147694
rect 84660 147688 84712 147694
rect 84528 147636 84608 147642
rect 84476 147630 84608 147636
rect 84660 147630 84712 147636
rect 84488 147614 84608 147630
rect 84580 140026 84608 147614
rect 84580 139998 84792 140026
rect 84764 137986 84792 139998
rect 84672 137958 84792 137986
rect 84672 128382 84700 137958
rect 84476 128376 84528 128382
rect 84660 128376 84712 128382
rect 84528 128324 84608 128330
rect 84476 128318 84608 128324
rect 84660 128318 84712 128324
rect 84488 128302 84608 128318
rect 84580 120714 84608 128302
rect 84580 120686 84792 120714
rect 84764 118674 84792 120686
rect 84672 118646 84792 118674
rect 84672 109070 84700 118646
rect 84476 109064 84528 109070
rect 84660 109064 84712 109070
rect 84528 109012 84608 109018
rect 84476 109006 84608 109012
rect 84660 109006 84712 109012
rect 84488 108990 84608 109006
rect 84580 101402 84608 108990
rect 84580 101374 84700 101402
rect 84672 89758 84700 101374
rect 84476 89752 84528 89758
rect 84660 89752 84712 89758
rect 84528 89700 84608 89706
rect 84476 89694 84608 89700
rect 84660 89694 84712 89700
rect 84488 89678 84608 89694
rect 84580 80084 84608 89678
rect 84580 80056 84700 80084
rect 84672 66298 84700 80056
rect 84568 66292 84620 66298
rect 84568 66234 84620 66240
rect 84660 66292 84712 66298
rect 84660 66234 84712 66240
rect 84580 60738 84608 66234
rect 84580 60710 84700 60738
rect 84672 48346 84700 60710
rect 84568 48340 84620 48346
rect 84568 48282 84620 48288
rect 84660 48340 84712 48346
rect 84660 48282 84712 48288
rect 84580 41426 84608 48282
rect 84580 41398 84700 41426
rect 84672 29102 84700 41398
rect 84660 29096 84712 29102
rect 84660 29038 84712 29044
rect 84568 29028 84620 29034
rect 84568 28970 84620 28976
rect 84580 22114 84608 28970
rect 84580 22086 84700 22114
rect 84672 12458 84700 22086
rect 84488 12430 84700 12458
rect 84384 4072 84436 4078
rect 84290 4040 84346 4049
rect 84384 4014 84436 4020
rect 84290 3975 84346 3984
rect 84488 3330 84516 12430
rect 84856 4146 84884 317784
rect 84936 317766 84988 317772
rect 85132 309194 85160 320062
rect 85868 318714 85896 320076
rect 85856 318708 85908 318714
rect 85856 318650 85908 318656
rect 86236 318102 86264 320076
rect 86420 320062 86710 320090
rect 86224 318096 86276 318102
rect 86224 318038 86276 318044
rect 86420 316010 86448 320062
rect 87064 318782 87092 320076
rect 87052 318776 87104 318782
rect 87052 318718 87104 318724
rect 87524 317966 87552 320076
rect 87708 320062 87906 320090
rect 87512 317960 87564 317966
rect 87512 317902 87564 317908
rect 87708 316010 87736 320062
rect 88248 318164 88300 318170
rect 88248 318106 88300 318112
rect 85684 315982 86448 316010
rect 87064 315982 87736 316010
rect 85120 309188 85172 309194
rect 85120 309130 85172 309136
rect 85684 5098 85712 315982
rect 87064 5166 87092 315982
rect 87052 5160 87104 5166
rect 87052 5102 87104 5108
rect 85672 5092 85724 5098
rect 85672 5034 85724 5040
rect 88260 4146 88288 318106
rect 88352 317490 88380 320076
rect 88536 320062 88734 320090
rect 88904 320062 89194 320090
rect 88340 317484 88392 317490
rect 88340 317426 88392 317432
rect 88432 315988 88484 315994
rect 88432 315930 88484 315936
rect 88444 5234 88472 315930
rect 88432 5228 88484 5234
rect 88432 5170 88484 5176
rect 84844 4140 84896 4146
rect 84844 4082 84896 4088
rect 87328 4140 87380 4146
rect 87328 4082 87380 4088
rect 88248 4140 88300 4146
rect 88248 4082 88300 4088
rect 86132 4072 86184 4078
rect 86132 4014 86184 4020
rect 84476 3324 84528 3330
rect 84476 3266 84528 3272
rect 84936 3324 84988 3330
rect 84936 3266 84988 3272
rect 83004 3256 83056 3262
rect 83004 3198 83056 3204
rect 83832 3256 83884 3262
rect 83832 3198 83884 3204
rect 83844 480 83872 3198
rect 84948 480 84976 3266
rect 86144 480 86172 4014
rect 87340 480 87368 4082
rect 88536 3482 88564 320062
rect 88904 315994 88932 320062
rect 88984 318436 89036 318442
rect 88984 318378 89036 318384
rect 88892 315988 88944 315994
rect 88892 315930 88944 315936
rect 88996 4010 89024 318378
rect 89076 318300 89128 318306
rect 89076 318242 89128 318248
rect 89088 4078 89116 318242
rect 89548 317898 89576 320076
rect 89536 317892 89588 317898
rect 89536 317834 89588 317840
rect 90008 317762 90036 320076
rect 90100 320062 90390 320090
rect 89996 317756 90048 317762
rect 89996 317698 90048 317704
rect 90100 316010 90128 320062
rect 89824 315982 90128 316010
rect 89824 5302 89852 315982
rect 90468 307873 90496 320198
rect 91218 320062 91324 320090
rect 91008 318640 91060 318646
rect 91008 318582 91060 318588
rect 90454 307864 90510 307873
rect 90454 307799 90510 307808
rect 90178 307728 90234 307737
rect 90178 307663 90234 307672
rect 90192 298246 90220 307663
rect 89996 298240 90048 298246
rect 89996 298182 90048 298188
rect 90180 298240 90232 298246
rect 90180 298182 90232 298188
rect 90008 296721 90036 298182
rect 89994 296712 90050 296721
rect 89994 296647 90050 296656
rect 90270 296712 90326 296721
rect 90270 296647 90326 296656
rect 90284 287094 90312 296647
rect 90088 287088 90140 287094
rect 90088 287030 90140 287036
rect 90272 287088 90324 287094
rect 90272 287030 90324 287036
rect 90100 273358 90128 287030
rect 90088 273352 90140 273358
rect 90088 273294 90140 273300
rect 89996 267776 90048 267782
rect 89996 267718 90048 267724
rect 90008 265690 90036 267718
rect 90008 265662 90128 265690
rect 90100 260846 90128 265662
rect 89996 260840 90048 260846
rect 89996 260782 90048 260788
rect 90088 260840 90140 260846
rect 90088 260782 90140 260788
rect 90008 253978 90036 260782
rect 89996 253972 90048 253978
rect 89996 253914 90048 253920
rect 90088 253836 90140 253842
rect 90088 253778 90140 253784
rect 90100 241482 90128 253778
rect 90008 241454 90128 241482
rect 90008 240145 90036 241454
rect 89994 240136 90050 240145
rect 89994 240071 90050 240080
rect 90178 240136 90234 240145
rect 91020 240122 91048 318582
rect 90178 240071 90234 240080
rect 90928 240094 91048 240122
rect 90192 230518 90220 240071
rect 90928 230518 90956 240094
rect 89996 230512 90048 230518
rect 89996 230454 90048 230460
rect 90180 230512 90232 230518
rect 90824 230512 90876 230518
rect 90180 230454 90232 230460
rect 90638 230480 90694 230489
rect 90008 227066 90036 230454
rect 90638 230415 90694 230424
rect 90822 230480 90824 230489
rect 90916 230512 90968 230518
rect 90876 230480 90878 230489
rect 90916 230454 90968 230460
rect 90822 230415 90878 230424
rect 90008 227038 90220 227066
rect 90192 224890 90220 227038
rect 90100 224862 90220 224890
rect 90100 217410 90128 224862
rect 90652 220862 90680 230415
rect 90640 220856 90692 220862
rect 90640 220798 90692 220804
rect 91008 220856 91060 220862
rect 91008 220798 91060 220804
rect 91020 220726 91048 220798
rect 91008 220720 91060 220726
rect 91008 220662 91060 220668
rect 90008 217382 90128 217410
rect 90008 205698 90036 217382
rect 91100 212492 91152 212498
rect 91100 212434 91152 212440
rect 91112 211154 91140 212434
rect 91112 211138 91232 211154
rect 91112 211132 91244 211138
rect 91112 211126 91192 211132
rect 91192 211074 91244 211080
rect 91204 211043 91232 211074
rect 89996 205692 90048 205698
rect 89996 205634 90048 205640
rect 90088 205556 90140 205562
rect 90088 205498 90140 205504
rect 90100 198098 90128 205498
rect 91008 202836 91060 202842
rect 91008 202778 91060 202784
rect 90008 198070 90128 198098
rect 90008 193225 90036 198070
rect 89994 193216 90050 193225
rect 89994 193151 90050 193160
rect 90178 193216 90234 193225
rect 90178 193151 90234 193160
rect 90192 174010 90220 193151
rect 91020 183598 91048 202778
rect 91008 183592 91060 183598
rect 91008 183534 91060 183540
rect 91008 180872 91060 180878
rect 91008 180814 91060 180820
rect 91020 178702 91048 180814
rect 91008 178696 91060 178702
rect 91008 178638 91060 178644
rect 89996 174004 90048 174010
rect 89996 173946 90048 173952
rect 90180 174004 90232 174010
rect 90180 173946 90232 173952
rect 90008 157486 90036 173946
rect 91192 171148 91244 171154
rect 91192 171090 91244 171096
rect 91204 162897 91232 171090
rect 91190 162888 91246 162897
rect 91190 162823 91246 162832
rect 91098 162616 91154 162625
rect 91098 162551 91154 162560
rect 89996 157480 90048 157486
rect 89996 157422 90048 157428
rect 89996 157344 90048 157350
rect 89996 157286 90048 157292
rect 90008 135425 90036 157286
rect 91112 153241 91140 162551
rect 91098 153232 91154 153241
rect 91098 153167 91154 153176
rect 91190 153096 91246 153105
rect 91190 153031 91246 153040
rect 89994 135416 90050 135425
rect 89994 135351 90050 135360
rect 89994 135280 90050 135289
rect 89994 135215 90050 135224
rect 90008 125610 90036 135215
rect 91204 133958 91232 153031
rect 91008 133952 91060 133958
rect 91008 133894 91060 133900
rect 91192 133952 91244 133958
rect 91192 133894 91244 133900
rect 90008 125594 90128 125610
rect 90008 125588 90140 125594
rect 90008 125582 90088 125588
rect 90088 125530 90140 125536
rect 90180 125588 90232 125594
rect 90180 125530 90232 125536
rect 90192 115977 90220 125530
rect 91020 124166 91048 133894
rect 91008 124160 91060 124166
rect 91008 124102 91060 124108
rect 91192 124160 91244 124166
rect 91192 124102 91244 124108
rect 89994 115968 90050 115977
rect 89994 115903 89996 115912
rect 90048 115903 90050 115912
rect 90178 115968 90234 115977
rect 90178 115903 90180 115912
rect 89996 115874 90048 115880
rect 90232 115903 90234 115912
rect 90180 115874 90232 115880
rect 90192 96665 90220 115874
rect 91204 114617 91232 124102
rect 91006 114608 91062 114617
rect 90928 114566 91006 114594
rect 90928 114510 90956 114566
rect 91006 114543 91062 114552
rect 91190 114608 91246 114617
rect 91190 114543 91246 114552
rect 90916 114504 90968 114510
rect 90916 114446 90968 114452
rect 91008 104916 91060 104922
rect 91008 104858 91060 104864
rect 91020 104802 91048 104858
rect 91020 104774 91140 104802
rect 89994 96656 90050 96665
rect 89994 96591 90050 96600
rect 90178 96656 90234 96665
rect 90178 96591 90234 96600
rect 90008 86902 90036 96591
rect 91112 95266 91140 104774
rect 91008 95260 91060 95266
rect 91008 95202 91060 95208
rect 91100 95260 91152 95266
rect 91100 95202 91152 95208
rect 89996 86896 90048 86902
rect 89996 86838 90048 86844
rect 91020 85513 91048 95202
rect 91006 85504 91062 85513
rect 91006 85439 91062 85448
rect 91098 85368 91154 85377
rect 91098 85303 91154 85312
rect 89996 77308 90048 77314
rect 89996 77250 90048 77256
rect 90008 67590 90036 77250
rect 89996 67584 90048 67590
rect 89996 67526 90048 67532
rect 91112 66366 91140 85303
rect 91100 66360 91152 66366
rect 91100 66302 91152 66308
rect 91008 66292 91060 66298
rect 91008 66234 91060 66240
rect 89996 58064 90048 58070
rect 89996 58006 90048 58012
rect 90008 41342 90036 58006
rect 91020 56710 91048 66234
rect 91008 56704 91060 56710
rect 91008 56646 91060 56652
rect 90916 55276 90968 55282
rect 90916 55218 90968 55224
rect 90928 46986 90956 55218
rect 90916 46980 90968 46986
rect 90916 46922 90968 46928
rect 91008 46980 91060 46986
rect 91008 46922 91060 46928
rect 91020 46850 91048 46922
rect 91008 46844 91060 46850
rect 91008 46786 91060 46792
rect 91192 46844 91244 46850
rect 91192 46786 91244 46792
rect 89996 41336 90048 41342
rect 89996 41278 90048 41284
rect 89996 41200 90048 41206
rect 89996 41142 90048 41148
rect 90008 28966 90036 41142
rect 91204 29034 91232 46786
rect 91008 29028 91060 29034
rect 91008 28970 91060 28976
rect 91192 29028 91244 29034
rect 91192 28970 91244 28976
rect 89996 28960 90048 28966
rect 89996 28902 90048 28908
rect 91020 27606 91048 28970
rect 91008 27600 91060 27606
rect 91008 27542 91060 27548
rect 89996 19372 90048 19378
rect 89996 19314 90048 19320
rect 89812 5296 89864 5302
rect 89812 5238 89864 5244
rect 89720 4140 89772 4146
rect 89720 4082 89772 4088
rect 89076 4072 89128 4078
rect 89076 4014 89128 4020
rect 88984 4004 89036 4010
rect 88984 3946 89036 3952
rect 88444 3454 88564 3482
rect 88444 3398 88472 3454
rect 88432 3392 88484 3398
rect 88432 3334 88484 3340
rect 88524 3392 88576 3398
rect 88524 3334 88576 3340
rect 88536 480 88564 3334
rect 89732 480 89760 4082
rect 90008 3058 90036 19314
rect 91008 18012 91060 18018
rect 91008 17954 91060 17960
rect 91020 12510 91048 17954
rect 91008 12504 91060 12510
rect 91008 12446 91060 12452
rect 90916 12436 90968 12442
rect 90916 12378 90968 12384
rect 90928 9654 90956 12378
rect 90916 9648 90968 9654
rect 90916 9590 90968 9596
rect 90916 9512 90968 9518
rect 90916 9454 90968 9460
rect 89996 3052 90048 3058
rect 89996 2994 90048 3000
rect 90928 480 90956 9454
rect 91296 3126 91324 320062
rect 91664 317694 91692 320076
rect 91744 318368 91796 318374
rect 91744 318310 91796 318316
rect 91652 317688 91704 317694
rect 91652 317630 91704 317636
rect 91756 4146 91784 318310
rect 92032 317558 92060 320076
rect 92492 317626 92520 320076
rect 92860 318034 92888 320076
rect 93044 320062 93242 320090
rect 93320 320062 93702 320090
rect 92848 318028 92900 318034
rect 92848 317970 92900 317976
rect 92480 317620 92532 317626
rect 92480 317562 92532 317568
rect 92020 317552 92072 317558
rect 92020 317494 92072 317500
rect 93044 317422 93072 320062
rect 93124 318572 93176 318578
rect 93124 318514 93176 318520
rect 93032 317416 93084 317422
rect 93032 317358 93084 317364
rect 92572 315988 92624 315994
rect 92572 315930 92624 315936
rect 91744 4140 91796 4146
rect 91744 4082 91796 4088
rect 92112 3732 92164 3738
rect 92112 3674 92164 3680
rect 91284 3120 91336 3126
rect 91284 3062 91336 3068
rect 92124 480 92152 3674
rect 92584 2854 92612 315930
rect 92848 307828 92900 307834
rect 92848 307770 92900 307776
rect 92860 299606 92888 307770
rect 92848 299600 92900 299606
rect 92848 299542 92900 299548
rect 92848 299464 92900 299470
rect 92848 299406 92900 299412
rect 92860 269142 92888 299406
rect 92756 269136 92808 269142
rect 92756 269078 92808 269084
rect 92848 269136 92900 269142
rect 92848 269078 92900 269084
rect 92768 260914 92796 269078
rect 92756 260908 92808 260914
rect 92756 260850 92808 260856
rect 92848 260772 92900 260778
rect 92848 260714 92900 260720
rect 92860 259434 92888 260714
rect 92676 259406 92888 259434
rect 92676 249830 92704 259406
rect 92664 249824 92716 249830
rect 92664 249766 92716 249772
rect 92848 249824 92900 249830
rect 92848 249766 92900 249772
rect 92860 236722 92888 249766
rect 92768 236694 92888 236722
rect 92768 227066 92796 236694
rect 92768 227038 92980 227066
rect 92952 224890 92980 227038
rect 92860 224862 92980 224890
rect 92860 217410 92888 224862
rect 92768 217382 92888 217410
rect 92768 212537 92796 217382
rect 92754 212528 92810 212537
rect 92754 212463 92810 212472
rect 92938 212528 92994 212537
rect 92938 212463 92994 212472
rect 92952 193322 92980 212463
rect 92756 193316 92808 193322
rect 92756 193258 92808 193264
rect 92940 193316 92992 193322
rect 92940 193258 92992 193264
rect 92768 157434 92796 193258
rect 92768 157406 92888 157434
rect 92860 157332 92888 157406
rect 92768 157304 92888 157332
rect 92768 135425 92796 157304
rect 92754 135416 92810 135425
rect 92754 135351 92810 135360
rect 92754 135280 92810 135289
rect 92754 135215 92810 135224
rect 92768 125610 92796 135215
rect 92768 125594 92888 125610
rect 92768 125588 92900 125594
rect 92768 125582 92848 125588
rect 92848 125530 92900 125536
rect 92940 125588 92992 125594
rect 92940 125530 92992 125536
rect 92952 115977 92980 125530
rect 92754 115968 92810 115977
rect 92754 115903 92756 115912
rect 92808 115903 92810 115912
rect 92938 115968 92994 115977
rect 92938 115903 92940 115912
rect 92756 115874 92808 115880
rect 92992 115903 92994 115912
rect 92940 115874 92992 115880
rect 92952 96665 92980 115874
rect 92754 96656 92810 96665
rect 92754 96591 92810 96600
rect 92938 96656 92994 96665
rect 92938 96591 92994 96600
rect 92768 86902 92796 96591
rect 92756 86896 92808 86902
rect 92756 86838 92808 86844
rect 92756 77308 92808 77314
rect 92756 77250 92808 77256
rect 92768 67590 92796 77250
rect 92756 67584 92808 67590
rect 92756 67526 92808 67532
rect 92756 58064 92808 58070
rect 92756 58006 92808 58012
rect 92768 48346 92796 58006
rect 92756 48340 92808 48346
rect 92756 48282 92808 48288
rect 92848 48204 92900 48210
rect 92848 48146 92900 48152
rect 92860 27742 92888 48146
rect 92848 27736 92900 27742
rect 92848 27678 92900 27684
rect 92756 27668 92808 27674
rect 92756 27610 92808 27616
rect 92768 2990 92796 27610
rect 93136 3330 93164 318514
rect 93320 315994 93348 320062
rect 93768 318504 93820 318510
rect 93768 318446 93820 318452
rect 93308 315988 93360 315994
rect 93308 315930 93360 315936
rect 93780 4146 93808 318446
rect 94056 317422 94084 320076
rect 94240 320062 94530 320090
rect 94608 320062 94898 320090
rect 94044 317416 94096 317422
rect 94044 317358 94096 317364
rect 93952 316056 94004 316062
rect 93952 315998 94004 316004
rect 93860 315988 93912 315994
rect 93860 315930 93912 315936
rect 93872 77246 93900 315930
rect 93964 77246 93992 315998
rect 94240 315994 94268 320062
rect 94608 316062 94636 320062
rect 95240 316124 95292 316130
rect 95240 316066 95292 316072
rect 94596 316056 94648 316062
rect 94596 315998 94648 316004
rect 94228 315988 94280 315994
rect 94228 315930 94280 315936
rect 94044 307896 94096 307902
rect 94044 307838 94096 307844
rect 94056 307766 94084 307838
rect 94044 307760 94096 307766
rect 94044 307702 94096 307708
rect 94044 298172 94096 298178
rect 94044 298114 94096 298120
rect 94056 288454 94084 298114
rect 94044 288448 94096 288454
rect 94044 288390 94096 288396
rect 94136 288448 94188 288454
rect 94136 288390 94188 288396
rect 94148 287065 94176 288390
rect 94134 287056 94190 287065
rect 94134 286991 94190 287000
rect 94318 287056 94374 287065
rect 94318 286991 94374 287000
rect 94332 277438 94360 286991
rect 94136 277432 94188 277438
rect 94136 277374 94188 277380
rect 94320 277432 94372 277438
rect 94320 277374 94372 277380
rect 94148 265690 94176 277374
rect 94056 265662 94176 265690
rect 94056 251258 94084 265662
rect 94044 251252 94096 251258
rect 94044 251194 94096 251200
rect 94136 251252 94188 251258
rect 94136 251194 94188 251200
rect 94148 245002 94176 251194
rect 94136 244996 94188 245002
rect 94136 244938 94188 244944
rect 94136 231872 94188 231878
rect 94136 231814 94188 231820
rect 94148 225078 94176 231814
rect 94136 225072 94188 225078
rect 94136 225014 94188 225020
rect 94044 224936 94096 224942
rect 94044 224878 94096 224884
rect 94056 222193 94084 224878
rect 94042 222184 94098 222193
rect 94042 222119 94098 222128
rect 94318 222184 94374 222193
rect 94318 222119 94374 222128
rect 94332 212566 94360 222119
rect 94136 212560 94188 212566
rect 94136 212502 94188 212508
rect 94320 212560 94372 212566
rect 94320 212502 94372 212508
rect 94148 205766 94176 212502
rect 94136 205760 94188 205766
rect 94136 205702 94188 205708
rect 94044 205624 94096 205630
rect 94044 205566 94096 205572
rect 94056 202842 94084 205566
rect 94044 202836 94096 202842
rect 94044 202778 94096 202784
rect 94136 193248 94188 193254
rect 94136 193190 94188 193196
rect 94148 188442 94176 193190
rect 94148 188414 94268 188442
rect 94240 173942 94268 188414
rect 94136 173936 94188 173942
rect 94136 173878 94188 173884
rect 94228 173936 94280 173942
rect 94228 173878 94280 173884
rect 94148 172514 94176 173878
rect 94136 172508 94188 172514
rect 94136 172450 94188 172456
rect 94320 172508 94372 172514
rect 94320 172450 94372 172456
rect 94332 162897 94360 172450
rect 94134 162888 94190 162897
rect 94134 162823 94190 162832
rect 94318 162888 94374 162897
rect 94318 162823 94374 162832
rect 94148 156670 94176 162823
rect 94136 156664 94188 156670
rect 94136 156606 94188 156612
rect 94320 147008 94372 147014
rect 94320 146950 94372 146956
rect 94332 133929 94360 146950
rect 94134 133920 94190 133929
rect 94134 133855 94190 133864
rect 94318 133920 94374 133929
rect 94318 133855 94374 133864
rect 94148 125610 94176 133855
rect 94056 125582 94176 125610
rect 94056 118454 94084 125582
rect 94044 118448 94096 118454
rect 94044 118390 94096 118396
rect 94136 118380 94188 118386
rect 94136 118322 94188 118328
rect 94148 106593 94176 118322
rect 94134 106584 94190 106593
rect 94134 106519 94190 106528
rect 94042 106312 94098 106321
rect 94042 106247 94098 106256
rect 94056 104854 94084 106247
rect 94044 104848 94096 104854
rect 94044 104790 94096 104796
rect 94044 95260 94096 95266
rect 94044 95202 94096 95208
rect 94056 87145 94084 95202
rect 94042 87136 94098 87145
rect 94042 87071 94098 87080
rect 94042 87000 94098 87009
rect 94042 86935 94098 86944
rect 94056 85542 94084 86935
rect 94044 85536 94096 85542
rect 94044 85478 94096 85484
rect 94320 80980 94372 80986
rect 94320 80922 94372 80928
rect 93860 77240 93912 77246
rect 93860 77182 93912 77188
rect 93952 77240 94004 77246
rect 93952 77182 94004 77188
rect 93952 77104 94004 77110
rect 93952 77046 94004 77052
rect 93860 77036 93912 77042
rect 93860 76978 93912 76984
rect 93308 4140 93360 4146
rect 93308 4082 93360 4088
rect 93768 4140 93820 4146
rect 93768 4082 93820 4088
rect 93124 3324 93176 3330
rect 93124 3266 93176 3272
rect 92756 2984 92808 2990
rect 92756 2926 92808 2932
rect 92572 2848 92624 2854
rect 92572 2790 92624 2796
rect 93320 480 93348 4082
rect 93872 3466 93900 76978
rect 93964 3806 93992 77046
rect 94332 74526 94360 80922
rect 94320 74520 94372 74526
rect 94320 74462 94372 74468
rect 94136 64932 94188 64938
rect 94136 64874 94188 64880
rect 94148 60042 94176 64874
rect 94136 60036 94188 60042
rect 94136 59978 94188 59984
rect 94136 50652 94188 50658
rect 94136 50594 94188 50600
rect 94148 31822 94176 50594
rect 94136 31816 94188 31822
rect 94136 31758 94188 31764
rect 94136 31612 94188 31618
rect 94136 31554 94188 31560
rect 94148 22114 94176 31554
rect 94056 22086 94176 22114
rect 94056 19394 94084 22086
rect 94056 19366 94176 19394
rect 94148 12510 94176 19366
rect 94136 12504 94188 12510
rect 94136 12446 94188 12452
rect 94228 12368 94280 12374
rect 94228 12310 94280 12316
rect 94240 9654 94268 12310
rect 94228 9648 94280 9654
rect 94228 9590 94280 9596
rect 94504 4140 94556 4146
rect 94504 4082 94556 4088
rect 93952 3800 94004 3806
rect 93952 3742 94004 3748
rect 93860 3460 93912 3466
rect 93860 3402 93912 3408
rect 94516 480 94544 4082
rect 95252 3670 95280 316066
rect 95240 3664 95292 3670
rect 95240 3606 95292 3612
rect 95344 3534 95372 320076
rect 95436 320062 95726 320090
rect 95896 320062 96186 320090
rect 96264 320062 96554 320090
rect 96724 320062 97014 320090
rect 97184 320062 97382 320090
rect 97552 320062 97842 320090
rect 95436 3602 95464 320062
rect 95896 316130 95924 320062
rect 95884 316124 95936 316130
rect 95884 316066 95936 316072
rect 96264 316010 96292 320062
rect 96528 317892 96580 317898
rect 96528 317834 96580 317840
rect 96344 317824 96396 317830
rect 96344 317766 96396 317772
rect 95620 315982 96292 316010
rect 95620 302274 95648 315982
rect 96356 314786 96384 317766
rect 95528 302246 95648 302274
rect 95896 314758 96384 314786
rect 95528 302138 95556 302246
rect 95528 302110 95740 302138
rect 95712 273306 95740 302110
rect 95528 273278 95740 273306
rect 95528 273170 95556 273278
rect 95528 273142 95648 273170
rect 95620 241482 95648 273142
rect 95620 241454 95740 241482
rect 95712 234666 95740 241454
rect 95700 234660 95752 234666
rect 95700 234602 95752 234608
rect 95608 234592 95660 234598
rect 95608 234534 95660 234540
rect 95620 222170 95648 234534
rect 95620 222142 95740 222170
rect 95712 215354 95740 222142
rect 95700 215348 95752 215354
rect 95700 215290 95752 215296
rect 95608 215280 95660 215286
rect 95608 215222 95660 215228
rect 95620 202858 95648 215222
rect 95620 202830 95740 202858
rect 95712 196042 95740 202830
rect 95700 196036 95752 196042
rect 95700 195978 95752 195984
rect 95608 195968 95660 195974
rect 95608 195910 95660 195916
rect 95620 183546 95648 195910
rect 95528 183518 95648 183546
rect 95528 176730 95556 183518
rect 95516 176724 95568 176730
rect 95516 176666 95568 176672
rect 95608 176656 95660 176662
rect 95608 176598 95660 176604
rect 95620 157434 95648 176598
rect 95528 157406 95648 157434
rect 95528 157298 95556 157406
rect 95528 157270 95648 157298
rect 95620 138122 95648 157270
rect 95528 138094 95648 138122
rect 95528 137850 95556 138094
rect 95528 137822 95648 137850
rect 95620 118794 95648 137822
rect 95608 118788 95660 118794
rect 95608 118730 95660 118736
rect 95608 118652 95660 118658
rect 95608 118594 95660 118600
rect 95620 62914 95648 118594
rect 95528 62886 95648 62914
rect 95528 62642 95556 62886
rect 95528 62614 95648 62642
rect 95620 41426 95648 62614
rect 95528 41398 95648 41426
rect 95528 41290 95556 41398
rect 95528 41262 95648 41290
rect 95620 21978 95648 41262
rect 95620 21950 95740 21978
rect 95712 3874 95740 21950
rect 95896 4146 95924 314758
rect 95884 4140 95936 4146
rect 95884 4082 95936 4088
rect 95700 3868 95752 3874
rect 95700 3810 95752 3816
rect 95424 3596 95476 3602
rect 95424 3538 95476 3544
rect 95332 3528 95384 3534
rect 95332 3470 95384 3476
rect 96540 3466 96568 317834
rect 96620 315988 96672 315994
rect 96620 315930 96672 315936
rect 96632 4010 96660 315930
rect 96724 4078 96752 320062
rect 97184 316010 97212 320062
rect 97264 318164 97316 318170
rect 97264 318106 97316 318112
rect 97000 315982 97212 316010
rect 97000 302410 97028 315982
rect 96908 302382 97028 302410
rect 96908 302274 96936 302382
rect 96816 302246 96936 302274
rect 96816 302138 96844 302246
rect 96816 302110 97028 302138
rect 97000 273306 97028 302110
rect 96816 273278 97028 273306
rect 96816 273170 96844 273278
rect 96816 273142 97028 273170
rect 97000 253994 97028 273142
rect 96816 253966 97028 253994
rect 96816 253858 96844 253966
rect 96816 253830 97028 253858
rect 97000 234682 97028 253830
rect 96816 234654 97028 234682
rect 96816 234546 96844 234654
rect 96816 234518 97028 234546
rect 97000 215370 97028 234518
rect 96816 215342 97028 215370
rect 96816 215234 96844 215342
rect 96816 215206 97028 215234
rect 97000 196058 97028 215206
rect 96816 196030 97028 196058
rect 96816 195922 96844 196030
rect 96816 195894 97028 195922
rect 97000 176746 97028 195894
rect 96816 176718 97028 176746
rect 96816 176610 96844 176718
rect 96816 176582 97028 176610
rect 97000 157434 97028 176582
rect 96816 157406 97028 157434
rect 96816 157298 96844 157406
rect 96816 157270 96936 157298
rect 96908 157162 96936 157270
rect 96908 157134 97028 157162
rect 97000 60761 97028 157134
rect 96986 60752 97042 60761
rect 96986 60687 97042 60696
rect 96986 56672 97042 56681
rect 96986 56607 97042 56616
rect 97000 56574 97028 56607
rect 96988 56568 97040 56574
rect 96988 56510 97040 56516
rect 96988 47048 97040 47054
rect 96988 46990 97040 46996
rect 97000 46918 97028 46990
rect 96988 46912 97040 46918
rect 96988 46854 97040 46860
rect 96988 37324 97040 37330
rect 96988 37266 97040 37272
rect 97000 28966 97028 37266
rect 96988 28960 97040 28966
rect 96988 28902 97040 28908
rect 96988 21956 97040 21962
rect 96988 21898 97040 21904
rect 96896 4140 96948 4146
rect 96896 4082 96948 4088
rect 96712 4072 96764 4078
rect 96712 4014 96764 4020
rect 96620 4004 96672 4010
rect 96620 3946 96672 3952
rect 95700 3460 95752 3466
rect 95700 3402 95752 3408
rect 96528 3460 96580 3466
rect 96528 3402 96580 3408
rect 95712 480 95740 3402
rect 96908 480 96936 4082
rect 97000 3942 97028 21898
rect 96988 3936 97040 3942
rect 96988 3878 97040 3884
rect 97276 3262 97304 318106
rect 97552 315994 97580 320062
rect 98196 318442 98224 320076
rect 98184 318436 98236 318442
rect 98184 318378 98236 318384
rect 98656 317762 98684 320076
rect 98840 320062 99038 320090
rect 98644 317756 98696 317762
rect 98644 317698 98696 317704
rect 97908 317688 97960 317694
rect 97908 317630 97960 317636
rect 97540 315988 97592 315994
rect 97540 315930 97592 315936
rect 97920 4146 97948 317630
rect 98840 316010 98868 320062
rect 99484 318578 99512 320076
rect 99472 318572 99524 318578
rect 99472 318514 99524 318520
rect 99852 318306 99880 320076
rect 99840 318300 99892 318306
rect 99840 318242 99892 318248
rect 100312 318238 100340 320076
rect 100300 318232 100352 318238
rect 100300 318174 100352 318180
rect 100680 318170 100708 320076
rect 101140 318374 101168 320076
rect 101508 318646 101536 320076
rect 101496 318640 101548 318646
rect 101496 318582 101548 318588
rect 101128 318368 101180 318374
rect 101128 318310 101180 318316
rect 100668 318164 100720 318170
rect 100668 318106 100720 318112
rect 100024 317620 100076 317626
rect 100024 317562 100076 317568
rect 98104 315982 98868 316010
rect 97908 4140 97960 4146
rect 97908 4082 97960 4088
rect 98104 3890 98132 315982
rect 98104 3862 98316 3890
rect 98092 3664 98144 3670
rect 98092 3606 98144 3612
rect 97264 3256 97316 3262
rect 97264 3198 97316 3204
rect 98104 480 98132 3606
rect 98288 3398 98316 3862
rect 100036 3534 100064 317562
rect 101968 317490 101996 320076
rect 102336 318510 102364 320076
rect 102324 318504 102376 318510
rect 102324 318446 102376 318452
rect 102796 317830 102824 320076
rect 103164 317898 103192 320076
rect 103152 317892 103204 317898
rect 103152 317834 103204 317840
rect 102784 317824 102836 317830
rect 102784 317766 102836 317772
rect 103624 317694 103652 320076
rect 103612 317688 103664 317694
rect 103612 317630 103664 317636
rect 103428 317552 103480 317558
rect 103428 317494 103480 317500
rect 100116 317484 100168 317490
rect 100116 317426 100168 317432
rect 101956 317484 102008 317490
rect 101956 317426 102008 317432
rect 102784 317484 102836 317490
rect 102784 317426 102836 317432
rect 100128 3738 100156 317426
rect 102796 4298 102824 317426
rect 102612 4270 102824 4298
rect 101588 4072 101640 4078
rect 101588 4014 101640 4020
rect 100484 3936 100536 3942
rect 100484 3878 100536 3884
rect 100116 3732 100168 3738
rect 100116 3674 100168 3680
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 100024 3528 100076 3534
rect 100024 3470 100076 3476
rect 98276 3392 98328 3398
rect 98276 3334 98328 3340
rect 99300 480 99328 3470
rect 100496 480 100524 3878
rect 101600 480 101628 4014
rect 102612 3670 102640 4270
rect 103440 4146 103468 317494
rect 103992 317490 104020 320076
rect 104360 317626 104388 320076
rect 104348 317620 104400 317626
rect 104348 317562 104400 317568
rect 103980 317484 104032 317490
rect 103980 317426 104032 317432
rect 104452 316010 104480 320198
rect 105004 319410 105032 320198
rect 105004 319382 105124 319410
rect 104808 317484 104860 317490
rect 104808 317426 104860 317432
rect 103716 315982 104480 316010
rect 102784 4140 102836 4146
rect 102784 4082 102836 4088
rect 103428 4140 103480 4146
rect 103428 4082 103480 4088
rect 102600 3664 102652 3670
rect 102600 3606 102652 3612
rect 102796 480 102824 4082
rect 103716 3942 103744 315982
rect 103704 3936 103756 3942
rect 103704 3878 103756 3884
rect 104820 3534 104848 317426
rect 105096 311982 105124 319382
rect 105648 317558 105676 320076
rect 105636 317552 105688 317558
rect 105636 317494 105688 317500
rect 106016 317490 106044 320076
rect 106292 320062 106490 320090
rect 106660 320062 106858 320090
rect 107028 320062 107318 320090
rect 107686 320062 107884 320090
rect 106004 317484 106056 317490
rect 106004 317426 106056 317432
rect 105084 311976 105136 311982
rect 105084 311918 105136 311924
rect 105176 311772 105228 311778
rect 105176 311714 105228 311720
rect 105188 302258 105216 311714
rect 105176 302252 105228 302258
rect 105176 302194 105228 302200
rect 105084 298172 105136 298178
rect 105084 298114 105136 298120
rect 105096 298058 105124 298114
rect 105174 298072 105230 298081
rect 105096 298030 105174 298058
rect 105174 298007 105230 298016
rect 105358 298072 105414 298081
rect 105358 298007 105414 298016
rect 105372 292466 105400 298007
rect 105176 292460 105228 292466
rect 105176 292402 105228 292408
rect 105360 292460 105412 292466
rect 105360 292402 105412 292408
rect 105188 283014 105216 292402
rect 105176 283008 105228 283014
rect 105176 282950 105228 282956
rect 105176 282804 105228 282810
rect 105176 282746 105228 282752
rect 105188 280158 105216 282746
rect 105176 280152 105228 280158
rect 105176 280094 105228 280100
rect 105176 273148 105228 273154
rect 105176 273090 105228 273096
rect 105188 270502 105216 273090
rect 105176 270496 105228 270502
rect 105176 270438 105228 270444
rect 105176 263492 105228 263498
rect 105176 263434 105228 263440
rect 105188 260846 105216 263434
rect 105176 260840 105228 260846
rect 105176 260782 105228 260788
rect 105176 253836 105228 253842
rect 105176 253778 105228 253784
rect 105188 251190 105216 253778
rect 105176 251184 105228 251190
rect 105176 251126 105228 251132
rect 105084 241528 105136 241534
rect 105084 241470 105136 241476
rect 105096 234666 105124 241470
rect 105084 234660 105136 234666
rect 105084 234602 105136 234608
rect 105176 234524 105228 234530
rect 105176 234466 105228 234472
rect 105188 231826 105216 234466
rect 105096 231798 105216 231826
rect 105096 225010 105124 231798
rect 105084 225004 105136 225010
rect 105084 224946 105136 224952
rect 105084 222216 105136 222222
rect 105084 222158 105136 222164
rect 105096 215354 105124 222158
rect 105084 215348 105136 215354
rect 105084 215290 105136 215296
rect 105176 215212 105228 215218
rect 105176 215154 105228 215160
rect 105188 212514 105216 215154
rect 105096 212486 105216 212514
rect 105096 205698 105124 212486
rect 105084 205692 105136 205698
rect 105084 205634 105136 205640
rect 105084 202904 105136 202910
rect 105084 202846 105136 202852
rect 105096 196042 105124 202846
rect 105084 196036 105136 196042
rect 105084 195978 105136 195984
rect 105176 195900 105228 195906
rect 105176 195842 105228 195848
rect 105188 193202 105216 195842
rect 105096 193174 105216 193202
rect 105096 186386 105124 193174
rect 105084 186380 105136 186386
rect 105084 186322 105136 186328
rect 105084 183592 105136 183598
rect 105084 183534 105136 183540
rect 105096 176730 105124 183534
rect 105084 176724 105136 176730
rect 105084 176666 105136 176672
rect 105176 176588 105228 176594
rect 105176 176530 105228 176536
rect 105188 173890 105216 176530
rect 105096 173862 105216 173890
rect 105096 169114 105124 173862
rect 104900 169108 104952 169114
rect 104900 169050 104952 169056
rect 105084 169108 105136 169114
rect 105084 169050 105136 169056
rect 104912 164257 104940 169050
rect 104898 164248 104954 164257
rect 104898 164183 104954 164192
rect 105082 164248 105138 164257
rect 105082 164183 105138 164192
rect 105096 157418 105124 164183
rect 105084 157412 105136 157418
rect 105084 157354 105136 157360
rect 105176 157276 105228 157282
rect 105176 157218 105228 157224
rect 105188 147762 105216 157218
rect 105176 147756 105228 147762
rect 105176 147698 105228 147704
rect 105084 147620 105136 147626
rect 105084 147562 105136 147568
rect 105096 143546 105124 147562
rect 105084 143540 105136 143546
rect 105084 143482 105136 143488
rect 105084 137964 105136 137970
rect 105084 137906 105136 137912
rect 105096 133906 105124 137906
rect 105096 133878 105216 133906
rect 105188 128450 105216 133878
rect 105176 128444 105228 128450
rect 105176 128386 105228 128392
rect 105084 128308 105136 128314
rect 105084 128250 105136 128256
rect 105096 124166 105124 128250
rect 105084 124160 105136 124166
rect 105084 124102 105136 124108
rect 105176 114572 105228 114578
rect 105176 114514 105228 114520
rect 105188 109138 105216 114514
rect 105176 109132 105228 109138
rect 105176 109074 105228 109080
rect 105084 108996 105136 109002
rect 105084 108938 105136 108944
rect 105096 104854 105124 108938
rect 105084 104848 105136 104854
rect 105084 104790 105136 104796
rect 105176 95260 105228 95266
rect 105176 95202 105228 95208
rect 105188 89826 105216 95202
rect 105176 89820 105228 89826
rect 105176 89762 105228 89768
rect 105084 89684 105136 89690
rect 105084 89626 105136 89632
rect 105096 85542 105124 89626
rect 105084 85536 105136 85542
rect 105084 85478 105136 85484
rect 104992 84108 105044 84114
rect 104992 84050 105044 84056
rect 105004 74594 105032 84050
rect 104992 74588 105044 74594
rect 104992 74530 105044 74536
rect 104992 66292 105044 66298
rect 104992 66234 105044 66240
rect 105004 64870 105032 66234
rect 104992 64864 105044 64870
rect 104992 64806 105044 64812
rect 105268 64864 105320 64870
rect 105268 64806 105320 64812
rect 105280 46986 105308 64806
rect 104900 46980 104952 46986
rect 104900 46922 104952 46928
rect 105268 46980 105320 46986
rect 105268 46922 105320 46928
rect 104912 41342 104940 46922
rect 104900 41336 104952 41342
rect 104900 41278 104952 41284
rect 105176 41336 105228 41342
rect 105176 41278 105228 41284
rect 105188 31822 105216 41278
rect 105176 31816 105228 31822
rect 105176 31758 105228 31764
rect 105084 31748 105136 31754
rect 105084 31690 105136 31696
rect 105096 28914 105124 31690
rect 105096 28886 105216 28914
rect 105188 4298 105216 28886
rect 105004 4270 105216 4298
rect 105004 4078 105032 4270
rect 106292 4146 106320 320062
rect 106660 316010 106688 320062
rect 107028 316010 107056 320062
rect 106384 315982 106688 316010
rect 106752 315982 107056 316010
rect 105176 4140 105228 4146
rect 105176 4082 105228 4088
rect 106280 4140 106332 4146
rect 106280 4082 106332 4088
rect 104992 4072 105044 4078
rect 104992 4014 105044 4020
rect 103980 3528 104032 3534
rect 103980 3470 104032 3476
rect 104808 3528 104860 3534
rect 104808 3470 104860 3476
rect 103992 480 104020 3470
rect 105188 480 105216 4082
rect 106384 480 106412 315982
rect 106752 302258 106780 315982
rect 106556 302252 106608 302258
rect 106556 302194 106608 302200
rect 106740 302252 106792 302258
rect 106740 302194 106792 302200
rect 106568 302138 106596 302194
rect 106568 302110 106688 302138
rect 106660 292618 106688 302110
rect 106660 292590 106780 292618
rect 106752 282946 106780 292590
rect 106556 282940 106608 282946
rect 106556 282882 106608 282888
rect 106740 282940 106792 282946
rect 106740 282882 106792 282888
rect 106568 282826 106596 282882
rect 106568 282798 106688 282826
rect 106660 280158 106688 282798
rect 106648 280152 106700 280158
rect 106648 280094 106700 280100
rect 106832 273284 106884 273290
rect 106832 273226 106884 273232
rect 106844 270502 106872 273226
rect 106832 270496 106884 270502
rect 106832 270438 106884 270444
rect 106924 260908 106976 260914
rect 106924 260850 106976 260856
rect 106936 254046 106964 260850
rect 106924 254040 106976 254046
rect 106924 253982 106976 253988
rect 106832 253904 106884 253910
rect 106832 253846 106884 253852
rect 106844 244202 106872 253846
rect 106660 244174 106872 244202
rect 106660 241505 106688 244174
rect 106646 241496 106702 241505
rect 106646 241431 106702 241440
rect 106554 235376 106610 235385
rect 106554 235311 106610 235320
rect 106568 230450 106596 235311
rect 106556 230444 106608 230450
rect 106556 230386 106608 230392
rect 106464 220924 106516 220930
rect 106464 220866 106516 220872
rect 106476 220794 106504 220866
rect 106464 220788 106516 220794
rect 106464 220730 106516 220736
rect 106648 220788 106700 220794
rect 106648 220730 106700 220736
rect 106660 215234 106688 220730
rect 106568 215206 106688 215234
rect 106568 202910 106596 215206
rect 106556 202904 106608 202910
rect 106556 202846 106608 202852
rect 106740 202904 106792 202910
rect 106740 202846 106792 202852
rect 106752 196042 106780 202846
rect 106740 196036 106792 196042
rect 106740 195978 106792 195984
rect 106832 195968 106884 195974
rect 106832 195910 106884 195916
rect 106844 193225 106872 195910
rect 106646 193216 106702 193225
rect 106646 193151 106702 193160
rect 106830 193216 106886 193225
rect 106830 193151 106886 193160
rect 106660 183598 106688 193151
rect 106648 183592 106700 183598
rect 106648 183534 106700 183540
rect 106924 183592 106976 183598
rect 106924 183534 106976 183540
rect 106936 173942 106964 183534
rect 106740 173936 106792 173942
rect 106462 173904 106518 173913
rect 106462 173839 106518 173848
rect 106738 173904 106740 173913
rect 106924 173936 106976 173942
rect 106792 173904 106794 173913
rect 106924 173878 106976 173884
rect 106738 173839 106794 173848
rect 106476 164257 106504 173839
rect 106462 164248 106518 164257
rect 106462 164183 106518 164192
rect 106646 164248 106702 164257
rect 106646 164183 106648 164192
rect 106700 164183 106702 164192
rect 106648 164154 106700 164160
rect 106648 157344 106700 157350
rect 106648 157286 106700 157292
rect 106660 154578 106688 157286
rect 106660 154550 106780 154578
rect 106752 147694 106780 154550
rect 106556 147688 106608 147694
rect 106740 147688 106792 147694
rect 106608 147636 106688 147642
rect 106556 147630 106688 147636
rect 106740 147630 106792 147636
rect 106568 147614 106688 147630
rect 106660 144906 106688 147614
rect 106648 144900 106700 144906
rect 106648 144842 106700 144848
rect 106648 137964 106700 137970
rect 106648 137906 106700 137912
rect 106660 135266 106688 137906
rect 106660 135238 106780 135266
rect 106752 124234 106780 135238
rect 106464 124228 106516 124234
rect 106464 124170 106516 124176
rect 106740 124228 106792 124234
rect 106740 124170 106792 124176
rect 106476 124098 106504 124170
rect 106464 124092 106516 124098
rect 106464 124034 106516 124040
rect 106556 114640 106608 114646
rect 106556 114582 106608 114588
rect 106568 109138 106596 114582
rect 106556 109132 106608 109138
rect 106556 109074 106608 109080
rect 106556 108996 106608 109002
rect 106556 108938 106608 108944
rect 106568 104938 106596 108938
rect 106568 104910 106688 104938
rect 106660 103494 106688 104910
rect 106648 103488 106700 103494
rect 106648 103430 106700 103436
rect 106556 93900 106608 93906
rect 106556 93842 106608 93848
rect 106568 89826 106596 93842
rect 106556 89820 106608 89826
rect 106556 89762 106608 89768
rect 106648 85604 106700 85610
rect 106648 85546 106700 85552
rect 106660 75970 106688 85546
rect 106568 75942 106688 75970
rect 106568 75886 106596 75942
rect 106556 75880 106608 75886
rect 106556 75822 106608 75828
rect 106464 66360 106516 66366
rect 106464 66302 106516 66308
rect 106476 66230 106504 66302
rect 106464 66224 106516 66230
rect 106464 66166 106516 66172
rect 106556 66224 106608 66230
rect 106556 66166 106608 66172
rect 106568 51066 106596 66166
rect 106556 51060 106608 51066
rect 106556 51002 106608 51008
rect 106740 51060 106792 51066
rect 106740 51002 106792 51008
rect 106752 43466 106780 51002
rect 106752 43438 106872 43466
rect 106844 38622 106872 43438
rect 106832 38616 106884 38622
rect 106832 38558 106884 38564
rect 106832 31612 106884 31618
rect 106832 31554 106884 31560
rect 106844 4146 106872 31554
rect 107856 4146 107884 320062
rect 108132 317490 108160 320076
rect 108514 320062 108804 320090
rect 108776 317642 108804 320062
rect 108960 318306 108988 320076
rect 108948 318300 109000 318306
rect 108948 318242 109000 318248
rect 109328 317966 109356 320076
rect 109802 320062 110000 320090
rect 109972 318050 110000 320062
rect 110156 318170 110184 320076
rect 110144 318164 110196 318170
rect 110144 318106 110196 318112
rect 109972 318022 110368 318050
rect 109316 317960 109368 317966
rect 109316 317902 109368 317908
rect 110236 317960 110288 317966
rect 110236 317902 110288 317908
rect 108776 317614 108988 317642
rect 108120 317484 108172 317490
rect 108120 317426 108172 317432
rect 108856 317484 108908 317490
rect 108856 317426 108908 317432
rect 106832 4140 106884 4146
rect 106832 4082 106884 4088
rect 107568 4140 107620 4146
rect 107568 4082 107620 4088
rect 107844 4140 107896 4146
rect 107844 4082 107896 4088
rect 108764 4140 108816 4146
rect 108764 4082 108816 4088
rect 107580 480 107608 4082
rect 108776 480 108804 4082
rect 108868 3262 108896 317426
rect 108960 3398 108988 317614
rect 110248 3466 110276 317902
rect 110340 4010 110368 318022
rect 110616 317490 110644 320076
rect 110984 318034 111012 320076
rect 111458 320062 111656 320090
rect 111064 318300 111116 318306
rect 111064 318242 111116 318248
rect 110972 318028 111024 318034
rect 110972 317970 111024 317976
rect 110604 317484 110656 317490
rect 110604 317426 110656 317432
rect 110328 4004 110380 4010
rect 110328 3946 110380 3952
rect 111076 3534 111104 318242
rect 111156 318164 111208 318170
rect 111156 318106 111208 318112
rect 111168 3670 111196 318106
rect 111628 3874 111656 320062
rect 111812 318102 111840 320076
rect 112272 318170 112300 320076
rect 112260 318164 112312 318170
rect 112260 318106 112312 318112
rect 111800 318096 111852 318102
rect 111800 318038 111852 318044
rect 112640 318034 112668 320076
rect 113100 318238 113128 320076
rect 113088 318232 113140 318238
rect 113088 318174 113140 318180
rect 113468 318034 113496 320076
rect 113928 318102 113956 320076
rect 113916 318096 113968 318102
rect 113916 318038 113968 318044
rect 111708 318028 111760 318034
rect 111708 317970 111760 317976
rect 112628 318028 112680 318034
rect 112628 317970 112680 317976
rect 113088 318028 113140 318034
rect 113088 317970 113140 317976
rect 113456 318028 113508 318034
rect 113456 317970 113508 317976
rect 111616 3868 111668 3874
rect 111616 3810 111668 3816
rect 111156 3664 111208 3670
rect 111156 3606 111208 3612
rect 111064 3528 111116 3534
rect 111064 3470 111116 3476
rect 111720 3466 111748 317970
rect 113100 3670 113128 317970
rect 113824 317484 113876 317490
rect 113824 317426 113876 317432
rect 113088 3664 113140 3670
rect 113088 3606 113140 3612
rect 113836 3602 113864 317426
rect 114296 4078 114324 320076
rect 114756 318102 114784 320076
rect 114376 318096 114428 318102
rect 114376 318038 114428 318044
rect 114744 318096 114796 318102
rect 114744 318038 114796 318044
rect 114284 4072 114336 4078
rect 114284 4014 114336 4020
rect 113824 3596 113876 3602
rect 113824 3538 113876 3544
rect 112352 3528 112404 3534
rect 112352 3470 112404 3476
rect 110236 3460 110288 3466
rect 110236 3402 110288 3408
rect 111708 3460 111760 3466
rect 111708 3402 111760 3408
rect 108948 3392 109000 3398
rect 108948 3334 109000 3340
rect 111156 3392 111208 3398
rect 111156 3334 111208 3340
rect 108856 3256 108908 3262
rect 108856 3198 108908 3204
rect 109960 3256 110012 3262
rect 109960 3198 110012 3204
rect 109972 480 110000 3198
rect 111168 480 111196 3334
rect 112364 480 112392 3470
rect 114388 3398 114416 318038
rect 114468 318028 114520 318034
rect 114468 317970 114520 317976
rect 113548 3392 113600 3398
rect 113548 3334 113600 3340
rect 114376 3392 114428 3398
rect 114376 3334 114428 3340
rect 113560 480 113588 3334
rect 114480 3194 114508 317970
rect 115124 317898 115152 320076
rect 115506 320062 115796 320090
rect 115664 318096 115716 318102
rect 115664 318038 115716 318044
rect 115112 317892 115164 317898
rect 115112 317834 115164 317840
rect 115676 4010 115704 318038
rect 114744 4004 114796 4010
rect 114744 3946 114796 3952
rect 115664 4004 115716 4010
rect 115664 3946 115716 3952
rect 114468 3188 114520 3194
rect 114468 3130 114520 3136
rect 114756 480 114784 3946
rect 115768 3738 115796 320062
rect 115952 318034 115980 320076
rect 116320 318102 116348 320076
rect 116794 320062 116900 320090
rect 116584 318164 116636 318170
rect 116584 318106 116636 318112
rect 116308 318096 116360 318102
rect 116308 318038 116360 318044
rect 115940 318028 115992 318034
rect 115940 317970 115992 317976
rect 115848 317892 115900 317898
rect 115848 317834 115900 317840
rect 115860 3806 115888 317834
rect 115848 3800 115900 3806
rect 115848 3742 115900 3748
rect 115756 3732 115808 3738
rect 115756 3674 115808 3680
rect 115940 3528 115992 3534
rect 115940 3470 115992 3476
rect 115952 480 115980 3470
rect 116596 3330 116624 318106
rect 116872 318050 116900 320062
rect 117148 318646 117176 320076
rect 117136 318640 117188 318646
rect 117136 318582 117188 318588
rect 117228 318096 117280 318102
rect 116872 318022 117084 318050
rect 117228 318038 117280 318044
rect 116952 5092 117004 5098
rect 116952 5034 117004 5040
rect 116584 3324 116636 3330
rect 116584 3266 116636 3272
rect 116964 2854 116992 5034
rect 117056 3058 117084 318022
rect 117136 318028 117188 318034
rect 117136 317970 117188 317976
rect 117148 4978 117176 317970
rect 117240 5098 117268 318038
rect 117608 317626 117636 320076
rect 117990 320062 118280 320090
rect 118252 318050 118280 320062
rect 118436 318782 118464 320076
rect 118424 318776 118476 318782
rect 118424 318718 118476 318724
rect 118252 318022 118648 318050
rect 118804 318034 118832 320076
rect 119264 318102 119292 320076
rect 119252 318096 119304 318102
rect 119252 318038 119304 318044
rect 117596 317620 117648 317626
rect 117596 317562 117648 317568
rect 118516 317620 118568 317626
rect 118516 317562 118568 317568
rect 117228 5092 117280 5098
rect 117228 5034 117280 5040
rect 117148 4950 117268 4978
rect 117136 3596 117188 3602
rect 117136 3538 117188 3544
rect 117044 3052 117096 3058
rect 117044 2994 117096 3000
rect 116952 2848 117004 2854
rect 116952 2790 117004 2796
rect 117148 480 117176 3538
rect 117240 2990 117268 4950
rect 118240 3460 118292 3466
rect 118240 3402 118292 3408
rect 117228 2984 117280 2990
rect 117228 2926 117280 2932
rect 118252 480 118280 3402
rect 118528 3398 118556 317562
rect 118620 3466 118648 318022
rect 118792 318028 118844 318034
rect 118792 317970 118844 317976
rect 119632 317898 119660 320076
rect 120092 318306 120120 320076
rect 120080 318300 120132 318306
rect 120080 318242 120132 318248
rect 119896 318096 119948 318102
rect 119896 318038 119948 318044
rect 119620 317892 119672 317898
rect 119620 317834 119672 317840
rect 119436 3868 119488 3874
rect 119436 3810 119488 3816
rect 118608 3460 118660 3466
rect 118608 3402 118660 3408
rect 118516 3392 118568 3398
rect 118516 3334 118568 3340
rect 119448 480 119476 3810
rect 119908 3126 119936 318038
rect 119988 318028 120040 318034
rect 119988 317970 120040 317976
rect 119896 3120 119948 3126
rect 119896 3062 119948 3068
rect 120000 2922 120028 317970
rect 120264 317960 120316 317966
rect 120264 317902 120316 317908
rect 119988 2916 120040 2922
rect 119988 2858 120040 2864
rect 120276 626 120304 317902
rect 120460 317626 120488 320076
rect 120920 318034 120948 320076
rect 121288 318170 121316 320076
rect 121276 318164 121328 318170
rect 121276 318106 121328 318112
rect 121748 318102 121776 320076
rect 121736 318096 121788 318102
rect 121736 318038 121788 318044
rect 120908 318028 120960 318034
rect 120908 317970 120960 317976
rect 122116 317830 122144 320076
rect 122590 320062 122696 320090
rect 122564 318096 122616 318102
rect 122564 318038 122616 318044
rect 122104 317824 122156 317830
rect 122104 317766 122156 317772
rect 120448 317620 120500 317626
rect 120448 317562 120500 317568
rect 121368 317620 121420 317626
rect 121368 317562 121420 317568
rect 121380 3942 121408 317562
rect 121368 3936 121420 3942
rect 121368 3878 121420 3884
rect 122576 3534 122604 318038
rect 122668 3874 122696 320062
rect 122944 317966 122972 320076
rect 122932 317960 122984 317966
rect 122932 317902 122984 317908
rect 122748 317824 122800 317830
rect 122748 317766 122800 317772
rect 122656 3868 122708 3874
rect 122656 3810 122708 3816
rect 122564 3528 122616 3534
rect 122564 3470 122616 3476
rect 121828 3324 121880 3330
rect 121828 3266 121880 3272
rect 120276 598 120672 626
rect 120644 480 120672 598
rect 121840 480 121868 3266
rect 122760 3194 122788 317766
rect 123404 317762 123432 320076
rect 123772 318442 123800 320076
rect 123760 318436 123812 318442
rect 123760 318378 123812 318384
rect 124232 318374 124260 320076
rect 124220 318368 124272 318374
rect 124220 318310 124272 318316
rect 123484 318232 123536 318238
rect 123484 318174 123536 318180
rect 123392 317756 123444 317762
rect 123392 317698 123444 317704
rect 123024 3664 123076 3670
rect 123024 3606 123076 3612
rect 122748 3188 122800 3194
rect 122748 3130 122800 3136
rect 123036 480 123064 3606
rect 123496 3534 123524 318174
rect 124600 317966 124628 320076
rect 125074 320062 125180 320090
rect 125152 318050 125180 320062
rect 125152 318022 125364 318050
rect 124128 317960 124180 317966
rect 124128 317902 124180 317908
rect 124588 317960 124640 317966
rect 124588 317902 124640 317908
rect 124036 317756 124088 317762
rect 124036 317698 124088 317704
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124048 3262 124076 317698
rect 124140 3618 124168 317902
rect 125336 4146 125364 318022
rect 125324 4140 125376 4146
rect 125324 4082 125376 4088
rect 125428 4026 125456 320076
rect 125508 317960 125560 317966
rect 125508 317902 125560 317908
rect 125336 3998 125456 4026
rect 124140 3590 124352 3618
rect 124324 3534 124352 3590
rect 124220 3528 124272 3534
rect 124220 3470 124272 3476
rect 124312 3528 124364 3534
rect 124312 3470 124364 3476
rect 124036 3256 124088 3262
rect 124036 3198 124088 3204
rect 124232 480 124260 3470
rect 125336 3233 125364 3998
rect 125520 3398 125548 317902
rect 125888 317898 125916 320076
rect 126256 317966 126284 320076
rect 126624 318714 126652 320076
rect 126612 318708 126664 318714
rect 126612 318650 126664 318656
rect 126244 317960 126296 317966
rect 126244 317902 126296 317908
rect 126888 317960 126940 317966
rect 126888 317902 126940 317908
rect 125876 317892 125928 317898
rect 125876 317834 125928 317840
rect 126900 3602 126928 317902
rect 127084 317762 127112 320076
rect 127452 317966 127480 320076
rect 127912 318578 127940 320076
rect 127900 318572 127952 318578
rect 127900 318514 127952 318520
rect 128280 318238 128308 320076
rect 128268 318232 128320 318238
rect 128268 318174 128320 318180
rect 128740 317966 128768 320076
rect 127440 317960 127492 317966
rect 127440 317902 127492 317908
rect 128268 317960 128320 317966
rect 128268 317902 128320 317908
rect 128728 317960 128780 317966
rect 128728 317902 128780 317908
rect 127072 317756 127124 317762
rect 127072 317698 127124 317704
rect 128176 317756 128228 317762
rect 128176 317698 128228 317704
rect 128188 4078 128216 317698
rect 127532 4072 127584 4078
rect 128176 4072 128228 4078
rect 127584 4020 127848 4026
rect 127532 4014 127848 4020
rect 128176 4014 128228 4020
rect 127544 3998 127848 4014
rect 126612 3596 126664 3602
rect 126612 3538 126664 3544
rect 126888 3596 126940 3602
rect 126888 3538 126940 3544
rect 125416 3392 125468 3398
rect 125416 3334 125468 3340
rect 125508 3392 125560 3398
rect 125508 3334 125560 3340
rect 125322 3224 125378 3233
rect 125322 3159 125378 3168
rect 125428 480 125456 3334
rect 126624 480 126652 3538
rect 127820 480 127848 3998
rect 128280 3505 128308 317902
rect 129108 317830 129136 320076
rect 129096 317824 129148 317830
rect 129096 317766 129148 317772
rect 129464 317824 129516 317830
rect 129464 317766 129516 317772
rect 129476 6594 129504 317766
rect 129464 6588 129516 6594
rect 129464 6530 129516 6536
rect 129568 4049 129596 320076
rect 129936 317966 129964 320076
rect 129648 317960 129700 317966
rect 129648 317902 129700 317908
rect 129924 317960 129976 317966
rect 129924 317902 129976 317908
rect 129554 4040 129610 4049
rect 129004 4004 129056 4010
rect 129660 4010 129688 317902
rect 130396 317830 130424 320076
rect 130778 320062 130976 320090
rect 130384 317824 130436 317830
rect 130384 317766 130436 317772
rect 130844 317824 130896 317830
rect 130844 317766 130896 317772
rect 130856 6526 130884 317766
rect 130844 6520 130896 6526
rect 130844 6462 130896 6468
rect 129554 3975 129610 3984
rect 129648 4004 129700 4010
rect 129004 3946 129056 3952
rect 129648 3946 129700 3952
rect 128266 3496 128322 3505
rect 128266 3431 128322 3440
rect 129016 480 129044 3946
rect 130948 3913 130976 320062
rect 131028 317960 131080 317966
rect 131028 317902 131080 317908
rect 130934 3904 130990 3913
rect 130934 3839 130990 3848
rect 131040 3806 131068 317902
rect 131224 317898 131252 320076
rect 131212 317892 131264 317898
rect 131212 317834 131264 317840
rect 131592 317830 131620 320076
rect 132066 320062 132264 320090
rect 132132 318504 132184 318510
rect 132132 318446 132184 318452
rect 131580 317824 131632 317830
rect 131580 317766 131632 317772
rect 132144 317694 132172 318446
rect 132236 318050 132264 320062
rect 132420 318510 132448 320076
rect 132408 318504 132460 318510
rect 132408 318446 132460 318452
rect 132236 318022 132356 318050
rect 132880 318034 132908 320076
rect 133262 320062 133552 320090
rect 133144 318776 133196 318782
rect 133144 318718 133196 318724
rect 132224 317824 132276 317830
rect 132224 317766 132276 317772
rect 132132 317688 132184 317694
rect 132132 317630 132184 317636
rect 132236 6458 132264 317766
rect 132224 6452 132276 6458
rect 132224 6394 132276 6400
rect 130200 3800 130252 3806
rect 130200 3742 130252 3748
rect 131028 3800 131080 3806
rect 132328 3777 132356 318022
rect 132868 318028 132920 318034
rect 132868 317970 132920 317976
rect 132408 317892 132460 317898
rect 132408 317834 132460 317840
rect 131028 3742 131080 3748
rect 132314 3768 132370 3777
rect 130212 480 130240 3742
rect 131396 3732 131448 3738
rect 132420 3738 132448 317834
rect 132314 3703 132370 3712
rect 132408 3732 132460 3738
rect 131396 3674 131448 3680
rect 132408 3674 132460 3680
rect 131408 480 131436 3674
rect 133156 3466 133184 318718
rect 133236 318640 133288 318646
rect 133236 318582 133288 318588
rect 133248 3534 133276 318582
rect 133524 318510 133552 320062
rect 133512 318504 133564 318510
rect 133512 318446 133564 318452
rect 133708 317490 133736 320076
rect 133788 318028 133840 318034
rect 133788 317970 133840 317976
rect 133696 317484 133748 317490
rect 133696 317426 133748 317432
rect 133800 6390 133828 317970
rect 134076 317830 134104 320076
rect 134536 318646 134564 320076
rect 134524 318640 134576 318646
rect 134524 318582 134576 318588
rect 134524 317960 134576 317966
rect 134524 317902 134576 317908
rect 134064 317824 134116 317830
rect 134064 317766 134116 317772
rect 133788 6384 133840 6390
rect 133788 6326 133840 6332
rect 134536 4214 134564 317902
rect 134904 317762 134932 320076
rect 135364 318034 135392 320076
rect 135732 318782 135760 320076
rect 135720 318776 135772 318782
rect 135720 318718 135772 318724
rect 135352 318028 135404 318034
rect 135352 317970 135404 317976
rect 136192 317898 136220 320076
rect 136560 318186 136588 320076
rect 136468 318158 136588 318186
rect 136180 317892 136232 317898
rect 136180 317834 136232 317840
rect 135168 317824 135220 317830
rect 135168 317766 135220 317772
rect 134892 317756 134944 317762
rect 134892 317698 134944 317704
rect 135180 6322 135208 317766
rect 135904 317688 135956 317694
rect 135904 317630 135956 317636
rect 135168 6316 135220 6322
rect 135168 6258 135220 6264
rect 134524 4208 134576 4214
rect 134524 4150 134576 4156
rect 133236 3528 133288 3534
rect 133236 3470 133288 3476
rect 133144 3460 133196 3466
rect 133144 3402 133196 3408
rect 135916 3058 135944 317630
rect 136468 6186 136496 318158
rect 137020 318034 137048 320076
rect 136548 318028 136600 318034
rect 136548 317970 136600 317976
rect 137008 318028 137060 318034
rect 137008 317970 137060 317976
rect 136560 6254 136588 317970
rect 137388 317830 137416 320076
rect 137376 317824 137428 317830
rect 137376 317766 137428 317772
rect 137756 317558 137784 320076
rect 137928 318028 137980 318034
rect 137928 317970 137980 317976
rect 137744 317552 137796 317558
rect 137744 317494 137796 317500
rect 136548 6248 136600 6254
rect 136548 6190 136600 6196
rect 136456 6180 136508 6186
rect 136456 6122 136508 6128
rect 136088 3528 136140 3534
rect 136088 3470 136140 3476
rect 134892 3052 134944 3058
rect 134892 2994 134944 3000
rect 135904 3052 135956 3058
rect 135904 2994 135956 3000
rect 132592 2984 132644 2990
rect 132592 2926 132644 2932
rect 132604 480 132632 2926
rect 133788 2848 133840 2854
rect 133788 2790 133840 2796
rect 133800 480 133828 2790
rect 134904 480 134932 2994
rect 136100 480 136128 3470
rect 137940 3058 137968 317970
rect 138216 317694 138244 320076
rect 138204 317688 138256 317694
rect 138204 317630 138256 317636
rect 138584 317490 138612 320076
rect 139058 320062 139256 320090
rect 138572 317484 138624 317490
rect 138572 317426 138624 317432
rect 139228 317422 139256 320062
rect 139412 317626 139440 320076
rect 139400 317620 139452 317626
rect 139400 317562 139452 317568
rect 139872 317490 139900 320076
rect 140254 320062 140544 320090
rect 139308 317484 139360 317490
rect 139308 317426 139360 317432
rect 139860 317484 139912 317490
rect 139860 317426 139912 317432
rect 139216 317416 139268 317422
rect 139216 317358 139268 317364
rect 139320 4282 139348 317426
rect 140516 8022 140544 320062
rect 140700 318306 140728 320076
rect 140688 318300 140740 318306
rect 140688 318242 140740 318248
rect 140688 317620 140740 317626
rect 140688 317562 140740 317568
rect 140596 317484 140648 317490
rect 140596 317426 140648 317432
rect 140504 8016 140556 8022
rect 140504 7958 140556 7964
rect 140608 4350 140636 317426
rect 140596 4344 140648 4350
rect 140596 4286 140648 4292
rect 139308 4276 139360 4282
rect 139308 4218 139360 4224
rect 140700 3466 140728 317562
rect 141068 317490 141096 320076
rect 141542 320062 141648 320090
rect 141910 320062 142108 320090
rect 141424 317960 141476 317966
rect 141424 317902 141476 317908
rect 141056 317484 141108 317490
rect 141056 317426 141108 317432
rect 141436 3534 141464 317902
rect 141620 316010 141648 320062
rect 142080 318850 142108 320062
rect 142068 318844 142120 318850
rect 142068 318786 142120 318792
rect 142356 317490 142384 320076
rect 142738 320062 142936 320090
rect 142068 317484 142120 317490
rect 142068 317426 142120 317432
rect 142344 317484 142396 317490
rect 142344 317426 142396 317432
rect 141620 315982 142016 316010
rect 141988 7954 142016 315982
rect 141976 7948 142028 7954
rect 141976 7890 142028 7896
rect 142080 4418 142108 317426
rect 142908 316010 142936 320062
rect 143184 318073 143212 320076
rect 143170 318064 143226 318073
rect 143170 317999 143226 318008
rect 143552 317490 143580 320076
rect 144026 320062 144132 320090
rect 143448 317484 143500 317490
rect 143448 317426 143500 317432
rect 143540 317484 143592 317490
rect 143540 317426 143592 317432
rect 142908 315982 143396 316010
rect 143368 7886 143396 315982
rect 143356 7880 143408 7886
rect 143356 7822 143408 7828
rect 143460 4486 143488 317426
rect 144104 316010 144132 320062
rect 144380 317626 144408 320076
rect 144840 317744 144868 320076
rect 144748 317716 144868 317744
rect 144368 317620 144420 317626
rect 144368 317562 144420 317568
rect 144644 317484 144696 317490
rect 144644 317426 144696 317432
rect 144104 315982 144592 316010
rect 144564 7818 144592 315982
rect 144552 7812 144604 7818
rect 144552 7754 144604 7760
rect 144656 4554 144684 317426
rect 144748 4622 144776 317716
rect 144828 317620 144880 317626
rect 144828 317562 144880 317568
rect 144736 4616 144788 4622
rect 144736 4558 144788 4564
rect 144644 4548 144696 4554
rect 144644 4490 144696 4496
rect 143448 4480 143500 4486
rect 143448 4422 143500 4428
rect 142068 4412 142120 4418
rect 142068 4354 142120 4360
rect 141424 3528 141476 3534
rect 141424 3470 141476 3476
rect 144460 3528 144512 3534
rect 144460 3470 144512 3476
rect 139676 3460 139728 3466
rect 139676 3402 139728 3408
rect 140688 3460 140740 3466
rect 140688 3402 140740 3408
rect 137928 3052 137980 3058
rect 137928 2994 137980 3000
rect 138480 2984 138532 2990
rect 138480 2926 138532 2932
rect 137284 2848 137336 2854
rect 137284 2790 137336 2796
rect 137296 480 137324 2790
rect 138492 480 138520 2926
rect 139688 480 139716 3402
rect 142068 3120 142120 3126
rect 142068 3062 142120 3068
rect 140872 2916 140924 2922
rect 140872 2858 140924 2864
rect 140884 480 140912 2858
rect 142080 480 142108 3062
rect 143264 3052 143316 3058
rect 143264 2994 143316 3000
rect 143276 480 143304 2994
rect 144472 480 144500 3470
rect 144840 3369 144868 317562
rect 145208 317490 145236 320076
rect 145668 318714 145696 320076
rect 146050 320062 146248 320090
rect 145656 318708 145708 318714
rect 145656 318650 145708 318656
rect 145656 318096 145708 318102
rect 145656 318038 145708 318044
rect 145564 317756 145616 317762
rect 145564 317698 145616 317704
rect 145196 317484 145248 317490
rect 145196 317426 145248 317432
rect 145576 4842 145604 317698
rect 145484 4814 145604 4842
rect 144826 3360 144882 3369
rect 144826 3295 144882 3304
rect 145484 3126 145512 4814
rect 145564 4140 145616 4146
rect 145564 4082 145616 4088
rect 145576 3346 145604 4082
rect 145668 3534 145696 318038
rect 146116 317484 146168 317490
rect 146116 317426 146168 317432
rect 146128 7750 146156 317426
rect 146116 7744 146168 7750
rect 146116 7686 146168 7692
rect 146220 4690 146248 320062
rect 146496 317490 146524 320076
rect 146864 318102 146892 320076
rect 147338 320062 147536 320090
rect 147404 318436 147456 318442
rect 147404 318378 147456 318384
rect 147416 318209 147444 318378
rect 147402 318200 147458 318209
rect 147402 318135 147458 318144
rect 146852 318096 146904 318102
rect 146852 318038 146904 318044
rect 146576 318028 146628 318034
rect 146576 317970 146628 317976
rect 146484 317484 146536 317490
rect 146484 317426 146536 317432
rect 146208 4684 146260 4690
rect 146208 4626 146260 4632
rect 145656 3528 145708 3534
rect 145656 3470 145708 3476
rect 145576 3318 145696 3346
rect 145472 3120 145524 3126
rect 145472 3062 145524 3068
rect 145668 480 145696 3318
rect 146588 610 146616 317970
rect 147404 317484 147456 317490
rect 147404 317426 147456 317432
rect 147416 315874 147444 317426
rect 147508 316010 147536 320062
rect 147692 317762 147720 320076
rect 148152 318714 148180 320076
rect 148140 318708 148192 318714
rect 148140 318650 148192 318656
rect 147862 318200 147918 318209
rect 147862 318135 147864 318144
rect 147916 318135 147918 318144
rect 147864 318106 147916 318112
rect 148324 317824 148376 317830
rect 148324 317766 148376 317772
rect 147680 317756 147732 317762
rect 147680 317698 147732 317704
rect 147508 315982 147628 316010
rect 147416 315846 147536 315874
rect 147508 7682 147536 315846
rect 147496 7676 147548 7682
rect 147496 7618 147548 7624
rect 147600 4758 147628 315982
rect 147588 4752 147640 4758
rect 147588 4694 147640 4700
rect 148336 4078 148364 317766
rect 148520 317490 148548 320076
rect 148784 317756 148836 317762
rect 148784 317698 148836 317704
rect 148508 317484 148560 317490
rect 148508 317426 148560 317432
rect 148796 7614 148824 317698
rect 148784 7608 148836 7614
rect 148784 7550 148836 7556
rect 148888 5438 148916 320076
rect 149348 318374 149376 320076
rect 149730 320062 149836 320090
rect 150190 320062 150388 320090
rect 150558 320062 150848 320090
rect 151018 320062 151216 320090
rect 151386 320062 151676 320090
rect 149808 318442 149836 320062
rect 149704 318436 149756 318442
rect 149704 318378 149756 318384
rect 149796 318436 149848 318442
rect 149796 318378 149848 318384
rect 150256 318436 150308 318442
rect 150256 318378 150308 318384
rect 149336 318368 149388 318374
rect 149336 318310 149388 318316
rect 148968 317484 149020 317490
rect 148968 317426 149020 317432
rect 148980 5506 149008 317426
rect 148968 5500 149020 5506
rect 148968 5442 149020 5448
rect 148876 5432 148928 5438
rect 148876 5374 148928 5380
rect 148324 4072 148376 4078
rect 148324 4014 148376 4020
rect 149244 3936 149296 3942
rect 149244 3878 149296 3884
rect 148048 3528 148100 3534
rect 148048 3470 148100 3476
rect 146576 604 146628 610
rect 146576 546 146628 552
rect 146852 604 146904 610
rect 146852 546 146904 552
rect 146864 480 146892 546
rect 148060 480 148088 3470
rect 149256 480 149284 3878
rect 149716 2854 149744 318378
rect 150268 5370 150296 318378
rect 150256 5364 150308 5370
rect 150256 5306 150308 5312
rect 150360 5302 150388 320062
rect 150820 318850 150848 320062
rect 150808 318844 150860 318850
rect 150808 318786 150860 318792
rect 150900 318164 150952 318170
rect 150900 318106 150952 318112
rect 150912 312662 150940 318106
rect 151084 317620 151136 317626
rect 151084 317562 151136 317568
rect 151096 312746 151124 317562
rect 151188 312882 151216 320062
rect 151648 316010 151676 320062
rect 151832 317490 151860 320076
rect 152200 317558 152228 320076
rect 152674 320062 152872 320090
rect 152464 318300 152516 318306
rect 152464 318242 152516 318248
rect 152188 317552 152240 317558
rect 152188 317494 152240 317500
rect 151820 317484 151872 317490
rect 151820 317426 151872 317432
rect 151648 315982 151768 316010
rect 151188 312854 151676 312882
rect 151096 312718 151308 312746
rect 150900 312656 150952 312662
rect 150900 312598 150952 312604
rect 151176 312656 151228 312662
rect 151176 312598 151228 312604
rect 151084 309188 151136 309194
rect 151084 309130 151136 309136
rect 151096 299470 151124 309130
rect 151084 299464 151136 299470
rect 151084 299406 151136 299412
rect 151084 289876 151136 289882
rect 151084 289818 151136 289824
rect 151096 280158 151124 289818
rect 151084 280152 151136 280158
rect 151084 280094 151136 280100
rect 151084 270564 151136 270570
rect 151084 270506 151136 270512
rect 151096 260846 151124 270506
rect 151084 260840 151136 260846
rect 151084 260782 151136 260788
rect 151084 251252 151136 251258
rect 151084 251194 151136 251200
rect 151096 241505 151124 251194
rect 151082 241496 151138 241505
rect 151082 241431 151138 241440
rect 150990 241360 151046 241369
rect 150990 241295 151046 241304
rect 151004 231878 151032 241295
rect 150992 231872 151044 231878
rect 150992 231814 151044 231820
rect 151084 231872 151136 231878
rect 151084 231814 151136 231820
rect 151096 222193 151124 231814
rect 151082 222184 151138 222193
rect 151082 222119 151138 222128
rect 150990 222048 151046 222057
rect 150990 221983 151046 221992
rect 151004 212566 151032 221983
rect 150992 212560 151044 212566
rect 150992 212502 151044 212508
rect 151084 212560 151136 212566
rect 151084 212502 151136 212508
rect 151096 202881 151124 212502
rect 151082 202872 151138 202881
rect 151082 202807 151138 202816
rect 150990 202736 151046 202745
rect 150990 202671 151046 202680
rect 151004 193254 151032 202671
rect 150992 193248 151044 193254
rect 150992 193190 151044 193196
rect 151084 193248 151136 193254
rect 151084 193190 151136 193196
rect 151096 183569 151124 193190
rect 151082 183560 151138 183569
rect 151082 183495 151138 183504
rect 150990 183424 151046 183433
rect 150990 183359 151046 183368
rect 151004 173942 151032 183359
rect 150992 173936 151044 173942
rect 150992 173878 151044 173884
rect 151084 173936 151136 173942
rect 151084 173878 151136 173884
rect 151096 164218 151124 173878
rect 151084 164212 151136 164218
rect 151084 164154 151136 164160
rect 151084 154624 151136 154630
rect 151084 154566 151136 154572
rect 151096 144906 151124 154566
rect 151084 144900 151136 144906
rect 151084 144842 151136 144848
rect 151084 135312 151136 135318
rect 151084 135254 151136 135260
rect 151096 125594 151124 135254
rect 151084 125588 151136 125594
rect 151084 125530 151136 125536
rect 151084 116000 151136 116006
rect 151084 115942 151136 115948
rect 151096 106282 151124 115942
rect 151084 106276 151136 106282
rect 151084 106218 151136 106224
rect 151084 96688 151136 96694
rect 151084 96630 151136 96636
rect 151096 86970 151124 96630
rect 151084 86964 151136 86970
rect 151084 86906 151136 86912
rect 151084 77308 151136 77314
rect 151084 77250 151136 77256
rect 151096 67590 151124 77250
rect 151084 67584 151136 67590
rect 151084 67526 151136 67532
rect 151084 57996 151136 58002
rect 151084 57938 151136 57944
rect 151096 48278 151124 57938
rect 151084 48272 151136 48278
rect 151084 48214 151136 48220
rect 151084 38684 151136 38690
rect 151084 38626 151136 38632
rect 151096 28966 151124 38626
rect 151084 28960 151136 28966
rect 151084 28902 151136 28908
rect 151084 19372 151136 19378
rect 151084 19314 151136 19320
rect 151096 9659 151124 19314
rect 151082 9650 151138 9659
rect 151082 9585 151138 9594
rect 150348 5296 150400 5302
rect 150348 5238 150400 5244
rect 151188 3942 151216 312598
rect 151176 3936 151228 3942
rect 151176 3878 151228 3884
rect 151280 3398 151308 312718
rect 151648 5234 151676 312854
rect 151636 5228 151688 5234
rect 151636 5170 151688 5176
rect 151740 5166 151768 315982
rect 151728 5160 151780 5166
rect 151728 5102 151780 5108
rect 152476 3874 152504 318242
rect 152648 317484 152700 317490
rect 152648 317426 152700 317432
rect 152660 315874 152688 317426
rect 152844 316010 152872 320062
rect 152844 315982 152964 316010
rect 152660 315846 152872 315874
rect 152844 8702 152872 315846
rect 152936 8770 152964 315982
rect 153028 8974 153056 320076
rect 153108 317552 153160 317558
rect 153108 317494 153160 317500
rect 153016 8968 153068 8974
rect 153016 8910 153068 8916
rect 152924 8764 152976 8770
rect 152924 8706 152976 8712
rect 152832 8696 152884 8702
rect 152832 8638 152884 8644
rect 153120 5098 153148 317494
rect 153488 317490 153516 320076
rect 153856 318374 153884 320076
rect 154330 320062 154436 320090
rect 153844 318368 153896 318374
rect 153844 318310 153896 318316
rect 154304 318368 154356 318374
rect 154304 318310 154356 318316
rect 153844 317960 153896 317966
rect 153844 317902 153896 317908
rect 153476 317484 153528 317490
rect 153476 317426 153528 317432
rect 153198 9480 153254 9489
rect 153198 9415 153254 9424
rect 153108 5092 153160 5098
rect 153108 5034 153160 5040
rect 151544 3868 151596 3874
rect 151544 3810 151596 3816
rect 152464 3868 152516 3874
rect 152464 3810 152516 3816
rect 151268 3392 151320 3398
rect 151268 3334 151320 3340
rect 150440 3188 150492 3194
rect 150440 3130 150492 3136
rect 149704 2848 149756 2854
rect 149704 2790 149756 2796
rect 150452 480 150480 3130
rect 151556 480 151584 3810
rect 153212 3058 153240 9415
rect 153856 4078 153884 317902
rect 153936 317620 153988 317626
rect 153936 317562 153988 317568
rect 153844 4072 153896 4078
rect 153844 4014 153896 4020
rect 153948 3890 153976 317562
rect 154316 8906 154344 318310
rect 154408 9654 154436 320062
rect 154684 317558 154712 320076
rect 154672 317552 154724 317558
rect 154672 317494 154724 317500
rect 155144 317490 155172 320076
rect 155526 320062 155724 320090
rect 155224 317756 155276 317762
rect 155224 317698 155276 317704
rect 154488 317484 154540 317490
rect 154488 317426 154540 317432
rect 155132 317484 155184 317490
rect 155132 317426 155184 317432
rect 154396 9648 154448 9654
rect 154396 9590 154448 9596
rect 154304 8900 154356 8906
rect 154304 8842 154356 8848
rect 154500 5030 154528 317426
rect 154488 5024 154540 5030
rect 154488 4966 154540 4972
rect 153856 3862 153976 3890
rect 155132 3936 155184 3942
rect 155132 3878 155184 3884
rect 153856 3126 153884 3862
rect 153936 3664 153988 3670
rect 153936 3606 153988 3612
rect 153844 3120 153896 3126
rect 153844 3062 153896 3068
rect 152740 3052 152792 3058
rect 152740 2994 152792 3000
rect 153200 3052 153252 3058
rect 153200 2994 153252 3000
rect 151726 2952 151782 2961
rect 151726 2887 151728 2896
rect 151780 2887 151782 2896
rect 151728 2858 151780 2864
rect 152752 480 152780 2994
rect 153948 480 153976 3606
rect 155144 480 155172 3878
rect 155236 3670 155264 317698
rect 155696 9518 155724 320062
rect 155972 317558 156000 320076
rect 155868 317552 155920 317558
rect 155868 317494 155920 317500
rect 155960 317552 156012 317558
rect 155960 317494 156012 317500
rect 155776 317484 155828 317490
rect 155776 317426 155828 317432
rect 155788 9586 155816 317426
rect 155776 9580 155828 9586
rect 155776 9522 155828 9528
rect 155684 9512 155736 9518
rect 155684 9454 155736 9460
rect 155880 4962 155908 317494
rect 156340 317490 156368 320076
rect 156814 320062 157012 320090
rect 156604 318164 156656 318170
rect 156604 318106 156656 318112
rect 156328 317484 156380 317490
rect 156328 317426 156380 317432
rect 156616 7478 156644 318106
rect 156984 9382 157012 320062
rect 157064 317484 157116 317490
rect 157064 317426 157116 317432
rect 157076 9450 157104 317426
rect 157064 9444 157116 9450
rect 157064 9386 157116 9392
rect 156972 9376 157024 9382
rect 156972 9318 157024 9324
rect 156604 7472 156656 7478
rect 156604 7414 156656 7420
rect 157168 5574 157196 320076
rect 157642 320062 157840 320090
rect 158010 320062 158300 320090
rect 158470 320062 158668 320090
rect 157248 317552 157300 317558
rect 157248 317494 157300 317500
rect 157156 5568 157208 5574
rect 157156 5510 157208 5516
rect 155868 4956 155920 4962
rect 155868 4898 155920 4904
rect 157260 4894 157288 317494
rect 157812 315926 157840 320062
rect 157984 318504 158036 318510
rect 157984 318446 158036 318452
rect 157800 315920 157852 315926
rect 157800 315862 157852 315868
rect 157248 4888 157300 4894
rect 157248 4830 157300 4836
rect 156328 4072 156380 4078
rect 156328 4014 156380 4020
rect 155224 3664 155276 3670
rect 155224 3606 155276 3612
rect 156340 480 156368 4014
rect 157996 3330 158024 318446
rect 158076 317688 158128 317694
rect 158076 317630 158128 317636
rect 158088 3641 158116 317630
rect 158272 316010 158300 320062
rect 158272 315982 158576 316010
rect 158444 315920 158496 315926
rect 158444 315862 158496 315868
rect 158456 9246 158484 315862
rect 158548 9314 158576 315982
rect 158536 9308 158588 9314
rect 158536 9250 158588 9256
rect 158444 9240 158496 9246
rect 158444 9182 158496 9188
rect 158640 5409 158668 320062
rect 158824 317558 158852 320076
rect 159284 318442 159312 320076
rect 159456 318776 159508 318782
rect 159456 318718 159508 318724
rect 159364 318640 159416 318646
rect 159364 318582 159416 318588
rect 159272 318436 159324 318442
rect 159272 318378 159324 318384
rect 158812 317552 158864 317558
rect 158812 317494 158864 317500
rect 158626 5400 158682 5409
rect 158626 5335 158682 5344
rect 158074 3632 158130 3641
rect 158074 3567 158130 3576
rect 159376 3398 159404 318582
rect 159364 3392 159416 3398
rect 159364 3334 159416 3340
rect 159468 3330 159496 318718
rect 159652 317490 159680 320076
rect 159836 320062 160034 320090
rect 159640 317484 159692 317490
rect 159640 317426 159692 317432
rect 159836 9110 159864 320062
rect 160480 318374 160508 320076
rect 160468 318368 160520 318374
rect 160468 318310 160520 318316
rect 160744 317824 160796 317830
rect 160744 317766 160796 317772
rect 159916 317552 159968 317558
rect 159916 317494 159968 317500
rect 159928 9178 159956 317494
rect 160008 317484 160060 317490
rect 160008 317426 160060 317432
rect 159916 9172 159968 9178
rect 159916 9114 159968 9120
rect 159824 9104 159876 9110
rect 159824 9046 159876 9052
rect 160020 5273 160048 317426
rect 160006 5264 160062 5273
rect 160006 5199 160062 5208
rect 157524 3324 157576 3330
rect 157524 3266 157576 3272
rect 157984 3324 158036 3330
rect 157984 3266 158036 3272
rect 159456 3324 159508 3330
rect 159456 3266 159508 3272
rect 157248 2984 157300 2990
rect 157246 2952 157248 2961
rect 157300 2952 157302 2961
rect 157246 2887 157302 2896
rect 157536 480 157564 3266
rect 158720 3256 158772 3262
rect 158720 3198 158772 3204
rect 159914 3224 159970 3233
rect 158732 480 158760 3198
rect 159914 3159 159970 3168
rect 159928 480 159956 3159
rect 160756 2854 160784 317766
rect 160848 317490 160876 320076
rect 160836 317484 160888 317490
rect 160836 317426 160888 317432
rect 161308 7002 161336 320076
rect 161676 318510 161704 320076
rect 161664 318504 161716 318510
rect 161664 318446 161716 318452
rect 162136 317490 162164 320076
rect 162518 320062 162716 320090
rect 161388 317484 161440 317490
rect 161388 317426 161440 317432
rect 162124 317484 162176 317490
rect 162124 317426 162176 317432
rect 161296 6996 161348 7002
rect 161296 6938 161348 6944
rect 161400 5137 161428 317426
rect 162124 309188 162176 309194
rect 162124 309130 162176 309136
rect 162136 9790 162164 309130
rect 162124 9784 162176 9790
rect 162124 9726 162176 9732
rect 161940 9716 161992 9722
rect 161940 9658 161992 9664
rect 161952 6662 161980 9658
rect 162688 9042 162716 320062
rect 162964 318646 162992 320076
rect 162952 318640 163004 318646
rect 162952 318582 163004 318588
rect 163332 317490 163360 320076
rect 163502 318064 163558 318073
rect 163502 317999 163558 318008
rect 162768 317484 162820 317490
rect 162768 317426 162820 317432
rect 163320 317484 163372 317490
rect 163320 317426 163372 317432
rect 162676 9036 162728 9042
rect 162676 8978 162728 8984
rect 161940 6656 161992 6662
rect 161940 6598 161992 6604
rect 161386 5128 161442 5137
rect 161386 5063 161442 5072
rect 162780 5001 162808 317426
rect 162766 4992 162822 5001
rect 162766 4927 162822 4936
rect 162308 3596 162360 3602
rect 162308 3538 162360 3544
rect 161112 3188 161164 3194
rect 161112 3130 161164 3136
rect 160744 2848 160796 2854
rect 160744 2790 160796 2796
rect 161124 480 161152 3130
rect 162320 480 162348 3538
rect 163516 3262 163544 317999
rect 163792 317558 163820 320076
rect 163976 319410 164004 320198
rect 230664 320146 230716 320152
rect 231492 320204 231794 320210
rect 231544 320198 231794 320204
rect 235566 320210 235672 320226
rect 240442 320210 240732 320226
rect 241730 320210 241928 320226
rect 235566 320204 235684 320210
rect 235566 320198 235632 320204
rect 231492 320146 231544 320152
rect 240442 320204 240744 320210
rect 240442 320198 240692 320204
rect 235632 320146 235684 320152
rect 240692 320146 240744 320152
rect 241336 320204 241388 320210
rect 241730 320204 241940 320210
rect 241730 320198 241888 320204
rect 241336 320146 241388 320152
rect 241888 320146 241940 320152
rect 242716 320204 242768 320210
rect 242716 320146 242768 320152
rect 244280 320204 244332 320210
rect 244280 320146 244332 320152
rect 244384 320198 244582 320226
rect 245120 320210 245410 320226
rect 246408 320210 246698 320226
rect 248064 320210 248354 320226
rect 245108 320204 245410 320210
rect 163976 319382 164096 319410
rect 164068 318730 164096 319382
rect 164240 318776 164292 318782
rect 163976 318702 164096 318730
rect 164238 318744 164240 318753
rect 164292 318744 164294 318753
rect 164148 318708 164200 318714
rect 163976 318238 164004 318702
rect 164238 318679 164294 318688
rect 164148 318650 164200 318656
rect 164056 318640 164108 318646
rect 164160 318594 164188 318650
rect 164108 318588 164188 318594
rect 164056 318582 164188 318588
rect 164068 318566 164188 318582
rect 163964 318232 164016 318238
rect 163964 318174 164016 318180
rect 163780 317552 163832 317558
rect 163780 317494 163832 317500
rect 164056 317552 164108 317558
rect 164056 317494 164108 317500
rect 164068 8974 164096 317494
rect 164620 317490 164648 320076
rect 164884 318572 164936 318578
rect 164884 318514 164936 318520
rect 164148 317484 164200 317490
rect 164148 317426 164200 317432
rect 164608 317484 164660 317490
rect 164608 317426 164660 317432
rect 164056 8968 164108 8974
rect 164056 8910 164108 8916
rect 164160 4865 164188 317426
rect 164146 4856 164202 4865
rect 164146 4791 164202 4800
rect 164700 4072 164752 4078
rect 164700 4014 164752 4020
rect 163504 3256 163556 3262
rect 163504 3198 163556 3204
rect 163504 2984 163556 2990
rect 163504 2926 163556 2932
rect 163596 2984 163648 2990
rect 163596 2926 163648 2932
rect 163516 480 163544 2926
rect 163608 2854 163636 2926
rect 163596 2848 163648 2854
rect 163596 2790 163648 2796
rect 164712 480 164740 4014
rect 164896 3602 164924 318514
rect 164988 317558 165016 320076
rect 164976 317552 165028 317558
rect 164976 317494 165028 317500
rect 165344 317484 165396 317490
rect 165344 317426 165396 317432
rect 165356 12510 165384 317426
rect 165344 12504 165396 12510
rect 165344 12446 165396 12452
rect 165448 11150 165476 320076
rect 165816 317558 165844 320076
rect 166172 317620 166224 317626
rect 166172 317562 166224 317568
rect 165528 317552 165580 317558
rect 165528 317494 165580 317500
rect 165804 317552 165856 317558
rect 165804 317494 165856 317500
rect 165436 11144 165488 11150
rect 165436 11086 165488 11092
rect 165540 8362 165568 317494
rect 166184 316418 166212 317562
rect 166276 317490 166304 320076
rect 166658 320062 166764 320090
rect 166264 317484 166316 317490
rect 166264 317426 166316 317432
rect 166184 316390 166304 316418
rect 165528 8356 165580 8362
rect 165528 8298 165580 8304
rect 164792 3596 164844 3602
rect 164792 3538 164844 3544
rect 164884 3596 164936 3602
rect 164884 3538 164936 3544
rect 164804 3482 164832 3538
rect 166276 3505 166304 316390
rect 166736 14074 166764 320062
rect 167000 318776 167052 318782
rect 166998 318744 167000 318753
rect 167052 318744 167054 318753
rect 166998 318679 167054 318688
rect 166908 317552 166960 317558
rect 166908 317494 166960 317500
rect 166816 317484 166868 317490
rect 166816 317426 166868 317432
rect 166724 14068 166776 14074
rect 166724 14010 166776 14016
rect 166828 13870 166856 317426
rect 166816 13864 166868 13870
rect 166816 13806 166868 13812
rect 166920 5545 166948 317494
rect 167104 317490 167132 320076
rect 167472 317558 167500 320076
rect 167946 320062 168052 320090
rect 167644 317892 167696 317898
rect 167644 317834 167696 317840
rect 167460 317552 167512 317558
rect 167460 317494 167512 317500
rect 167092 317484 167144 317490
rect 167092 317426 167144 317432
rect 166906 5536 166962 5545
rect 166906 5471 166962 5480
rect 167656 3602 167684 317834
rect 168024 14142 168052 320062
rect 168300 317642 168328 320076
rect 168208 317614 168328 317642
rect 168104 317484 168156 317490
rect 168104 317426 168156 317432
rect 168012 14136 168064 14142
rect 168012 14078 168064 14084
rect 168116 13938 168144 317426
rect 168208 14210 168236 317614
rect 168288 317552 168340 317558
rect 168288 317494 168340 317500
rect 168196 14204 168248 14210
rect 168196 14146 168248 14152
rect 168300 14006 168328 317494
rect 168760 317490 168788 320076
rect 169142 320062 169340 320090
rect 169602 320062 169708 320090
rect 168748 317484 168800 317490
rect 168748 317426 168800 317432
rect 169312 316010 169340 320062
rect 169576 317484 169628 317490
rect 169576 317426 169628 317432
rect 169312 315982 169524 316010
rect 169496 16454 169524 315982
rect 169484 16448 169536 16454
rect 169484 16390 169536 16396
rect 169588 14278 169616 317426
rect 169576 14272 169628 14278
rect 169576 14214 169628 14220
rect 168288 14000 168340 14006
rect 168288 13942 168340 13948
rect 168104 13932 168156 13938
rect 168104 13874 168156 13880
rect 169680 5574 169708 320062
rect 169956 317490 169984 320076
rect 170430 320062 170536 320090
rect 170798 320062 171088 320090
rect 169944 317484 169996 317490
rect 169944 317426 169996 317432
rect 170508 316010 170536 320062
rect 170956 317484 171008 317490
rect 170956 317426 171008 317432
rect 170508 315982 170904 316010
rect 170876 16386 170904 315982
rect 170864 16380 170916 16386
rect 170864 16322 170916 16328
rect 170968 14346 170996 317426
rect 170956 14340 171008 14346
rect 170956 14282 171008 14288
rect 170588 6588 170640 6594
rect 170588 6530 170640 6536
rect 169668 5568 169720 5574
rect 169668 5510 169720 5516
rect 169392 4004 169444 4010
rect 169392 3946 169444 3952
rect 167092 3596 167144 3602
rect 167092 3538 167144 3544
rect 167644 3596 167696 3602
rect 167644 3538 167696 3544
rect 168288 3596 168340 3602
rect 168288 3538 168340 3544
rect 165894 3496 165950 3505
rect 164804 3454 164924 3482
rect 164896 3398 164924 3454
rect 165894 3431 165950 3440
rect 166262 3496 166318 3505
rect 166262 3431 166318 3440
rect 164884 3392 164936 3398
rect 164884 3334 164936 3340
rect 165908 480 165936 3431
rect 167104 480 167132 3538
rect 168300 3194 168328 3538
rect 168196 3188 168248 3194
rect 168196 3130 168248 3136
rect 168288 3188 168340 3194
rect 168288 3130 168340 3136
rect 168208 480 168236 3130
rect 169404 480 169432 3946
rect 170600 480 170628 6530
rect 171060 5642 171088 320062
rect 171244 317490 171272 320076
rect 171612 317626 171640 320076
rect 171600 317620 171652 317626
rect 171600 317562 171652 317568
rect 171980 317558 172008 320076
rect 172440 317642 172468 320076
rect 172152 317620 172204 317626
rect 172152 317562 172204 317568
rect 172348 317614 172468 317642
rect 171968 317552 172020 317558
rect 171968 317494 172020 317500
rect 171232 317484 171284 317490
rect 171232 317426 171284 317432
rect 172164 16318 172192 317562
rect 172244 317484 172296 317490
rect 172244 317426 172296 317432
rect 172152 16312 172204 16318
rect 172152 16254 172204 16260
rect 172256 9722 172284 317426
rect 172348 9790 172376 317614
rect 172428 317552 172480 317558
rect 172428 317494 172480 317500
rect 172336 9784 172388 9790
rect 172336 9726 172388 9732
rect 172244 9716 172296 9722
rect 172244 9658 172296 9664
rect 172440 5710 172468 317494
rect 172808 317490 172836 320076
rect 173268 317558 173296 320076
rect 173650 320062 173756 320090
rect 173256 317552 173308 317558
rect 173256 317494 173308 317500
rect 172796 317484 172848 317490
rect 172796 317426 172848 317432
rect 173624 317484 173676 317490
rect 173624 317426 173676 317432
rect 173636 16250 173664 317426
rect 173624 16244 173676 16250
rect 173624 16186 173676 16192
rect 173728 9858 173756 320062
rect 174096 317558 174124 320076
rect 173808 317552 173860 317558
rect 173808 317494 173860 317500
rect 174084 317552 174136 317558
rect 174084 317494 174136 317500
rect 173716 9852 173768 9858
rect 173716 9794 173768 9800
rect 173820 5778 173848 317494
rect 174464 317490 174492 320076
rect 174938 320062 175044 320090
rect 174452 317484 174504 317490
rect 174452 317426 174504 317432
rect 175016 9926 175044 320062
rect 175188 317552 175240 317558
rect 175188 317494 175240 317500
rect 175096 317484 175148 317490
rect 175096 317426 175148 317432
rect 175004 9920 175056 9926
rect 175004 9862 175056 9868
rect 174176 6520 174228 6526
rect 174176 6462 174228 6468
rect 173808 5772 173860 5778
rect 173808 5714 173860 5720
rect 172428 5704 172480 5710
rect 172428 5646 172480 5652
rect 171048 5636 171100 5642
rect 171048 5578 171100 5584
rect 171782 4040 171838 4049
rect 171782 3975 171838 3984
rect 171796 480 171824 3975
rect 172980 3800 173032 3806
rect 172980 3742 173032 3748
rect 172992 480 173020 3742
rect 174188 480 174216 6462
rect 175108 5846 175136 317426
rect 175096 5840 175148 5846
rect 175096 5782 175148 5788
rect 175200 3330 175228 317494
rect 175292 317490 175320 320076
rect 175752 317558 175780 320076
rect 176134 320062 176424 320090
rect 175740 317552 175792 317558
rect 175740 317494 175792 317500
rect 175280 317484 175332 317490
rect 175280 317426 175332 317432
rect 176292 317484 176344 317490
rect 176292 317426 176344 317432
rect 176304 16182 176332 317426
rect 176292 16176 176344 16182
rect 176292 16118 176344 16124
rect 176396 9994 176424 320062
rect 176580 317642 176608 320076
rect 176488 317614 176608 317642
rect 176384 9988 176436 9994
rect 176384 9930 176436 9936
rect 176488 8498 176516 317614
rect 176568 317552 176620 317558
rect 176568 317494 176620 317500
rect 176476 8492 176528 8498
rect 176476 8434 176528 8440
rect 176580 5914 176608 317494
rect 176948 317490 176976 320076
rect 177408 317558 177436 320076
rect 177776 317762 177804 320076
rect 177764 317756 177816 317762
rect 177764 317698 177816 317704
rect 177396 317552 177448 317558
rect 177396 317494 177448 317500
rect 177856 317552 177908 317558
rect 177856 317494 177908 317500
rect 176936 317484 176988 317490
rect 176936 317426 176988 317432
rect 177868 10062 177896 317494
rect 178236 317490 178264 320076
rect 178604 317558 178632 320076
rect 179078 320062 179276 320090
rect 178592 317552 178644 317558
rect 178592 317494 178644 317500
rect 179052 317552 179104 317558
rect 179052 317494 179104 317500
rect 177948 317484 178000 317490
rect 177948 317426 178000 317432
rect 178224 317484 178276 317490
rect 178224 317426 178276 317432
rect 177856 10056 177908 10062
rect 177856 9998 177908 10004
rect 177764 6452 177816 6458
rect 177764 6394 177816 6400
rect 176568 5908 176620 5914
rect 176568 5850 176620 5856
rect 175370 3904 175426 3913
rect 175370 3839 175426 3848
rect 175188 3324 175240 3330
rect 175188 3266 175240 3272
rect 175384 480 175412 3839
rect 176568 3732 176620 3738
rect 176568 3674 176620 3680
rect 176580 480 176608 3674
rect 177776 480 177804 6394
rect 177960 5982 177988 317426
rect 179064 315738 179092 317494
rect 179144 317484 179196 317490
rect 179144 317426 179196 317432
rect 179156 315874 179184 317426
rect 179248 316010 179276 320062
rect 179432 317558 179460 320076
rect 179420 317552 179472 317558
rect 179420 317494 179472 317500
rect 179892 317490 179920 320076
rect 180260 317694 180288 320076
rect 180248 317688 180300 317694
rect 180720 317642 180748 320076
rect 180248 317630 180300 317636
rect 180628 317614 180748 317642
rect 179880 317484 179932 317490
rect 179880 317426 179932 317432
rect 180524 317484 180576 317490
rect 180524 317426 180576 317432
rect 179248 315982 179368 316010
rect 179156 315846 179276 315874
rect 179064 315710 179184 315738
rect 179156 10130 179184 315710
rect 179144 10124 179196 10130
rect 179144 10066 179196 10072
rect 179248 6050 179276 315846
rect 179236 6044 179288 6050
rect 179236 5986 179288 5992
rect 177948 5976 178000 5982
rect 177948 5918 178000 5924
rect 178958 3768 179014 3777
rect 179340 3738 179368 315982
rect 180536 10198 180564 317426
rect 180524 10192 180576 10198
rect 180524 10134 180576 10140
rect 180628 6866 180656 317614
rect 180708 317552 180760 317558
rect 180708 317494 180760 317500
rect 180616 6860 180668 6866
rect 180616 6802 180668 6808
rect 180720 6118 180748 317494
rect 181088 317490 181116 320076
rect 181562 320062 181760 320090
rect 181930 320062 182128 320090
rect 181076 317484 181128 317490
rect 181076 317426 181128 317432
rect 181628 317484 181680 317490
rect 181628 317426 181680 317432
rect 181640 315874 181668 317426
rect 181732 316010 181760 320062
rect 181732 315982 182036 316010
rect 181640 315846 181944 315874
rect 181916 10266 181944 315846
rect 181904 10260 181956 10266
rect 181904 10202 181956 10208
rect 182008 8566 182036 315982
rect 181996 8560 182048 8566
rect 181996 8502 182048 8508
rect 182100 6798 182128 320062
rect 182376 317490 182404 320076
rect 182744 317830 182772 320076
rect 183126 320062 183416 320090
rect 182732 317824 182784 317830
rect 182732 317766 182784 317772
rect 182364 317484 182416 317490
rect 182364 317426 182416 317432
rect 183192 317484 183244 317490
rect 183192 317426 183244 317432
rect 183204 315874 183232 317426
rect 183388 316010 183416 320062
rect 183572 317558 183600 320076
rect 183940 317626 183968 320076
rect 183928 317620 183980 317626
rect 183928 317562 183980 317568
rect 183560 317552 183612 317558
rect 183560 317494 183612 317500
rect 184400 317490 184428 320076
rect 184584 320062 184782 320090
rect 184388 317484 184440 317490
rect 184388 317426 184440 317432
rect 183388 315982 183508 316010
rect 183204 315846 183416 315874
rect 183388 11014 183416 315846
rect 183376 11008 183428 11014
rect 183376 10950 183428 10956
rect 182088 6792 182140 6798
rect 182088 6734 182140 6740
rect 183480 6730 183508 315982
rect 184584 10878 184612 320062
rect 185228 318578 185256 320076
rect 185216 318572 185268 318578
rect 185216 318514 185268 318520
rect 184848 317620 184900 317626
rect 184848 317562 184900 317568
rect 184664 317552 184716 317558
rect 184664 317494 184716 317500
rect 184676 10946 184704 317494
rect 184756 317484 184808 317490
rect 184756 317426 184808 317432
rect 184664 10940 184716 10946
rect 184664 10882 184716 10888
rect 184572 10872 184624 10878
rect 184572 10814 184624 10820
rect 183468 6724 183520 6730
rect 183468 6666 183520 6672
rect 184768 6662 184796 317426
rect 184756 6656 184808 6662
rect 184756 6598 184808 6604
rect 184860 6474 184888 317562
rect 185596 317490 185624 320076
rect 186070 320062 186176 320090
rect 185584 317484 185636 317490
rect 185584 317426 185636 317432
rect 186148 10810 186176 320062
rect 186424 317694 186452 320076
rect 186412 317688 186464 317694
rect 186412 317630 186464 317636
rect 186884 317490 186912 320076
rect 187266 320062 187464 320090
rect 186228 317484 186280 317490
rect 186228 317426 186280 317432
rect 186872 317484 186924 317490
rect 186872 317426 186924 317432
rect 186136 10804 186188 10810
rect 186136 10746 186188 10752
rect 186240 6594 186268 317426
rect 187436 10742 187464 320062
rect 187712 317762 187740 320076
rect 187700 317756 187752 317762
rect 187700 317698 187752 317704
rect 187608 317688 187660 317694
rect 187608 317630 187660 317636
rect 187516 317484 187568 317490
rect 187516 317426 187568 317432
rect 187424 10736 187476 10742
rect 187424 10678 187476 10684
rect 186228 6588 186280 6594
rect 186228 6530 186280 6536
rect 187528 6526 187556 317426
rect 184768 6446 184888 6474
rect 187516 6520 187568 6526
rect 187516 6462 187568 6468
rect 181352 6384 181404 6390
rect 181352 6326 181404 6332
rect 180708 6112 180760 6118
rect 180708 6054 180760 6060
rect 178958 3703 179014 3712
rect 179328 3732 179380 3738
rect 178972 480 179000 3703
rect 179328 3674 179380 3680
rect 180156 2916 180208 2922
rect 180156 2858 180208 2864
rect 180168 480 180196 2858
rect 181364 480 181392 6326
rect 184768 4146 184796 6446
rect 184848 6316 184900 6322
rect 184848 6258 184900 6264
rect 183744 4140 183796 4146
rect 183744 4082 183796 4088
rect 184756 4140 184808 4146
rect 184756 4082 184808 4088
rect 182548 3392 182600 3398
rect 182548 3334 182600 3340
rect 182560 480 182588 3334
rect 183756 480 183784 4082
rect 184860 480 184888 6258
rect 187620 4078 187648 317630
rect 188080 317490 188108 320076
rect 188554 320062 188660 320090
rect 188922 320062 189028 320090
rect 188068 317484 188120 317490
rect 188068 317426 188120 317432
rect 188632 316010 188660 320062
rect 188896 317484 188948 317490
rect 188896 317426 188948 317432
rect 188632 315982 188844 316010
rect 188816 10674 188844 315982
rect 188804 10668 188856 10674
rect 188804 10610 188856 10616
rect 188908 6458 188936 317426
rect 188896 6452 188948 6458
rect 188896 6394 188948 6400
rect 188436 6248 188488 6254
rect 188436 6190 188488 6196
rect 186044 4072 186096 4078
rect 186044 4014 186096 4020
rect 187608 4072 187660 4078
rect 187608 4014 187660 4020
rect 186056 480 186084 4014
rect 187240 3052 187292 3058
rect 187240 2994 187292 3000
rect 187252 480 187280 2994
rect 188448 480 188476 6190
rect 189000 3058 189028 320062
rect 189368 317490 189396 320076
rect 189736 317694 189764 320076
rect 190196 317966 190224 320076
rect 190184 317960 190236 317966
rect 190184 317902 190236 317908
rect 189724 317688 189776 317694
rect 189724 317630 189776 317636
rect 190276 317688 190328 317694
rect 190276 317630 190328 317636
rect 189356 317484 189408 317490
rect 189356 317426 189408 317432
rect 190288 10606 190316 317630
rect 190564 317490 190592 320076
rect 191024 317694 191052 320076
rect 191406 320062 191696 320090
rect 191012 317688 191064 317694
rect 191012 317630 191064 317636
rect 191564 317688 191616 317694
rect 191564 317630 191616 317636
rect 190368 317484 190420 317490
rect 190368 317426 190420 317432
rect 190552 317484 190604 317490
rect 190552 317426 190604 317432
rect 190276 10600 190328 10606
rect 190276 10542 190328 10548
rect 190380 6390 190408 317426
rect 191576 10538 191604 317630
rect 191564 10532 191616 10538
rect 191564 10474 191616 10480
rect 191668 8430 191696 320062
rect 191852 317694 191880 320076
rect 191840 317688 191892 317694
rect 191840 317630 191892 317636
rect 192220 317490 192248 320076
rect 192680 318782 192708 320076
rect 193062 320062 193168 320090
rect 192668 318776 192720 318782
rect 192668 318718 192720 318724
rect 193036 317688 193088 317694
rect 193036 317630 193088 317636
rect 191748 317484 191800 317490
rect 191748 317426 191800 317432
rect 192208 317484 192260 317490
rect 192208 317426 192260 317432
rect 192944 317484 192996 317490
rect 192944 317426 192996 317432
rect 191656 8424 191708 8430
rect 191656 8366 191708 8372
rect 190368 6384 190420 6390
rect 190368 6326 190420 6332
rect 191760 6322 191788 317426
rect 192956 10470 192984 317426
rect 192944 10464 192996 10470
rect 192944 10406 192996 10412
rect 191748 6316 191800 6322
rect 191748 6258 191800 6264
rect 193048 6254 193076 317630
rect 193036 6248 193088 6254
rect 193036 6190 193088 6196
rect 193140 6186 193168 320062
rect 193508 317490 193536 320076
rect 193772 317824 193824 317830
rect 193772 317766 193824 317772
rect 193784 317506 193812 317766
rect 193876 317694 193904 320076
rect 194258 320062 194456 320090
rect 193864 317688 193916 317694
rect 193864 317630 193916 317636
rect 193496 317484 193548 317490
rect 193784 317478 193996 317506
rect 193496 317426 193548 317432
rect 193968 309262 193996 317478
rect 194324 317484 194376 317490
rect 194324 317426 194376 317432
rect 193956 309256 194008 309262
rect 193956 309198 194008 309204
rect 193864 307828 193916 307834
rect 193864 307770 193916 307776
rect 193876 298110 193904 307770
rect 193864 298104 193916 298110
rect 193864 298046 193916 298052
rect 193864 288448 193916 288454
rect 193864 288390 193916 288396
rect 193876 278769 193904 288390
rect 193678 278760 193734 278769
rect 193678 278695 193734 278704
rect 193862 278760 193918 278769
rect 193862 278695 193918 278704
rect 193692 269142 193720 278695
rect 193680 269136 193732 269142
rect 193680 269078 193732 269084
rect 193864 269136 193916 269142
rect 193864 269078 193916 269084
rect 193876 259457 193904 269078
rect 193678 259448 193734 259457
rect 193678 259383 193734 259392
rect 193862 259448 193918 259457
rect 193862 259383 193918 259392
rect 193692 249830 193720 259383
rect 193680 249824 193732 249830
rect 193680 249766 193732 249772
rect 193864 249824 193916 249830
rect 193864 249766 193916 249772
rect 193876 241777 193904 249766
rect 193862 241768 193918 241777
rect 193862 241703 193918 241712
rect 193862 241632 193918 241641
rect 193862 241567 193918 241576
rect 193876 240145 193904 241567
rect 193678 240136 193734 240145
rect 193678 240071 193734 240080
rect 193862 240136 193918 240145
rect 193862 240071 193918 240080
rect 193692 230518 193720 240071
rect 193680 230512 193732 230518
rect 193680 230454 193732 230460
rect 193864 230512 193916 230518
rect 193864 230454 193916 230460
rect 193876 220833 193904 230454
rect 193678 220824 193734 220833
rect 193678 220759 193734 220768
rect 193862 220824 193918 220833
rect 193862 220759 193918 220768
rect 193692 211177 193720 220759
rect 193678 211168 193734 211177
rect 193678 211103 193734 211112
rect 193862 211168 193918 211177
rect 193862 211103 193918 211112
rect 193876 201482 193904 211103
rect 193680 201476 193732 201482
rect 193680 201418 193732 201424
rect 193864 201476 193916 201482
rect 193864 201418 193916 201424
rect 193692 191865 193720 201418
rect 193678 191856 193734 191865
rect 193678 191791 193734 191800
rect 193862 191856 193918 191865
rect 193862 191791 193918 191800
rect 193876 182170 193904 191791
rect 193680 182164 193732 182170
rect 193680 182106 193732 182112
rect 193864 182164 193916 182170
rect 193864 182106 193916 182112
rect 193692 172553 193720 182106
rect 193678 172544 193734 172553
rect 193678 172479 193734 172488
rect 193862 172544 193918 172553
rect 193862 172479 193918 172488
rect 193876 162858 193904 172479
rect 193864 162852 193916 162858
rect 193864 162794 193916 162800
rect 193864 153264 193916 153270
rect 193864 153206 193916 153212
rect 193876 143546 193904 153206
rect 193864 143540 193916 143546
rect 193864 143482 193916 143488
rect 193864 133952 193916 133958
rect 193864 133894 193916 133900
rect 193876 124166 193904 133894
rect 193864 124160 193916 124166
rect 193864 124102 193916 124108
rect 193864 114572 193916 114578
rect 193864 114514 193916 114520
rect 193876 104854 193904 114514
rect 193864 104848 193916 104854
rect 193864 104790 193916 104796
rect 193864 95260 193916 95266
rect 193864 95202 193916 95208
rect 193876 85542 193904 95202
rect 193864 85536 193916 85542
rect 193864 85478 193916 85484
rect 193864 75948 193916 75954
rect 193864 75890 193916 75896
rect 193876 66230 193904 75890
rect 193864 66224 193916 66230
rect 193864 66166 193916 66172
rect 193864 56636 193916 56642
rect 193864 56578 193916 56584
rect 193876 46918 193904 56578
rect 193864 46912 193916 46918
rect 193864 46854 193916 46860
rect 193956 29028 194008 29034
rect 193956 28970 194008 28976
rect 193968 22114 193996 28970
rect 193784 22086 193996 22114
rect 193784 19310 193812 22086
rect 193772 19304 193824 19310
rect 193772 19246 193824 19252
rect 193772 12436 193824 12442
rect 193772 12378 193824 12384
rect 193784 9738 193812 12378
rect 194336 10402 194364 317426
rect 194324 10396 194376 10402
rect 194324 10338 194376 10344
rect 193784 9710 193904 9738
rect 192024 6180 192076 6186
rect 192024 6122 192076 6128
rect 193128 6180 193180 6186
rect 193128 6122 193180 6128
rect 190828 3936 190880 3942
rect 190828 3878 190880 3884
rect 188988 3052 189040 3058
rect 188988 2994 189040 3000
rect 189632 2848 189684 2854
rect 189632 2790 189684 2796
rect 189644 480 189672 2790
rect 190840 480 190868 3878
rect 192036 480 192064 6122
rect 193876 4214 193904 9710
rect 194428 6769 194456 320062
rect 194704 317694 194732 320076
rect 195072 318646 195100 320076
rect 195060 318640 195112 318646
rect 195060 318582 195112 318588
rect 194508 317688 194560 317694
rect 194508 317630 194560 317636
rect 194692 317688 194744 317694
rect 194692 317630 194744 317636
rect 194414 6760 194470 6769
rect 194414 6695 194470 6704
rect 193864 4208 193916 4214
rect 193864 4150 193916 4156
rect 194520 3942 194548 317630
rect 195532 317490 195560 320076
rect 195716 320062 195914 320090
rect 195520 317484 195572 317490
rect 195520 317426 195572 317432
rect 195716 10849 195744 320062
rect 196360 317762 196388 320076
rect 196348 317756 196400 317762
rect 196348 317698 196400 317704
rect 195796 317688 195848 317694
rect 195796 317630 195848 317636
rect 195702 10840 195758 10849
rect 195702 10775 195758 10784
rect 195808 10334 195836 317630
rect 196728 317490 196756 320076
rect 197188 317914 197216 320076
rect 197556 318714 197584 320076
rect 197544 318708 197596 318714
rect 197544 318650 197596 318656
rect 197096 317886 197216 317914
rect 195888 317484 195940 317490
rect 195888 317426 195940 317432
rect 196716 317484 196768 317490
rect 196716 317426 196768 317432
rect 195796 10328 195848 10334
rect 195796 10270 195848 10276
rect 195900 6633 195928 317426
rect 197096 10713 197124 317886
rect 197176 317756 197228 317762
rect 197176 317698 197228 317704
rect 197082 10704 197138 10713
rect 197082 10639 197138 10648
rect 197188 8634 197216 317698
rect 198016 317490 198044 320076
rect 198398 320062 198596 320090
rect 197268 317484 197320 317490
rect 197268 317426 197320 317432
rect 198004 317484 198056 317490
rect 198004 317426 198056 317432
rect 197176 8628 197228 8634
rect 197176 8570 197228 8576
rect 195886 6624 195942 6633
rect 195886 6559 195942 6568
rect 197280 6497 197308 317426
rect 198004 309188 198056 309194
rect 198004 309130 198056 309136
rect 198016 7070 198044 309130
rect 198568 10577 198596 320062
rect 198844 317762 198872 320076
rect 198832 317756 198884 317762
rect 198832 317698 198884 317704
rect 199212 317490 199240 320076
rect 199686 320062 199884 320090
rect 198648 317484 198700 317490
rect 198648 317426 198700 317432
rect 199200 317484 199252 317490
rect 199200 317426 199252 317432
rect 198554 10568 198610 10577
rect 198554 10503 198610 10512
rect 198004 7064 198056 7070
rect 198004 7006 198056 7012
rect 197266 6488 197322 6497
rect 197266 6423 197322 6432
rect 198660 6361 198688 317426
rect 199856 10441 199884 320062
rect 200040 318306 200068 320076
rect 200028 318300 200080 318306
rect 200028 318242 200080 318248
rect 200028 317756 200080 317762
rect 200028 317698 200080 317704
rect 199936 317484 199988 317490
rect 199936 317426 199988 317432
rect 199842 10432 199898 10441
rect 199842 10367 199898 10376
rect 198646 6352 198702 6361
rect 198646 6287 198702 6296
rect 199948 6225 199976 317426
rect 199934 6216 199990 6225
rect 199934 6151 199990 6160
rect 198004 4276 198056 4282
rect 198004 4218 198056 4224
rect 194508 3936 194560 3942
rect 194508 3878 194560 3884
rect 194416 3868 194468 3874
rect 194416 3810 194468 3816
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 193232 480 193260 3470
rect 194428 480 194456 3810
rect 195612 3120 195664 3126
rect 195612 3062 195664 3068
rect 195624 480 195652 3062
rect 196808 2984 196860 2990
rect 196808 2926 196860 2932
rect 196820 480 196848 2926
rect 198016 480 198044 4218
rect 200040 3874 200068 317698
rect 200500 317490 200528 320076
rect 200882 320062 201172 320090
rect 201342 320062 201448 320090
rect 201144 317642 201172 320062
rect 201144 317614 201356 317642
rect 200488 317484 200540 317490
rect 200488 317426 200540 317432
rect 201224 317484 201276 317490
rect 201224 317426 201276 317432
rect 201236 14414 201264 317426
rect 201224 14408 201276 14414
rect 201224 14350 201276 14356
rect 201328 10305 201356 317614
rect 201314 10296 201370 10305
rect 201314 10231 201370 10240
rect 200028 3868 200080 3874
rect 200028 3810 200080 3816
rect 201420 3806 201448 320062
rect 201696 317490 201724 320076
rect 202156 318714 202184 320076
rect 202144 318708 202196 318714
rect 202144 318650 202196 318656
rect 202524 318374 202552 320076
rect 202696 318708 202748 318714
rect 202696 318650 202748 318656
rect 202512 318368 202564 318374
rect 202512 318310 202564 318316
rect 202144 318028 202196 318034
rect 202144 317970 202196 317976
rect 201684 317484 201736 317490
rect 201684 317426 201736 317432
rect 201500 4344 201552 4350
rect 201500 4286 201552 4292
rect 201408 3800 201460 3806
rect 201408 3742 201460 3748
rect 199200 3664 199252 3670
rect 199200 3606 199252 3612
rect 199212 480 199240 3606
rect 200396 3460 200448 3466
rect 200396 3402 200448 3408
rect 200408 480 200436 3402
rect 201512 480 201540 4286
rect 202156 4282 202184 317970
rect 202708 15026 202736 318650
rect 202984 317762 203012 320076
rect 203352 318034 203380 320076
rect 203340 318028 203392 318034
rect 203340 317970 203392 317976
rect 202972 317756 203024 317762
rect 202972 317698 203024 317704
rect 203812 317490 203840 320076
rect 203996 320062 204194 320090
rect 203892 318028 203944 318034
rect 203892 317970 203944 317976
rect 202788 317484 202840 317490
rect 202788 317426 202840 317432
rect 203800 317484 203852 317490
rect 203800 317426 203852 317432
rect 202800 15162 202828 317426
rect 202788 15156 202840 15162
rect 202788 15098 202840 15104
rect 202696 15020 202748 15026
rect 202696 14962 202748 14968
rect 203904 14958 203932 317970
rect 203892 14952 203944 14958
rect 203892 14894 203944 14900
rect 203996 14822 204024 320062
rect 204076 317756 204128 317762
rect 204076 317698 204128 317704
rect 204088 15094 204116 317698
rect 204640 317490 204668 320076
rect 205008 318782 205036 320076
rect 205390 320062 205588 320090
rect 204996 318776 205048 318782
rect 204996 318718 205048 318724
rect 204168 317484 204220 317490
rect 204168 317426 204220 317432
rect 204628 317484 204680 317490
rect 204628 317426 204680 317432
rect 205456 317484 205508 317490
rect 205456 317426 205508 317432
rect 204076 15088 204128 15094
rect 204076 15030 204128 15036
rect 203984 14816 204036 14822
rect 203984 14758 204036 14764
rect 202696 8016 202748 8022
rect 202696 7958 202748 7964
rect 202144 4276 202196 4282
rect 202144 4218 202196 4224
rect 202708 480 202736 7958
rect 204180 3738 204208 317426
rect 204904 309188 204956 309194
rect 204904 309130 204956 309136
rect 204916 183666 204944 309130
rect 204904 183660 204956 183666
rect 204904 183602 204956 183608
rect 204720 183592 204772 183598
rect 204720 183534 204772 183540
rect 204732 173942 204760 183534
rect 204720 173936 204772 173942
rect 204720 173878 204772 173884
rect 204904 173936 204956 173942
rect 204904 173878 204956 173884
rect 204916 164150 204944 173878
rect 204812 164144 204864 164150
rect 204812 164086 204864 164092
rect 204904 164144 204956 164150
rect 204904 164086 204956 164092
rect 204824 154737 204852 164086
rect 204810 154728 204866 154737
rect 204810 154663 204866 154672
rect 204902 154592 204958 154601
rect 204902 154527 204958 154536
rect 204916 144838 204944 154527
rect 204812 144832 204864 144838
rect 204812 144774 204864 144780
rect 204904 144832 204956 144838
rect 204904 144774 204956 144780
rect 204824 135425 204852 144774
rect 204810 135416 204866 135425
rect 204810 135351 204866 135360
rect 204902 135280 204958 135289
rect 204902 135215 204958 135224
rect 204916 130370 204944 135215
rect 204916 130342 205036 130370
rect 205008 125610 205036 130342
rect 205008 125582 205128 125610
rect 205100 116006 205128 125582
rect 204904 116000 204956 116006
rect 204904 115942 204956 115948
rect 205088 116000 205140 116006
rect 205088 115942 205140 115948
rect 204916 106350 204944 115942
rect 204720 106344 204772 106350
rect 204720 106286 204772 106292
rect 204904 106344 204956 106350
rect 204904 106286 204956 106292
rect 204732 96694 204760 106286
rect 204720 96688 204772 96694
rect 204720 96630 204772 96636
rect 204904 96688 204956 96694
rect 204904 96630 204956 96636
rect 204916 87038 204944 96630
rect 204720 87032 204772 87038
rect 204720 86974 204772 86980
rect 204904 87032 204956 87038
rect 204904 86974 204956 86980
rect 204732 85542 204760 86974
rect 204720 85536 204772 85542
rect 204720 85478 204772 85484
rect 204904 75948 204956 75954
rect 204904 75890 204956 75896
rect 204916 66230 204944 75890
rect 204904 66224 204956 66230
rect 204904 66166 204956 66172
rect 204904 56636 204956 56642
rect 204904 56578 204956 56584
rect 204916 46918 204944 56578
rect 204904 46912 204956 46918
rect 204904 46854 204956 46860
rect 204904 37324 204956 37330
rect 204904 37266 204956 37272
rect 204916 27606 204944 37266
rect 204904 27600 204956 27606
rect 204904 27542 204956 27548
rect 204904 18012 204956 18018
rect 204904 17954 204956 17960
rect 204916 9738 204944 17954
rect 205468 14890 205496 317426
rect 205456 14884 205508 14890
rect 205456 14826 205508 14832
rect 204824 9710 204944 9738
rect 204824 7070 204852 9710
rect 205560 7070 205588 320062
rect 205836 317490 205864 320076
rect 206204 318034 206232 320076
rect 206678 320062 206876 320090
rect 206192 318028 206244 318034
rect 206192 317970 206244 317976
rect 206652 318028 206704 318034
rect 206652 317970 206704 317976
rect 205824 317484 205876 317490
rect 205824 317426 205876 317432
rect 206664 315738 206692 317970
rect 206744 317484 206796 317490
rect 206744 317426 206796 317432
rect 206756 315874 206784 317426
rect 206848 316010 206876 320062
rect 207032 317490 207060 320076
rect 207492 318034 207520 320076
rect 207874 320062 208164 320090
rect 207848 318096 207900 318102
rect 207848 318038 207900 318044
rect 207480 318028 207532 318034
rect 207480 317970 207532 317976
rect 207020 317484 207072 317490
rect 207020 317426 207072 317432
rect 206848 315982 206968 316010
rect 206756 315846 206876 315874
rect 206664 315710 206784 315738
rect 206756 16114 206784 315710
rect 206744 16108 206796 16114
rect 206744 16050 206796 16056
rect 206848 14754 206876 315846
rect 206836 14748 206888 14754
rect 206836 14690 206888 14696
rect 205640 8832 205692 8838
rect 205638 8800 205640 8809
rect 205692 8800 205694 8809
rect 205638 8735 205694 8744
rect 206284 7948 206336 7954
rect 206284 7890 206336 7896
rect 204812 7064 204864 7070
rect 204812 7006 204864 7012
rect 205548 7064 205600 7070
rect 205548 7006 205600 7012
rect 205088 4412 205140 4418
rect 205088 4354 205140 4360
rect 204168 3732 204220 3738
rect 204168 3674 204220 3680
rect 203892 3188 203944 3194
rect 203892 3130 203944 3136
rect 203904 480 203932 3130
rect 205100 480 205128 4354
rect 206296 480 206324 7890
rect 206940 7138 206968 315982
rect 207860 315738 207888 318038
rect 208032 317484 208084 317490
rect 208032 317426 208084 317432
rect 208044 315874 208072 317426
rect 208136 316010 208164 320062
rect 208320 318102 208348 320076
rect 208688 318782 208716 320076
rect 208676 318776 208728 318782
rect 208676 318718 208728 318724
rect 209044 318436 209096 318442
rect 209044 318378 209096 318384
rect 208308 318096 208360 318102
rect 208308 318038 208360 318044
rect 208216 318028 208268 318034
rect 208216 317970 208268 317976
rect 208228 316146 208256 317970
rect 208228 316118 208348 316146
rect 208136 315982 208256 316010
rect 208044 315846 208164 315874
rect 207860 315710 208072 315738
rect 208044 11286 208072 315710
rect 208032 11280 208084 11286
rect 208032 11222 208084 11228
rect 208136 11218 208164 315846
rect 208124 11212 208176 11218
rect 208124 11154 208176 11160
rect 208228 7206 208256 315982
rect 208216 7200 208268 7206
rect 208216 7142 208268 7148
rect 206928 7132 206980 7138
rect 206928 7074 206980 7080
rect 208320 3670 208348 316118
rect 209056 4486 209084 318378
rect 209148 317490 209176 320076
rect 209530 320062 209636 320090
rect 209136 317484 209188 317490
rect 209136 317426 209188 317432
rect 209608 11354 209636 320062
rect 209976 318442 210004 320076
rect 209964 318436 210016 318442
rect 209964 318378 210016 318384
rect 210344 317490 210372 320076
rect 210818 320062 211016 320090
rect 209688 317484 209740 317490
rect 209688 317426 209740 317432
rect 210332 317484 210384 317490
rect 210332 317426 210384 317432
rect 209596 11348 209648 11354
rect 209596 11290 209648 11296
rect 209700 7274 209728 317426
rect 210988 11422 211016 320062
rect 211172 317490 211200 320076
rect 211632 318034 211660 320076
rect 212014 320062 212304 320090
rect 211988 318164 212040 318170
rect 211988 318106 212040 318112
rect 211620 318028 211672 318034
rect 211620 317970 211672 317976
rect 211068 317484 211120 317490
rect 211068 317426 211120 317432
rect 211160 317484 211212 317490
rect 211160 317426 211212 317432
rect 210976 11416 211028 11422
rect 210976 11358 211028 11364
rect 209872 7880 209924 7886
rect 209872 7822 209924 7828
rect 209688 7268 209740 7274
rect 209688 7210 209740 7216
rect 208676 4480 208728 4486
rect 208676 4422 208728 4428
rect 209044 4480 209096 4486
rect 209044 4422 209096 4428
rect 208308 3664 208360 3670
rect 207478 3632 207534 3641
rect 208308 3606 208360 3612
rect 207478 3567 207534 3576
rect 207492 480 207520 3567
rect 208688 480 208716 4422
rect 209884 480 209912 7822
rect 211080 7342 211108 317426
rect 212000 302258 212028 318106
rect 212080 317484 212132 317490
rect 212080 317426 212132 317432
rect 212092 315874 212120 317426
rect 212276 316010 212304 320062
rect 212460 318442 212488 320076
rect 212448 318436 212500 318442
rect 212448 318378 212500 318384
rect 212448 318028 212500 318034
rect 212448 317970 212500 317976
rect 212276 315982 212396 316010
rect 212092 315846 212304 315874
rect 211804 302252 211856 302258
rect 211804 302194 211856 302200
rect 211988 302252 212040 302258
rect 211988 302194 212040 302200
rect 211816 302138 211844 302194
rect 211816 302110 211936 302138
rect 211908 292618 211936 302110
rect 211908 292590 212028 292618
rect 212000 282946 212028 292590
rect 211804 282940 211856 282946
rect 211804 282882 211856 282888
rect 211988 282940 212040 282946
rect 211988 282882 212040 282888
rect 211816 282826 211844 282882
rect 211816 282798 211936 282826
rect 211908 273306 211936 282798
rect 211908 273278 212028 273306
rect 212000 263634 212028 273278
rect 211804 263628 211856 263634
rect 211804 263570 211856 263576
rect 211988 263628 212040 263634
rect 211988 263570 212040 263576
rect 211816 263514 211844 263570
rect 211816 263486 211936 263514
rect 211908 253994 211936 263486
rect 211908 253966 212028 253994
rect 212000 244322 212028 253966
rect 211804 244316 211856 244322
rect 211804 244258 211856 244264
rect 211988 244316 212040 244322
rect 211988 244258 212040 244264
rect 211816 244202 211844 244258
rect 211816 244174 211936 244202
rect 211908 234682 211936 244174
rect 211908 234654 212028 234682
rect 212000 225010 212028 234654
rect 211804 225004 211856 225010
rect 211804 224946 211856 224952
rect 211988 225004 212040 225010
rect 211988 224946 212040 224952
rect 211816 224890 211844 224946
rect 211816 224862 211936 224890
rect 211908 215370 211936 224862
rect 211908 215342 212028 215370
rect 212000 205698 212028 215342
rect 211804 205692 211856 205698
rect 211804 205634 211856 205640
rect 211988 205692 212040 205698
rect 211988 205634 212040 205640
rect 211816 205578 211844 205634
rect 211816 205550 211936 205578
rect 211908 196058 211936 205550
rect 211908 196030 212028 196058
rect 212000 186386 212028 196030
rect 211804 186380 211856 186386
rect 211804 186322 211856 186328
rect 211988 186380 212040 186386
rect 211988 186322 212040 186328
rect 211816 186266 211844 186322
rect 211816 186238 211936 186266
rect 211908 183569 211936 186238
rect 211710 183560 211766 183569
rect 211710 183495 211766 183504
rect 211894 183560 211950 183569
rect 211894 183495 211950 183504
rect 211724 173942 211752 183495
rect 211712 173936 211764 173942
rect 211712 173878 211764 173884
rect 211988 173936 212040 173942
rect 211988 173878 212040 173884
rect 212000 167074 212028 173878
rect 211804 167068 211856 167074
rect 211804 167010 211856 167016
rect 211988 167068 212040 167074
rect 211988 167010 212040 167016
rect 211816 166954 211844 167010
rect 211816 166926 211936 166954
rect 211908 164218 211936 166926
rect 211896 164212 211948 164218
rect 211896 164154 211948 164160
rect 211896 157344 211948 157350
rect 211896 157286 211948 157292
rect 211908 154578 211936 157286
rect 211908 154550 212028 154578
rect 212000 147694 212028 154550
rect 211804 147688 211856 147694
rect 211988 147688 212040 147694
rect 211856 147636 211936 147642
rect 211804 147630 211936 147636
rect 211988 147630 212040 147636
rect 211816 147614 211936 147630
rect 211908 144906 211936 147614
rect 211896 144900 211948 144906
rect 211896 144842 211948 144848
rect 211896 137964 211948 137970
rect 211896 137906 211948 137912
rect 211908 135266 211936 137906
rect 211908 135238 212028 135266
rect 212000 128382 212028 135238
rect 211804 128376 211856 128382
rect 211988 128376 212040 128382
rect 211856 128324 211936 128330
rect 211804 128318 211936 128324
rect 211988 128318 212040 128324
rect 211816 128302 211936 128318
rect 211908 125594 211936 128302
rect 211896 125588 211948 125594
rect 211896 125530 211948 125536
rect 211896 118652 211948 118658
rect 211896 118594 211948 118600
rect 211908 115954 211936 118594
rect 211908 115926 212028 115954
rect 212000 109070 212028 115926
rect 211804 109064 211856 109070
rect 211988 109064 212040 109070
rect 211856 109012 211936 109018
rect 211804 109006 211936 109012
rect 211988 109006 212040 109012
rect 211816 108990 211936 109006
rect 211908 106282 211936 108990
rect 211896 106276 211948 106282
rect 211896 106218 211948 106224
rect 211896 99340 211948 99346
rect 211896 99282 211948 99288
rect 211908 96642 211936 99282
rect 211908 96614 212028 96642
rect 212000 89758 212028 96614
rect 211804 89752 211856 89758
rect 211988 89752 212040 89758
rect 211856 89700 211936 89706
rect 211804 89694 211936 89700
rect 211988 89694 212040 89700
rect 211816 89678 211936 89694
rect 211908 86970 211936 89678
rect 211896 86964 211948 86970
rect 211896 86906 211948 86912
rect 211988 77308 212040 77314
rect 211988 77250 212040 77256
rect 212000 75886 212028 77250
rect 211988 75880 212040 75886
rect 211988 75822 212040 75828
rect 211896 70372 211948 70378
rect 211896 70314 211948 70320
rect 211908 60738 211936 70314
rect 211908 60710 212028 60738
rect 212000 57934 212028 60710
rect 211988 57928 212040 57934
rect 211988 57870 212040 57876
rect 211896 50720 211948 50726
rect 211896 50662 211948 50668
rect 211908 41426 211936 50662
rect 211908 41398 212028 41426
rect 212000 38622 212028 41398
rect 211988 38616 212040 38622
rect 211988 38558 212040 38564
rect 211896 29028 211948 29034
rect 211896 28970 211948 28976
rect 211908 22114 211936 28970
rect 211908 22086 212028 22114
rect 212000 12458 212028 22086
rect 212276 16046 212304 315846
rect 212264 16040 212316 16046
rect 212264 15982 212316 15988
rect 211816 12430 212028 12458
rect 211068 7336 211120 7342
rect 211068 7278 211120 7284
rect 211816 4486 211844 12430
rect 212368 11490 212396 315982
rect 212356 11484 212408 11490
rect 212356 11426 212408 11432
rect 212460 7410 212488 317970
rect 212828 317490 212856 320076
rect 213288 318034 213316 320076
rect 213670 320062 213868 320090
rect 213276 318028 213328 318034
rect 213276 317970 213328 317976
rect 213644 318028 213696 318034
rect 213644 317970 213696 317976
rect 212816 317484 212868 317490
rect 212816 317426 212868 317432
rect 213656 11558 213684 317970
rect 213736 317484 213788 317490
rect 213736 317426 213788 317432
rect 213644 11552 213696 11558
rect 213644 11494 213696 11500
rect 213460 7812 213512 7818
rect 213460 7754 213512 7760
rect 212448 7404 212500 7410
rect 212448 7346 212500 7352
rect 212264 4548 212316 4554
rect 212264 4490 212316 4496
rect 211804 4480 211856 4486
rect 211804 4422 211856 4428
rect 211068 3596 211120 3602
rect 211068 3538 211120 3544
rect 211080 480 211108 3538
rect 212276 480 212304 4490
rect 213472 480 213500 7754
rect 213748 7478 213776 317426
rect 213736 7472 213788 7478
rect 213736 7414 213788 7420
rect 213840 3602 213868 320062
rect 214116 318034 214144 320076
rect 214484 318714 214512 320076
rect 214944 318782 214972 320076
rect 214932 318776 214984 318782
rect 214932 318718 214984 318724
rect 214472 318708 214524 318714
rect 214472 318650 214524 318656
rect 215116 318708 215168 318714
rect 215116 318650 215168 318656
rect 214104 318028 214156 318034
rect 214104 317970 214156 317976
rect 215128 11626 215156 318650
rect 215312 318170 215340 320076
rect 215300 318164 215352 318170
rect 215300 318106 215352 318112
rect 215772 318034 215800 320076
rect 216154 320062 216352 320090
rect 216522 320062 216628 320090
rect 215944 318504 215996 318510
rect 215944 318446 215996 318452
rect 215208 318028 215260 318034
rect 215208 317970 215260 317976
rect 215760 318028 215812 318034
rect 215760 317970 215812 317976
rect 215116 11620 215168 11626
rect 215116 11562 215168 11568
rect 215116 8832 215168 8838
rect 215114 8800 215116 8809
rect 215168 8800 215170 8809
rect 215114 8735 215170 8744
rect 215220 7546 215248 317970
rect 215208 7540 215260 7546
rect 215208 7482 215260 7488
rect 215116 4820 215168 4826
rect 215116 4762 215168 4768
rect 215576 4820 215628 4826
rect 215576 4762 215628 4768
rect 215128 4729 215156 4762
rect 215588 4729 215616 4762
rect 215114 4720 215170 4729
rect 215114 4655 215170 4664
rect 215574 4720 215630 4729
rect 215574 4655 215630 4664
rect 215852 4616 215904 4622
rect 215852 4558 215904 4564
rect 215116 4548 215168 4554
rect 215116 4490 215168 4496
rect 215128 4457 215156 4490
rect 215300 4480 215352 4486
rect 215114 4448 215170 4457
rect 215114 4383 215170 4392
rect 215298 4448 215300 4457
rect 215352 4448 215354 4457
rect 215298 4383 215354 4392
rect 213828 3596 213880 3602
rect 213828 3538 213880 3544
rect 214654 3360 214710 3369
rect 214654 3295 214710 3304
rect 214668 480 214696 3295
rect 215864 480 215892 4558
rect 215956 4536 215984 318446
rect 216324 15978 216352 320062
rect 216496 318164 216548 318170
rect 216496 318106 216548 318112
rect 216404 318028 216456 318034
rect 216404 317970 216456 317976
rect 216312 15972 216364 15978
rect 216312 15914 216364 15920
rect 216416 11694 216444 317970
rect 216404 11688 216456 11694
rect 216404 11630 216456 11636
rect 216508 8294 216536 318106
rect 216496 8288 216548 8294
rect 216496 8230 216548 8236
rect 216600 8226 216628 320062
rect 216968 318034 216996 320076
rect 217336 318510 217364 320076
rect 217810 320062 218008 320090
rect 217324 318504 217376 318510
rect 217324 318446 217376 318452
rect 216956 318028 217008 318034
rect 216956 317970 217008 317976
rect 217876 318028 217928 318034
rect 217876 317970 217928 317976
rect 217888 12442 217916 317970
rect 217876 12436 217928 12442
rect 217876 12378 217928 12384
rect 216588 8220 216640 8226
rect 216588 8162 216640 8168
rect 217980 8158 218008 320062
rect 218164 318034 218192 320076
rect 218624 318170 218652 320076
rect 219006 320062 219296 320090
rect 218704 318232 218756 318238
rect 218704 318174 218756 318180
rect 218612 318164 218664 318170
rect 218612 318106 218664 318112
rect 218152 318028 218204 318034
rect 218152 317970 218204 317976
rect 217968 8152 218020 8158
rect 217968 8094 218020 8100
rect 218716 7954 218744 318174
rect 219164 318028 219216 318034
rect 219164 317970 219216 317976
rect 219072 16584 219124 16590
rect 219072 16526 219124 16532
rect 218704 7948 218756 7954
rect 218704 7890 218756 7896
rect 219084 7834 219112 16526
rect 219176 12374 219204 317970
rect 219164 12368 219216 12374
rect 219164 12310 219216 12316
rect 219268 8090 219296 320062
rect 219348 318164 219400 318170
rect 219348 318106 219400 318112
rect 219360 16590 219388 318106
rect 219452 318034 219480 320076
rect 219834 320062 220124 320090
rect 220096 318764 220124 320062
rect 220176 318776 220228 318782
rect 220096 318736 220176 318764
rect 220176 318718 220228 318724
rect 220280 318170 220308 320076
rect 220268 318164 220320 318170
rect 220268 318106 220320 318112
rect 219440 318028 219492 318034
rect 219440 317970 219492 317976
rect 220544 318028 220596 318034
rect 220544 317970 220596 317976
rect 219348 16584 219400 16590
rect 219348 16526 219400 16532
rect 220556 12306 220584 317970
rect 220544 12300 220596 12306
rect 220544 12242 220596 12248
rect 220648 12238 220676 320076
rect 221108 318170 221136 320076
rect 220728 318164 220780 318170
rect 220728 318106 220780 318112
rect 221096 318164 221148 318170
rect 221096 318106 221148 318112
rect 220636 12232 220688 12238
rect 220636 12174 220688 12180
rect 219256 8084 219308 8090
rect 219256 8026 219308 8032
rect 220740 8022 220768 318106
rect 221476 318034 221504 320076
rect 221464 318028 221516 318034
rect 221464 317970 221516 317976
rect 221936 12170 221964 320076
rect 222304 318714 222332 320076
rect 222292 318708 222344 318714
rect 222292 318650 222344 318656
rect 222108 318164 222160 318170
rect 222108 318106 222160 318112
rect 222016 318028 222068 318034
rect 222016 317970 222068 317976
rect 221924 12164 221976 12170
rect 221924 12106 221976 12112
rect 220728 8016 220780 8022
rect 220728 7958 220780 7964
rect 222028 7954 222056 317970
rect 219256 7948 219308 7954
rect 219256 7890 219308 7896
rect 222016 7948 222068 7954
rect 222016 7890 222068 7896
rect 219084 7806 219204 7834
rect 217048 7744 217100 7750
rect 217048 7686 217100 7692
rect 216036 4548 216088 4554
rect 215956 4508 216036 4536
rect 216036 4490 216088 4496
rect 217060 480 217088 7686
rect 218980 4684 219032 4690
rect 218980 4626 219032 4632
rect 218150 3496 218206 3505
rect 218150 3431 218206 3440
rect 218164 480 218192 3431
rect 218992 3346 219020 4626
rect 219176 3534 219204 7806
rect 219268 4690 219296 7890
rect 220544 7676 220596 7682
rect 220544 7618 220596 7624
rect 219256 4684 219308 4690
rect 219256 4626 219308 4632
rect 219164 3528 219216 3534
rect 219164 3470 219216 3476
rect 218992 3318 219388 3346
rect 219360 480 219388 3318
rect 220556 480 220584 7618
rect 222120 3466 222148 318106
rect 222764 318034 222792 320076
rect 223146 320062 223436 320090
rect 223606 320062 223712 320090
rect 222752 318028 222804 318034
rect 222752 317970 222804 317976
rect 223408 12102 223436 320062
rect 223488 318028 223540 318034
rect 223488 317970 223540 317976
rect 223396 12096 223448 12102
rect 223396 12038 223448 12044
rect 223500 7886 223528 317970
rect 223684 311234 223712 320062
rect 223960 318034 223988 320076
rect 224434 320062 224540 320090
rect 223948 318028 224000 318034
rect 223948 317970 224000 317976
rect 224512 316010 224540 320062
rect 224788 318238 224816 320076
rect 224972 320062 225262 320090
rect 225630 320062 225828 320090
rect 226090 320062 226288 320090
rect 224776 318232 224828 318238
rect 224776 318174 224828 318180
rect 224776 318028 224828 318034
rect 224776 317970 224828 317976
rect 224512 315982 224724 316010
rect 223672 311228 223724 311234
rect 223672 311170 223724 311176
rect 224696 12034 224724 315982
rect 224684 12028 224736 12034
rect 224684 11970 224736 11976
rect 223488 7880 223540 7886
rect 223488 7822 223540 7828
rect 224788 7818 224816 317970
rect 224868 311228 224920 311234
rect 224868 311170 224920 311176
rect 224776 7812 224828 7818
rect 224776 7754 224828 7760
rect 224132 7608 224184 7614
rect 224132 7550 224184 7556
rect 222936 4616 222988 4622
rect 222936 4558 222988 4564
rect 222108 3460 222160 3466
rect 222108 3402 222160 3408
rect 221740 3256 221792 3262
rect 221740 3198 221792 3204
rect 221752 480 221780 3198
rect 222948 480 222976 4558
rect 224144 480 224172 7550
rect 224880 3913 224908 311170
rect 224972 307086 225000 320062
rect 225800 316010 225828 320062
rect 225800 315982 226104 316010
rect 224960 307080 225012 307086
rect 224960 307022 225012 307028
rect 226076 11966 226104 315982
rect 226156 307080 226208 307086
rect 226156 307022 226208 307028
rect 226064 11960 226116 11966
rect 226064 11902 226116 11908
rect 224960 8832 225012 8838
rect 224958 8800 224960 8809
rect 225012 8800 225014 8809
rect 224958 8735 225014 8744
rect 226168 7750 226196 307022
rect 226156 7744 226208 7750
rect 226156 7686 226208 7692
rect 225328 4208 225380 4214
rect 225328 4150 225380 4156
rect 224866 3904 224922 3913
rect 224866 3839 224922 3848
rect 225340 480 225368 4150
rect 226260 3777 226288 320062
rect 226444 318034 226472 320076
rect 226918 320062 227024 320090
rect 226432 318028 226484 318034
rect 226432 317970 226484 317976
rect 226996 313970 227024 320062
rect 227272 318209 227300 320076
rect 227258 318200 227314 318209
rect 227640 318186 227668 320076
rect 227258 318135 227314 318144
rect 227548 318158 227668 318186
rect 226996 313942 227300 313970
rect 227272 302138 227300 313942
rect 227272 302110 227392 302138
rect 227364 299470 227392 302110
rect 227352 299464 227404 299470
rect 227352 299406 227404 299412
rect 227444 289876 227496 289882
rect 227444 289818 227496 289824
rect 227456 282946 227484 289818
rect 227260 282940 227312 282946
rect 227260 282882 227312 282888
rect 227444 282940 227496 282946
rect 227444 282882 227496 282888
rect 227272 282826 227300 282882
rect 227272 282798 227392 282826
rect 227364 273306 227392 282798
rect 227364 273278 227484 273306
rect 227456 263634 227484 273278
rect 227260 263628 227312 263634
rect 227260 263570 227312 263576
rect 227444 263628 227496 263634
rect 227444 263570 227496 263576
rect 227272 263514 227300 263570
rect 227272 263486 227392 263514
rect 227364 253994 227392 263486
rect 227364 253966 227484 253994
rect 227456 244322 227484 253966
rect 227260 244316 227312 244322
rect 227260 244258 227312 244264
rect 227444 244316 227496 244322
rect 227444 244258 227496 244264
rect 227272 244202 227300 244258
rect 227272 244174 227392 244202
rect 227364 234682 227392 244174
rect 227364 234654 227484 234682
rect 227456 225010 227484 234654
rect 227260 225004 227312 225010
rect 227260 224946 227312 224952
rect 227444 225004 227496 225010
rect 227444 224946 227496 224952
rect 227272 224890 227300 224946
rect 227272 224862 227392 224890
rect 227364 215370 227392 224862
rect 227364 215342 227484 215370
rect 227456 205698 227484 215342
rect 227260 205692 227312 205698
rect 227260 205634 227312 205640
rect 227444 205692 227496 205698
rect 227444 205634 227496 205640
rect 227272 205578 227300 205634
rect 227272 205550 227392 205578
rect 227364 196058 227392 205550
rect 227364 196030 227484 196058
rect 227456 186386 227484 196030
rect 227260 186380 227312 186386
rect 227260 186322 227312 186328
rect 227444 186380 227496 186386
rect 227444 186322 227496 186328
rect 227272 186266 227300 186322
rect 227272 186238 227392 186266
rect 227364 183569 227392 186238
rect 227166 183560 227222 183569
rect 227166 183495 227222 183504
rect 227350 183560 227406 183569
rect 227350 183495 227406 183504
rect 227180 173942 227208 183495
rect 227168 173936 227220 173942
rect 227168 173878 227220 173884
rect 227444 173936 227496 173942
rect 227444 173878 227496 173884
rect 227456 167074 227484 173878
rect 227260 167068 227312 167074
rect 227260 167010 227312 167016
rect 227444 167068 227496 167074
rect 227444 167010 227496 167016
rect 227272 166954 227300 167010
rect 227272 166926 227392 166954
rect 227364 164218 227392 166926
rect 227352 164212 227404 164218
rect 227352 164154 227404 164160
rect 227352 157344 227404 157350
rect 227352 157286 227404 157292
rect 227364 154578 227392 157286
rect 227364 154550 227484 154578
rect 227456 147694 227484 154550
rect 227260 147688 227312 147694
rect 227444 147688 227496 147694
rect 227312 147636 227392 147642
rect 227260 147630 227392 147636
rect 227444 147630 227496 147636
rect 227272 147614 227392 147630
rect 227364 144906 227392 147614
rect 227352 144900 227404 144906
rect 227352 144842 227404 144848
rect 227352 137964 227404 137970
rect 227352 137906 227404 137912
rect 227364 135266 227392 137906
rect 227364 135238 227484 135266
rect 227456 128382 227484 135238
rect 227260 128376 227312 128382
rect 227444 128376 227496 128382
rect 227312 128324 227392 128330
rect 227260 128318 227392 128324
rect 227444 128318 227496 128324
rect 227272 128302 227392 128318
rect 227364 125594 227392 128302
rect 227352 125588 227404 125594
rect 227352 125530 227404 125536
rect 227352 118652 227404 118658
rect 227352 118594 227404 118600
rect 227364 115954 227392 118594
rect 227364 115926 227484 115954
rect 227456 109070 227484 115926
rect 227260 109064 227312 109070
rect 227444 109064 227496 109070
rect 227312 109012 227392 109018
rect 227260 109006 227392 109012
rect 227444 109006 227496 109012
rect 227272 108990 227392 109006
rect 227364 106282 227392 108990
rect 227352 106276 227404 106282
rect 227352 106218 227404 106224
rect 227352 99340 227404 99346
rect 227352 99282 227404 99288
rect 227364 96642 227392 99282
rect 227364 96614 227484 96642
rect 227456 89758 227484 96614
rect 227260 89752 227312 89758
rect 227444 89752 227496 89758
rect 227312 89700 227392 89706
rect 227260 89694 227392 89700
rect 227444 89694 227496 89700
rect 227272 89678 227392 89694
rect 227364 86970 227392 89678
rect 227352 86964 227404 86970
rect 227352 86906 227404 86912
rect 227444 77308 227496 77314
rect 227444 77250 227496 77256
rect 227456 70258 227484 77250
rect 227364 70230 227484 70258
rect 227364 60738 227392 70230
rect 227364 60710 227484 60738
rect 227456 57934 227484 60710
rect 227444 57928 227496 57934
rect 227444 57870 227496 57876
rect 227352 51060 227404 51066
rect 227352 51002 227404 51008
rect 227364 41426 227392 51002
rect 227364 41398 227484 41426
rect 227456 31770 227484 41398
rect 227272 31754 227484 31770
rect 227260 31748 227496 31754
rect 227312 31742 227444 31748
rect 227260 31690 227312 31696
rect 227444 31690 227496 31696
rect 227272 31659 227300 31690
rect 227456 22137 227484 31690
rect 227442 22128 227498 22137
rect 227442 22063 227498 22072
rect 227350 19408 227406 19417
rect 227350 19343 227406 19352
rect 227364 19310 227392 19343
rect 227352 19304 227404 19310
rect 227352 19246 227404 19252
rect 227548 7614 227576 318158
rect 228100 318034 228128 320076
rect 228482 320062 228772 320090
rect 227628 318028 227680 318034
rect 227628 317970 227680 317976
rect 228088 318028 228140 318034
rect 228088 317970 228140 317976
rect 227640 7682 227668 317970
rect 228744 315994 228772 320062
rect 228824 318028 228876 318034
rect 228824 317970 228876 317976
rect 228732 315988 228784 315994
rect 228732 315930 228784 315936
rect 228836 11830 228864 317970
rect 228824 11824 228876 11830
rect 228824 11766 228876 11772
rect 228928 8265 228956 320076
rect 229296 318034 229324 320076
rect 229756 318617 229784 320076
rect 230138 320062 230428 320090
rect 229742 318608 229798 318617
rect 229742 318543 229798 318552
rect 229284 318028 229336 318034
rect 229284 317970 229336 317976
rect 230296 318028 230348 318034
rect 230296 317970 230348 317976
rect 229008 315988 229060 315994
rect 229008 315930 229060 315936
rect 228914 8256 228970 8265
rect 228914 8191 228970 8200
rect 227628 7676 227680 7682
rect 227628 7618 227680 7624
rect 227536 7608 227588 7614
rect 227536 7550 227588 7556
rect 226524 5500 226576 5506
rect 226524 5442 226576 5448
rect 226246 3768 226302 3777
rect 226246 3703 226302 3712
rect 226536 480 226564 5442
rect 227720 5432 227772 5438
rect 227720 5374 227772 5380
rect 227732 480 227760 5374
rect 228916 4208 228968 4214
rect 228916 4150 228968 4156
rect 228928 480 228956 4150
rect 229020 3641 229048 315930
rect 230308 11762 230336 317970
rect 230296 11756 230348 11762
rect 230296 11698 230348 11704
rect 230400 8129 230428 320062
rect 230584 315382 230612 320076
rect 230572 315376 230624 315382
rect 230572 315318 230624 315324
rect 230676 313834 230704 320146
rect 230584 313806 230704 313834
rect 230768 320062 230966 320090
rect 231426 320062 231532 320090
rect 230584 307086 230612 313806
rect 230572 307080 230624 307086
rect 230572 307022 230624 307028
rect 230768 307018 230796 320062
rect 231504 318186 231532 320062
rect 231504 318158 231624 318186
rect 231596 315874 231624 318158
rect 232240 318073 232268 320076
rect 232424 320062 232622 320090
rect 232226 318064 232282 318073
rect 231860 318028 231912 318034
rect 232226 317999 232282 318008
rect 231860 317970 231912 317976
rect 231596 315846 231716 315874
rect 231492 315376 231544 315382
rect 231492 315318 231544 315324
rect 230756 307012 230808 307018
rect 230756 306954 230808 306960
rect 231504 12345 231532 315318
rect 231584 307080 231636 307086
rect 231584 307022 231636 307028
rect 231490 12336 231546 12345
rect 231490 12271 231546 12280
rect 231596 12209 231624 307022
rect 231582 12200 231638 12209
rect 231582 12135 231638 12144
rect 230386 8120 230442 8129
rect 230386 8055 230442 8064
rect 231688 7993 231716 315846
rect 231872 307086 231900 317970
rect 232424 316010 232452 320062
rect 233068 318034 233096 320076
rect 233252 320062 233450 320090
rect 233620 320062 233910 320090
rect 233056 318028 233108 318034
rect 233056 317970 233108 317976
rect 232056 315982 232452 316010
rect 231860 307080 231912 307086
rect 231860 307022 231912 307028
rect 231768 307012 231820 307018
rect 231768 306954 231820 306960
rect 231674 7984 231730 7993
rect 231674 7919 231730 7928
rect 230112 5364 230164 5370
rect 230112 5306 230164 5312
rect 229006 3632 229062 3641
rect 229006 3567 229062 3576
rect 230124 480 230152 5306
rect 231308 5296 231360 5302
rect 231308 5238 231360 5244
rect 231320 480 231348 5238
rect 231780 3505 231808 306954
rect 232056 302258 232084 315982
rect 233252 307086 233280 320062
rect 233332 318028 233384 318034
rect 233332 317970 233384 317976
rect 233344 311846 233372 317970
rect 233620 316010 233648 320062
rect 234264 318034 234292 320076
rect 234724 318345 234752 320076
rect 235106 320062 235396 320090
rect 234710 318336 234766 318345
rect 234710 318271 234766 318280
rect 234252 318028 234304 318034
rect 234252 317970 234304 317976
rect 233436 315982 233648 316010
rect 234896 316056 234948 316062
rect 234896 315998 234948 316004
rect 234620 315988 234672 315994
rect 233332 311840 233384 311846
rect 233332 311782 233384 311788
rect 233056 307080 233108 307086
rect 233056 307022 233108 307028
rect 233240 307080 233292 307086
rect 233240 307022 233292 307028
rect 232044 302252 232096 302258
rect 232044 302194 232096 302200
rect 233068 12073 233096 307022
rect 233436 302326 233464 315982
rect 234620 315930 234672 315936
rect 234344 311840 234396 311846
rect 234344 311782 234396 311788
rect 233424 302320 233476 302326
rect 233424 302262 233476 302268
rect 233148 302252 233200 302258
rect 233148 302194 233200 302200
rect 233054 12064 233110 12073
rect 233054 11999 233110 12008
rect 233160 7857 233188 302194
rect 234356 299538 234384 311782
rect 234632 307086 234660 315930
rect 234528 307080 234580 307086
rect 234528 307022 234580 307028
rect 234620 307080 234672 307086
rect 234620 307022 234672 307028
rect 234436 302252 234488 302258
rect 234436 302194 234488 302200
rect 234252 299532 234304 299538
rect 234252 299474 234304 299480
rect 234344 299532 234396 299538
rect 234344 299474 234396 299480
rect 234264 296721 234292 299474
rect 233974 296712 234030 296721
rect 233974 296647 234030 296656
rect 234250 296712 234306 296721
rect 234250 296647 234306 296656
rect 233988 287094 234016 296647
rect 233976 287088 234028 287094
rect 233976 287030 234028 287036
rect 234068 287088 234120 287094
rect 234068 287030 234120 287036
rect 234080 283642 234108 287030
rect 234080 283614 234200 283642
rect 234172 270434 234200 283614
rect 234160 270428 234212 270434
rect 234160 270370 234212 270376
rect 234068 260908 234120 260914
rect 234068 260850 234120 260856
rect 234080 251258 234108 260850
rect 234068 251252 234120 251258
rect 234068 251194 234120 251200
rect 234160 251252 234212 251258
rect 234160 251194 234212 251200
rect 234172 240174 234200 251194
rect 234068 240168 234120 240174
rect 234068 240110 234120 240116
rect 234160 240168 234212 240174
rect 234160 240110 234212 240116
rect 234080 234666 234108 240110
rect 234068 234660 234120 234666
rect 234068 234602 234120 234608
rect 234160 234524 234212 234530
rect 234160 234466 234212 234472
rect 234172 225078 234200 234466
rect 234160 225072 234212 225078
rect 234160 225014 234212 225020
rect 234068 224936 234120 224942
rect 234068 224878 234120 224884
rect 234080 217977 234108 224878
rect 233790 217968 233846 217977
rect 233790 217903 233846 217912
rect 234066 217968 234122 217977
rect 234066 217903 234122 217912
rect 233804 216646 233832 217903
rect 233792 216640 233844 216646
rect 233792 216582 233844 216588
rect 233792 208412 233844 208418
rect 233792 208354 233844 208360
rect 233804 203590 233832 208354
rect 233792 203584 233844 203590
rect 233792 203526 233844 203532
rect 234344 203584 234396 203590
rect 234344 203526 234396 203532
rect 234356 178650 234384 203526
rect 234172 178622 234384 178650
rect 234172 173913 234200 178622
rect 234158 173904 234214 173913
rect 234158 173839 234214 173848
rect 234342 173904 234398 173913
rect 234342 173839 234398 173848
rect 234356 162858 234384 173839
rect 234160 162852 234212 162858
rect 234160 162794 234212 162800
rect 234344 162852 234396 162858
rect 234344 162794 234396 162800
rect 234172 161430 234200 162794
rect 234160 161424 234212 161430
rect 234160 161366 234212 161372
rect 234160 151836 234212 151842
rect 234160 151778 234212 151784
rect 234172 144974 234200 151778
rect 234160 144968 234212 144974
rect 234160 144910 234212 144916
rect 234252 144832 234304 144838
rect 234252 144774 234304 144780
rect 234264 142118 234292 144774
rect 234252 142112 234304 142118
rect 234252 142054 234304 142060
rect 234252 124228 234304 124234
rect 234252 124170 234304 124176
rect 234264 119406 234292 124170
rect 234252 119400 234304 119406
rect 234252 119342 234304 119348
rect 234068 114640 234120 114646
rect 234120 114588 234200 114594
rect 234068 114582 234200 114588
rect 234080 114566 234200 114582
rect 234172 114510 234200 114566
rect 234160 114504 234212 114510
rect 234160 114446 234212 114452
rect 234252 104916 234304 104922
rect 234252 104858 234304 104864
rect 234264 100094 234292 104858
rect 234252 100088 234304 100094
rect 234252 100030 234304 100036
rect 234160 95260 234212 95266
rect 234160 95202 234212 95208
rect 234172 91798 234200 95202
rect 234160 91792 234212 91798
rect 234160 91734 234212 91740
rect 234344 87100 234396 87106
rect 234344 87042 234396 87048
rect 234356 86986 234384 87042
rect 234264 86958 234384 86986
rect 234264 85542 234292 86958
rect 234252 85536 234304 85542
rect 234252 85478 234304 85484
rect 234160 75948 234212 75954
rect 234160 75890 234212 75896
rect 234172 70530 234200 75890
rect 234172 70502 234292 70530
rect 234264 67658 234292 70502
rect 234068 67652 234120 67658
rect 234068 67594 234120 67600
rect 234252 67652 234304 67658
rect 234252 67594 234304 67600
rect 234080 66230 234108 67594
rect 234068 66224 234120 66230
rect 234068 66166 234120 66172
rect 234252 57860 234304 57866
rect 234252 57802 234304 57808
rect 234264 48346 234292 57802
rect 234068 48340 234120 48346
rect 234068 48282 234120 48288
rect 234252 48340 234304 48346
rect 234252 48282 234304 48288
rect 234080 46918 234108 48282
rect 234068 46912 234120 46918
rect 234068 46854 234120 46860
rect 234068 38684 234120 38690
rect 234068 38626 234120 38632
rect 234080 31634 234108 38626
rect 234080 31606 234292 31634
rect 234264 22114 234292 31606
rect 234264 22086 234384 22114
rect 234356 19310 234384 22086
rect 234344 19304 234396 19310
rect 234344 19246 234396 19252
rect 234448 10010 234476 302194
rect 234356 9982 234476 10010
rect 233146 7848 233202 7857
rect 233146 7783 233202 7792
rect 234356 7721 234384 9982
rect 234436 8424 234488 8430
rect 234434 8392 234436 8401
rect 234488 8392 234490 8401
rect 234434 8327 234490 8336
rect 234342 7712 234398 7721
rect 234342 7647 234398 7656
rect 233700 5228 233752 5234
rect 233700 5170 233752 5176
rect 231860 4412 231912 4418
rect 231860 4354 231912 4360
rect 231872 4298 231900 4354
rect 232504 4344 232556 4350
rect 231872 4282 231992 4298
rect 232504 4286 232556 4292
rect 231872 4276 232004 4282
rect 231872 4270 231952 4276
rect 231952 4218 232004 4224
rect 231766 3496 231822 3505
rect 231766 3431 231822 3440
rect 232516 480 232544 4286
rect 233712 480 233740 5170
rect 234540 3369 234568 307022
rect 234908 296818 234936 315998
rect 235368 315874 235396 320062
rect 235644 320062 235934 320090
rect 236196 320062 236394 320090
rect 236472 320062 236762 320090
rect 235448 319932 235500 319938
rect 235448 319874 235500 319880
rect 235460 315994 235488 319874
rect 235644 316062 235672 320062
rect 236196 317422 236224 320062
rect 236184 317416 236236 317422
rect 236184 317358 236236 317364
rect 235632 316056 235684 316062
rect 235632 315998 235684 316004
rect 236472 315994 236500 320062
rect 237208 318617 237236 320076
rect 237392 320062 237590 320090
rect 237194 318608 237250 318617
rect 237194 318543 237250 318552
rect 235448 315988 235500 315994
rect 235448 315930 235500 315936
rect 236000 315988 236052 315994
rect 236000 315930 236052 315936
rect 236460 315988 236512 315994
rect 236460 315930 236512 315936
rect 235368 315846 235948 315874
rect 235816 307080 235868 307086
rect 235816 307022 235868 307028
rect 234896 296812 234948 296818
rect 234896 296754 234948 296760
rect 235724 296812 235776 296818
rect 235724 296754 235776 296760
rect 235736 296682 235764 296754
rect 235724 296676 235776 296682
rect 235724 296618 235776 296624
rect 235724 287156 235776 287162
rect 235724 287098 235776 287104
rect 235736 209778 235764 287098
rect 235724 209772 235776 209778
rect 235724 209714 235776 209720
rect 235540 200184 235592 200190
rect 235540 200126 235592 200132
rect 235552 180849 235580 200126
rect 235538 180840 235594 180849
rect 235538 180775 235594 180784
rect 235722 180840 235778 180849
rect 235722 180775 235724 180784
rect 235776 180775 235778 180784
rect 235724 180746 235776 180752
rect 235632 171148 235684 171154
rect 235632 171090 235684 171096
rect 235644 169266 235672 171090
rect 235552 169238 235672 169266
rect 235552 154601 235580 169238
rect 235538 154592 235594 154601
rect 235538 154527 235594 154536
rect 235722 154592 235778 154601
rect 235722 154527 235778 154536
rect 235736 96626 235764 154527
rect 235724 96620 235776 96626
rect 235724 96562 235776 96568
rect 235724 87032 235776 87038
rect 235724 86974 235776 86980
rect 235736 77246 235764 86974
rect 235724 77240 235776 77246
rect 235724 77182 235776 77188
rect 235724 67652 235776 67658
rect 235724 67594 235776 67600
rect 235736 57934 235764 67594
rect 235724 57928 235776 57934
rect 235724 57870 235776 57876
rect 235724 48340 235776 48346
rect 235724 48282 235776 48288
rect 235736 38622 235764 48282
rect 235724 38616 235776 38622
rect 235724 38558 235776 38564
rect 235724 29028 235776 29034
rect 235724 28970 235776 28976
rect 235736 19310 235764 28970
rect 234620 19304 234672 19310
rect 234620 19246 234672 19252
rect 235724 19304 235776 19310
rect 235724 19246 235776 19252
rect 234632 11937 234660 19246
rect 234618 11928 234674 11937
rect 234618 11863 234674 11872
rect 235828 11801 235856 307022
rect 235814 11792 235870 11801
rect 235814 11727 235870 11736
rect 235920 7585 235948 315846
rect 236012 307086 236040 315930
rect 236184 307828 236236 307834
rect 236184 307770 236236 307776
rect 236000 307080 236052 307086
rect 236000 307022 236052 307028
rect 236196 306746 236224 307770
rect 237392 307086 237420 320062
rect 238036 318850 238064 320076
rect 238128 320062 238418 320090
rect 238786 320062 238892 320090
rect 237656 318844 237708 318850
rect 237656 318786 237708 318792
rect 238024 318844 238076 318850
rect 238024 318786 238076 318792
rect 237668 317422 237696 318786
rect 237656 317416 237708 317422
rect 237656 317358 237708 317364
rect 238128 315994 238156 320062
rect 238576 317416 238628 317422
rect 238576 317358 238628 317364
rect 237472 315988 237524 315994
rect 237472 315930 237524 315936
rect 238116 315988 238168 315994
rect 238116 315930 238168 315936
rect 237288 307080 237340 307086
rect 237288 307022 237340 307028
rect 237380 307080 237432 307086
rect 237380 307022 237432 307028
rect 236184 306740 236236 306746
rect 236184 306682 236236 306688
rect 237104 306740 237156 306746
rect 237104 306682 237156 306688
rect 237116 289762 237144 306682
rect 237116 289734 237236 289762
rect 237208 26874 237236 289734
rect 237116 26846 237236 26874
rect 237116 14686 237144 26846
rect 237104 14680 237156 14686
rect 237104 14622 237156 14628
rect 237300 11665 237328 307022
rect 237484 302190 237512 315930
rect 237472 302184 237524 302190
rect 237472 302126 237524 302132
rect 238392 302184 238444 302190
rect 238392 302126 238444 302132
rect 238404 289762 238432 302126
rect 238404 289734 238524 289762
rect 238496 26874 238524 289734
rect 238404 26846 238524 26874
rect 238404 14550 238432 26846
rect 238588 14618 238616 317358
rect 238864 316198 238892 320062
rect 239048 320062 239246 320090
rect 239324 320062 239614 320090
rect 239784 320062 240074 320090
rect 239048 318866 239076 320062
rect 238956 318838 239076 318866
rect 238956 317422 238984 318838
rect 238944 317416 238996 317422
rect 238944 317358 238996 317364
rect 238852 316192 238904 316198
rect 238852 316134 238904 316140
rect 238852 316056 238904 316062
rect 238852 315998 238904 316004
rect 238760 315988 238812 315994
rect 238760 315930 238812 315936
rect 238668 307080 238720 307086
rect 238668 307022 238720 307028
rect 238576 14612 238628 14618
rect 238576 14554 238628 14560
rect 238392 14544 238444 14550
rect 238392 14486 238444 14492
rect 238680 12578 238708 307022
rect 238772 307018 238800 315930
rect 238864 307086 238892 315998
rect 239324 315994 239352 320062
rect 239784 316062 239812 320062
rect 240888 318850 240916 320076
rect 240980 320062 241270 320090
rect 240508 318844 240560 318850
rect 240508 318786 240560 318792
rect 240876 318844 240928 318850
rect 240876 318786 240928 318792
rect 240520 317422 240548 318786
rect 240508 317416 240560 317422
rect 240508 317358 240560 317364
rect 239956 316192 240008 316198
rect 239956 316134 240008 316140
rect 239772 316056 239824 316062
rect 239772 315998 239824 316004
rect 239312 315988 239364 315994
rect 239312 315930 239364 315936
rect 238944 307828 238996 307834
rect 238944 307770 238996 307776
rect 238852 307080 238904 307086
rect 238852 307022 238904 307028
rect 238760 307012 238812 307018
rect 238760 306954 238812 306960
rect 238956 302258 238984 307770
rect 239864 307080 239916 307086
rect 239864 307022 239916 307028
rect 238944 302252 238996 302258
rect 238944 302194 238996 302200
rect 239772 302184 239824 302190
rect 239772 302126 239824 302132
rect 239784 278066 239812 302126
rect 239692 278038 239812 278066
rect 239692 14482 239720 278038
rect 239876 15201 239904 307022
rect 239862 15192 239918 15201
rect 239862 15127 239918 15136
rect 239680 14476 239732 14482
rect 239680 14418 239732 14424
rect 239968 12646 239996 316134
rect 240980 315994 241008 320062
rect 241244 317416 241296 317422
rect 241244 317358 241296 317364
rect 240140 315988 240192 315994
rect 240140 315930 240192 315936
rect 240968 315988 241020 315994
rect 240968 315930 241020 315936
rect 240152 307086 240180 315930
rect 240140 307080 240192 307086
rect 240140 307022 240192 307028
rect 240048 307012 240100 307018
rect 240048 306954 240100 306960
rect 240060 12714 240088 306954
rect 241256 278066 241284 317358
rect 241164 278038 241284 278066
rect 241164 12782 241192 278038
rect 241152 12776 241204 12782
rect 241152 12718 241204 12724
rect 240048 12708 240100 12714
rect 240048 12650 240100 12656
rect 239956 12640 240008 12646
rect 239956 12582 240008 12588
rect 238668 12572 238720 12578
rect 238668 12514 238720 12520
rect 237286 11656 237342 11665
rect 237286 11591 237342 11600
rect 239586 8800 239642 8809
rect 238392 8764 238444 8770
rect 239586 8735 239642 8744
rect 238392 8706 238444 8712
rect 236000 8696 236052 8702
rect 236000 8638 236052 8644
rect 235906 7576 235962 7585
rect 235906 7511 235962 7520
rect 234804 5160 234856 5166
rect 234804 5102 234856 5108
rect 234526 3360 234582 3369
rect 234526 3295 234582 3304
rect 234816 480 234844 5102
rect 236012 480 236040 8638
rect 237196 5092 237248 5098
rect 237196 5034 237248 5040
rect 237208 480 237236 5034
rect 238404 480 238432 8706
rect 239600 480 239628 8735
rect 239772 8492 239824 8498
rect 239772 8434 239824 8440
rect 239784 8401 239812 8434
rect 241348 8430 241376 320146
rect 242084 318850 242112 320076
rect 242176 320062 242558 320090
rect 241612 318844 241664 318850
rect 241612 318786 241664 318792
rect 242072 318844 242124 318850
rect 242072 318786 242124 318792
rect 241520 315988 241572 315994
rect 241520 315930 241572 315936
rect 241532 307086 241560 315930
rect 241624 314158 241652 318786
rect 242176 315994 242204 320062
rect 242164 315988 242216 315994
rect 242164 315930 242216 315936
rect 241612 314152 241664 314158
rect 241612 314094 241664 314100
rect 242624 314152 242676 314158
rect 242624 314094 242676 314100
rect 241428 307080 241480 307086
rect 241428 307022 241480 307028
rect 241520 307080 241572 307086
rect 241520 307022 241572 307028
rect 241336 8424 241388 8430
rect 239770 8392 239826 8401
rect 241336 8366 241388 8372
rect 239770 8327 239826 8336
rect 241440 6934 241468 307022
rect 242636 298110 242664 314094
rect 242624 298104 242676 298110
rect 242624 298046 242676 298052
rect 242624 288448 242676 288454
rect 242624 288390 242676 288396
rect 242636 270502 242664 288390
rect 242532 270496 242584 270502
rect 242532 270438 242584 270444
rect 242624 270496 242676 270502
rect 242624 270438 242676 270444
rect 242544 249801 242572 270438
rect 242346 249792 242402 249801
rect 242346 249727 242402 249736
rect 242530 249792 242586 249801
rect 242530 249727 242586 249736
rect 242360 240174 242388 249727
rect 242348 240168 242400 240174
rect 242348 240110 242400 240116
rect 242532 240168 242584 240174
rect 242532 240110 242584 240116
rect 242544 230489 242572 240110
rect 242346 230480 242402 230489
rect 242346 230415 242402 230424
rect 242530 230480 242586 230489
rect 242530 230415 242586 230424
rect 242360 220862 242388 230415
rect 242348 220856 242400 220862
rect 242348 220798 242400 220804
rect 242532 220856 242584 220862
rect 242532 220798 242584 220804
rect 242544 211138 242572 220798
rect 242348 211132 242400 211138
rect 242348 211074 242400 211080
rect 242532 211132 242584 211138
rect 242532 211074 242584 211080
rect 242360 201521 242388 211074
rect 242346 201512 242402 201521
rect 242346 201447 242402 201456
rect 242530 201512 242586 201521
rect 242530 201447 242586 201456
rect 242544 191826 242572 201447
rect 242348 191820 242400 191826
rect 242348 191762 242400 191768
rect 242532 191820 242584 191826
rect 242532 191762 242584 191768
rect 242360 182209 242388 191762
rect 242346 182200 242402 182209
rect 242346 182135 242402 182144
rect 242530 182200 242586 182209
rect 242530 182135 242586 182144
rect 242544 172514 242572 182135
rect 242532 172508 242584 172514
rect 242532 172450 242584 172456
rect 242532 162920 242584 162926
rect 242532 162862 242584 162868
rect 242544 153202 242572 162862
rect 242532 153196 242584 153202
rect 242532 153138 242584 153144
rect 242532 143608 242584 143614
rect 242532 143550 242584 143556
rect 242544 133890 242572 143550
rect 242532 133884 242584 133890
rect 242532 133826 242584 133832
rect 242532 124228 242584 124234
rect 242532 124170 242584 124176
rect 242544 114510 242572 124170
rect 242532 114504 242584 114510
rect 242532 114446 242584 114452
rect 242532 104916 242584 104922
rect 242532 104858 242584 104864
rect 242544 95198 242572 104858
rect 242532 95192 242584 95198
rect 242532 95134 242584 95140
rect 242532 85604 242584 85610
rect 242532 85546 242584 85552
rect 242544 75886 242572 85546
rect 242532 75880 242584 75886
rect 242532 75822 242584 75828
rect 242532 66292 242584 66298
rect 242532 66234 242584 66240
rect 242544 56574 242572 66234
rect 242532 56568 242584 56574
rect 242532 56510 242584 56516
rect 242532 46980 242584 46986
rect 242532 46922 242584 46928
rect 242544 37262 242572 46922
rect 242532 37256 242584 37262
rect 242532 37198 242584 37204
rect 242532 27668 242584 27674
rect 242532 27610 242584 27616
rect 242544 22794 242572 27610
rect 242360 22766 242572 22794
rect 242360 19258 242388 22766
rect 242360 19230 242480 19258
rect 242452 12850 242480 19230
rect 242440 12844 242492 12850
rect 242440 12786 242492 12792
rect 242728 8838 242756 320146
rect 242926 320062 243032 320090
rect 242900 315988 242952 315994
rect 242900 315930 242952 315936
rect 242808 307080 242860 307086
rect 242808 307022 242860 307028
rect 242716 8832 242768 8838
rect 242716 8774 242768 8780
rect 241980 8764 242032 8770
rect 241980 8706 242032 8712
rect 241428 6928 241480 6934
rect 241428 6870 241480 6876
rect 240784 5024 240836 5030
rect 240784 4966 240836 4972
rect 240796 480 240824 4966
rect 241992 480 242020 8706
rect 242820 5098 242848 307022
rect 242912 306882 242940 315930
rect 243004 307068 243032 320062
rect 243096 320062 243386 320090
rect 243754 320062 244044 320090
rect 243096 315994 243124 320062
rect 244016 316010 244044 320062
rect 244200 319444 244228 320076
rect 244108 319416 244228 319444
rect 244108 316130 244136 319416
rect 244096 316124 244148 316130
rect 244096 316066 244148 316072
rect 243084 315988 243136 315994
rect 244016 315982 244228 316010
rect 243084 315930 243136 315936
rect 244096 315920 244148 315926
rect 244096 315862 244148 315868
rect 243004 307040 244044 307068
rect 242900 306876 242952 306882
rect 242900 306818 242952 306824
rect 243912 306876 243964 306882
rect 243912 306818 243964 306824
rect 243924 298110 243952 306818
rect 243912 298104 243964 298110
rect 243912 298046 243964 298052
rect 243820 288448 243872 288454
rect 243820 288390 243872 288396
rect 243832 278866 243860 288390
rect 243820 278860 243872 278866
rect 243820 278802 243872 278808
rect 243820 277432 243872 277438
rect 243820 277374 243872 277380
rect 243832 269210 243860 277374
rect 243820 269204 243872 269210
rect 243820 269146 243872 269152
rect 243728 269068 243780 269074
rect 243728 269010 243780 269016
rect 243740 264466 243768 269010
rect 243648 264438 243768 264466
rect 243648 249830 243676 264438
rect 243636 249824 243688 249830
rect 243636 249766 243688 249772
rect 243820 249824 243872 249830
rect 243820 249766 243872 249772
rect 243832 245018 243860 249766
rect 243648 244990 243860 245018
rect 243648 230518 243676 244990
rect 243636 230512 243688 230518
rect 243636 230454 243688 230460
rect 243820 230512 243872 230518
rect 243820 230454 243872 230460
rect 243832 220810 243860 230454
rect 243740 220782 243860 220810
rect 243740 211206 243768 220782
rect 243728 211200 243780 211206
rect 243728 211142 243780 211148
rect 243820 211200 243872 211206
rect 243820 211142 243872 211148
rect 243832 206258 243860 211142
rect 243740 206230 243860 206258
rect 243740 191894 243768 206230
rect 243728 191888 243780 191894
rect 243728 191830 243780 191836
rect 243820 191888 243872 191894
rect 243820 191830 243872 191836
rect 243832 182186 243860 191830
rect 243740 182158 243860 182186
rect 243740 172582 243768 182158
rect 243728 172576 243780 172582
rect 243728 172518 243780 172524
rect 243820 172576 243872 172582
rect 243820 172518 243872 172524
rect 243832 172446 243860 172518
rect 243820 172440 243872 172446
rect 243820 172382 243872 172388
rect 243912 172440 243964 172446
rect 243912 172382 243964 172388
rect 243924 162874 243952 172382
rect 243832 162846 243952 162874
rect 243832 161430 243860 162846
rect 243820 161424 243872 161430
rect 243820 161366 243872 161372
rect 243820 151836 243872 151842
rect 243820 151778 243872 151784
rect 243832 143614 243860 151778
rect 243636 143608 243688 143614
rect 243636 143550 243688 143556
rect 243820 143608 243872 143614
rect 243820 143550 243872 143556
rect 243648 133958 243676 143550
rect 243636 133952 243688 133958
rect 243636 133894 243688 133900
rect 243820 133952 243872 133958
rect 243820 133894 243872 133900
rect 243832 133822 243860 133894
rect 243820 133816 243872 133822
rect 243820 133758 243872 133764
rect 243820 124228 243872 124234
rect 243820 124170 243872 124176
rect 243832 122806 243860 124170
rect 243820 122800 243872 122806
rect 243820 122742 243872 122748
rect 243820 113212 243872 113218
rect 243820 113154 243872 113160
rect 243832 104990 243860 113154
rect 243820 104984 243872 104990
rect 243820 104926 243872 104932
rect 243636 104916 243688 104922
rect 243636 104858 243688 104864
rect 243648 95266 243676 104858
rect 243636 95260 243688 95266
rect 243636 95202 243688 95208
rect 243820 95260 243872 95266
rect 243820 95202 243872 95208
rect 243832 90250 243860 95202
rect 243648 90222 243860 90250
rect 243648 75954 243676 90222
rect 243636 75948 243688 75954
rect 243636 75890 243688 75896
rect 243820 75948 243872 75954
rect 243820 75890 243872 75896
rect 243832 71074 243860 75890
rect 243648 71046 243860 71074
rect 243648 56642 243676 71046
rect 243636 56636 243688 56642
rect 243636 56578 243688 56584
rect 243820 56636 243872 56642
rect 243820 56578 243872 56584
rect 243832 46889 243860 56578
rect 243634 46880 243690 46889
rect 243634 46815 243690 46824
rect 243818 46880 243874 46889
rect 243818 46815 243874 46824
rect 243648 37330 243676 46815
rect 243636 37324 243688 37330
rect 243636 37266 243688 37272
rect 243820 37324 243872 37330
rect 243820 37266 243872 37272
rect 243832 27554 243860 37266
rect 243740 27526 243860 27554
rect 243740 18018 243768 27526
rect 243728 18012 243780 18018
rect 243728 17954 243780 17960
rect 243820 18012 243872 18018
rect 243820 17954 243872 17960
rect 243832 12918 243860 17954
rect 243820 12912 243872 12918
rect 243820 12854 243872 12860
rect 244016 9382 244044 307040
rect 244004 9376 244056 9382
rect 244004 9318 244056 9324
rect 244108 9217 244136 315862
rect 244094 9208 244150 9217
rect 244094 9143 244150 9152
rect 243176 8696 243228 8702
rect 243176 8638 243228 8644
rect 242900 8560 242952 8566
rect 242900 8502 242952 8508
rect 242808 5092 242860 5098
rect 242808 5034 242860 5040
rect 242912 2990 242940 8502
rect 242900 2984 242952 2990
rect 242900 2926 242952 2932
rect 243188 480 243216 8638
rect 244200 5030 244228 315982
rect 244292 307086 244320 320146
rect 244280 307080 244332 307086
rect 244280 307022 244332 307028
rect 244384 296342 244412 320198
rect 245160 320198 245410 320204
rect 245660 320204 245712 320210
rect 245108 320146 245160 320152
rect 245660 320146 245712 320152
rect 246396 320204 246698 320210
rect 246448 320198 246698 320204
rect 247132 320204 247184 320210
rect 246396 320146 246448 320152
rect 247132 320146 247184 320152
rect 248052 320204 248354 320210
rect 248104 320198 248354 320204
rect 252862 320210 253060 320226
rect 252862 320204 253072 320210
rect 252862 320198 253020 320204
rect 248052 320146 248104 320152
rect 253020 320146 253072 320152
rect 253756 320204 253808 320210
rect 253756 320146 253808 320152
rect 253860 320198 254058 320226
rect 255714 320210 256004 320226
rect 255714 320204 256016 320210
rect 255714 320198 255964 320204
rect 245028 318850 245056 320076
rect 245016 318844 245068 318850
rect 245016 318786 245068 318792
rect 245568 318844 245620 318850
rect 245568 318786 245620 318792
rect 245580 309126 245608 318786
rect 245568 309120 245620 309126
rect 245568 309062 245620 309068
rect 245672 307086 245700 320146
rect 245856 318850 245884 320076
rect 246238 320062 246528 320090
rect 245752 318844 245804 318850
rect 245752 318786 245804 318792
rect 245844 318844 245896 318850
rect 245844 318786 245896 318792
rect 245476 307080 245528 307086
rect 245476 307022 245528 307028
rect 245660 307080 245712 307086
rect 245660 307022 245712 307028
rect 244372 296336 244424 296342
rect 244372 296278 244424 296284
rect 245384 296336 245436 296342
rect 245384 296278 245436 296284
rect 245292 19304 245344 19310
rect 245292 19246 245344 19252
rect 245304 12866 245332 19246
rect 245396 12986 245424 296278
rect 245384 12980 245436 12986
rect 245384 12922 245436 12928
rect 245304 12838 245424 12866
rect 245396 5506 245424 12838
rect 245488 9450 245516 307022
rect 245568 299532 245620 299538
rect 245568 299474 245620 299480
rect 245580 19310 245608 299474
rect 245764 294642 245792 318786
rect 246500 315246 246528 320062
rect 246488 315240 246540 315246
rect 246488 315182 246540 315188
rect 246948 315240 247000 315246
rect 246948 315182 247000 315188
rect 246856 307080 246908 307086
rect 246856 307022 246908 307028
rect 245752 294636 245804 294642
rect 245752 294578 245804 294584
rect 246764 294636 246816 294642
rect 246764 294578 246816 294584
rect 245568 19304 245620 19310
rect 245568 19246 245620 19252
rect 246776 13054 246804 294578
rect 246764 13048 246816 13054
rect 246764 12990 246816 12996
rect 246764 9580 246816 9586
rect 246764 9522 246816 9528
rect 245568 9512 245620 9518
rect 245568 9454 245620 9460
rect 245476 9444 245528 9450
rect 245476 9386 245528 9392
rect 245384 5500 245436 5506
rect 245384 5442 245436 5448
rect 244188 5024 244240 5030
rect 244188 4966 244240 4972
rect 244372 4956 244424 4962
rect 244372 4898 244424 4904
rect 244186 4584 244242 4593
rect 244186 4519 244242 4528
rect 244200 4486 244228 4519
rect 244188 4480 244240 4486
rect 244188 4422 244240 4428
rect 244384 480 244412 4898
rect 245580 480 245608 9454
rect 246776 480 246804 9522
rect 246868 9314 246896 307022
rect 246960 298110 246988 315182
rect 247052 307358 247080 320076
rect 247040 307352 247092 307358
rect 247040 307294 247092 307300
rect 247144 307034 247172 320146
rect 247236 320062 247526 320090
rect 247894 320062 248184 320090
rect 247236 309806 247264 320062
rect 248156 317422 248184 320062
rect 248432 320062 248722 320090
rect 249182 320062 249288 320090
rect 248144 317416 248196 317422
rect 248144 317358 248196 317364
rect 248328 317416 248380 317422
rect 248328 317358 248380 317364
rect 248340 311658 248368 317358
rect 248248 311630 248368 311658
rect 247224 309800 247276 309806
rect 247224 309742 247276 309748
rect 248144 307352 248196 307358
rect 248144 307294 248196 307300
rect 247144 307006 247264 307034
rect 246948 298104 247000 298110
rect 246948 298046 247000 298052
rect 247236 294642 247264 307006
rect 247224 294636 247276 294642
rect 247224 294578 247276 294584
rect 248052 294636 248104 294642
rect 248052 294578 248104 294584
rect 246948 288448 247000 288454
rect 246948 288390 247000 288396
rect 246960 259457 246988 288390
rect 246946 259448 247002 259457
rect 246946 259383 247002 259392
rect 247130 259448 247186 259457
rect 247130 259383 247186 259392
rect 247144 249830 247172 259383
rect 246948 249824 247000 249830
rect 246948 249766 247000 249772
rect 247132 249824 247184 249830
rect 247132 249766 247184 249772
rect 246960 240145 246988 249766
rect 246946 240136 247002 240145
rect 246946 240071 247002 240080
rect 247130 240136 247186 240145
rect 247130 240071 247186 240080
rect 247144 230518 247172 240071
rect 246948 230512 247000 230518
rect 246948 230454 247000 230460
rect 247132 230512 247184 230518
rect 247132 230454 247184 230460
rect 246960 220833 246988 230454
rect 246946 220824 247002 220833
rect 246946 220759 247002 220768
rect 247130 220824 247186 220833
rect 247130 220759 247186 220768
rect 247144 211177 247172 220759
rect 246946 211168 247002 211177
rect 246946 211103 247002 211112
rect 247130 211168 247186 211177
rect 247130 211103 247186 211112
rect 246960 201482 246988 211103
rect 246948 201476 247000 201482
rect 246948 201418 247000 201424
rect 247132 201476 247184 201482
rect 247132 201418 247184 201424
rect 247144 191865 247172 201418
rect 246946 191856 247002 191865
rect 246946 191791 247002 191800
rect 247130 191856 247186 191865
rect 247130 191791 247186 191800
rect 246960 182170 246988 191791
rect 246948 182164 247000 182170
rect 246948 182106 247000 182112
rect 247132 182164 247184 182170
rect 247132 182106 247184 182112
rect 247144 172553 247172 182106
rect 246946 172544 247002 172553
rect 246946 172479 247002 172488
rect 247130 172544 247186 172553
rect 247130 172479 247186 172488
rect 246960 143546 246988 172479
rect 246948 143540 247000 143546
rect 246948 143482 247000 143488
rect 247132 143540 247184 143546
rect 247132 143482 247184 143488
rect 247144 133929 247172 143482
rect 246946 133920 247002 133929
rect 246946 133855 247002 133864
rect 247130 133920 247186 133929
rect 247130 133855 247186 133864
rect 246960 104854 246988 133855
rect 246948 104848 247000 104854
rect 246948 104790 247000 104796
rect 246948 95260 247000 95266
rect 246948 95202 247000 95208
rect 246960 85542 246988 95202
rect 246948 85536 247000 85542
rect 246948 85478 247000 85484
rect 246948 75948 247000 75954
rect 246948 75890 247000 75896
rect 246960 66230 246988 75890
rect 246948 66224 247000 66230
rect 246948 66166 247000 66172
rect 246948 56636 247000 56642
rect 246948 56578 247000 56584
rect 246960 46918 246988 56578
rect 246948 46912 247000 46918
rect 246948 46854 247000 46860
rect 246948 37324 247000 37330
rect 246948 37266 247000 37272
rect 246960 9897 246988 37266
rect 248064 13734 248092 294578
rect 248156 13802 248184 307294
rect 248248 298110 248276 311630
rect 248328 309800 248380 309806
rect 248328 309742 248380 309748
rect 248236 298104 248288 298110
rect 248236 298046 248288 298052
rect 248236 288448 248288 288454
rect 248236 288390 248288 288396
rect 248248 143546 248276 288390
rect 248236 143540 248288 143546
rect 248236 143482 248288 143488
rect 248234 133920 248290 133929
rect 248234 133855 248290 133864
rect 248248 27606 248276 133855
rect 248236 27600 248288 27606
rect 248236 27542 248288 27548
rect 248236 18012 248288 18018
rect 248236 17954 248288 17960
rect 248248 17134 248276 17954
rect 248236 17128 248288 17134
rect 248236 17070 248288 17076
rect 248144 13796 248196 13802
rect 248144 13738 248196 13744
rect 248052 13728 248104 13734
rect 248052 13670 248104 13676
rect 246946 9888 247002 9897
rect 246946 9823 247002 9832
rect 246856 9308 246908 9314
rect 246856 9250 246908 9256
rect 248144 8764 248196 8770
rect 248144 8706 248196 8712
rect 248156 8673 248184 8706
rect 248142 8664 248198 8673
rect 248142 8599 248198 8608
rect 248340 6934 248368 309742
rect 248432 307086 248460 320062
rect 249260 318866 249288 320062
rect 249536 319444 249564 320076
rect 249904 319444 249932 320076
rect 250378 320062 250576 320090
rect 249444 319416 249564 319444
rect 249812 319416 249932 319444
rect 249260 318838 249380 318866
rect 248512 311636 248564 311642
rect 248512 311578 248564 311584
rect 248420 307080 248472 307086
rect 248420 307022 248472 307028
rect 248524 294642 248552 311578
rect 249352 311522 249380 318838
rect 249444 311642 249472 319416
rect 249432 311636 249484 311642
rect 249432 311578 249484 311584
rect 249352 311494 249472 311522
rect 248512 294636 248564 294642
rect 248512 294578 248564 294584
rect 249444 289882 249472 311494
rect 249812 307086 249840 319416
rect 250548 313954 250576 320062
rect 250732 319444 250760 320076
rect 251206 320062 251404 320090
rect 251574 320062 251680 320090
rect 250640 319416 250760 319444
rect 250536 313948 250588 313954
rect 250536 313890 250588 313896
rect 250640 311642 250668 319416
rect 251376 316198 251404 320062
rect 251652 319462 251680 320062
rect 251744 320062 252034 320090
rect 251456 319456 251508 319462
rect 251456 319398 251508 319404
rect 251640 319456 251692 319462
rect 251640 319398 251692 319404
rect 251364 316192 251416 316198
rect 251364 316134 251416 316140
rect 250996 313948 251048 313954
rect 250996 313890 251048 313896
rect 249892 311636 249944 311642
rect 249892 311578 249944 311584
rect 250628 311636 250680 311642
rect 250628 311578 250680 311584
rect 249708 307080 249760 307086
rect 249708 307022 249760 307028
rect 249800 307080 249852 307086
rect 249800 307022 249852 307028
rect 249524 294636 249576 294642
rect 249524 294578 249576 294584
rect 249432 289876 249484 289882
rect 249432 289818 249484 289824
rect 248420 143540 248472 143546
rect 248420 143482 248472 143488
rect 249432 143540 249484 143546
rect 249432 143482 249484 143488
rect 248432 133929 248460 143482
rect 249444 133929 249472 143482
rect 248418 133920 248474 133929
rect 248418 133855 248474 133864
rect 249430 133920 249486 133929
rect 249430 133855 249486 133864
rect 248420 17128 248472 17134
rect 248420 17070 248472 17076
rect 248432 8770 248460 17070
rect 249536 13666 249564 294578
rect 249616 289876 249668 289882
rect 249616 289818 249668 289824
rect 249628 270502 249656 289818
rect 249616 270496 249668 270502
rect 249616 270438 249668 270444
rect 249616 260908 249668 260914
rect 249616 260850 249668 260856
rect 249628 143546 249656 260850
rect 249616 143540 249668 143546
rect 249616 143482 249668 143488
rect 249614 133920 249670 133929
rect 249614 133855 249670 133864
rect 249628 27606 249656 133855
rect 249616 27600 249668 27606
rect 249616 27542 249668 27548
rect 249616 18012 249668 18018
rect 249616 17954 249668 17960
rect 249524 13660 249576 13666
rect 249524 13602 249576 13608
rect 249628 13546 249656 17954
rect 249444 13518 249656 13546
rect 249444 12322 249472 13518
rect 249444 12294 249564 12322
rect 249246 9480 249302 9489
rect 249246 9415 249302 9424
rect 248800 8906 249012 8922
rect 248788 8900 249012 8906
rect 248840 8894 249012 8900
rect 248788 8842 248840 8848
rect 248420 8764 248472 8770
rect 248420 8706 248472 8712
rect 248984 8514 249012 8894
rect 248984 8486 249196 8514
rect 248328 6928 248380 6934
rect 248328 6870 248380 6876
rect 247960 4888 248012 4894
rect 247960 4830 248012 4836
rect 247972 480 248000 4830
rect 249064 4752 249116 4758
rect 249064 4694 249116 4700
rect 249076 4593 249104 4694
rect 249062 4584 249118 4593
rect 249062 4519 249118 4528
rect 249168 480 249196 8486
rect 249260 4486 249288 9415
rect 249536 9382 249564 12294
rect 249524 9376 249576 9382
rect 249524 9318 249576 9324
rect 249338 9208 249394 9217
rect 249338 9143 249394 9152
rect 249352 8634 249380 9143
rect 249340 8628 249392 8634
rect 249340 8570 249392 8576
rect 249720 5370 249748 307022
rect 249904 296342 249932 311578
rect 251008 299538 251036 313890
rect 251468 309194 251496 319398
rect 251744 309602 251772 320062
rect 251732 309596 251784 309602
rect 251732 309538 251784 309544
rect 251272 309188 251324 309194
rect 251272 309130 251324 309136
rect 251456 309188 251508 309194
rect 251456 309130 251508 309136
rect 251088 307080 251140 307086
rect 251088 307022 251140 307028
rect 251284 307034 251312 309130
rect 250812 299532 250864 299538
rect 250812 299474 250864 299480
rect 250996 299532 251048 299538
rect 250996 299474 251048 299480
rect 249892 296336 249944 296342
rect 249892 296278 249944 296284
rect 250824 289882 250852 299474
rect 250904 296336 250956 296342
rect 250904 296278 250956 296284
rect 250812 289876 250864 289882
rect 250812 289818 250864 289824
rect 250810 240136 250866 240145
rect 250810 240071 250866 240080
rect 250824 230518 250852 240071
rect 250812 230512 250864 230518
rect 250812 230454 250864 230460
rect 250810 220824 250866 220833
rect 250810 220759 250866 220768
rect 250824 211177 250852 220759
rect 250810 211168 250866 211177
rect 250810 211103 250866 211112
rect 250812 182164 250864 182170
rect 250812 182106 250864 182112
rect 250824 172553 250852 182106
rect 250810 172544 250866 172553
rect 250810 172479 250866 172488
rect 250812 162852 250864 162858
rect 250812 162794 250864 162800
rect 250824 153241 250852 162794
rect 250810 153232 250866 153241
rect 250810 153167 250866 153176
rect 250812 19916 250864 19922
rect 250812 19858 250864 19864
rect 250824 12322 250852 19858
rect 250916 13598 250944 296278
rect 250996 289876 251048 289882
rect 250996 289818 251048 289824
rect 251008 270502 251036 289818
rect 250996 270496 251048 270502
rect 250996 270438 251048 270444
rect 250996 260908 251048 260914
rect 250996 260850 251048 260856
rect 251008 240145 251036 260850
rect 250994 240136 251050 240145
rect 250994 240071 251050 240080
rect 250996 230512 251048 230518
rect 250996 230454 251048 230460
rect 251008 220833 251036 230454
rect 250994 220824 251050 220833
rect 250994 220759 251050 220768
rect 250994 211168 251050 211177
rect 250994 211103 251050 211112
rect 251008 182170 251036 211103
rect 250996 182164 251048 182170
rect 250996 182106 251048 182112
rect 250994 172544 251050 172553
rect 250994 172479 251050 172488
rect 251008 162858 251036 172479
rect 250996 162852 251048 162858
rect 250996 162794 251048 162800
rect 250994 153232 251050 153241
rect 250994 153167 251050 153176
rect 251008 143546 251036 153167
rect 250996 143540 251048 143546
rect 250996 143482 251048 143488
rect 250994 133920 251050 133929
rect 250994 133855 251050 133864
rect 251008 46918 251036 133855
rect 250996 46912 251048 46918
rect 250996 46854 251048 46860
rect 250996 37324 251048 37330
rect 250996 37266 251048 37272
rect 251008 19922 251036 37266
rect 250996 19916 251048 19922
rect 250996 19858 251048 19864
rect 250904 13592 250956 13598
rect 250904 13534 250956 13540
rect 250824 12294 250944 12322
rect 250916 9654 250944 12294
rect 250352 9648 250404 9654
rect 250352 9590 250404 9596
rect 250904 9648 250956 9654
rect 250904 9590 250956 9596
rect 249798 8664 249854 8673
rect 249798 8599 249854 8608
rect 249708 5364 249760 5370
rect 249708 5306 249760 5312
rect 249248 4480 249300 4486
rect 249248 4422 249300 4428
rect 249812 3058 249840 8599
rect 249800 3052 249852 3058
rect 249800 2994 249852 3000
rect 250364 480 250392 9590
rect 251100 4690 251128 307022
rect 251284 307006 251404 307034
rect 251272 306944 251324 306950
rect 251272 306886 251324 306892
rect 251284 299470 251312 306886
rect 251272 299464 251324 299470
rect 251272 299406 251324 299412
rect 251376 297378 251404 307006
rect 251376 297350 252324 297378
rect 252192 297288 252244 297294
rect 252192 297230 252244 297236
rect 252098 240136 252154 240145
rect 252098 240071 252154 240080
rect 252112 230518 252140 240071
rect 252100 230512 252152 230518
rect 252100 230454 252152 230460
rect 252098 220824 252154 220833
rect 252098 220759 252154 220768
rect 252112 211177 252140 220759
rect 252098 211168 252154 211177
rect 252098 211103 252154 211112
rect 252100 182164 252152 182170
rect 252100 182106 252152 182112
rect 252112 172553 252140 182106
rect 252098 172544 252154 172553
rect 252098 172479 252154 172488
rect 252100 162852 252152 162858
rect 252100 162794 252152 162800
rect 252112 153241 252140 162794
rect 252098 153232 252154 153241
rect 252098 153167 252154 153176
rect 251180 143540 251232 143546
rect 251180 143482 251232 143488
rect 252100 143540 252152 143546
rect 252100 143482 252152 143488
rect 251192 133929 251220 143482
rect 252112 133929 252140 143482
rect 251178 133920 251234 133929
rect 251178 133855 251234 133864
rect 252098 133920 252154 133929
rect 252098 133855 252154 133864
rect 252100 95260 252152 95266
rect 252100 95202 252152 95208
rect 252112 87009 252140 95202
rect 252098 87000 252154 87009
rect 252098 86935 252154 86944
rect 252204 13530 252232 297230
rect 252296 270502 252324 297350
rect 252284 270496 252336 270502
rect 252284 270438 252336 270444
rect 252284 260908 252336 260914
rect 252284 260850 252336 260856
rect 252296 251190 252324 260850
rect 252284 251184 252336 251190
rect 252284 251126 252336 251132
rect 252284 241528 252336 241534
rect 252284 241470 252336 241476
rect 252296 240145 252324 241470
rect 252282 240136 252338 240145
rect 252282 240071 252338 240080
rect 252284 230512 252336 230518
rect 252284 230454 252336 230460
rect 252296 220833 252324 230454
rect 252282 220824 252338 220833
rect 252282 220759 252338 220768
rect 252282 211168 252338 211177
rect 252282 211103 252338 211112
rect 252296 201482 252324 211103
rect 252284 201476 252336 201482
rect 252284 201418 252336 201424
rect 252284 191888 252336 191894
rect 252284 191830 252336 191836
rect 252296 182170 252324 191830
rect 252284 182164 252336 182170
rect 252284 182106 252336 182112
rect 252282 172544 252338 172553
rect 252282 172479 252338 172488
rect 252296 162858 252324 172479
rect 252284 162852 252336 162858
rect 252284 162794 252336 162800
rect 252282 153232 252338 153241
rect 252282 153167 252338 153176
rect 252296 143546 252324 153167
rect 252284 143540 252336 143546
rect 252284 143482 252336 143488
rect 252282 133920 252338 133929
rect 252282 133855 252338 133864
rect 252296 124166 252324 133855
rect 252284 124160 252336 124166
rect 252284 124102 252336 124108
rect 252284 114572 252336 114578
rect 252284 114514 252336 114520
rect 252296 104854 252324 114514
rect 252284 104848 252336 104854
rect 252284 104790 252336 104796
rect 252282 87000 252338 87009
rect 252282 86935 252338 86944
rect 252296 85542 252324 86935
rect 252284 85536 252336 85542
rect 252284 85478 252336 85484
rect 252284 75948 252336 75954
rect 252284 75890 252336 75896
rect 252296 66230 252324 75890
rect 252284 66224 252336 66230
rect 252284 66166 252336 66172
rect 252284 56636 252336 56642
rect 252284 56578 252336 56584
rect 252296 46918 252324 56578
rect 252284 46912 252336 46918
rect 252284 46854 252336 46860
rect 252284 37324 252336 37330
rect 252284 37266 252336 37272
rect 252192 13524 252244 13530
rect 252192 13466 252244 13472
rect 252296 12458 252324 37266
rect 252112 12430 252324 12458
rect 252112 12322 252140 12430
rect 252112 12294 252232 12322
rect 252204 9586 252232 12294
rect 252192 9580 252244 9586
rect 252192 9522 252244 9528
rect 252388 5506 252416 320076
rect 252940 320062 253230 320090
rect 253400 320062 253690 320090
rect 252468 316192 252520 316198
rect 252468 316134 252520 316140
rect 252376 5500 252428 5506
rect 252376 5442 252428 5448
rect 251456 5160 251508 5166
rect 251456 5102 251508 5108
rect 251088 4684 251140 4690
rect 251088 4626 251140 4632
rect 251468 480 251496 5102
rect 252480 5030 252508 316134
rect 252560 315988 252612 315994
rect 252560 315930 252612 315936
rect 252572 307086 252600 315930
rect 252940 309233 252968 320062
rect 253400 315994 253428 320062
rect 253388 315988 253440 315994
rect 253388 315930 253440 315936
rect 252926 309224 252982 309233
rect 252926 309159 252982 309168
rect 252742 309088 252798 309097
rect 252742 309023 252798 309032
rect 252560 307080 252612 307086
rect 252560 307022 252612 307028
rect 252756 294642 252784 309023
rect 252744 294636 252796 294642
rect 252744 294578 252796 294584
rect 253664 294636 253716 294642
rect 253664 294578 253716 294584
rect 253676 13462 253704 294578
rect 253664 13456 253716 13462
rect 253664 13398 253716 13404
rect 253664 11076 253716 11082
rect 253664 11018 253716 11024
rect 252652 9308 252704 9314
rect 252652 9250 252704 9256
rect 252468 5024 252520 5030
rect 252468 4966 252520 4972
rect 252664 480 252692 9250
rect 253676 5438 253704 11018
rect 253768 9518 253796 320146
rect 253860 319410 253888 320198
rect 255964 320146 256016 320152
rect 256332 320204 256384 320210
rect 256332 320146 256384 320152
rect 258000 320198 258198 320226
rect 260484 320198 260682 320226
rect 261588 320210 261878 320226
rect 260840 320204 260892 320210
rect 254136 320062 254518 320090
rect 254886 320062 255176 320090
rect 255346 320062 255452 320090
rect 253860 319382 253980 319410
rect 253952 307086 253980 319382
rect 254136 309210 254164 320062
rect 255148 316010 255176 320062
rect 255148 315982 255268 316010
rect 254044 309182 254164 309210
rect 254044 309126 254072 309182
rect 254032 309120 254084 309126
rect 254032 309062 254084 309068
rect 253848 307080 253900 307086
rect 253848 307022 253900 307028
rect 253940 307080 253992 307086
rect 253940 307022 253992 307028
rect 255136 307080 255188 307086
rect 255136 307022 255188 307028
rect 253860 11082 253888 307022
rect 255044 299532 255096 299538
rect 255044 299474 255096 299480
rect 255056 13394 255084 299474
rect 255044 13388 255096 13394
rect 255044 13330 255096 13336
rect 255148 13122 255176 307022
rect 255240 299538 255268 315982
rect 255320 315036 255372 315042
rect 255320 314978 255372 314984
rect 255332 307154 255360 314978
rect 255320 307148 255372 307154
rect 255320 307090 255372 307096
rect 255424 307086 255452 320062
rect 255792 320062 256174 320090
rect 255792 316010 255820 320062
rect 255516 315982 255820 316010
rect 255412 307080 255464 307086
rect 255412 307022 255464 307028
rect 255516 307018 255544 315982
rect 255504 307012 255556 307018
rect 255504 306954 255556 306960
rect 255228 299532 255280 299538
rect 255228 299474 255280 299480
rect 255228 298172 255280 298178
rect 255228 298114 255280 298120
rect 255240 298042 255268 298114
rect 255228 298036 255280 298042
rect 255228 297978 255280 297984
rect 255228 288448 255280 288454
rect 255228 288390 255280 288396
rect 255240 278769 255268 288390
rect 255226 278760 255282 278769
rect 255226 278695 255282 278704
rect 255318 278624 255374 278633
rect 255318 278559 255374 278568
rect 255332 269142 255360 278559
rect 255228 269136 255280 269142
rect 255228 269078 255280 269084
rect 255320 269136 255372 269142
rect 255320 269078 255372 269084
rect 255240 240174 255268 269078
rect 255228 240168 255280 240174
rect 255228 240110 255280 240116
rect 255320 240168 255372 240174
rect 255320 240110 255372 240116
rect 255332 230518 255360 240110
rect 255228 230512 255280 230518
rect 255228 230454 255280 230460
rect 255320 230512 255372 230518
rect 255320 230454 255372 230460
rect 255240 229090 255268 230454
rect 255228 229084 255280 229090
rect 255228 229026 255280 229032
rect 255504 229084 255556 229090
rect 255504 229026 255556 229032
rect 255516 219473 255544 229026
rect 255318 219464 255374 219473
rect 255318 219399 255374 219408
rect 255502 219464 255558 219473
rect 255502 219399 255558 219408
rect 255332 211206 255360 219399
rect 255320 211200 255372 211206
rect 255320 211142 255372 211148
rect 255596 211064 255648 211070
rect 255596 211006 255648 211012
rect 255608 206242 255636 211006
rect 255412 206236 255464 206242
rect 255412 206178 255464 206184
rect 255596 206236 255648 206242
rect 255596 206178 255648 206184
rect 255424 190534 255452 206178
rect 255320 190528 255372 190534
rect 255320 190470 255372 190476
rect 255412 190528 255464 190534
rect 255412 190470 255464 190476
rect 255332 182186 255360 190470
rect 255332 182158 255452 182186
rect 255424 171154 255452 182158
rect 255320 171148 255372 171154
rect 255320 171090 255372 171096
rect 255412 171148 255464 171154
rect 255412 171090 255464 171096
rect 255332 162874 255360 171090
rect 255332 162846 255452 162874
rect 255424 153241 255452 162846
rect 255226 153232 255282 153241
rect 255226 153167 255282 153176
rect 255410 153232 255466 153241
rect 255410 153167 255466 153176
rect 255240 143449 255268 153167
rect 255226 143440 255282 143449
rect 255226 143375 255282 143384
rect 255410 133920 255466 133929
rect 255410 133855 255466 133864
rect 255424 125633 255452 133855
rect 255226 125624 255282 125633
rect 255226 125559 255282 125568
rect 255410 125624 255466 125633
rect 255410 125559 255466 125568
rect 255240 124166 255268 125559
rect 255228 124160 255280 124166
rect 255228 124102 255280 124108
rect 255228 106344 255280 106350
rect 255228 106286 255280 106292
rect 255240 104854 255268 106286
rect 255228 104848 255280 104854
rect 255228 104790 255280 104796
rect 255228 87032 255280 87038
rect 255228 86974 255280 86980
rect 255240 85542 255268 86974
rect 255228 85536 255280 85542
rect 255228 85478 255280 85484
rect 255228 75948 255280 75954
rect 255228 75890 255280 75896
rect 255240 66230 255268 75890
rect 255228 66224 255280 66230
rect 255228 66166 255280 66172
rect 255228 56636 255280 56642
rect 255228 56578 255280 56584
rect 255240 46918 255268 56578
rect 255228 46912 255280 46918
rect 255228 46854 255280 46860
rect 255228 37324 255280 37330
rect 255228 37266 255280 37272
rect 255240 27606 255268 37266
rect 255228 27600 255280 27606
rect 255228 27542 255280 27548
rect 255228 18012 255280 18018
rect 255228 17954 255280 17960
rect 255136 13116 255188 13122
rect 255136 13058 255188 13064
rect 255240 12458 255268 17954
rect 256344 13326 256372 320146
rect 256542 320062 256648 320090
rect 256620 318850 256648 320062
rect 256424 318844 256476 318850
rect 256424 318786 256476 318792
rect 256608 318844 256660 318850
rect 256608 318786 256660 318792
rect 256436 315042 256464 318786
rect 256988 316130 257016 320076
rect 257080 320062 257370 320090
rect 257448 320062 257830 320090
rect 256976 316124 257028 316130
rect 256976 316066 257028 316072
rect 257080 316010 257108 320062
rect 256712 315982 257108 316010
rect 256424 315036 256476 315042
rect 256424 314978 256476 314984
rect 256516 307148 256568 307154
rect 256516 307090 256568 307096
rect 256424 307080 256476 307086
rect 256424 307022 256476 307028
rect 256332 13320 256384 13326
rect 256332 13262 256384 13268
rect 255240 12430 255360 12458
rect 255332 12322 255360 12430
rect 255056 12294 255360 12322
rect 253848 11076 253900 11082
rect 253848 11018 253900 11024
rect 253756 9512 253808 9518
rect 253756 9454 253808 9460
rect 253848 9444 253900 9450
rect 253848 9386 253900 9392
rect 253664 5432 253716 5438
rect 253664 5374 253716 5380
rect 253860 480 253888 9386
rect 255056 9058 255084 12294
rect 255136 11076 255188 11082
rect 255136 11018 255188 11024
rect 255148 9178 255176 11018
rect 256436 9450 256464 307022
rect 256424 9444 256476 9450
rect 256424 9386 256476 9392
rect 256528 9314 256556 307090
rect 256712 307086 256740 315982
rect 257448 315042 257476 320062
rect 258000 319410 258028 320198
rect 258658 320062 258856 320090
rect 259026 320062 259224 320090
rect 259486 320062 259592 320090
rect 258000 319382 258120 319410
rect 257804 316124 257856 316130
rect 257804 316066 257856 316072
rect 257436 315036 257488 315042
rect 257436 314978 257488 314984
rect 256700 307080 256752 307086
rect 256700 307022 256752 307028
rect 256608 307012 256660 307018
rect 256608 306954 256660 306960
rect 256516 9308 256568 9314
rect 256516 9250 256568 9256
rect 256240 9240 256292 9246
rect 256240 9182 256292 9188
rect 255136 9172 255188 9178
rect 255136 9114 255188 9120
rect 255056 9030 255176 9058
rect 255042 5400 255098 5409
rect 255042 5335 255098 5344
rect 255056 480 255084 5335
rect 255148 5166 255176 9030
rect 255136 5160 255188 5166
rect 255136 5102 255188 5108
rect 256252 480 256280 9182
rect 256620 5302 256648 306954
rect 256698 15192 256754 15201
rect 256698 15127 256754 15136
rect 256712 14793 256740 15127
rect 256698 14784 256754 14793
rect 256698 14719 256754 14728
rect 257816 13258 257844 316066
rect 257896 315036 257948 315042
rect 257896 314978 257948 314984
rect 257804 13252 257856 13258
rect 257804 13194 257856 13200
rect 257908 9246 257936 314978
rect 257988 307080 258040 307086
rect 258092 307068 258120 319382
rect 258828 315994 258856 320062
rect 259196 318730 259224 320062
rect 259196 318702 259316 318730
rect 258816 315988 258868 315994
rect 258816 315930 258868 315936
rect 259288 309194 259316 318702
rect 259368 315988 259420 315994
rect 259368 315930 259420 315936
rect 259460 315988 259512 315994
rect 259460 315930 259512 315936
rect 259184 309188 259236 309194
rect 259184 309130 259236 309136
rect 259276 309188 259328 309194
rect 259276 309130 259328 309136
rect 258092 307040 258212 307068
rect 257988 307022 258040 307028
rect 257804 9240 257856 9246
rect 257804 9182 257856 9188
rect 257896 9240 257948 9246
rect 257896 9182 257948 9188
rect 256608 5296 256660 5302
rect 256608 5238 256660 5244
rect 257436 4616 257488 4622
rect 257436 4558 257488 4564
rect 257448 480 257476 4558
rect 257816 3126 257844 9182
rect 258000 5234 258028 307022
rect 258184 297378 258212 307040
rect 259196 302326 259224 309130
rect 259184 302320 259236 302326
rect 259184 302262 259236 302268
rect 259184 302184 259236 302190
rect 259184 302126 259236 302132
rect 259196 297498 259224 302126
rect 259184 297492 259236 297498
rect 259184 297434 259236 297440
rect 258184 297350 259224 297378
rect 259090 240136 259146 240145
rect 259090 240071 259146 240080
rect 259104 230518 259132 240071
rect 259092 230512 259144 230518
rect 259092 230454 259144 230460
rect 259090 220824 259146 220833
rect 259090 220759 259146 220768
rect 259104 211177 259132 220759
rect 259090 211168 259146 211177
rect 259090 211103 259146 211112
rect 259092 182164 259144 182170
rect 259092 182106 259144 182112
rect 259104 172553 259132 182106
rect 259090 172544 259146 172553
rect 259090 172479 259146 172488
rect 259092 162852 259144 162858
rect 259092 162794 259144 162800
rect 259104 153241 259132 162794
rect 259090 153232 259146 153241
rect 259090 153167 259146 153176
rect 259092 143540 259144 143546
rect 259092 143482 259144 143488
rect 259104 125633 259132 143482
rect 259090 125624 259146 125633
rect 259090 125559 259146 125568
rect 259092 114572 259144 114578
rect 259092 114514 259144 114520
rect 259104 106321 259132 114514
rect 259090 106312 259146 106321
rect 259090 106247 259146 106256
rect 259196 22778 259224 297350
rect 259276 289876 259328 289882
rect 259276 289818 259328 289824
rect 259288 270502 259316 289818
rect 259276 270496 259328 270502
rect 259276 270438 259328 270444
rect 259276 260908 259328 260914
rect 259276 260850 259328 260856
rect 259288 240145 259316 260850
rect 259274 240136 259330 240145
rect 259274 240071 259330 240080
rect 259276 230512 259328 230518
rect 259276 230454 259328 230460
rect 259288 220833 259316 230454
rect 259274 220824 259330 220833
rect 259274 220759 259330 220768
rect 259274 211168 259330 211177
rect 259274 211103 259330 211112
rect 259288 182170 259316 211103
rect 259276 182164 259328 182170
rect 259276 182106 259328 182112
rect 259274 172544 259330 172553
rect 259274 172479 259330 172488
rect 259288 162858 259316 172479
rect 259276 162852 259328 162858
rect 259276 162794 259328 162800
rect 259274 153232 259330 153241
rect 259274 153167 259330 153176
rect 259288 143546 259316 153167
rect 259276 143540 259328 143546
rect 259276 143482 259328 143488
rect 259274 125624 259330 125633
rect 259274 125559 259330 125568
rect 259288 114578 259316 125559
rect 259276 114572 259328 114578
rect 259276 114514 259328 114520
rect 259274 106312 259330 106321
rect 259274 106247 259330 106256
rect 259288 104854 259316 106247
rect 259276 104848 259328 104854
rect 259276 104790 259328 104796
rect 259276 95260 259328 95266
rect 259276 95202 259328 95208
rect 259288 85542 259316 95202
rect 259276 85536 259328 85542
rect 259276 85478 259328 85484
rect 259276 75948 259328 75954
rect 259276 75890 259328 75896
rect 259288 66230 259316 75890
rect 259276 66224 259328 66230
rect 259276 66166 259328 66172
rect 259276 56636 259328 56642
rect 259276 56578 259328 56584
rect 259288 46918 259316 56578
rect 259276 46912 259328 46918
rect 259276 46854 259328 46860
rect 259276 37324 259328 37330
rect 259276 37266 259328 37272
rect 259184 22772 259236 22778
rect 259184 22714 259236 22720
rect 259288 13002 259316 37266
rect 259196 12974 259316 13002
rect 259196 9625 259224 12974
rect 259380 12322 259408 315930
rect 259472 307018 259500 315930
rect 259460 307012 259512 307018
rect 259460 306954 259512 306960
rect 259564 302122 259592 320062
rect 259656 320062 259854 320090
rect 260024 320062 260314 320090
rect 259656 307086 259684 320062
rect 260024 315994 260052 320062
rect 260484 319410 260512 320198
rect 260840 320146 260892 320152
rect 261576 320204 261878 320210
rect 261628 320198 261878 320204
rect 263336 320198 263534 320226
rect 264072 320210 264362 320226
rect 263600 320204 263652 320210
rect 261576 320146 261628 320152
rect 260484 319382 260604 319410
rect 260012 315988 260064 315994
rect 260012 315930 260064 315936
rect 259644 307080 259696 307086
rect 259644 307022 259696 307028
rect 259552 302116 259604 302122
rect 259552 302058 259604 302064
rect 260472 302116 260524 302122
rect 260472 302058 260524 302064
rect 260484 190466 260512 302058
rect 260288 190460 260340 190466
rect 260288 190402 260340 190408
rect 260472 190460 260524 190466
rect 260472 190402 260524 190408
rect 260300 180849 260328 190402
rect 260286 180840 260342 180849
rect 260286 180775 260342 180784
rect 260470 180840 260526 180849
rect 260470 180775 260526 180784
rect 260484 26246 260512 180775
rect 260472 26240 260524 26246
rect 260472 26182 260524 26188
rect 260576 13705 260604 319382
rect 260748 307080 260800 307086
rect 260852 307068 260880 320146
rect 261050 320062 261340 320090
rect 261510 320062 261616 320090
rect 261312 315994 261340 320062
rect 261588 318850 261616 320062
rect 261576 318844 261628 318850
rect 261576 318786 261628 318792
rect 261668 318844 261720 318850
rect 261668 318786 261720 318792
rect 261300 315988 261352 315994
rect 261300 315930 261352 315936
rect 261680 313936 261708 318786
rect 262324 315994 262352 320076
rect 262508 320062 262706 320090
rect 262784 320062 263166 320090
rect 262128 315988 262180 315994
rect 262128 315930 262180 315936
rect 262312 315988 262364 315994
rect 262312 315930 262364 315936
rect 261680 313908 261800 313936
rect 261772 309074 261800 313908
rect 261772 309046 262076 309074
rect 260852 307040 260972 307068
rect 260748 307022 260800 307028
rect 260656 307012 260708 307018
rect 260656 306954 260708 306960
rect 260562 13696 260618 13705
rect 260562 13631 260618 13640
rect 259288 12294 259408 12322
rect 259182 9616 259238 9625
rect 259182 9551 259238 9560
rect 258630 5264 258686 5273
rect 257988 5228 258040 5234
rect 258630 5199 258686 5208
rect 257988 5170 258040 5176
rect 257804 3120 257856 3126
rect 257804 3062 257856 3068
rect 258644 480 258672 5199
rect 259288 4894 259316 12294
rect 260668 9178 260696 306954
rect 259828 9172 259880 9178
rect 259828 9114 259880 9120
rect 260656 9172 260708 9178
rect 260656 9114 260708 9120
rect 259276 4888 259328 4894
rect 259276 4830 259328 4836
rect 259840 480 259868 9114
rect 260760 5166 260788 307022
rect 260944 297378 260972 307040
rect 260944 297350 261984 297378
rect 261956 13569 261984 297350
rect 262048 66230 262076 309046
rect 262036 66224 262088 66230
rect 262036 66166 262088 66172
rect 262036 49428 262088 49434
rect 262036 49370 262088 49376
rect 262048 33250 262076 49370
rect 262036 33244 262088 33250
rect 262036 33186 262088 33192
rect 262036 29708 262088 29714
rect 262036 29650 262088 29656
rect 262048 23390 262076 29650
rect 262036 23384 262088 23390
rect 262036 23326 262088 23332
rect 261942 13560 261998 13569
rect 261942 13495 261998 13504
rect 260748 5160 260800 5166
rect 260748 5102 260800 5108
rect 262140 5030 262168 315930
rect 262404 315784 262456 315790
rect 262404 315726 262456 315732
rect 262312 312792 262364 312798
rect 262312 312734 262364 312740
rect 262220 312724 262272 312730
rect 262220 312666 262272 312672
rect 262232 307086 262260 312666
rect 262220 307080 262272 307086
rect 262220 307022 262272 307028
rect 262324 306066 262352 312734
rect 262416 307018 262444 315726
rect 262508 312730 262536 320062
rect 262784 312798 262812 320062
rect 263336 319410 263364 320198
rect 263600 320146 263652 320152
rect 264060 320204 264362 320210
rect 264112 320198 264362 320204
rect 266478 320210 266676 320226
rect 266478 320204 266688 320210
rect 266478 320198 266636 320204
rect 264060 320146 264112 320152
rect 266636 320146 266688 320152
rect 263336 319382 263456 319410
rect 262772 312792 262824 312798
rect 262772 312734 262824 312740
rect 262496 312724 262548 312730
rect 262496 312666 262548 312672
rect 263324 307080 263376 307086
rect 263324 307022 263376 307028
rect 262404 307012 262456 307018
rect 262404 306954 262456 306960
rect 262312 306060 262364 306066
rect 262312 306002 262364 306008
rect 263232 306060 263284 306066
rect 263232 306002 263284 306008
rect 262220 66224 262272 66230
rect 262220 66166 262272 66172
rect 262232 49434 262260 66166
rect 262220 49428 262272 49434
rect 262220 49370 262272 49376
rect 262220 23384 262272 23390
rect 262220 23326 262272 23332
rect 262232 13841 262260 23326
rect 262218 13832 262274 13841
rect 262218 13767 262274 13776
rect 262402 13832 262458 13841
rect 262402 13767 262458 13776
rect 262416 9489 262444 13767
rect 263244 13433 263272 306002
rect 263230 13424 263286 13433
rect 263230 13359 263286 13368
rect 263336 13274 263364 307022
rect 263244 13246 263364 13274
rect 262402 9480 262458 9489
rect 262402 9415 262458 9424
rect 263244 9353 263272 13246
rect 263230 9344 263286 9353
rect 263230 9279 263286 9288
rect 263428 8786 263456 319382
rect 263612 307034 263640 320146
rect 263994 320062 264192 320090
rect 264822 320062 264928 320090
rect 265190 320062 265296 320090
rect 264164 313954 264192 320062
rect 264152 313948 264204 313954
rect 264152 313890 264204 313896
rect 264704 313948 264756 313954
rect 264704 313890 264756 313896
rect 264716 309126 264744 313890
rect 264704 309120 264756 309126
rect 264704 309062 264756 309068
rect 264796 309052 264848 309058
rect 264796 308994 264848 309000
rect 263508 307012 263560 307018
rect 263612 307006 263732 307034
rect 263508 306954 263560 306960
rect 263244 8758 263456 8786
rect 263244 5273 263272 8758
rect 263416 6996 263468 7002
rect 263416 6938 263468 6944
rect 263230 5264 263286 5273
rect 263230 5199 263286 5208
rect 262218 5128 262274 5137
rect 262218 5063 262274 5072
rect 261024 5024 261076 5030
rect 261024 4966 261076 4972
rect 262128 5024 262180 5030
rect 262128 4966 262180 4972
rect 261036 480 261064 4966
rect 262232 480 262260 5063
rect 263428 480 263456 6938
rect 263520 5409 263548 306954
rect 263704 294001 263732 307006
rect 263690 293992 263746 294001
rect 263690 293927 263746 293936
rect 264702 293992 264758 294001
rect 264702 293927 264758 293936
rect 264716 284306 264744 293927
rect 264520 284300 264572 284306
rect 264520 284242 264572 284248
rect 264704 284300 264756 284306
rect 264704 284242 264756 284248
rect 264532 274689 264560 284242
rect 264518 274680 264574 274689
rect 264518 274615 264574 274624
rect 264702 274680 264758 274689
rect 264702 274615 264704 274624
rect 264756 274615 264758 274624
rect 264704 274586 264756 274592
rect 264612 264988 264664 264994
rect 264612 264930 264664 264936
rect 264624 192574 264652 264930
rect 264612 192568 264664 192574
rect 264612 192510 264664 192516
rect 264612 185700 264664 185706
rect 264612 185642 264664 185648
rect 264624 180826 264652 185642
rect 264624 180798 264744 180826
rect 264716 169810 264744 180798
rect 264624 169782 264744 169810
rect 264624 169726 264652 169782
rect 264612 169720 264664 169726
rect 264612 169662 264664 169668
rect 264612 160132 264664 160138
rect 264612 160074 264664 160080
rect 264624 160018 264652 160074
rect 264532 159990 264652 160018
rect 264532 150482 264560 159990
rect 264520 150476 264572 150482
rect 264520 150418 264572 150424
rect 264612 150476 264664 150482
rect 264612 150418 264664 150424
rect 264624 150362 264652 150418
rect 264532 150334 264652 150362
rect 264532 140826 264560 150334
rect 264808 143546 264836 308994
rect 264796 143540 264848 143546
rect 264796 143482 264848 143488
rect 264520 140820 264572 140826
rect 264520 140762 264572 140768
rect 264612 140820 264664 140826
rect 264612 140762 264664 140768
rect 264624 140706 264652 140762
rect 264532 140678 264652 140706
rect 264532 131170 264560 140678
rect 264794 133920 264850 133929
rect 264794 133855 264850 133864
rect 264520 131164 264572 131170
rect 264520 131106 264572 131112
rect 264612 131164 264664 131170
rect 264612 131106 264664 131112
rect 264624 131050 264652 131106
rect 264532 131022 264652 131050
rect 264532 121514 264560 131022
rect 264520 121508 264572 121514
rect 264520 121450 264572 121456
rect 264612 121508 264664 121514
rect 264612 121450 264664 121456
rect 264624 121394 264652 121450
rect 264532 121366 264652 121394
rect 264532 111858 264560 121366
rect 264520 111852 264572 111858
rect 264520 111794 264572 111800
rect 264612 111852 264664 111858
rect 264612 111794 264664 111800
rect 264624 111722 264652 111794
rect 264612 111716 264664 111722
rect 264612 111658 264664 111664
rect 264612 102196 264664 102202
rect 264612 102138 264664 102144
rect 264624 102082 264652 102138
rect 264532 102054 264652 102082
rect 264532 92546 264560 102054
rect 264520 92540 264572 92546
rect 264520 92482 264572 92488
rect 264612 92540 264664 92546
rect 264612 92482 264664 92488
rect 264624 92410 264652 92482
rect 264612 92404 264664 92410
rect 264612 92346 264664 92352
rect 264612 82884 264664 82890
rect 264612 82826 264664 82832
rect 264624 82770 264652 82826
rect 264532 82742 264652 82770
rect 264532 73234 264560 82742
rect 264520 73228 264572 73234
rect 264520 73170 264572 73176
rect 264612 73228 264664 73234
rect 264612 73170 264664 73176
rect 264624 53786 264652 73170
rect 264612 53780 264664 53786
rect 264612 53722 264664 53728
rect 264612 44328 264664 44334
rect 264612 44270 264664 44276
rect 264624 33250 264652 44270
rect 264428 33244 264480 33250
rect 264428 33186 264480 33192
rect 264612 33244 264664 33250
rect 264612 33186 264664 33192
rect 264440 24886 264468 33186
rect 264428 24880 264480 24886
rect 264428 24822 264480 24828
rect 264704 24880 264756 24886
rect 264704 24822 264756 24828
rect 264716 15201 264744 24822
rect 264702 15192 264758 15201
rect 264702 15127 264758 15136
rect 264808 9217 264836 133855
rect 264794 9208 264850 9217
rect 264794 9143 264850 9152
rect 263506 5400 263562 5409
rect 263506 5335 263562 5344
rect 264900 5098 264928 320062
rect 265268 315994 265296 320062
rect 265360 320062 265650 320090
rect 266018 320062 266308 320090
rect 265256 315988 265308 315994
rect 265256 315930 265308 315936
rect 265360 314673 265388 320062
rect 266084 315988 266136 315994
rect 266084 315930 266136 315936
rect 265346 314664 265402 314673
rect 265346 314599 265402 314608
rect 265806 314664 265862 314673
rect 265806 314599 265862 314608
rect 265820 302190 265848 314599
rect 265808 302184 265860 302190
rect 265808 302126 265860 302132
rect 266096 299538 266124 315930
rect 266084 299532 266136 299538
rect 266084 299474 266136 299480
rect 266176 299532 266228 299538
rect 266176 299474 266228 299480
rect 265900 292664 265952 292670
rect 265900 292606 265952 292612
rect 265912 292534 265940 292606
rect 265900 292528 265952 292534
rect 265900 292470 265952 292476
rect 265992 292460 266044 292466
rect 265992 292402 266044 292408
rect 266004 230518 266032 292402
rect 265992 230512 266044 230518
rect 265992 230454 266044 230460
rect 265992 218068 266044 218074
rect 265992 218010 266044 218016
rect 266004 181014 266032 218010
rect 265992 181008 266044 181014
rect 265992 180950 266044 180956
rect 265992 180872 266044 180878
rect 265992 180814 266044 180820
rect 266004 179382 266032 180814
rect 265992 179376 266044 179382
rect 265992 179318 266044 179324
rect 265992 169788 266044 169794
rect 265992 169730 266044 169736
rect 266004 160070 266032 169730
rect 265992 160064 266044 160070
rect 265992 160006 266044 160012
rect 265992 150476 266044 150482
rect 265992 150418 266044 150424
rect 264980 143540 265032 143546
rect 264980 143482 265032 143488
rect 264992 133929 265020 143482
rect 266004 140758 266032 150418
rect 265992 140752 266044 140758
rect 265992 140694 266044 140700
rect 264978 133920 265034 133929
rect 264978 133855 265034 133864
rect 265992 131164 266044 131170
rect 265992 131106 266044 131112
rect 266004 121446 266032 131106
rect 265992 121440 266044 121446
rect 265992 121382 266044 121388
rect 265992 111852 266044 111858
rect 265992 111794 266044 111800
rect 266004 102134 266032 111794
rect 265992 102128 266044 102134
rect 265992 102070 266044 102076
rect 265992 92540 266044 92546
rect 265992 92482 266044 92488
rect 266004 82822 266032 92482
rect 265992 82816 266044 82822
rect 265992 82758 266044 82764
rect 265992 73228 266044 73234
rect 265992 73170 266044 73176
rect 266004 35850 266032 73170
rect 266004 35822 266124 35850
rect 265162 15056 265218 15065
rect 265162 14991 265218 15000
rect 265176 13297 265204 14991
rect 265162 13288 265218 13297
rect 265162 13223 265218 13232
rect 266096 13161 266124 35822
rect 266082 13152 266138 13161
rect 266082 13087 266138 13096
rect 266188 13002 266216 299474
rect 266096 12974 266216 13002
rect 266096 9602 266124 12974
rect 266096 9574 266216 9602
rect 266188 9081 266216 9574
rect 266174 9072 266230 9081
rect 266174 9007 266230 9016
rect 266280 5137 266308 320062
rect 266556 320062 266846 320090
rect 266924 320062 267306 320090
rect 266452 315920 266504 315926
rect 266452 315862 266504 315868
rect 266464 307018 266492 315862
rect 266452 307012 266504 307018
rect 266452 306954 266504 306960
rect 266556 306406 266584 320062
rect 266924 317422 266952 320062
rect 267384 319462 267412 320334
rect 269868 320210 270158 320226
rect 267464 320204 267516 320210
rect 267464 320146 267516 320152
rect 269120 320204 269172 320210
rect 269120 320146 269172 320152
rect 269856 320204 270158 320210
rect 269908 320198 270158 320204
rect 269856 320146 269908 320152
rect 267372 319456 267424 319462
rect 267372 319398 267424 319404
rect 266912 317416 266964 317422
rect 266912 317358 266964 317364
rect 266544 306400 266596 306406
rect 266544 306342 266596 306348
rect 267096 306400 267148 306406
rect 267096 306342 267148 306348
rect 267108 303618 267136 306342
rect 267096 303612 267148 303618
rect 267096 303554 267148 303560
rect 267096 299464 267148 299470
rect 267096 299406 267148 299412
rect 267108 293978 267136 299406
rect 267108 293950 267228 293978
rect 267200 287774 267228 293950
rect 267188 287768 267240 287774
rect 267188 287710 267240 287716
rect 267280 282940 267332 282946
rect 267280 282882 267332 282888
rect 267292 186454 267320 282882
rect 267280 186448 267332 186454
rect 267280 186390 267332 186396
rect 267096 186380 267148 186386
rect 267096 186322 267148 186328
rect 267108 180849 267136 186322
rect 267094 180840 267150 180849
rect 267094 180775 267150 180784
rect 267278 180840 267334 180849
rect 267278 180775 267334 180784
rect 267292 179382 267320 180775
rect 267280 179376 267332 179382
rect 267280 179318 267332 179324
rect 267280 169788 267332 169794
rect 267280 169730 267332 169736
rect 267292 160070 267320 169730
rect 267280 160064 267332 160070
rect 267280 160006 267332 160012
rect 267280 150476 267332 150482
rect 267280 150418 267332 150424
rect 267292 140758 267320 150418
rect 267280 140752 267332 140758
rect 267280 140694 267332 140700
rect 267280 131164 267332 131170
rect 267280 131106 267332 131112
rect 267292 121446 267320 131106
rect 267280 121440 267332 121446
rect 267280 121382 267332 121388
rect 267280 111852 267332 111858
rect 267280 111794 267332 111800
rect 267292 102134 267320 111794
rect 267280 102128 267332 102134
rect 267280 102070 267332 102076
rect 267280 92540 267332 92546
rect 267280 92482 267332 92488
rect 267292 82822 267320 92482
rect 267280 82816 267332 82822
rect 267280 82758 267332 82764
rect 267280 73228 267332 73234
rect 267280 73170 267332 73176
rect 267292 63510 267320 73170
rect 267280 63504 267332 63510
rect 267280 63446 267332 63452
rect 267280 53848 267332 53854
rect 267280 53790 267332 53796
rect 267292 44130 267320 53790
rect 267280 44124 267332 44130
rect 267280 44066 267332 44072
rect 267372 35828 267424 35834
rect 267372 35770 267424 35776
rect 267384 13025 267412 35770
rect 267370 13016 267426 13025
rect 267370 12951 267426 12960
rect 267476 9110 267504 320146
rect 267556 319456 267608 319462
rect 267556 319398 267608 319404
rect 267568 315926 267596 319398
rect 267648 317416 267700 317422
rect 267648 317358 267700 317364
rect 267740 317416 267792 317422
rect 267740 317358 267792 317364
rect 267556 315920 267608 315926
rect 267556 315862 267608 315868
rect 267556 307012 267608 307018
rect 267556 306954 267608 306960
rect 267372 9104 267424 9110
rect 267372 9046 267424 9052
rect 267464 9104 267516 9110
rect 267464 9046 267516 9052
rect 267004 9036 267056 9042
rect 267004 8978 267056 8984
rect 266266 5128 266322 5137
rect 264612 5092 264664 5098
rect 264612 5034 264664 5040
rect 264888 5092 264940 5098
rect 266266 5063 266322 5072
rect 264888 5034 264940 5040
rect 264624 480 264652 5034
rect 265806 4992 265862 5001
rect 265806 4927 265862 4936
rect 265820 480 265848 4927
rect 267016 480 267044 8978
rect 267384 3194 267412 9046
rect 267568 9042 267596 306954
rect 267556 9036 267608 9042
rect 267556 8978 267608 8984
rect 267660 5001 267688 317358
rect 267752 307086 267780 317358
rect 268120 314702 268148 320076
rect 268502 320062 268792 320090
rect 268764 316010 268792 320062
rect 268948 317422 268976 320076
rect 268936 317416 268988 317422
rect 268936 317358 268988 317364
rect 268764 315982 269068 316010
rect 267832 314696 267884 314702
rect 267832 314638 267884 314644
rect 268108 314696 268160 314702
rect 268108 314638 268160 314644
rect 267740 307080 267792 307086
rect 267740 307022 267792 307028
rect 267844 299538 267872 314638
rect 269040 307170 269068 315982
rect 268856 307142 269068 307170
rect 267832 299532 267884 299538
rect 267832 299474 267884 299480
rect 268752 299532 268804 299538
rect 268752 299474 268804 299480
rect 268764 277386 268792 299474
rect 268856 297430 268884 307142
rect 268936 307080 268988 307086
rect 268936 307022 268988 307028
rect 268844 297424 268896 297430
rect 268844 297366 268896 297372
rect 268844 287768 268896 287774
rect 268844 287710 268896 287716
rect 268856 278118 268884 287710
rect 268844 278112 268896 278118
rect 268844 278054 268896 278060
rect 268672 277358 268792 277386
rect 268672 273290 268700 277358
rect 268660 273284 268712 273290
rect 268660 273226 268712 273232
rect 268752 268252 268804 268258
rect 268752 268194 268804 268200
rect 268660 267776 268712 267782
rect 268660 267718 268712 267724
rect 268672 258482 268700 267718
rect 268764 258806 268792 268194
rect 268752 258800 268804 258806
rect 268752 258742 268804 258748
rect 268672 258454 268884 258482
rect 268752 244724 268804 244730
rect 268752 244666 268804 244672
rect 268660 244316 268712 244322
rect 268660 244258 268712 244264
rect 268672 239170 268700 244258
rect 268764 239494 268792 244666
rect 268856 244322 268884 258454
rect 268844 244316 268896 244322
rect 268844 244258 268896 244264
rect 268752 239488 268804 239494
rect 268752 239430 268804 239436
rect 268672 239142 268884 239170
rect 268752 229764 268804 229770
rect 268752 229706 268804 229712
rect 268660 225004 268712 225010
rect 268660 224946 268712 224952
rect 268672 219994 268700 224946
rect 268764 224534 268792 229706
rect 268856 225010 268884 239142
rect 268844 225004 268896 225010
rect 268844 224946 268896 224952
rect 268752 224528 268804 224534
rect 268752 224470 268804 224476
rect 268672 219966 268884 219994
rect 268752 210452 268804 210458
rect 268752 210394 268804 210400
rect 268660 205692 268712 205698
rect 268660 205634 268712 205640
rect 268672 200682 268700 205634
rect 268764 201006 268792 210394
rect 268856 205698 268884 219966
rect 268844 205692 268896 205698
rect 268844 205634 268896 205640
rect 268752 201000 268804 201006
rect 268752 200942 268804 200948
rect 268672 200654 268884 200682
rect 268752 191140 268804 191146
rect 268752 191082 268804 191088
rect 268660 186380 268712 186386
rect 268660 186322 268712 186328
rect 268672 176746 268700 186322
rect 268764 181490 268792 191082
rect 268856 186386 268884 200654
rect 268844 186380 268896 186386
rect 268844 186322 268896 186328
rect 268752 181484 268804 181490
rect 268752 181426 268804 181432
rect 268672 176718 268792 176746
rect 268764 176610 268792 176718
rect 268580 176582 268792 176610
rect 268580 162194 268608 176582
rect 268752 171624 268804 171630
rect 268752 171566 268804 171572
rect 268764 162382 268792 171566
rect 268752 162376 268804 162382
rect 268752 162318 268804 162324
rect 268580 162166 268884 162194
rect 268752 152516 268804 152522
rect 268752 152458 268804 152464
rect 268660 147688 268712 147694
rect 268660 147630 268712 147636
rect 268672 138666 268700 147630
rect 268764 142866 268792 152458
rect 268856 147694 268884 162166
rect 268844 147688 268896 147694
rect 268844 147630 268896 147636
rect 268752 142860 268804 142866
rect 268752 142802 268804 142808
rect 268672 138638 268792 138666
rect 268764 137986 268792 138638
rect 268764 137958 268884 137986
rect 268752 133204 268804 133210
rect 268752 133146 268804 133152
rect 268660 128376 268712 128382
rect 268660 128318 268712 128324
rect 268672 122806 268700 128318
rect 268764 123554 268792 133146
rect 268856 128382 268884 137958
rect 268844 128376 268896 128382
rect 268844 128318 268896 128324
rect 268752 123548 268804 123554
rect 268752 123490 268804 123496
rect 268660 122800 268712 122806
rect 268660 122742 268712 122748
rect 268752 113892 268804 113898
rect 268752 113834 268804 113840
rect 268660 109064 268712 109070
rect 268660 109006 268712 109012
rect 268672 103494 268700 109006
rect 268764 108594 268792 113834
rect 268844 113212 268896 113218
rect 268844 113154 268896 113160
rect 268856 109070 268884 113154
rect 268844 109064 268896 109070
rect 268844 109006 268896 109012
rect 268752 108588 268804 108594
rect 268752 108530 268804 108536
rect 268660 103488 268712 103494
rect 268660 103430 268712 103436
rect 268752 94376 268804 94382
rect 268752 94318 268804 94324
rect 268568 93900 268620 93906
rect 268568 93842 268620 93848
rect 268580 84810 268608 93842
rect 268764 84930 268792 94318
rect 268752 84924 268804 84930
rect 268752 84866 268804 84872
rect 268580 84782 268884 84810
rect 268752 75132 268804 75138
rect 268752 75074 268804 75080
rect 268660 70440 268712 70446
rect 268660 70382 268712 70388
rect 268672 56624 268700 70382
rect 268764 65550 268792 75074
rect 268856 70446 268884 84782
rect 268844 70440 268896 70446
rect 268844 70382 268896 70388
rect 268752 65544 268804 65550
rect 268752 65486 268804 65492
rect 268580 56596 268700 56624
rect 268580 26738 268608 56596
rect 268752 55888 268804 55894
rect 268752 55830 268804 55836
rect 268764 46238 268792 55830
rect 268752 46232 268804 46238
rect 268752 46174 268804 46180
rect 268752 32224 268804 32230
rect 268752 32166 268804 32172
rect 268764 26926 268792 32166
rect 268752 26920 268804 26926
rect 268752 26862 268804 26868
rect 268580 26710 268884 26738
rect 268752 17264 268804 17270
rect 268752 17206 268804 17212
rect 267646 4992 267702 5001
rect 267646 4927 267702 4936
rect 268108 4956 268160 4962
rect 268108 4898 268160 4904
rect 267372 3188 267424 3194
rect 267372 3130 267424 3136
rect 268120 480 268148 4898
rect 268764 4894 268792 17206
rect 268856 15065 268884 26710
rect 268842 15056 268898 15065
rect 268842 14991 268898 15000
rect 268948 8945 268976 307022
rect 269132 305794 269160 320146
rect 269330 320062 269436 320090
rect 269790 320062 269988 320090
rect 270618 320062 270816 320090
rect 270986 320062 271276 320090
rect 271446 320062 271644 320090
rect 271814 320062 271920 320090
rect 269408 318850 269436 320062
rect 269212 318844 269264 318850
rect 269212 318786 269264 318792
rect 269396 318844 269448 318850
rect 269396 318786 269448 318792
rect 269224 311794 269252 318786
rect 269960 316010 269988 320062
rect 270500 316056 270552 316062
rect 269960 315982 270448 316010
rect 270500 315998 270552 316004
rect 269224 311766 270356 311794
rect 269120 305788 269172 305794
rect 269120 305730 269172 305736
rect 270224 305788 270276 305794
rect 270224 305730 270276 305736
rect 269028 297424 269080 297430
rect 269028 297366 269080 297372
rect 269040 287774 269068 297366
rect 269028 287768 269080 287774
rect 269028 287710 269080 287716
rect 269028 278112 269080 278118
rect 269028 278054 269080 278060
rect 269040 268258 269068 278054
rect 269028 268252 269080 268258
rect 269028 268194 269080 268200
rect 269028 258800 269080 258806
rect 269028 258742 269080 258748
rect 269040 244730 269068 258742
rect 269028 244724 269080 244730
rect 269028 244666 269080 244672
rect 269028 239488 269080 239494
rect 269028 239430 269080 239436
rect 269040 229770 269068 239430
rect 269028 229764 269080 229770
rect 269028 229706 269080 229712
rect 269028 224528 269080 224534
rect 269028 224470 269080 224476
rect 269040 210458 269068 224470
rect 269028 210452 269080 210458
rect 269028 210394 269080 210400
rect 269028 201000 269080 201006
rect 269028 200942 269080 200948
rect 269040 191146 269068 200942
rect 269028 191140 269080 191146
rect 269028 191082 269080 191088
rect 269028 181484 269080 181490
rect 269028 181426 269080 181432
rect 269040 171630 269068 181426
rect 269028 171624 269080 171630
rect 269028 171566 269080 171572
rect 269028 162376 269080 162382
rect 269028 162318 269080 162324
rect 269040 152522 269068 162318
rect 269028 152516 269080 152522
rect 269028 152458 269080 152464
rect 269028 142860 269080 142866
rect 269028 142802 269080 142808
rect 269040 133210 269068 142802
rect 269028 133204 269080 133210
rect 269028 133146 269080 133152
rect 269028 123548 269080 123554
rect 269028 123490 269080 123496
rect 269040 113898 269068 123490
rect 269028 113892 269080 113898
rect 269028 113834 269080 113840
rect 269028 108588 269080 108594
rect 269028 108530 269080 108536
rect 269040 94382 269068 108530
rect 269028 94376 269080 94382
rect 269028 94318 269080 94324
rect 269028 84924 269080 84930
rect 269028 84866 269080 84872
rect 269040 75138 269068 84866
rect 269028 75132 269080 75138
rect 269028 75074 269080 75080
rect 269028 65544 269080 65550
rect 269028 65486 269080 65492
rect 269040 55894 269068 65486
rect 269028 55888 269080 55894
rect 269028 55830 269080 55836
rect 269028 46232 269080 46238
rect 269028 46174 269080 46180
rect 269040 32230 269068 46174
rect 269028 32224 269080 32230
rect 269028 32166 269080 32172
rect 269028 26920 269080 26926
rect 269028 26862 269080 26868
rect 269040 17270 269068 26862
rect 269028 17264 269080 17270
rect 269028 17206 269080 17212
rect 270236 14793 270264 305730
rect 270328 14929 270356 311766
rect 270314 14920 270370 14929
rect 270314 14855 270370 14864
rect 270222 14784 270278 14793
rect 270222 14719 270278 14728
rect 268934 8936 268990 8945
rect 268934 8871 268990 8880
rect 268752 4888 268804 4894
rect 270420 4865 270448 315982
rect 270512 307086 270540 315998
rect 270788 309194 270816 320062
rect 271248 315994 271276 320062
rect 271236 315988 271288 315994
rect 271236 315930 271288 315936
rect 271616 315874 271644 320062
rect 271892 319462 271920 320062
rect 271696 319456 271748 319462
rect 271696 319398 271748 319404
rect 271880 319456 271932 319462
rect 271880 319398 271932 319404
rect 271708 316062 271736 319398
rect 353944 318776 353996 318782
rect 353944 318718 353996 318724
rect 329104 318640 329156 318646
rect 329104 318582 329156 318588
rect 322204 317960 322256 317966
rect 322204 317902 322256 317908
rect 318064 317824 318116 317830
rect 318064 317766 318116 317772
rect 313924 317688 313976 317694
rect 313924 317630 313976 317636
rect 307024 317620 307076 317626
rect 307024 317562 307076 317568
rect 311164 317620 311216 317626
rect 311164 317562 311216 317568
rect 300124 317552 300176 317558
rect 300124 317494 300176 317500
rect 276664 317484 276716 317490
rect 276664 317426 276716 317432
rect 271696 316056 271748 316062
rect 271696 315998 271748 316004
rect 271788 315988 271840 315994
rect 271788 315930 271840 315936
rect 271616 315846 271736 315874
rect 270776 309188 270828 309194
rect 270776 309130 270828 309136
rect 271512 309188 271564 309194
rect 271512 309130 271564 309136
rect 270500 307080 270552 307086
rect 270500 307022 270552 307028
rect 271524 299470 271552 309130
rect 271604 307080 271656 307086
rect 271604 307022 271656 307028
rect 271512 299464 271564 299470
rect 271512 299406 271564 299412
rect 271512 293548 271564 293554
rect 271512 293490 271564 293496
rect 271524 14657 271552 293490
rect 271510 14648 271566 14657
rect 271510 14583 271566 14592
rect 271616 14521 271644 307022
rect 271602 14512 271658 14521
rect 271602 14447 271658 14456
rect 271708 8974 271736 315846
rect 270500 8968 270552 8974
rect 270500 8910 270552 8916
rect 271696 8968 271748 8974
rect 271696 8910 271748 8916
rect 268752 4830 268804 4836
rect 269302 4856 269358 4865
rect 269302 4791 269358 4800
rect 270406 4856 270462 4865
rect 270406 4791 270462 4800
rect 269316 480 269344 4791
rect 270512 480 270540 8910
rect 271800 4826 271828 315930
rect 271880 12504 271932 12510
rect 271880 12446 271932 12452
rect 271696 4820 271748 4826
rect 271696 4762 271748 4768
rect 271788 4820 271840 4826
rect 271788 4762 271840 4768
rect 271708 480 271736 4762
rect 271892 610 271920 12446
rect 274640 11144 274692 11150
rect 274640 11086 274692 11092
rect 274088 8356 274140 8362
rect 274088 8298 274140 8304
rect 271880 604 271932 610
rect 271880 546 271932 552
rect 272892 604 272944 610
rect 272892 546 272944 552
rect 272904 480 272932 546
rect 274100 480 274128 8298
rect 274652 610 274680 11086
rect 276478 5536 276534 5545
rect 276478 5471 276534 5480
rect 274640 604 274692 610
rect 274640 546 274692 552
rect 275284 604 275336 610
rect 275284 546 275336 552
rect 275296 480 275324 546
rect 276492 480 276520 5471
rect 276676 3262 276704 317426
rect 285680 16448 285732 16454
rect 285680 16390 285732 16396
rect 284300 14272 284352 14278
rect 284300 14214 284352 14220
rect 282920 14204 282972 14210
rect 282920 14146 282972 14152
rect 281540 14136 281592 14142
rect 281540 14078 281592 14084
rect 278872 14068 278924 14074
rect 278872 14010 278924 14016
rect 278780 13932 278832 13938
rect 278780 13874 278832 13880
rect 277400 13864 277452 13870
rect 277400 13806 277452 13812
rect 276664 3256 276716 3262
rect 276664 3198 276716 3204
rect 277412 610 277440 13806
rect 278792 3398 278820 13874
rect 278780 3392 278832 3398
rect 278780 3334 278832 3340
rect 277400 604 277452 610
rect 277400 546 277452 552
rect 277676 604 277728 610
rect 277676 546 277728 552
rect 277688 480 277716 546
rect 278884 480 278912 14010
rect 280160 14000 280212 14006
rect 280160 13942 280212 13948
rect 280068 3392 280120 3398
rect 280068 3334 280120 3340
rect 280080 480 280108 3334
rect 280172 610 280200 13942
rect 281552 610 281580 14078
rect 282932 610 282960 14146
rect 284312 626 284340 14214
rect 280160 604 280212 610
rect 280160 546 280212 552
rect 281264 604 281316 610
rect 281264 546 281316 552
rect 281540 604 281592 610
rect 281540 546 281592 552
rect 282460 604 282512 610
rect 282460 546 282512 552
rect 282920 604 282972 610
rect 282920 546 282972 552
rect 283656 604 283708 610
rect 284312 598 284800 626
rect 285692 610 285720 16390
rect 288440 16380 288492 16386
rect 288440 16322 288492 16328
rect 287060 14340 287112 14346
rect 287060 14282 287112 14288
rect 287072 5574 287100 14282
rect 286968 5568 287020 5574
rect 286968 5510 287020 5516
rect 287060 5568 287112 5574
rect 287060 5510 287112 5516
rect 288348 5568 288400 5574
rect 288348 5510 288400 5516
rect 286980 5386 287008 5510
rect 286980 5358 287192 5386
rect 283656 546 283708 552
rect 281276 480 281304 546
rect 282472 480 282500 546
rect 283668 480 283696 546
rect 284772 480 284800 598
rect 285680 604 285732 610
rect 285680 546 285732 552
rect 285956 604 286008 610
rect 285956 546 286008 552
rect 285968 480 285996 546
rect 287164 480 287192 5358
rect 288360 480 288388 5510
rect 288452 610 288480 16322
rect 292580 16312 292632 16318
rect 292580 16254 292632 16260
rect 291200 9716 291252 9722
rect 291200 9658 291252 9664
rect 290740 5636 290792 5642
rect 290740 5578 290792 5584
rect 288440 604 288492 610
rect 288440 546 288492 552
rect 289544 604 289596 610
rect 289544 546 289596 552
rect 289556 480 289584 546
rect 290752 480 290780 5578
rect 291212 610 291240 9658
rect 292592 610 292620 16254
rect 296720 16244 296772 16250
rect 296720 16186 296772 16192
rect 295340 9784 295392 9790
rect 295340 9726 295392 9732
rect 294328 5704 294380 5710
rect 294328 5646 294380 5652
rect 291200 604 291252 610
rect 291200 546 291252 552
rect 291936 604 291988 610
rect 291936 546 291988 552
rect 292580 604 292632 610
rect 292580 546 292632 552
rect 293132 604 293184 610
rect 293132 546 293184 552
rect 291948 480 291976 546
rect 293144 480 293172 546
rect 294340 480 294368 5646
rect 295352 610 295380 9726
rect 295340 604 295392 610
rect 295340 546 295392 552
rect 295524 604 295576 610
rect 295524 546 295576 552
rect 295536 480 295564 546
rect 296732 480 296760 16186
rect 298100 9852 298152 9858
rect 298100 9794 298152 9800
rect 297916 5772 297968 5778
rect 297916 5714 297968 5720
rect 297928 480 297956 5714
rect 298112 610 298140 9794
rect 300136 3398 300164 317494
rect 303620 16176 303672 16182
rect 303620 16118 303672 16124
rect 302240 9920 302292 9926
rect 302240 9862 302292 9868
rect 301412 5840 301464 5846
rect 301412 5782 301464 5788
rect 300124 3392 300176 3398
rect 300124 3334 300176 3340
rect 300308 3324 300360 3330
rect 300308 3266 300360 3272
rect 298100 604 298152 610
rect 298100 546 298152 552
rect 299112 604 299164 610
rect 299112 546 299164 552
rect 299124 480 299152 546
rect 300320 480 300348 3266
rect 301424 480 301452 5782
rect 302252 626 302280 9862
rect 302252 598 302648 626
rect 303632 610 303660 16118
rect 305000 9988 305052 9994
rect 305000 9930 305052 9936
rect 305012 3398 305040 9930
rect 305092 5908 305144 5914
rect 305092 5850 305144 5856
rect 305000 3392 305052 3398
rect 305000 3334 305052 3340
rect 305104 3210 305132 5850
rect 307036 3398 307064 317562
rect 309140 10056 309192 10062
rect 309140 9998 309192 10004
rect 308588 5976 308640 5982
rect 308588 5918 308640 5924
rect 306196 3392 306248 3398
rect 306196 3334 306248 3340
rect 307024 3392 307076 3398
rect 307024 3334 307076 3340
rect 305012 3182 305132 3210
rect 302620 480 302648 598
rect 303620 604 303672 610
rect 303620 546 303672 552
rect 303804 604 303856 610
rect 303804 546 303856 552
rect 303816 480 303844 546
rect 305012 480 305040 3182
rect 306208 480 306236 3334
rect 307392 2984 307444 2990
rect 307392 2926 307444 2932
rect 307404 480 307432 2926
rect 308600 480 308628 5918
rect 309152 610 309180 9998
rect 311176 3330 311204 317562
rect 313372 10124 313424 10130
rect 313372 10066 313424 10072
rect 312176 6044 312228 6050
rect 312176 5986 312228 5992
rect 310980 3324 311032 3330
rect 310980 3266 311032 3272
rect 311164 3324 311216 3330
rect 311164 3266 311216 3272
rect 309140 604 309192 610
rect 309140 546 309192 552
rect 309784 604 309836 610
rect 309784 546 309836 552
rect 309796 480 309824 546
rect 310992 480 311020 3266
rect 312188 480 312216 5986
rect 313384 480 313412 10066
rect 313936 2990 313964 317630
rect 316040 10192 316092 10198
rect 316040 10134 316092 10140
rect 315764 6112 315816 6118
rect 315764 6054 315816 6060
rect 313924 2984 313976 2990
rect 313924 2926 313976 2932
rect 314568 2916 314620 2922
rect 314568 2858 314620 2864
rect 314580 480 314608 2858
rect 315776 480 315804 6054
rect 316052 610 316080 10134
rect 318076 4978 318104 317766
rect 320180 10260 320232 10266
rect 320180 10202 320232 10208
rect 319260 6860 319312 6866
rect 319260 6802 319312 6808
rect 318076 4950 318196 4978
rect 318168 2990 318196 4950
rect 318064 2984 318116 2990
rect 318064 2926 318116 2932
rect 318156 2984 318208 2990
rect 318156 2926 318208 2932
rect 316040 604 316092 610
rect 316040 546 316092 552
rect 316960 604 317012 610
rect 316960 546 317012 552
rect 316972 480 317000 546
rect 318076 480 318104 2926
rect 319272 480 319300 6802
rect 320192 626 320220 10202
rect 322216 3058 322244 317902
rect 325056 317892 325108 317898
rect 325056 317834 325108 317840
rect 325068 309126 325096 317834
rect 325056 309120 325108 309126
rect 325056 309062 325108 309068
rect 324964 299532 325016 299538
rect 324964 299474 325016 299480
rect 324976 292618 325004 299474
rect 324976 292590 325096 292618
rect 325068 289814 325096 292590
rect 325056 289808 325108 289814
rect 325056 289750 325108 289756
rect 324964 280220 325016 280226
rect 324964 280162 325016 280168
rect 324976 273306 325004 280162
rect 324976 273278 325096 273306
rect 325068 270502 325096 273278
rect 325056 270496 325108 270502
rect 325056 270438 325108 270444
rect 324964 260908 325016 260914
rect 324964 260850 325016 260856
rect 324976 251258 325004 260850
rect 324780 251252 324832 251258
rect 324780 251194 324832 251200
rect 324964 251252 325016 251258
rect 324964 251194 325016 251200
rect 324792 251122 324820 251194
rect 324780 251116 324832 251122
rect 324780 251058 324832 251064
rect 324872 241596 324924 241602
rect 324872 241538 324924 241544
rect 324884 241466 324912 241538
rect 324872 241460 324924 241466
rect 324872 241402 324924 241408
rect 325056 234660 325108 234666
rect 325056 234602 325108 234608
rect 325068 231849 325096 234602
rect 324870 231840 324926 231849
rect 324870 231775 324926 231784
rect 325054 231840 325110 231849
rect 325054 231775 325110 231784
rect 324884 222222 324912 231775
rect 324872 222216 324924 222222
rect 324872 222158 324924 222164
rect 325148 222216 325200 222222
rect 325148 222158 325200 222164
rect 325160 215422 325188 222158
rect 325148 215416 325200 215422
rect 325148 215358 325200 215364
rect 325056 215280 325108 215286
rect 325056 215222 325108 215228
rect 325068 212537 325096 215222
rect 324870 212528 324926 212537
rect 324870 212463 324926 212472
rect 325054 212528 325110 212537
rect 325054 212463 325110 212472
rect 324884 202910 324912 212463
rect 324872 202904 324924 202910
rect 324872 202846 324924 202852
rect 325148 202904 325200 202910
rect 325148 202846 325200 202852
rect 325160 196110 325188 202846
rect 325148 196104 325200 196110
rect 325148 196046 325200 196052
rect 325056 195968 325108 195974
rect 325056 195910 325108 195916
rect 325068 193225 325096 195910
rect 324870 193216 324926 193225
rect 324870 193151 324926 193160
rect 325054 193216 325110 193225
rect 325054 193151 325110 193160
rect 324884 183598 324912 193151
rect 324872 183592 324924 183598
rect 324872 183534 324924 183540
rect 325148 183592 325200 183598
rect 325148 183534 325200 183540
rect 325160 176798 325188 183534
rect 325148 176792 325200 176798
rect 325148 176734 325200 176740
rect 325056 176656 325108 176662
rect 325056 176598 325108 176604
rect 325068 173913 325096 176598
rect 324870 173904 324926 173913
rect 324870 173839 324926 173848
rect 325054 173904 325110 173913
rect 325054 173839 325110 173848
rect 324884 167006 324912 173839
rect 324872 167000 324924 167006
rect 324872 166942 324924 166948
rect 325056 167000 325108 167006
rect 325056 166942 325108 166948
rect 325068 164234 325096 166942
rect 325068 164206 325188 164234
rect 325160 157486 325188 164206
rect 325148 157480 325200 157486
rect 325148 157422 325200 157428
rect 325056 157276 325108 157282
rect 325056 157218 325108 157224
rect 325068 154562 325096 157218
rect 325056 154556 325108 154562
rect 325056 154498 325108 154504
rect 325240 154556 325292 154562
rect 325240 154498 325292 154504
rect 325252 144945 325280 154498
rect 324962 144936 325018 144945
rect 324962 144871 325018 144880
rect 325238 144936 325294 144945
rect 325238 144871 325294 144880
rect 324976 138038 325004 144871
rect 324964 138032 325016 138038
rect 324964 137974 325016 137980
rect 325056 137964 325108 137970
rect 325056 137906 325108 137912
rect 325068 135250 325096 137906
rect 325056 135244 325108 135250
rect 325056 135186 325108 135192
rect 325240 135244 325292 135250
rect 325240 135186 325292 135192
rect 325252 125633 325280 135186
rect 324962 125624 325018 125633
rect 324962 125559 325018 125568
rect 325238 125624 325294 125633
rect 325238 125559 325294 125568
rect 324976 118726 325004 125559
rect 324964 118720 325016 118726
rect 324964 118662 325016 118668
rect 325056 118652 325108 118658
rect 325056 118594 325108 118600
rect 325068 115938 325096 118594
rect 325056 115932 325108 115938
rect 325056 115874 325108 115880
rect 325240 115932 325292 115938
rect 325240 115874 325292 115880
rect 325252 106321 325280 115874
rect 324962 106312 325018 106321
rect 324962 106247 325018 106256
rect 325238 106312 325294 106321
rect 325238 106247 325294 106256
rect 324976 101454 325004 106247
rect 324780 101448 324832 101454
rect 324780 101390 324832 101396
rect 324964 101448 325016 101454
rect 324964 101390 325016 101396
rect 324792 89706 324820 101390
rect 324792 89678 325004 89706
rect 324976 80102 325004 89678
rect 324964 80096 325016 80102
rect 324964 80038 325016 80044
rect 325056 79960 325108 79966
rect 325056 79902 325108 79908
rect 325068 77246 325096 79902
rect 325056 77240 325108 77246
rect 325056 77182 325108 77188
rect 324964 67652 325016 67658
rect 324964 67594 325016 67600
rect 324976 60738 325004 67594
rect 324792 60710 325004 60738
rect 324792 48278 324820 60710
rect 324596 48272 324648 48278
rect 324596 48214 324648 48220
rect 324780 48272 324832 48278
rect 324780 48214 324832 48220
rect 324608 46918 324636 48214
rect 324596 46912 324648 46918
rect 324596 46854 324648 46860
rect 324872 38548 324924 38554
rect 324872 38490 324924 38496
rect 324884 31822 324912 38490
rect 324872 31816 324924 31822
rect 324872 31758 324924 31764
rect 324872 31680 324924 31686
rect 324872 31622 324924 31628
rect 324884 22114 324912 31622
rect 324884 22086 325188 22114
rect 325160 21978 325188 22086
rect 325160 21950 325372 21978
rect 322940 11008 322992 11014
rect 322940 10950 322992 10956
rect 322848 6792 322900 6798
rect 322848 6734 322900 6740
rect 321652 3052 321704 3058
rect 321652 2994 321704 3000
rect 322204 3052 322256 3058
rect 322204 2994 322256 3000
rect 320192 598 320496 626
rect 320468 480 320496 598
rect 321664 480 321692 2994
rect 322860 480 322888 6734
rect 322952 610 322980 10950
rect 325344 3330 325372 21950
rect 327080 10940 327132 10946
rect 327080 10882 327132 10888
rect 326436 6724 326488 6730
rect 326436 6666 326488 6672
rect 325240 3324 325292 3330
rect 325240 3266 325292 3272
rect 325332 3324 325384 3330
rect 325332 3266 325384 3272
rect 322940 604 322992 610
rect 322940 546 322992 552
rect 324044 604 324096 610
rect 324044 546 324096 552
rect 324056 480 324084 546
rect 325252 480 325280 3266
rect 326448 480 326476 6666
rect 327092 610 327120 10882
rect 328828 4140 328880 4146
rect 328828 4082 328880 4088
rect 327080 604 327132 610
rect 327080 546 327132 552
rect 327632 604 327684 610
rect 327632 546 327684 552
rect 327644 480 327672 546
rect 328840 480 328868 4082
rect 329116 3398 329144 318582
rect 331864 318572 331916 318578
rect 331864 318514 331916 318520
rect 331312 10872 331364 10878
rect 331312 10814 331364 10820
rect 330024 6656 330076 6662
rect 330024 6598 330076 6604
rect 329104 3392 329156 3398
rect 329104 3334 329156 3340
rect 330036 480 330064 6598
rect 331324 626 331352 10814
rect 331876 4010 331904 318514
rect 348424 318504 348476 318510
rect 348424 318446 348476 318452
rect 347044 318436 347096 318442
rect 347044 318378 347096 318384
rect 345664 318368 345716 318374
rect 345664 318310 345716 318316
rect 336004 318300 336056 318306
rect 336004 318242 336056 318248
rect 333980 10804 334032 10810
rect 333980 10746 334032 10752
rect 333612 6588 333664 6594
rect 333612 6530 333664 6536
rect 331864 4004 331916 4010
rect 331864 3946 331916 3952
rect 332416 2916 332468 2922
rect 332416 2858 332468 2864
rect 331232 598 331352 626
rect 331232 480 331260 598
rect 332428 480 332456 2858
rect 333624 480 333652 6530
rect 333992 610 334020 10746
rect 336016 4078 336044 318242
rect 342904 318164 342956 318170
rect 342904 318106 342956 318112
rect 340144 318096 340196 318102
rect 340144 318038 340196 318044
rect 338120 10736 338172 10742
rect 338120 10678 338172 10684
rect 337108 6520 337160 6526
rect 337108 6462 337160 6468
rect 335912 4072 335964 4078
rect 335912 4014 335964 4020
rect 336004 4072 336056 4078
rect 336004 4014 336056 4020
rect 333980 604 334032 610
rect 333980 546 334032 552
rect 334716 604 334768 610
rect 334716 546 334768 552
rect 334728 480 334756 546
rect 335924 480 335952 4014
rect 337120 480 337148 6462
rect 338132 626 338160 10678
rect 340156 5386 340184 318038
rect 340880 10668 340932 10674
rect 340880 10610 340932 10616
rect 340696 6452 340748 6458
rect 340696 6394 340748 6400
rect 340156 5358 340276 5386
rect 340248 4010 340276 5358
rect 340236 4004 340288 4010
rect 340236 3946 340288 3952
rect 339500 2984 339552 2990
rect 339500 2926 339552 2932
rect 338132 598 338344 626
rect 338316 480 338344 598
rect 339512 480 339540 2926
rect 340708 480 340736 6394
rect 340892 610 340920 10610
rect 342916 2922 342944 318106
rect 345020 10600 345072 10606
rect 345020 10542 345072 10548
rect 344284 6384 344336 6390
rect 344284 6326 344336 6332
rect 342904 2916 342956 2922
rect 342904 2858 342956 2864
rect 343088 2848 343140 2854
rect 343088 2790 343140 2796
rect 340880 604 340932 610
rect 340880 546 340932 552
rect 341892 604 341944 610
rect 341892 546 341944 552
rect 341904 480 341932 546
rect 343100 480 343128 2790
rect 344296 480 344324 6326
rect 345032 4298 345060 10542
rect 345032 4270 345428 4298
rect 345018 4176 345074 4185
rect 345018 4111 345020 4120
rect 345072 4111 345074 4120
rect 345020 4082 345072 4088
rect 345400 626 345428 4270
rect 345676 2990 345704 318310
rect 346676 3052 346728 3058
rect 346676 2994 346728 3000
rect 345664 2984 345716 2990
rect 345664 2926 345716 2932
rect 345400 598 345520 626
rect 345492 480 345520 598
rect 346688 480 346716 2994
rect 347056 2922 347084 318378
rect 347780 10532 347832 10538
rect 347780 10474 347832 10480
rect 347792 3330 347820 10474
rect 347872 6316 347924 6322
rect 347872 6258 347924 6264
rect 347780 3324 347832 3330
rect 347780 3266 347832 3272
rect 347044 2916 347096 2922
rect 347044 2858 347096 2864
rect 347884 480 347912 6258
rect 348436 2990 348464 318446
rect 349804 318028 349856 318034
rect 349804 317970 349856 317976
rect 349068 3324 349120 3330
rect 349068 3266 349120 3272
rect 348424 2984 348476 2990
rect 348424 2926 348476 2932
rect 349080 480 349108 3266
rect 349816 2990 349844 317970
rect 351920 10464 351972 10470
rect 351920 10406 351972 10412
rect 351368 6248 351420 6254
rect 351368 6190 351420 6196
rect 350264 3120 350316 3126
rect 350264 3062 350316 3068
rect 349804 2984 349856 2990
rect 349804 2926 349856 2932
rect 350276 480 350304 3062
rect 351380 480 351408 6190
rect 351932 610 351960 10406
rect 353956 3126 353984 318718
rect 356704 318708 356756 318714
rect 356704 318650 356756 318656
rect 356152 10396 356204 10402
rect 356152 10338 356204 10344
rect 354956 6180 355008 6186
rect 354956 6122 355008 6128
rect 354586 4176 354642 4185
rect 354586 4111 354588 4120
rect 354640 4111 354642 4120
rect 354588 4082 354640 4088
rect 353944 3120 353996 3126
rect 353944 3062 353996 3068
rect 353760 3052 353812 3058
rect 353760 2994 353812 3000
rect 351920 604 351972 610
rect 351920 546 351972 552
rect 352564 604 352616 610
rect 352564 546 352616 552
rect 352576 480 352604 546
rect 353772 480 353800 2994
rect 354968 480 354996 6122
rect 356164 480 356192 10338
rect 356716 3233 356744 318650
rect 374642 318608 374698 318617
rect 374642 318543 374698 318552
rect 367742 318472 367798 318481
rect 367742 318407 367798 318416
rect 360844 318232 360896 318238
rect 360844 318174 360896 318180
rect 364982 318200 365038 318209
rect 358820 10328 358872 10334
rect 358820 10270 358872 10276
rect 358542 6760 358598 6769
rect 358542 6695 358598 6704
rect 357348 3936 357400 3942
rect 357348 3878 357400 3884
rect 356702 3224 356758 3233
rect 356702 3159 356758 3168
rect 357360 480 357388 3878
rect 358556 480 358584 6695
rect 358832 610 358860 10270
rect 360856 5386 360884 318174
rect 364982 318135 365038 318144
rect 362958 10840 363014 10849
rect 362958 10775 363014 10784
rect 362130 6624 362186 6633
rect 362130 6559 362186 6568
rect 360856 5358 361068 5386
rect 361040 3942 361068 5358
rect 360936 3936 360988 3942
rect 360936 3878 360988 3884
rect 361028 3936 361080 3942
rect 361028 3878 361080 3884
rect 359648 3392 359700 3398
rect 359648 3334 359700 3340
rect 359660 3233 359688 3334
rect 359646 3224 359702 3233
rect 359646 3159 359702 3168
rect 358820 604 358872 610
rect 358820 546 358872 552
rect 359740 604 359792 610
rect 359740 546 359792 552
rect 359752 480 359780 546
rect 360948 480 360976 3878
rect 362144 480 362172 6559
rect 362972 626 363000 10775
rect 364996 4078 365024 318135
rect 365718 10704 365774 10713
rect 365718 10639 365774 10648
rect 364892 4072 364944 4078
rect 364890 4040 364892 4049
rect 364984 4072 365036 4078
rect 364944 4040 364946 4049
rect 364984 4014 365036 4020
rect 364890 3975 364946 3984
rect 365732 3194 365760 10639
rect 365810 6488 365866 6497
rect 365810 6423 365866 6432
rect 364524 3188 364576 3194
rect 364524 3130 364576 3136
rect 365720 3188 365772 3194
rect 365720 3130 365772 3136
rect 362972 598 363368 626
rect 363340 480 363368 598
rect 364536 480 364564 3130
rect 365824 3074 365852 6423
rect 367756 5574 367784 318407
rect 373262 318336 373318 318345
rect 373262 318271 373318 318280
rect 371882 318064 371938 318073
rect 371882 317999 371938 318008
rect 369858 10568 369914 10577
rect 369858 10503 369914 10512
rect 369214 6352 369270 6361
rect 369214 6287 369270 6296
rect 367744 5568 367796 5574
rect 367744 5510 367796 5516
rect 368204 5568 368256 5574
rect 368204 5510 368256 5516
rect 368216 4146 368244 5510
rect 368020 4140 368072 4146
rect 368020 4082 368072 4088
rect 368204 4140 368256 4146
rect 368204 4082 368256 4088
rect 369124 4140 369176 4146
rect 369124 4082 369176 4088
rect 367006 4040 367062 4049
rect 367006 3975 367062 3984
rect 367020 3194 367048 3975
rect 366916 3188 366968 3194
rect 366916 3130 366968 3136
rect 367008 3188 367060 3194
rect 367008 3130 367060 3136
rect 365732 3046 365852 3074
rect 365732 480 365760 3046
rect 366928 480 366956 3130
rect 368032 480 368060 4082
rect 369136 3942 369164 4082
rect 369124 3936 369176 3942
rect 369124 3878 369176 3884
rect 369228 480 369256 6287
rect 369872 610 369900 10503
rect 371896 3942 371924 317999
rect 372802 6216 372858 6225
rect 372802 6151 372858 6160
rect 371884 3936 371936 3942
rect 371884 3878 371936 3884
rect 371608 3868 371660 3874
rect 371608 3810 371660 3816
rect 369860 604 369912 610
rect 369860 546 369912 552
rect 370412 604 370464 610
rect 370412 546 370464 552
rect 370424 480 370452 546
rect 371620 480 371648 3810
rect 372816 480 372844 6151
rect 373276 4049 373304 318271
rect 374090 10432 374146 10441
rect 374090 10367 374146 10376
rect 373262 4040 373318 4049
rect 373262 3975 373318 3984
rect 374104 626 374132 10367
rect 374656 5386 374684 318543
rect 391940 16108 391992 16114
rect 391940 16050 391992 16056
rect 379520 15156 379572 15162
rect 379520 15098 379572 15104
rect 375380 14408 375432 14414
rect 375380 14350 375432 14356
rect 374656 5358 375328 5386
rect 375300 3194 375328 5358
rect 375196 3188 375248 3194
rect 375196 3130 375248 3136
rect 375288 3188 375340 3194
rect 375288 3130 375340 3136
rect 374012 598 374132 626
rect 374012 480 374040 598
rect 375208 480 375236 3130
rect 375392 610 375420 14350
rect 376758 10296 376814 10305
rect 376758 10231 376814 10240
rect 376772 610 376800 10231
rect 378784 3800 378836 3806
rect 378784 3742 378836 3748
rect 375380 604 375432 610
rect 375380 546 375432 552
rect 376392 604 376444 610
rect 376392 546 376444 552
rect 376760 604 376812 610
rect 376760 546 376812 552
rect 377588 604 377640 610
rect 377588 546 377640 552
rect 376404 480 376432 546
rect 377600 480 377628 546
rect 378796 480 378824 3742
rect 379532 610 379560 15098
rect 382372 15088 382424 15094
rect 382372 15030 382424 15036
rect 380900 15020 380952 15026
rect 380900 14962 380952 14968
rect 380912 626 380940 14962
rect 382280 4004 382332 4010
rect 382280 3946 382332 3952
rect 382292 3618 382320 3946
rect 382384 3806 382412 15030
rect 383660 14952 383712 14958
rect 383660 14894 383712 14900
rect 382372 3800 382424 3806
rect 382372 3742 382424 3748
rect 383568 3800 383620 3806
rect 383568 3742 383620 3748
rect 382292 3590 382412 3618
rect 379520 604 379572 610
rect 379520 546 379572 552
rect 379980 604 380032 610
rect 380912 598 381216 626
rect 379980 546 380032 552
rect 379992 480 380020 546
rect 381188 480 381216 598
rect 382384 480 382412 3590
rect 383580 480 383608 3742
rect 383672 3346 383700 14894
rect 387800 14884 387852 14890
rect 387800 14826 387852 14832
rect 386420 14816 386472 14822
rect 386420 14758 386472 14764
rect 385868 3732 385920 3738
rect 385868 3674 385920 3680
rect 383672 3318 384712 3346
rect 384684 480 384712 3318
rect 385880 480 385908 3674
rect 386432 3346 386460 14758
rect 387812 3346 387840 14826
rect 390560 14748 390612 14754
rect 390560 14690 390612 14696
rect 390572 3738 390600 14690
rect 390652 7064 390704 7070
rect 390652 7006 390704 7012
rect 390560 3732 390612 3738
rect 390560 3674 390612 3680
rect 386432 3318 387104 3346
rect 387812 3318 388300 3346
rect 387076 480 387104 3318
rect 388272 480 388300 3318
rect 389456 2848 389508 2854
rect 389456 2790 389508 2796
rect 389468 480 389496 2790
rect 390664 480 390692 7006
rect 391848 3732 391900 3738
rect 391848 3674 391900 3680
rect 391860 480 391888 3674
rect 391952 3346 391980 16050
rect 407120 16040 407172 16046
rect 407120 15982 407172 15988
rect 405740 11416 405792 11422
rect 405740 11358 405792 11364
rect 401600 11348 401652 11354
rect 401600 11290 401652 11296
rect 398840 11280 398892 11286
rect 398840 11222 398892 11228
rect 394700 11212 394752 11218
rect 394700 11154 394752 11160
rect 394240 7132 394292 7138
rect 394240 7074 394292 7080
rect 391952 3318 393084 3346
rect 393056 480 393084 3318
rect 394252 480 394280 7074
rect 394712 610 394740 11154
rect 397828 7200 397880 7206
rect 397828 7142 397880 7148
rect 396632 3664 396684 3670
rect 396632 3606 396684 3612
rect 394700 604 394752 610
rect 394700 546 394752 552
rect 395436 604 395488 610
rect 395436 546 395488 552
rect 395448 480 395476 546
rect 396644 480 396672 3606
rect 397840 480 397868 7142
rect 398852 626 398880 11222
rect 401324 7268 401376 7274
rect 401324 7210 401376 7216
rect 400220 3256 400272 3262
rect 400220 3198 400272 3204
rect 398852 598 399064 626
rect 399036 480 399064 598
rect 400232 480 400260 3198
rect 401336 480 401364 7210
rect 401612 610 401640 11290
rect 404912 7336 404964 7342
rect 404912 7278 404964 7284
rect 403716 2916 403768 2922
rect 403716 2858 403768 2864
rect 401600 604 401652 610
rect 401600 546 401652 552
rect 402520 604 402572 610
rect 402520 546 402572 552
rect 402532 480 402560 546
rect 403728 480 403756 2858
rect 404924 480 404952 7278
rect 405752 610 405780 11358
rect 407132 3482 407160 15982
rect 420920 15972 420972 15978
rect 420920 15914 420972 15920
rect 419540 11688 419592 11694
rect 419540 11630 419592 11636
rect 416872 11620 416924 11626
rect 416872 11562 416924 11568
rect 412640 11552 412692 11558
rect 412640 11494 412692 11500
rect 408500 11484 408552 11490
rect 408500 11426 408552 11432
rect 408512 3670 408540 11426
rect 412088 7472 412140 7478
rect 412088 7414 412140 7420
rect 408592 7404 408644 7410
rect 408592 7346 408644 7352
rect 408500 3664 408552 3670
rect 408500 3606 408552 3612
rect 408604 3482 408632 7346
rect 409696 3664 409748 3670
rect 409696 3606 409748 3612
rect 407132 3454 407344 3482
rect 405740 604 405792 610
rect 405740 546 405792 552
rect 406108 604 406160 610
rect 406108 546 406160 552
rect 406120 480 406148 546
rect 407316 480 407344 3454
rect 408512 3454 408632 3482
rect 408512 480 408540 3454
rect 409708 480 409736 3606
rect 410892 2984 410944 2990
rect 410892 2926 410944 2932
rect 410904 480 410932 2926
rect 412100 480 412128 7414
rect 412652 610 412680 11494
rect 415676 7540 415728 7546
rect 415676 7482 415728 7488
rect 414480 3596 414532 3602
rect 414480 3538 414532 3544
rect 412640 604 412692 610
rect 412640 546 412692 552
rect 413284 604 413336 610
rect 413284 546 413336 552
rect 413296 480 413324 546
rect 414492 480 414520 3538
rect 415688 480 415716 7482
rect 416884 480 416912 11562
rect 419172 8288 419224 8294
rect 419172 8230 419224 8236
rect 417976 3052 418028 3058
rect 417976 2994 418028 3000
rect 417988 480 418016 2994
rect 419184 480 419212 8230
rect 419552 610 419580 11630
rect 420932 610 420960 15914
rect 477500 15904 477552 15910
rect 477500 15846 477552 15852
rect 423680 12436 423732 12442
rect 423680 12378 423732 12384
rect 422760 8220 422812 8226
rect 422760 8162 422812 8168
rect 419540 604 419592 610
rect 419540 546 419592 552
rect 420368 604 420420 610
rect 420368 546 420420 552
rect 420920 604 420972 610
rect 420920 546 420972 552
rect 421564 604 421616 610
rect 421564 546 421616 552
rect 420380 480 420408 546
rect 421576 480 421604 546
rect 422772 480 422800 8162
rect 423692 610 423720 12378
rect 426440 12368 426492 12374
rect 426440 12310 426492 12316
rect 462318 12336 462374 12345
rect 426348 8152 426400 8158
rect 426348 8094 426400 8100
rect 425152 3120 425204 3126
rect 425152 3062 425204 3068
rect 423680 604 423732 610
rect 423680 546 423732 552
rect 423956 604 424008 610
rect 423956 546 424008 552
rect 423968 480 423996 546
rect 425164 480 425192 3062
rect 426360 480 426388 8094
rect 426452 610 426480 12310
rect 430580 12300 430632 12306
rect 462318 12271 462374 12280
rect 430580 12242 430632 12248
rect 429936 8084 429988 8090
rect 429936 8026 429988 8032
rect 428740 3528 428792 3534
rect 428740 3470 428792 3476
rect 426440 604 426492 610
rect 426440 546 426492 552
rect 427544 604 427596 610
rect 427544 546 427596 552
rect 427556 480 427584 546
rect 428752 480 428780 3470
rect 429948 480 429976 8026
rect 430592 610 430620 12242
rect 433340 12232 433392 12238
rect 433340 12174 433392 12180
rect 433352 3534 433380 12174
rect 437480 12164 437532 12170
rect 437480 12106 437532 12112
rect 433524 8016 433576 8022
rect 433524 7958 433576 7964
rect 433340 3528 433392 3534
rect 433340 3470 433392 3476
rect 432328 3324 432380 3330
rect 432328 3266 432380 3272
rect 430580 604 430632 610
rect 430580 546 430632 552
rect 431132 604 431184 610
rect 431132 546 431184 552
rect 431144 480 431172 546
rect 432340 480 432368 3266
rect 433536 480 433564 7958
rect 437020 7948 437072 7954
rect 437020 7890 437072 7896
rect 434628 3528 434680 3534
rect 434628 3470 434680 3476
rect 434640 480 434668 3470
rect 435824 3460 435876 3466
rect 435824 3402 435876 3408
rect 435836 480 435864 3402
rect 437032 480 437060 7890
rect 437492 610 437520 12106
rect 441620 12096 441672 12102
rect 441620 12038 441672 12044
rect 440608 7880 440660 7886
rect 440608 7822 440660 7828
rect 439412 3392 439464 3398
rect 439412 3334 439464 3340
rect 437480 604 437532 610
rect 437480 546 437532 552
rect 438216 604 438268 610
rect 438216 546 438268 552
rect 438228 480 438256 546
rect 439424 480 439452 3334
rect 440620 480 440648 7822
rect 441632 3482 441660 12038
rect 444380 12028 444432 12034
rect 444380 11970 444432 11976
rect 444196 7812 444248 7818
rect 444196 7754 444248 7760
rect 442998 3904 443054 3913
rect 442998 3839 443054 3848
rect 441632 3454 441844 3482
rect 441816 480 441844 3454
rect 443012 480 443040 3839
rect 444208 480 444236 7754
rect 444392 3482 444420 11970
rect 448520 11960 448572 11966
rect 448520 11902 448572 11908
rect 447784 7744 447836 7750
rect 447784 7686 447836 7692
rect 446588 4140 446640 4146
rect 446588 4082 446640 4088
rect 444392 3454 445432 3482
rect 445404 480 445432 3454
rect 446600 480 446628 4082
rect 447796 480 447824 7686
rect 448532 3482 448560 11902
rect 451280 11892 451332 11898
rect 451280 11834 451332 11840
rect 450174 3768 450230 3777
rect 450174 3703 450230 3712
rect 448532 3454 449020 3482
rect 448992 480 449020 3454
rect 450188 480 450216 3703
rect 451292 3534 451320 11834
rect 455420 11824 455472 11830
rect 455420 11766 455472 11772
rect 451372 7676 451424 7682
rect 451372 7618 451424 7624
rect 451280 3528 451332 3534
rect 451280 3470 451332 3476
rect 451384 1442 451412 7618
rect 454868 7608 454920 7614
rect 454868 7550 454920 7556
rect 453672 4072 453724 4078
rect 453672 4014 453724 4020
rect 452476 3528 452528 3534
rect 452476 3470 452528 3476
rect 451292 1414 451412 1442
rect 451292 480 451320 1414
rect 452488 480 452516 3470
rect 453684 480 453712 4014
rect 454880 480 454908 7550
rect 455432 610 455460 11766
rect 459652 11756 459704 11762
rect 459652 11698 459704 11704
rect 458454 8256 458510 8265
rect 458454 8191 458510 8200
rect 457258 3632 457314 3641
rect 457258 3567 457314 3576
rect 455420 604 455472 610
rect 455420 546 455472 552
rect 456064 604 456116 610
rect 456064 546 456116 552
rect 456076 480 456104 546
rect 457272 480 457300 3567
rect 458468 480 458496 8191
rect 459664 480 459692 11698
rect 462042 8120 462098 8129
rect 462042 8055 462098 8064
rect 460848 3188 460900 3194
rect 460848 3130 460900 3136
rect 460860 480 460888 3130
rect 462056 480 462084 8055
rect 462332 610 462360 12271
rect 466458 12200 466514 12209
rect 466458 12135 466514 12144
rect 465630 7984 465686 7993
rect 465630 7919 465686 7928
rect 464434 3496 464490 3505
rect 464434 3431 464490 3440
rect 462320 604 462372 610
rect 462320 546 462372 552
rect 463240 604 463292 610
rect 463240 546 463292 552
rect 463252 480 463280 546
rect 464448 480 464476 3431
rect 465644 480 465672 7919
rect 466472 610 466500 12135
rect 469218 12064 469274 12073
rect 469218 11999 469274 12008
rect 469126 7848 469182 7857
rect 469126 7783 469182 7792
rect 467932 3936 467984 3942
rect 467932 3878 467984 3884
rect 466460 604 466512 610
rect 466460 546 466512 552
rect 466828 604 466880 610
rect 466828 546 466880 552
rect 466840 480 466868 546
rect 467944 480 467972 3878
rect 469140 480 469168 7783
rect 469232 610 469260 11999
rect 473358 11928 473414 11937
rect 473358 11863 473414 11872
rect 472714 7712 472770 7721
rect 472714 7647 472770 7656
rect 471518 3360 471574 3369
rect 471518 3295 471574 3304
rect 469220 604 469272 610
rect 469220 546 469272 552
rect 470324 604 470376 610
rect 470324 546 470376 552
rect 470336 480 470364 546
rect 471532 480 471560 3295
rect 472728 480 472756 7647
rect 473372 626 473400 11863
rect 476302 7576 476358 7585
rect 476302 7511 476358 7520
rect 475106 4040 475162 4049
rect 475106 3975 475162 3984
rect 473372 598 473860 626
rect 473832 592 473860 598
rect 473832 564 473952 592
rect 473924 480 473952 564
rect 475120 480 475148 3975
rect 476316 480 476344 7511
rect 477512 3602 477540 15846
rect 489918 15192 489974 15201
rect 489918 15127 489974 15136
rect 478880 14680 478932 14686
rect 478880 14622 478932 14628
rect 477590 11792 477646 11801
rect 477590 11727 477646 11736
rect 477500 3596 477552 3602
rect 477500 3538 477552 3544
rect 477604 3482 477632 11727
rect 478696 3596 478748 3602
rect 478696 3538 478748 3544
rect 477512 3454 477632 3482
rect 477512 480 477540 3454
rect 478708 480 478736 3538
rect 478892 610 478920 14622
rect 484400 14612 484452 14618
rect 484400 14554 484452 14560
rect 483020 12572 483072 12578
rect 483020 12514 483072 12520
rect 480258 11656 480314 11665
rect 480258 11591 480314 11600
rect 480272 3482 480300 11591
rect 482284 3868 482336 3874
rect 482284 3810 482336 3816
rect 480272 3454 481128 3482
rect 478880 604 478932 610
rect 478880 546 478932 552
rect 479892 604 479944 610
rect 479892 546 479944 552
rect 479904 480 479932 546
rect 481100 480 481128 3454
rect 482296 480 482324 3810
rect 483032 3482 483060 12514
rect 484412 3482 484440 14554
rect 485780 14544 485832 14550
rect 485780 14486 485832 14492
rect 483032 3454 483520 3482
rect 484412 3454 484624 3482
rect 483492 480 483520 3454
rect 484596 480 484624 3454
rect 485792 480 485820 14486
rect 487160 14476 487212 14482
rect 487160 14418 487212 14424
rect 485872 12640 485924 12646
rect 485872 12582 485924 12588
rect 485884 3482 485912 12582
rect 487172 3482 487200 14418
rect 488540 12708 488592 12714
rect 488540 12650 488592 12656
rect 488552 3482 488580 12650
rect 485884 3454 487016 3482
rect 487172 3454 488212 3482
rect 488552 3454 489408 3482
rect 486988 480 487016 3454
rect 488184 480 488212 3454
rect 489380 480 489408 3454
rect 489932 610 489960 15127
rect 571338 15056 571394 15065
rect 571338 14991 571394 15000
rect 510620 13796 510672 13802
rect 510620 13738 510672 13744
rect 506480 13048 506532 13054
rect 506480 12990 506532 12996
rect 502340 12980 502392 12986
rect 502340 12922 502392 12928
rect 499580 12912 499632 12918
rect 499580 12854 499632 12860
rect 495440 12844 495492 12850
rect 495440 12786 495492 12792
rect 492680 12776 492732 12782
rect 492680 12718 492732 12724
rect 491760 8424 491812 8430
rect 491760 8366 491812 8372
rect 489920 604 489972 610
rect 489920 546 489972 552
rect 490564 604 490616 610
rect 490564 546 490616 552
rect 490576 480 490604 546
rect 491772 480 491800 8366
rect 492692 626 492720 12718
rect 495348 8492 495400 8498
rect 495348 8434 495400 8440
rect 494152 4208 494204 4214
rect 494152 4150 494204 4156
rect 492692 598 492904 626
rect 492876 592 492904 598
rect 492876 564 492996 592
rect 492968 480 492996 564
rect 494164 480 494192 4150
rect 495360 480 495388 8434
rect 495452 610 495480 12786
rect 498936 8560 498988 8566
rect 498936 8502 498988 8508
rect 497740 4276 497792 4282
rect 497740 4218 497792 4224
rect 495440 604 495492 610
rect 495440 546 495492 552
rect 496544 604 496596 610
rect 496544 546 496596 552
rect 496556 480 496584 546
rect 497752 480 497780 4218
rect 498948 480 498976 8502
rect 499592 610 499620 12854
rect 501236 4344 501288 4350
rect 501236 4286 501288 4292
rect 499580 604 499632 610
rect 499580 546 499632 552
rect 500132 604 500184 610
rect 500132 546 500184 552
rect 500144 480 500172 546
rect 501248 480 501276 4286
rect 502352 3534 502380 12922
rect 506020 8696 506072 8702
rect 506020 8638 506072 8644
rect 502432 8628 502484 8634
rect 502432 8570 502484 8576
rect 502340 3528 502392 3534
rect 502340 3470 502392 3476
rect 502444 480 502472 8570
rect 504824 4412 504876 4418
rect 504824 4354 504876 4360
rect 503628 3528 503680 3534
rect 503628 3470 503680 3476
rect 503640 480 503668 3470
rect 504836 480 504864 4354
rect 506032 480 506060 8638
rect 506492 610 506520 12990
rect 509608 8764 509660 8770
rect 509608 8706 509660 8712
rect 508412 4480 508464 4486
rect 508412 4422 508464 4428
rect 506480 604 506532 610
rect 506480 546 506532 552
rect 507216 604 507268 610
rect 507216 546 507268 552
rect 507228 480 507256 546
rect 508424 480 508452 4422
rect 509620 480 509648 8706
rect 510632 610 510660 13738
rect 513380 13728 513432 13734
rect 513380 13670 513432 13676
rect 549258 13696 549314 13705
rect 513196 8832 513248 8838
rect 513196 8774 513248 8780
rect 512000 4548 512052 4554
rect 512000 4490 512052 4496
rect 510620 604 510672 610
rect 510620 546 510672 552
rect 510804 604 510856 610
rect 510804 546 510856 552
rect 510816 480 510844 546
rect 512012 480 512040 4490
rect 513208 480 513236 8774
rect 513392 610 513420 13670
rect 517520 13660 517572 13666
rect 549258 13631 549314 13640
rect 517520 13602 517572 13608
rect 516784 8900 516836 8906
rect 516784 8842 516836 8848
rect 515588 4616 515640 4622
rect 515588 4558 515640 4564
rect 513380 604 513432 610
rect 513380 546 513432 552
rect 514392 604 514444 610
rect 514392 546 514444 552
rect 514404 480 514432 546
rect 515600 480 515628 4558
rect 516796 480 516824 8842
rect 517532 626 517560 13602
rect 520280 13592 520332 13598
rect 520280 13534 520332 13540
rect 519084 4684 519136 4690
rect 519084 4626 519136 4632
rect 517532 598 517928 626
rect 517900 480 517928 598
rect 519096 480 519124 4626
rect 520292 3534 520320 13534
rect 524420 13524 524472 13530
rect 524420 13466 524472 13472
rect 520372 9648 520424 9654
rect 520372 9590 520424 9596
rect 520280 3528 520332 3534
rect 520280 3470 520332 3476
rect 520384 1442 520412 9590
rect 523868 9580 523920 9586
rect 523868 9522 523920 9528
rect 522672 4752 522724 4758
rect 522672 4694 522724 4700
rect 521476 3528 521528 3534
rect 521476 3470 521528 3476
rect 520292 1414 520412 1442
rect 520292 480 520320 1414
rect 521488 480 521516 3470
rect 522684 480 522712 4694
rect 523880 480 523908 9522
rect 524432 610 524460 13466
rect 528560 13456 528612 13462
rect 528560 13398 528612 13404
rect 527456 9512 527508 9518
rect 527456 9454 527508 9460
rect 526260 5500 526312 5506
rect 526260 5442 526312 5448
rect 524420 604 524472 610
rect 524420 546 524472 552
rect 525064 604 525116 610
rect 525064 546 525116 552
rect 525076 480 525104 546
rect 526272 480 526300 5442
rect 527468 480 527496 9454
rect 528572 592 528600 13398
rect 531320 13388 531372 13394
rect 531320 13330 531372 13336
rect 531044 9444 531096 9450
rect 531044 9386 531096 9392
rect 529848 5432 529900 5438
rect 529848 5374 529900 5380
rect 528572 564 528692 592
rect 528664 480 528692 564
rect 529860 480 529888 5374
rect 531056 480 531084 9386
rect 531332 610 531360 13330
rect 535460 13320 535512 13326
rect 535460 13262 535512 13268
rect 534540 9376 534592 9382
rect 534540 9318 534592 9324
rect 533436 5364 533488 5370
rect 533436 5306 533488 5312
rect 531320 604 531372 610
rect 531320 546 531372 552
rect 532240 604 532292 610
rect 532240 546 532292 552
rect 532252 480 532280 546
rect 533448 480 533476 5306
rect 534552 480 534580 9318
rect 535472 626 535500 13262
rect 538220 13252 538272 13258
rect 538220 13194 538272 13200
rect 538128 9308 538180 9314
rect 538128 9250 538180 9256
rect 536932 5296 536984 5302
rect 536932 5238 536984 5244
rect 535472 598 535684 626
rect 535656 592 535684 598
rect 535656 564 535776 592
rect 535748 480 535776 564
rect 536944 480 536972 5238
rect 538140 480 538168 9250
rect 538232 610 538260 13194
rect 542360 13184 542412 13190
rect 542360 13126 542412 13132
rect 541716 9240 541768 9246
rect 541716 9182 541768 9188
rect 540520 5228 540572 5234
rect 540520 5170 540572 5176
rect 538220 604 538272 610
rect 538220 546 538272 552
rect 539324 604 539376 610
rect 539324 546 539376 552
rect 539336 480 539364 546
rect 540532 480 540560 5170
rect 541728 480 541756 9182
rect 542372 610 542400 13126
rect 546500 13116 546552 13122
rect 546500 13058 546552 13064
rect 545302 9616 545358 9625
rect 545302 9551 545358 9560
rect 544108 5160 544160 5166
rect 544108 5102 544160 5108
rect 542360 604 542412 610
rect 542360 546 542412 552
rect 542912 604 542964 610
rect 542912 546 542964 552
rect 542924 480 542952 546
rect 544120 480 544148 5102
rect 545316 480 545344 9551
rect 546512 480 546540 13058
rect 548892 9172 548944 9178
rect 548892 9114 548944 9120
rect 547696 5092 547748 5098
rect 547696 5034 547748 5040
rect 547708 480 547736 5034
rect 548904 480 548932 9114
rect 549272 610 549300 13631
rect 553398 13560 553454 13569
rect 553398 13495 553454 13504
rect 552386 9480 552442 9489
rect 552386 9415 552442 9424
rect 551192 5024 551244 5030
rect 551192 4966 551244 4972
rect 549260 604 549312 610
rect 549260 546 549312 552
rect 550088 604 550140 610
rect 550088 546 550140 552
rect 550100 480 550128 546
rect 551204 480 551232 4966
rect 552400 480 552428 9415
rect 553412 626 553440 13495
rect 556158 13424 556214 13433
rect 556158 13359 556214 13368
rect 555974 9344 556030 9353
rect 555974 9279 556030 9288
rect 554778 5400 554834 5409
rect 554778 5335 554834 5344
rect 553412 598 553624 626
rect 553596 480 553624 598
rect 554792 480 554820 5335
rect 555988 480 556016 9279
rect 556172 610 556200 13359
rect 560298 13288 560354 13297
rect 560298 13223 560354 13232
rect 559562 9208 559618 9217
rect 559562 9143 559618 9152
rect 558366 5264 558422 5273
rect 558366 5199 558422 5208
rect 556160 604 556212 610
rect 556160 546 556212 552
rect 557172 604 557224 610
rect 557172 546 557224 552
rect 557184 480 557212 546
rect 558380 480 558408 5199
rect 559576 480 559604 9143
rect 560312 626 560340 13223
rect 563058 13152 563114 13161
rect 563058 13087 563114 13096
rect 561956 4956 562008 4962
rect 561956 4898 562008 4904
rect 560312 598 560800 626
rect 560772 480 560800 598
rect 561968 480 561996 4898
rect 563072 3534 563100 13087
rect 567198 13016 567254 13025
rect 567198 12951 567254 12960
rect 566740 9104 566792 9110
rect 563150 9072 563206 9081
rect 566740 9046 566792 9052
rect 563150 9007 563206 9016
rect 563060 3528 563112 3534
rect 563060 3470 563112 3476
rect 563164 480 563192 9007
rect 565542 5128 565598 5137
rect 565542 5063 565598 5072
rect 564348 3528 564400 3534
rect 564348 3470 564400 3476
rect 564360 480 564388 3470
rect 565556 480 565584 5063
rect 566752 480 566780 9046
rect 567212 3482 567240 12951
rect 570236 9036 570288 9042
rect 570236 8978 570288 8984
rect 569038 4992 569094 5001
rect 569038 4927 569094 4936
rect 567212 3454 567884 3482
rect 567856 480 567884 3454
rect 569052 480 569080 4927
rect 570248 480 570276 8978
rect 571352 3482 571380 14991
rect 574098 14920 574154 14929
rect 574098 14855 574154 14864
rect 573822 8936 573878 8945
rect 573822 8871 573878 8880
rect 572628 4888 572680 4894
rect 572628 4830 572680 4836
rect 571352 3454 571472 3482
rect 571444 480 571472 3454
rect 572640 480 572668 4830
rect 573836 480 573864 8871
rect 574112 3482 574140 14855
rect 576858 14784 576914 14793
rect 576858 14719 576914 14728
rect 576214 4856 576270 4865
rect 576214 4791 576270 4800
rect 574112 3454 575060 3482
rect 575032 480 575060 3454
rect 576228 480 576256 4791
rect 576872 610 576900 14719
rect 578238 14648 578294 14657
rect 578238 14583 578294 14592
rect 578252 626 578280 14583
rect 580998 14512 581054 14521
rect 580998 14447 581054 14456
rect 579804 4820 579856 4826
rect 579804 4762 579856 4768
rect 576860 604 576912 610
rect 576860 546 576912 552
rect 577412 604 577464 610
rect 578252 598 578648 626
rect 577412 546 577464 552
rect 577424 480 577452 546
rect 578620 480 578648 598
rect 579816 480 579844 4762
rect 581012 3534 581040 14447
rect 581092 8968 581144 8974
rect 581092 8910 581144 8916
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581104 1442 581132 8910
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 581012 1414 581132 1442
rect 581012 480 581040 1414
rect 582208 480 582236 3470
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 78586 655968 78642 656024
rect 187698 655968 187754 656024
rect 78494 654880 78550 654936
rect 78402 653112 78458 653168
rect 78310 652024 78366 652080
rect 78218 647536 78274 647592
rect 75826 568112 75882 568168
rect 73066 567840 73122 567896
rect 70950 523640 71006 523696
rect 77206 567976 77262 568032
rect 78678 650392 78734 650448
rect 78770 649168 78826 649224
rect 78862 589600 78918 589656
rect 103334 570288 103390 570344
rect 94870 570152 94926 570208
rect 98366 570152 98422 570208
rect 101770 570152 101826 570208
rect 86774 568520 86830 568576
rect 93766 568248 93822 568304
rect 95146 568540 95202 568576
rect 95146 568520 95148 568540
rect 95148 568520 95200 568540
rect 95200 568520 95202 568540
rect 95146 568384 95202 568440
rect 91098 567724 91154 567760
rect 91098 567704 91100 567724
rect 91100 567704 91152 567724
rect 91152 567704 91154 567724
rect 96526 568248 96582 568304
rect 97906 568248 97962 568304
rect 100666 568268 100722 568304
rect 100666 568248 100668 568268
rect 100668 568248 100720 568268
rect 100720 568248 100722 568268
rect 101954 568520 102010 568576
rect 102966 568520 103022 568576
rect 103150 568540 103206 568576
rect 103150 568520 103152 568540
rect 103152 568520 103204 568540
rect 103204 568520 103206 568540
rect 97906 567704 97962 567760
rect 100666 567724 100722 567760
rect 100666 567704 100668 567724
rect 100668 567704 100720 567724
rect 100720 567704 100722 567724
rect 88338 567432 88394 567488
rect 86958 567296 87014 567352
rect 89994 567316 90050 567352
rect 89994 567296 89996 567316
rect 89996 567296 90048 567316
rect 90048 567296 90050 567316
rect 93674 567160 93730 567216
rect 95054 567160 95110 567216
rect 96434 567160 96490 567216
rect 99194 567160 99250 567216
rect 102046 568248 102102 568304
rect 109038 570152 109094 570208
rect 112258 570152 112314 570208
rect 117962 570152 118018 570208
rect 119986 570152 120042 570208
rect 104070 568520 104126 568576
rect 104806 568520 104862 568576
rect 105266 568520 105322 568576
rect 106186 568520 106242 568576
rect 106646 568520 106702 568576
rect 107566 568520 107622 568576
rect 107750 568520 107806 568576
rect 108946 568520 109002 568576
rect 110326 568520 110382 568576
rect 110694 568520 110750 568576
rect 111706 568520 111762 568576
rect 109866 568384 109922 568440
rect 110326 567704 110382 567760
rect 113638 569744 113694 569800
rect 114466 569608 114522 569664
rect 117134 569608 117190 569664
rect 114742 568656 114798 568712
rect 115846 568520 115902 568576
rect 118330 569744 118386 569800
rect 118054 568656 118110 568712
rect 119434 569064 119490 569120
rect 119250 568928 119306 568984
rect 118514 566480 118570 566536
rect 120722 569744 120778 569800
rect 120078 569608 120134 569664
rect 120630 567332 120632 567352
rect 120632 567332 120684 567352
rect 120684 567332 120686 567352
rect 120630 567296 120686 567332
rect 120998 569064 121054 569120
rect 122746 568792 122802 568848
rect 122102 566072 122158 566128
rect 126610 568520 126666 568576
rect 128450 568540 128506 568576
rect 128450 568520 128452 568540
rect 128452 568520 128504 568540
rect 128504 568520 128506 568540
rect 124126 568248 124182 568304
rect 124310 568268 124366 568304
rect 124310 568248 124312 568268
rect 124312 568248 124364 568268
rect 124364 568248 124366 568268
rect 125506 568248 125562 568304
rect 124862 567704 124918 567760
rect 123482 567160 123538 567216
rect 125046 567296 125102 567352
rect 125322 567160 125378 567216
rect 125322 523912 125378 523968
rect 126886 567160 126942 567216
rect 127622 567160 127678 567216
rect 128174 567160 128230 567216
rect 126886 523776 126942 523832
rect 145562 568248 145618 568304
rect 145562 524048 145618 524104
rect 188342 654880 188398 654936
rect 152462 524184 152518 524240
rect 188434 653112 188490 653168
rect 188526 652024 188582 652080
rect 188618 650392 188674 650448
rect 188710 649168 188766 649224
rect 188802 647536 188858 647592
rect 188894 589600 188950 589656
rect 202786 570152 202842 570208
rect 220726 570152 220782 570208
rect 238758 570152 238814 570208
rect 195978 568520 196034 568576
rect 197450 568520 197506 568576
rect 202234 568520 202290 568576
rect 194414 568384 194470 568440
rect 194414 567588 194470 567624
rect 194414 567568 194416 567588
rect 194416 567568 194468 567588
rect 194468 567568 194470 567588
rect 202418 523912 202474 523968
rect 217874 569608 217930 569664
rect 204166 568520 204222 568576
rect 204810 568520 204866 568576
rect 205546 568520 205602 568576
rect 207018 568520 207074 568576
rect 209594 568540 209650 568576
rect 209594 568520 209596 568540
rect 209596 568520 209648 568540
rect 209648 568520 209650 568540
rect 203706 568384 203762 568440
rect 204350 524184 204406 524240
rect 197450 523640 197506 523696
rect 211894 568520 211950 568576
rect 213090 568520 213146 568576
rect 214102 568520 214158 568576
rect 215574 568520 215630 568576
rect 217138 568520 217194 568576
rect 209042 567332 209044 567352
rect 209044 567332 209096 567352
rect 209096 567332 209098 567352
rect 209042 567296 209098 567332
rect 206282 567196 206284 567216
rect 206284 567196 206336 567216
rect 206336 567196 206338 567216
rect 206282 567160 206338 567196
rect 206926 567160 206982 567216
rect 208306 567160 208362 567216
rect 206190 523776 206246 523832
rect 211066 567296 211122 567352
rect 209686 567160 209742 567216
rect 210422 567160 210478 567216
rect 210974 567160 211030 567216
rect 210054 524048 210110 524104
rect 218978 568520 219034 568576
rect 220082 568384 220138 568440
rect 217966 567296 218022 567352
rect 212446 567160 212502 567216
rect 213826 567160 213882 567216
rect 215206 567160 215262 567216
rect 216586 567160 216642 567216
rect 217874 567160 217930 567216
rect 219346 567160 219402 567216
rect 221462 568520 221518 568576
rect 222382 568520 222438 568576
rect 223670 568520 223726 568576
rect 225878 568520 225934 568576
rect 226246 568520 226302 568576
rect 227166 568520 227222 568576
rect 227626 568520 227682 568576
rect 228362 568520 228418 568576
rect 229006 568520 229062 568576
rect 229374 568520 229430 568576
rect 230386 568520 230442 568576
rect 231766 568520 231822 568576
rect 233054 568520 233110 568576
rect 234526 568520 234582 568576
rect 235906 568520 235962 568576
rect 237286 568520 237342 568576
rect 238666 568520 238722 568576
rect 226154 568384 226210 568440
rect 224774 568268 224830 568304
rect 224774 568248 224776 568268
rect 224776 568248 224828 568268
rect 224828 568248 224830 568268
rect 222106 567160 222162 567216
rect 223486 567160 223542 567216
rect 224866 567160 224922 567216
rect 230478 568112 230534 568168
rect 231950 568112 232006 568168
rect 231858 567996 231914 568032
rect 231858 567976 231860 567996
rect 231860 567976 231912 567996
rect 231912 567976 231914 567996
rect 233146 568384 233202 568440
rect 233238 568268 233294 568304
rect 233238 568248 233240 568268
rect 233240 568248 233292 568268
rect 233292 568248 233294 568268
rect 234618 568384 234674 568440
rect 235998 568132 236054 568168
rect 235998 568112 236000 568132
rect 236000 568112 236052 568132
rect 236052 568112 236054 568132
rect 237378 568248 237434 568304
rect 240046 568520 240102 568576
rect 273994 520920 274050 520976
rect 273626 515208 273682 515264
rect 273534 511400 273590 511456
rect 273718 507592 273774 507648
rect 273534 505688 273590 505744
rect 273534 503784 273590 503840
rect 273626 501880 273682 501936
rect 273718 499976 273774 500032
rect 273718 498072 273774 498128
rect 273718 496168 273774 496224
rect 273626 494264 273682 494320
rect 273626 492360 273682 492416
rect 273442 490456 273498 490512
rect 273626 488552 273682 488608
rect 273534 486648 273590 486704
rect 273626 484744 273682 484800
rect 273626 482840 273682 482896
rect 273626 480936 273682 480992
rect 273626 479032 273682 479088
rect 273626 477128 273682 477184
rect 273626 475224 273682 475280
rect 273626 473356 273628 473376
rect 273628 473356 273680 473376
rect 273680 473356 273682 473376
rect 273626 473320 273682 473356
rect 273258 463800 273314 463856
rect 273258 461896 273314 461952
rect 273258 460028 273260 460048
rect 273260 460028 273312 460048
rect 273312 460028 273314 460048
rect 273258 459992 273314 460028
rect 273258 458124 273260 458144
rect 273260 458124 273312 458144
rect 273312 458124 273314 458144
rect 273258 458088 273314 458124
rect 273258 456220 273260 456240
rect 273260 456220 273312 456240
rect 273312 456220 273314 456240
rect 273258 456184 273314 456220
rect 273258 454316 273260 454336
rect 273260 454316 273312 454336
rect 273312 454316 273314 454336
rect 273258 454280 273314 454316
rect 273258 452412 273260 452432
rect 273260 452412 273312 452432
rect 273312 452412 273314 452432
rect 273258 452376 273314 452412
rect 273350 450472 273406 450528
rect 273534 471416 273590 471472
rect 273534 469512 273590 469568
rect 273534 467608 273590 467664
rect 273534 465704 273590 465760
rect 273442 448568 273498 448624
rect 273442 446664 273498 446720
rect 273442 444796 273444 444816
rect 273444 444796 273496 444816
rect 273496 444796 273498 444816
rect 273442 444760 273498 444796
rect 273442 442892 273444 442912
rect 273444 442892 273496 442912
rect 273496 442892 273498 442912
rect 273442 442856 273498 442892
rect 273442 440952 273498 441008
rect 273442 439048 273498 439104
rect 273258 433372 273260 433392
rect 273260 433372 273312 433392
rect 273312 433372 273314 433392
rect 273258 433336 273314 433372
rect 273258 431468 273260 431488
rect 273260 431468 273312 431488
rect 273312 431468 273314 431488
rect 273258 431432 273314 431468
rect 273258 429564 273260 429584
rect 273260 429564 273312 429584
rect 273312 429564 273314 429584
rect 273258 429528 273314 429564
rect 273258 427660 273260 427680
rect 273260 427660 273312 427680
rect 273312 427660 273314 427680
rect 273258 427624 273314 427660
rect 273258 425756 273260 425776
rect 273260 425756 273312 425776
rect 273312 425756 273314 425776
rect 273258 425720 273314 425756
rect 273442 423816 273498 423872
rect 273442 421912 273498 421968
rect 273442 420044 273444 420064
rect 273444 420044 273496 420064
rect 273496 420044 273498 420064
rect 273442 420008 273498 420044
rect 273442 418124 273498 418160
rect 273442 418104 273444 418124
rect 273444 418104 273496 418124
rect 273496 418104 273498 418124
rect 273442 416236 273444 416256
rect 273444 416236 273496 416256
rect 273496 416236 273498 416256
rect 273442 416200 273498 416236
rect 273442 414332 273444 414352
rect 273444 414332 273496 414352
rect 273496 414332 273498 414352
rect 273442 414296 273498 414332
rect 273442 412428 273444 412448
rect 273444 412428 273496 412448
rect 273496 412428 273498 412448
rect 273442 412392 273498 412428
rect 273442 410524 273444 410544
rect 273444 410524 273496 410544
rect 273496 410524 273498 410544
rect 273442 410488 273498 410524
rect 273442 408620 273444 408640
rect 273444 408620 273496 408640
rect 273496 408620 273498 408640
rect 273442 408584 273498 408620
rect 273442 406716 273444 406736
rect 273444 406716 273496 406736
rect 273496 406716 273498 406736
rect 273442 406680 273498 406716
rect 273442 402908 273444 402928
rect 273444 402908 273496 402928
rect 273496 402908 273498 402928
rect 273442 402872 273498 402908
rect 273442 401004 273444 401024
rect 273444 401004 273496 401024
rect 273496 401004 273498 401024
rect 273442 400968 273498 401004
rect 273442 399064 273498 399120
rect 273442 397160 273498 397216
rect 273442 395256 273498 395312
rect 273442 393352 273498 393408
rect 273442 391448 273498 391504
rect 273534 389544 273590 389600
rect 273626 387640 273682 387696
rect 273534 385736 273590 385792
rect 273258 336232 273314 336288
rect 273350 330520 273406 330576
rect 273534 381928 273590 381984
rect 273626 380296 273682 380352
rect 273626 368600 273682 368656
rect 273810 364792 273866 364848
rect 273534 361020 273536 361040
rect 273536 361020 273588 361040
rect 273588 361020 273590 361040
rect 273534 360984 273590 361020
rect 273810 359080 273866 359136
rect 273810 353404 273812 353424
rect 273812 353404 273864 353424
rect 273864 353404 273866 353424
rect 273810 353368 273866 353404
rect 273534 349596 273536 349616
rect 273536 349596 273588 349616
rect 273588 349596 273590 349616
rect 273534 349560 273590 349596
rect 273534 347692 273536 347712
rect 273536 347692 273588 347712
rect 273588 347692 273590 347712
rect 273534 347656 273590 347692
rect 273534 345752 273590 345808
rect 273626 343848 273682 343904
rect 273534 341944 273590 342000
rect 273534 340076 273536 340096
rect 273536 340076 273588 340096
rect 273588 340076 273590 340096
rect 273534 340040 273590 340076
rect 274270 519016 274326 519072
rect 274086 517112 274142 517168
rect 274178 513304 274234 513360
rect 274270 509496 274326 509552
rect 274454 378120 274510 378176
rect 274454 376216 274510 376272
rect 274454 374312 274510 374368
rect 274454 372408 274510 372464
rect 274454 370524 274510 370560
rect 274454 370504 274456 370524
rect 274456 370504 274508 370524
rect 274508 370504 274510 370524
rect 274638 437144 274694 437200
rect 274730 435240 274786 435296
rect 274638 383832 274694 383888
rect 274546 366696 274602 366752
rect 274362 362888 274418 362944
rect 274362 355272 274418 355328
rect 274546 351464 274602 351520
rect 273902 338136 273958 338192
rect 273810 334328 273866 334384
rect 274270 332460 274272 332480
rect 274272 332460 274324 332480
rect 274324 332460 274326 332480
rect 274270 332424 274326 332460
rect 273994 328616 274050 328672
rect 273534 326712 273590 326768
rect 273442 324808 273498 324864
rect 273534 322904 273590 322960
rect 280066 396072 280122 396128
rect 337750 517384 337806 517440
rect 320178 516704 320234 516760
rect 398838 516724 398894 516760
rect 398838 516704 398840 516724
rect 398840 516704 398892 516724
rect 398892 516704 398894 516724
rect 400218 516604 400220 516624
rect 400220 516604 400272 516624
rect 400272 516604 400274 516624
rect 400218 516568 400274 516604
rect 401598 516588 401654 516624
rect 401598 516568 401600 516588
rect 401600 516568 401652 516588
rect 401652 516568 401654 516588
rect 338394 516432 338450 516488
rect 340878 516432 340934 516488
rect 403346 516468 403348 516488
rect 403348 516468 403400 516488
rect 403400 516468 403402 516488
rect 403346 516432 403402 516468
rect 404358 516452 404414 516488
rect 404358 516432 404360 516452
rect 404360 516432 404412 516452
rect 404412 516432 404414 516452
rect 406014 516452 406070 516488
rect 406014 516432 406016 516452
rect 406016 516432 406068 516452
rect 406068 516432 406070 516452
rect 320178 512080 320234 512136
rect 316682 509088 316738 509144
rect 319442 507864 319498 507920
rect 318798 363432 318854 363488
rect 320362 507456 320418 507512
rect 319810 506232 319866 506288
rect 320178 506232 320234 506288
rect 319810 500964 319812 500984
rect 319812 500964 319864 500984
rect 319864 500964 319866 500984
rect 319810 500928 319866 500964
rect 320730 504736 320786 504792
rect 320546 503648 320602 503704
rect 320178 503104 320234 503160
rect 319994 500792 320050 500848
rect 320362 502424 320418 502480
rect 320270 499568 320326 499624
rect 319810 497936 319866 497992
rect 320270 497800 320326 497856
rect 320178 497256 320234 497312
rect 319810 495216 319866 495272
rect 319810 493720 319866 493776
rect 320178 494944 320234 495000
rect 319994 492632 320050 492688
rect 319810 491136 319866 491192
rect 320178 490320 320234 490376
rect 320086 489812 320088 489832
rect 320088 489812 320140 489832
rect 320140 489812 320142 489832
rect 320086 489776 320142 489812
rect 320454 496576 320510 496632
rect 320362 493448 320418 493504
rect 320270 488416 320326 488472
rect 319810 487872 319866 487928
rect 320178 487872 320234 487928
rect 320270 487328 320326 487384
rect 319718 486648 319774 486704
rect 319810 485560 319866 485616
rect 320178 484472 320234 484528
rect 319810 483012 319812 483032
rect 319812 483012 319864 483032
rect 319864 483012 319866 483032
rect 319810 482976 319866 483012
rect 320178 482024 320234 482080
rect 320638 500112 320694 500168
rect 320822 501336 320878 501392
rect 320730 498888 320786 498944
rect 320546 494536 320602 494592
rect 320454 487328 320510 487384
rect 320822 495488 320878 495544
rect 320638 492224 320694 492280
rect 320638 490900 320640 490920
rect 320640 490900 320692 490920
rect 320692 490900 320694 490920
rect 320638 490864 320694 490900
rect 320730 488416 320786 488472
rect 320454 486104 320510 486160
rect 320362 484064 320418 484120
rect 319810 479712 319866 479768
rect 320178 479712 320234 479768
rect 320178 476720 320234 476776
rect 320546 484880 320602 484936
rect 320730 482704 320786 482760
rect 320638 482568 320694 482624
rect 320454 481480 320510 481536
rect 320638 482296 320694 482352
rect 320546 480256 320602 480312
rect 320362 476720 320418 476776
rect 320178 474408 320234 474464
rect 320454 475904 320510 475960
rect 320270 473320 320326 473376
rect 320270 473184 320326 473240
rect 320178 471008 320234 471064
rect 320638 479032 320694 479088
rect 320638 477944 320694 478000
rect 320730 475904 320786 475960
rect 320638 475768 320694 475824
rect 320362 472232 320418 472288
rect 320362 472096 320418 472152
rect 320270 470056 320326 470112
rect 320270 469784 320326 469840
rect 320178 468560 320234 468616
rect 320546 473184 320602 473240
rect 320454 471008 320510 471064
rect 320454 470872 320510 470928
rect 320362 469104 320418 469160
rect 320822 475788 320878 475824
rect 320822 475768 320824 475788
rect 320824 475768 320876 475788
rect 320876 475768 320878 475788
rect 320822 475496 320878 475552
rect 320730 474408 320786 474464
rect 320638 468832 320694 468888
rect 320178 465160 320234 465216
rect 320178 464888 320234 464944
rect 320638 467608 320694 467664
rect 320178 392028 320180 392048
rect 320180 392028 320232 392048
rect 320232 392028 320234 392048
rect 320178 391992 320234 392028
rect 320454 442312 320510 442368
rect 320730 442312 320786 442368
rect 320270 389816 320326 389872
rect 320086 389000 320142 389056
rect 338670 396788 338672 396808
rect 338672 396788 338724 396808
rect 338724 396788 338726 396808
rect 338670 396752 338726 396788
rect 397458 396772 397514 396808
rect 397458 396752 397460 396772
rect 397460 396752 397512 396772
rect 397512 396752 397514 396772
rect 398838 396652 398840 396672
rect 398840 396652 398892 396672
rect 398892 396652 398894 396672
rect 398838 396616 398894 396652
rect 400218 396636 400274 396672
rect 400218 396616 400220 396636
rect 400220 396616 400272 396636
rect 400272 396616 400274 396636
rect 401598 396516 401600 396536
rect 401600 396516 401652 396536
rect 401652 396516 401654 396536
rect 401598 396480 401654 396516
rect 403346 396500 403402 396536
rect 403346 396480 403348 396500
rect 403348 396480 403400 396500
rect 403400 396480 403402 396500
rect 404358 396480 404414 396536
rect 406014 396480 406070 396536
rect 320270 387504 320326 387560
rect 320362 386416 320418 386472
rect 320178 386280 320234 386336
rect 320178 383696 320234 383752
rect 320270 383152 320326 383208
rect 320638 384784 320694 384840
rect 320362 380840 320418 380896
rect 320270 379616 320326 379672
rect 320178 379480 320234 379536
rect 320178 377712 320234 377768
rect 319810 375128 319866 375184
rect 320178 376760 320234 376816
rect 320454 378936 320510 378992
rect 320362 376624 320418 376680
rect 320270 376080 320326 376136
rect 320178 375400 320234 375456
rect 319994 373768 320050 373824
rect 320086 373088 320142 373144
rect 320178 372680 320234 372736
rect 320362 372544 320418 372600
rect 320270 371456 320326 371512
rect 320178 368464 320234 368520
rect 320730 383560 320786 383616
rect 320638 381248 320694 381304
rect 320822 382472 320878 382528
rect 320822 380160 320878 380216
rect 320546 378392 320602 378448
rect 320546 374312 320602 374368
rect 320822 377712 320878 377768
rect 320730 376760 320786 376816
rect 320638 372272 320694 372328
rect 320822 371184 320878 371240
rect 320454 369688 320510 369744
rect 320362 369144 320418 369200
rect 320270 367920 320326 367976
rect 319810 365608 319866 365664
rect 320178 364928 320234 364984
rect 319994 363740 319996 363760
rect 319996 363740 320048 363760
rect 320048 363740 320050 363760
rect 319994 363704 320050 363740
rect 319810 361392 319866 361448
rect 320086 362652 320088 362672
rect 320088 362652 320140 362672
rect 320140 362652 320142 362672
rect 320086 362616 320142 362652
rect 320178 361392 320234 361448
rect 320730 369416 320786 369472
rect 320638 366152 320694 366208
rect 320454 364384 320510 364440
rect 320362 362072 320418 362128
rect 320270 360984 320326 361040
rect 320270 360304 320326 360360
rect 320454 359760 320510 359816
rect 320362 358536 320418 358592
rect 320270 357856 320326 357912
rect 320178 356768 320234 356824
rect 320178 355544 320234 355600
rect 320178 354456 320234 354512
rect 320638 364928 320694 364984
rect 320546 357040 320602 357096
rect 320270 353368 320326 353424
rect 320270 353232 320326 353288
rect 320178 352552 320234 352608
rect 320822 368464 320878 368520
rect 320822 367240 320878 367296
rect 320730 359760 320786 359816
rect 320638 355952 320694 356008
rect 320362 352416 320418 352472
rect 320638 351192 320694 351248
rect 320362 350920 320418 350976
rect 320178 349696 320234 349752
rect 320822 354592 320878 354648
rect 320822 353232 320878 353288
rect 320730 350104 320786 350160
rect 320178 348608 320234 348664
rect 320178 346332 320180 346352
rect 320180 346332 320232 346352
rect 320232 346332 320234 346352
rect 320178 346296 320234 346332
rect 273442 321000 273498 321056
rect 70306 320592 70362 320648
rect 23386 318552 23442 318608
rect 17866 318416 17922 318472
rect 16486 318280 16542 318336
rect 15106 318144 15162 318200
rect 13726 318008 13782 318064
rect 5262 3304 5318 3360
rect 10046 3440 10102 3496
rect 19522 3712 19578 3768
rect 18326 3576 18382 3632
rect 29090 3848 29146 3904
rect 42154 3984 42210 4040
rect 69018 318688 69074 318744
rect 70214 318688 70270 318744
rect 70766 135224 70822 135280
rect 70950 135224 71006 135280
rect 70766 77288 70822 77344
rect 70950 77288 71006 77344
rect 71686 3304 71742 3360
rect 72330 287000 72386 287056
rect 72514 287000 72570 287056
rect 72330 277380 72332 277400
rect 72332 277380 72384 277400
rect 72384 277380 72386 277400
rect 72330 277344 72386 277380
rect 72606 277344 72662 277400
rect 72054 182144 72110 182200
rect 72330 182144 72386 182200
rect 72238 87080 72294 87136
rect 72146 86944 72202 87000
rect 75918 318416 75974 318472
rect 75550 318280 75606 318336
rect 75090 318144 75146 318200
rect 74722 318008 74778 318064
rect 73434 277344 73490 277400
rect 73618 277344 73674 277400
rect 73434 231820 73436 231840
rect 73436 231820 73488 231840
rect 73488 231820 73490 231840
rect 73434 231784 73490 231820
rect 73710 231820 73712 231840
rect 73712 231820 73764 231840
rect 73764 231820 73766 231840
rect 73710 231784 73766 231820
rect 73434 212508 73436 212528
rect 73436 212508 73488 212528
rect 73488 212508 73490 212528
rect 73434 212472 73490 212508
rect 73710 212508 73712 212528
rect 73712 212508 73764 212528
rect 73764 212508 73766 212528
rect 73710 212472 73766 212508
rect 73342 182144 73398 182200
rect 73618 182144 73674 182200
rect 73342 162832 73398 162888
rect 73618 162832 73674 162888
rect 73434 86944 73490 87000
rect 73618 86944 73674 87000
rect 75918 3712 75974 3768
rect 78034 318552 78090 318608
rect 78678 267688 78734 267744
rect 78954 267688 79010 267744
rect 77482 248376 77538 248432
rect 77850 248376 77906 248432
rect 77482 202852 77484 202872
rect 77484 202852 77536 202872
rect 77536 202852 77538 202872
rect 77482 202816 77538 202852
rect 78770 202816 78826 202872
rect 78862 202680 78918 202736
rect 77574 195744 77630 195800
rect 77482 125568 77538 125624
rect 77666 125568 77722 125624
rect 78770 125568 78826 125624
rect 78954 125568 79010 125624
rect 77574 87080 77630 87136
rect 77482 86944 77538 87000
rect 81622 287000 81678 287056
rect 81806 287000 81862 287056
rect 81714 258032 81770 258088
rect 81898 258032 81954 258088
rect 81714 222164 81716 222184
rect 81716 222164 81768 222184
rect 81768 222164 81770 222184
rect 81714 222128 81770 222164
rect 81806 221992 81862 222048
rect 81714 183504 81770 183560
rect 81898 183504 81954 183560
rect 81898 133864 81954 133920
rect 82082 133864 82138 133920
rect 81714 125568 81770 125624
rect 81898 125568 81954 125624
rect 81806 87080 81862 87136
rect 81714 86944 81770 87000
rect 81806 66272 81862 66328
rect 81806 66000 81862 66056
rect 73342 3440 73398 3496
rect 76102 3576 76158 3632
rect 80150 3848 80206 3904
rect 80150 3304 80206 3360
rect 79782 3168 79838 3224
rect 80058 3168 80114 3224
rect 82542 3340 82544 3360
rect 82544 3340 82596 3360
rect 82596 3340 82598 3360
rect 82542 3304 82598 3340
rect 84290 3984 84346 4040
rect 90454 307808 90510 307864
rect 90178 307672 90234 307728
rect 89994 296656 90050 296712
rect 90270 296656 90326 296712
rect 89994 240080 90050 240136
rect 90178 240080 90234 240136
rect 90638 230424 90694 230480
rect 90822 230460 90824 230480
rect 90824 230460 90876 230480
rect 90876 230460 90878 230480
rect 90822 230424 90878 230460
rect 89994 193160 90050 193216
rect 90178 193160 90234 193216
rect 91190 162832 91246 162888
rect 91098 162560 91154 162616
rect 91098 153176 91154 153232
rect 91190 153040 91246 153096
rect 89994 135360 90050 135416
rect 89994 135224 90050 135280
rect 89994 115932 90050 115968
rect 89994 115912 89996 115932
rect 89996 115912 90048 115932
rect 90048 115912 90050 115932
rect 90178 115932 90234 115968
rect 90178 115912 90180 115932
rect 90180 115912 90232 115932
rect 90232 115912 90234 115932
rect 91006 114552 91062 114608
rect 91190 114552 91246 114608
rect 89994 96600 90050 96656
rect 90178 96600 90234 96656
rect 91006 85448 91062 85504
rect 91098 85312 91154 85368
rect 92754 212472 92810 212528
rect 92938 212472 92994 212528
rect 92754 135360 92810 135416
rect 92754 135224 92810 135280
rect 92754 115932 92810 115968
rect 92754 115912 92756 115932
rect 92756 115912 92808 115932
rect 92808 115912 92810 115932
rect 92938 115932 92994 115968
rect 92938 115912 92940 115932
rect 92940 115912 92992 115932
rect 92992 115912 92994 115932
rect 92754 96600 92810 96656
rect 92938 96600 92994 96656
rect 94134 287000 94190 287056
rect 94318 287000 94374 287056
rect 94042 222128 94098 222184
rect 94318 222128 94374 222184
rect 94134 162832 94190 162888
rect 94318 162832 94374 162888
rect 94134 133864 94190 133920
rect 94318 133864 94374 133920
rect 94134 106528 94190 106584
rect 94042 106256 94098 106312
rect 94042 87080 94098 87136
rect 94042 86944 94098 87000
rect 96986 60696 97042 60752
rect 96986 56616 97042 56672
rect 105174 298016 105230 298072
rect 105358 298016 105414 298072
rect 104898 164192 104954 164248
rect 105082 164192 105138 164248
rect 106646 241440 106702 241496
rect 106554 235320 106610 235376
rect 106646 193160 106702 193216
rect 106830 193160 106886 193216
rect 106462 173848 106518 173904
rect 106738 173884 106740 173904
rect 106740 173884 106792 173904
rect 106792 173884 106794 173904
rect 106738 173848 106794 173884
rect 106462 164192 106518 164248
rect 106646 164212 106702 164248
rect 106646 164192 106648 164212
rect 106648 164192 106700 164212
rect 106700 164192 106702 164212
rect 125322 3168 125378 3224
rect 129554 3984 129610 4040
rect 128266 3440 128322 3496
rect 130934 3848 130990 3904
rect 132314 3712 132370 3768
rect 143170 318008 143226 318064
rect 144826 3304 144882 3360
rect 147402 318144 147458 318200
rect 147862 318164 147918 318200
rect 147862 318144 147864 318164
rect 147864 318144 147916 318164
rect 147916 318144 147918 318164
rect 151082 241440 151138 241496
rect 150990 241304 151046 241360
rect 151082 222128 151138 222184
rect 150990 221992 151046 222048
rect 151082 202816 151138 202872
rect 150990 202680 151046 202736
rect 151082 183504 151138 183560
rect 150990 183368 151046 183424
rect 151082 9594 151138 9650
rect 153198 9424 153254 9480
rect 151726 2916 151782 2952
rect 151726 2896 151728 2916
rect 151728 2896 151780 2916
rect 151780 2896 151782 2916
rect 158626 5344 158682 5400
rect 158074 3576 158130 3632
rect 160006 5208 160062 5264
rect 157246 2932 157248 2952
rect 157248 2932 157300 2952
rect 157300 2932 157302 2952
rect 157246 2896 157302 2932
rect 159914 3168 159970 3224
rect 163502 318008 163558 318064
rect 161386 5072 161442 5128
rect 162766 4936 162822 4992
rect 164238 318724 164240 318744
rect 164240 318724 164292 318744
rect 164292 318724 164294 318744
rect 164238 318688 164294 318724
rect 164146 4800 164202 4856
rect 166998 318724 167000 318744
rect 167000 318724 167052 318744
rect 167052 318724 167054 318744
rect 166998 318688 167054 318724
rect 166906 5480 166962 5536
rect 165894 3440 165950 3496
rect 166262 3440 166318 3496
rect 171782 3984 171838 4040
rect 175370 3848 175426 3904
rect 178958 3712 179014 3768
rect 193678 278704 193734 278760
rect 193862 278704 193918 278760
rect 193678 259392 193734 259448
rect 193862 259392 193918 259448
rect 193862 241712 193918 241768
rect 193862 241576 193918 241632
rect 193678 240080 193734 240136
rect 193862 240080 193918 240136
rect 193678 220768 193734 220824
rect 193862 220768 193918 220824
rect 193678 211112 193734 211168
rect 193862 211112 193918 211168
rect 193678 191800 193734 191856
rect 193862 191800 193918 191856
rect 193678 172488 193734 172544
rect 193862 172488 193918 172544
rect 194414 6704 194470 6760
rect 195702 10784 195758 10840
rect 197082 10648 197138 10704
rect 195886 6568 195942 6624
rect 198554 10512 198610 10568
rect 197266 6432 197322 6488
rect 199842 10376 199898 10432
rect 198646 6296 198702 6352
rect 199934 6160 199990 6216
rect 201314 10240 201370 10296
rect 204810 154672 204866 154728
rect 204902 154536 204958 154592
rect 204810 135360 204866 135416
rect 204902 135224 204958 135280
rect 205638 8780 205640 8800
rect 205640 8780 205692 8800
rect 205692 8780 205694 8800
rect 205638 8744 205694 8780
rect 207478 3576 207534 3632
rect 211710 183504 211766 183560
rect 211894 183504 211950 183560
rect 215114 8780 215116 8800
rect 215116 8780 215168 8800
rect 215168 8780 215170 8800
rect 215114 8744 215170 8780
rect 215114 4664 215170 4720
rect 215574 4664 215630 4720
rect 215114 4392 215170 4448
rect 215298 4428 215300 4448
rect 215300 4428 215352 4448
rect 215352 4428 215354 4448
rect 215298 4392 215354 4428
rect 214654 3304 214710 3360
rect 218150 3440 218206 3496
rect 224958 8780 224960 8800
rect 224960 8780 225012 8800
rect 225012 8780 225014 8800
rect 224958 8744 225014 8780
rect 224866 3848 224922 3904
rect 227258 318144 227314 318200
rect 227166 183504 227222 183560
rect 227350 183504 227406 183560
rect 227442 22072 227498 22128
rect 227350 19352 227406 19408
rect 229742 318552 229798 318608
rect 228914 8200 228970 8256
rect 226246 3712 226302 3768
rect 232226 318008 232282 318064
rect 231490 12280 231546 12336
rect 231582 12144 231638 12200
rect 230386 8064 230442 8120
rect 231674 7928 231730 7984
rect 229006 3576 229062 3632
rect 234710 318280 234766 318336
rect 233054 12008 233110 12064
rect 233974 296656 234030 296712
rect 234250 296656 234306 296712
rect 233790 217912 233846 217968
rect 234066 217912 234122 217968
rect 234158 173848 234214 173904
rect 234342 173848 234398 173904
rect 233146 7792 233202 7848
rect 234434 8372 234436 8392
rect 234436 8372 234488 8392
rect 234488 8372 234490 8392
rect 234434 8336 234490 8372
rect 234342 7656 234398 7712
rect 231766 3440 231822 3496
rect 237194 318552 237250 318608
rect 235538 180784 235594 180840
rect 235722 180804 235778 180840
rect 235722 180784 235724 180804
rect 235724 180784 235776 180804
rect 235776 180784 235778 180804
rect 235538 154536 235594 154592
rect 235722 154536 235778 154592
rect 234618 11872 234674 11928
rect 235814 11736 235870 11792
rect 239862 15136 239918 15192
rect 237286 11600 237342 11656
rect 239586 8744 239642 8800
rect 235906 7520 235962 7576
rect 234526 3304 234582 3360
rect 239770 8336 239826 8392
rect 242346 249736 242402 249792
rect 242530 249736 242586 249792
rect 242346 230424 242402 230480
rect 242530 230424 242586 230480
rect 242346 201456 242402 201512
rect 242530 201456 242586 201512
rect 242346 182144 242402 182200
rect 242530 182144 242586 182200
rect 243634 46824 243690 46880
rect 243818 46824 243874 46880
rect 244094 9152 244150 9208
rect 244186 4528 244242 4584
rect 246946 259392 247002 259448
rect 247130 259392 247186 259448
rect 246946 240080 247002 240136
rect 247130 240080 247186 240136
rect 246946 220768 247002 220824
rect 247130 220768 247186 220824
rect 246946 211112 247002 211168
rect 247130 211112 247186 211168
rect 246946 191800 247002 191856
rect 247130 191800 247186 191856
rect 246946 172488 247002 172544
rect 247130 172488 247186 172544
rect 246946 133864 247002 133920
rect 247130 133864 247186 133920
rect 248234 133864 248290 133920
rect 246946 9832 247002 9888
rect 248142 8608 248198 8664
rect 248418 133864 248474 133920
rect 249430 133864 249486 133920
rect 249614 133864 249670 133920
rect 249246 9424 249302 9480
rect 249062 4528 249118 4584
rect 249338 9152 249394 9208
rect 250810 240080 250866 240136
rect 250810 220768 250866 220824
rect 250810 211112 250866 211168
rect 250810 172488 250866 172544
rect 250810 153176 250866 153232
rect 250994 240080 251050 240136
rect 250994 220768 251050 220824
rect 250994 211112 251050 211168
rect 250994 172488 251050 172544
rect 250994 153176 251050 153232
rect 250994 133864 251050 133920
rect 249798 8608 249854 8664
rect 252098 240080 252154 240136
rect 252098 220768 252154 220824
rect 252098 211112 252154 211168
rect 252098 172488 252154 172544
rect 252098 153176 252154 153232
rect 251178 133864 251234 133920
rect 252098 133864 252154 133920
rect 252098 86944 252154 87000
rect 252282 240080 252338 240136
rect 252282 220768 252338 220824
rect 252282 211112 252338 211168
rect 252282 172488 252338 172544
rect 252282 153176 252338 153232
rect 252282 133864 252338 133920
rect 252282 86944 252338 87000
rect 252926 309168 252982 309224
rect 252742 309032 252798 309088
rect 255226 278704 255282 278760
rect 255318 278568 255374 278624
rect 255318 219408 255374 219464
rect 255502 219408 255558 219464
rect 255226 153176 255282 153232
rect 255410 153176 255466 153232
rect 255226 143384 255282 143440
rect 255410 133864 255466 133920
rect 255226 125568 255282 125624
rect 255410 125568 255466 125624
rect 255042 5344 255098 5400
rect 256698 15136 256754 15192
rect 256698 14728 256754 14784
rect 259090 240080 259146 240136
rect 259090 220768 259146 220824
rect 259090 211112 259146 211168
rect 259090 172488 259146 172544
rect 259090 153176 259146 153232
rect 259090 125568 259146 125624
rect 259090 106256 259146 106312
rect 259274 240080 259330 240136
rect 259274 220768 259330 220824
rect 259274 211112 259330 211168
rect 259274 172488 259330 172544
rect 259274 153176 259330 153232
rect 259274 125568 259330 125624
rect 259274 106256 259330 106312
rect 260286 180784 260342 180840
rect 260470 180784 260526 180840
rect 260562 13640 260618 13696
rect 259182 9560 259238 9616
rect 258630 5208 258686 5264
rect 261942 13504 261998 13560
rect 262218 13776 262274 13832
rect 262402 13776 262458 13832
rect 263230 13368 263286 13424
rect 262402 9424 262458 9480
rect 263230 9288 263286 9344
rect 263230 5208 263286 5264
rect 262218 5072 262274 5128
rect 263690 293936 263746 293992
rect 264702 293936 264758 293992
rect 264518 274624 264574 274680
rect 264702 274644 264758 274680
rect 264702 274624 264704 274644
rect 264704 274624 264756 274644
rect 264756 274624 264758 274644
rect 264794 133864 264850 133920
rect 264702 15136 264758 15192
rect 264794 9152 264850 9208
rect 263506 5344 263562 5400
rect 265346 314608 265402 314664
rect 265806 314608 265862 314664
rect 264978 133864 265034 133920
rect 265162 15000 265218 15056
rect 265162 13232 265218 13288
rect 266082 13096 266138 13152
rect 266174 9016 266230 9072
rect 267094 180784 267150 180840
rect 267278 180784 267334 180840
rect 267370 12960 267426 13016
rect 266266 5072 266322 5128
rect 265806 4936 265862 4992
rect 267646 4936 267702 4992
rect 268842 15000 268898 15056
rect 270314 14864 270370 14920
rect 270222 14728 270278 14784
rect 268934 8880 268990 8936
rect 271510 14592 271566 14648
rect 271602 14456 271658 14512
rect 269302 4800 269358 4856
rect 270406 4800 270462 4856
rect 276478 5480 276534 5536
rect 324870 231784 324926 231840
rect 325054 231784 325110 231840
rect 324870 212472 324926 212528
rect 325054 212472 325110 212528
rect 324870 193160 324926 193216
rect 325054 193160 325110 193216
rect 324870 173848 324926 173904
rect 325054 173848 325110 173904
rect 324962 144880 325018 144936
rect 325238 144880 325294 144936
rect 324962 125568 325018 125624
rect 325238 125568 325294 125624
rect 324962 106256 325018 106312
rect 325238 106256 325294 106312
rect 345018 4140 345074 4176
rect 345018 4120 345020 4140
rect 345020 4120 345072 4140
rect 345072 4120 345074 4140
rect 354586 4140 354642 4176
rect 354586 4120 354588 4140
rect 354588 4120 354640 4140
rect 354640 4120 354642 4140
rect 374642 318552 374698 318608
rect 367742 318416 367798 318472
rect 358542 6704 358598 6760
rect 356702 3168 356758 3224
rect 364982 318144 365038 318200
rect 362958 10784 363014 10840
rect 362130 6568 362186 6624
rect 359646 3168 359702 3224
rect 365718 10648 365774 10704
rect 364890 4020 364892 4040
rect 364892 4020 364944 4040
rect 364944 4020 364946 4040
rect 364890 3984 364946 4020
rect 365810 6432 365866 6488
rect 373262 318280 373318 318336
rect 371882 318008 371938 318064
rect 369858 10512 369914 10568
rect 369214 6296 369270 6352
rect 367006 3984 367062 4040
rect 372802 6160 372858 6216
rect 374090 10376 374146 10432
rect 373262 3984 373318 4040
rect 376758 10240 376814 10296
rect 462318 12280 462374 12336
rect 442998 3848 443054 3904
rect 450174 3712 450230 3768
rect 458454 8200 458510 8256
rect 457258 3576 457314 3632
rect 462042 8064 462098 8120
rect 466458 12144 466514 12200
rect 465630 7928 465686 7984
rect 464434 3440 464490 3496
rect 469218 12008 469274 12064
rect 469126 7792 469182 7848
rect 473358 11872 473414 11928
rect 472714 7656 472770 7712
rect 471518 3304 471574 3360
rect 476302 7520 476358 7576
rect 475106 3984 475162 4040
rect 489918 15136 489974 15192
rect 477590 11736 477646 11792
rect 480258 11600 480314 11656
rect 571338 15000 571394 15056
rect 549258 13640 549314 13696
rect 545302 9560 545358 9616
rect 553398 13504 553454 13560
rect 552386 9424 552442 9480
rect 556158 13368 556214 13424
rect 555974 9288 556030 9344
rect 554778 5344 554834 5400
rect 560298 13232 560354 13288
rect 559562 9152 559618 9208
rect 558366 5208 558422 5264
rect 563058 13096 563114 13152
rect 567198 12960 567254 13016
rect 563150 9016 563206 9072
rect 565542 5072 565598 5128
rect 569038 4936 569094 4992
rect 574098 14864 574154 14920
rect 573822 8880 573878 8936
rect 576858 14728 576914 14784
rect 576214 4800 576270 4856
rect 578238 14592 578294 14648
rect 580998 14456 581054 14512
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696540 480 696780
rect 583520 686204 584960 686444
rect -960 682124 480 682364
rect 583520 674508 584960 674748
rect -960 667844 480 668084
rect 583520 662676 584960 662916
rect 78581 656026 78647 656029
rect 80102 656026 80162 656587
rect 78581 656024 80162 656026
rect 78581 655968 78586 656024
rect 78642 655968 80162 656024
rect 78581 655966 80162 655968
rect 187693 656026 187759 656029
rect 190134 656026 190194 656587
rect 187693 656024 190194 656026
rect 187693 655968 187698 656024
rect 187754 655968 190194 656024
rect 187693 655966 190194 655968
rect 78581 655963 78647 655966
rect 187693 655963 187759 655966
rect 78489 654938 78555 654941
rect 80102 654938 80162 655459
rect 78489 654936 80162 654938
rect 78489 654880 78494 654936
rect 78550 654880 80162 654936
rect 78489 654878 80162 654880
rect 188337 654938 188403 654941
rect 190134 654938 190194 655459
rect 188337 654936 190194 654938
rect 188337 654880 188342 654936
rect 188398 654880 190194 654936
rect 188337 654878 190194 654880
rect 78489 654875 78555 654878
rect 188337 654875 188403 654878
rect -960 653428 480 653668
rect 78397 653170 78463 653173
rect 80102 653170 80162 653759
rect 78397 653168 80162 653170
rect 78397 653112 78402 653168
rect 78458 653112 80162 653168
rect 78397 653110 80162 653112
rect 188429 653170 188495 653173
rect 190134 653170 190194 653759
rect 188429 653168 190194 653170
rect 188429 653112 188434 653168
rect 188490 653112 190194 653168
rect 188429 653110 190194 653112
rect 78397 653107 78463 653110
rect 188429 653107 188495 653110
rect 78305 652082 78371 652085
rect 80102 652082 80162 652631
rect 78305 652080 80162 652082
rect 78305 652024 78310 652080
rect 78366 652024 80162 652080
rect 78305 652022 80162 652024
rect 188521 652082 188587 652085
rect 190134 652082 190194 652631
rect 188521 652080 190194 652082
rect 188521 652024 188526 652080
rect 188582 652024 190194 652080
rect 188521 652022 190194 652024
rect 78305 652019 78371 652022
rect 188521 652019 188587 652022
rect 583520 650980 584960 651220
rect 78673 650450 78739 650453
rect 80102 650450 80162 650931
rect 78673 650448 80162 650450
rect 78673 650392 78678 650448
rect 78734 650392 80162 650448
rect 78673 650390 80162 650392
rect 188613 650450 188679 650453
rect 190134 650450 190194 650931
rect 188613 650448 190194 650450
rect 188613 650392 188618 650448
rect 188674 650392 190194 650448
rect 188613 650390 190194 650392
rect 78673 650387 78739 650390
rect 188613 650387 188679 650390
rect 78765 649226 78831 649229
rect 80102 649226 80162 649803
rect 78765 649224 80162 649226
rect 78765 649168 78770 649224
rect 78826 649168 80162 649224
rect 78765 649166 80162 649168
rect 188705 649226 188771 649229
rect 190134 649226 190194 649803
rect 188705 649224 190194 649226
rect 188705 649168 188710 649224
rect 188766 649168 190194 649224
rect 188705 649166 190194 649168
rect 78765 649163 78831 649166
rect 188705 649163 188771 649166
rect 78213 647594 78279 647597
rect 80102 647594 80162 648103
rect 78213 647592 80162 647594
rect 78213 647536 78218 647592
rect 78274 647536 80162 647592
rect 78213 647534 80162 647536
rect 188797 647594 188863 647597
rect 190134 647594 190194 648103
rect 188797 647592 190194 647594
rect 188797 647536 188802 647592
rect 188858 647536 190194 647592
rect 188797 647534 190194 647536
rect 78213 647531 78279 647534
rect 188797 647531 188863 647534
rect 583520 639284 584960 639524
rect -960 639012 480 639252
rect 583520 627588 584960 627828
rect -960 624732 480 624972
rect 583520 615756 584960 615996
rect -960 610316 480 610556
rect 583520 604060 584960 604300
rect -960 595900 480 596140
rect 583520 592364 584960 592604
rect 78857 589658 78923 589661
rect 80102 589658 80162 590255
rect 78857 589656 80162 589658
rect 78857 589600 78862 589656
rect 78918 589600 80162 589656
rect 78857 589598 80162 589600
rect 188889 589658 188955 589661
rect 190134 589658 190194 590255
rect 188889 589656 190194 589658
rect 188889 589600 188894 589656
rect 188950 589600 190194 589656
rect 188889 589598 190194 589600
rect 78857 589595 78923 589598
rect 188889 589595 188955 589598
rect -960 581620 480 581860
rect 583520 580668 584960 580908
rect 103329 570346 103395 570349
rect 103462 570346 103468 570348
rect 103329 570344 103468 570346
rect 103329 570288 103334 570344
rect 103390 570288 103468 570344
rect 103329 570286 103468 570288
rect 103329 570283 103395 570286
rect 103462 570284 103468 570286
rect 103532 570284 103538 570348
rect 94865 570212 94931 570213
rect 98361 570212 98427 570213
rect 94814 570148 94820 570212
rect 94884 570210 94931 570212
rect 94884 570208 94976 570210
rect 94926 570152 94976 570208
rect 94884 570150 94976 570152
rect 94884 570148 94931 570150
rect 98310 570148 98316 570212
rect 98380 570210 98427 570212
rect 101765 570212 101831 570213
rect 98380 570208 98472 570210
rect 98422 570152 98472 570208
rect 98380 570150 98472 570152
rect 101765 570208 101812 570212
rect 101876 570210 101882 570212
rect 101765 570152 101770 570208
rect 98380 570148 98427 570150
rect 94865 570147 94931 570148
rect 98361 570147 98427 570148
rect 101765 570148 101812 570152
rect 101876 570150 101922 570210
rect 101876 570148 101882 570150
rect 108798 570148 108804 570212
rect 108868 570210 108874 570212
rect 109033 570210 109099 570213
rect 108868 570208 109099 570210
rect 108868 570152 109038 570208
rect 109094 570152 109099 570208
rect 108868 570150 109099 570152
rect 108868 570148 108874 570150
rect 101765 570147 101831 570148
rect 109033 570147 109099 570150
rect 112253 570212 112319 570213
rect 112253 570208 112300 570212
rect 112364 570210 112370 570212
rect 112253 570152 112258 570208
rect 112253 570148 112300 570152
rect 112364 570150 112410 570210
rect 112364 570148 112370 570150
rect 113214 570148 113220 570212
rect 113284 570210 113290 570212
rect 117957 570210 118023 570213
rect 113284 570208 118023 570210
rect 113284 570152 117962 570208
rect 118018 570152 118023 570208
rect 113284 570150 118023 570152
rect 113284 570148 113290 570150
rect 112253 570147 112319 570148
rect 117957 570147 118023 570150
rect 119838 570148 119844 570212
rect 119908 570210 119914 570212
rect 119981 570210 120047 570213
rect 119908 570208 120047 570210
rect 119908 570152 119986 570208
rect 120042 570152 120047 570208
rect 119908 570150 120047 570152
rect 119908 570148 119914 570150
rect 119981 570147 120047 570150
rect 202781 570210 202847 570213
rect 220721 570212 220787 570213
rect 238753 570212 238819 570213
rect 203006 570210 203012 570212
rect 202781 570208 203012 570210
rect 202781 570152 202786 570208
rect 202842 570152 203012 570208
rect 202781 570150 203012 570152
rect 202781 570147 202847 570150
rect 203006 570148 203012 570150
rect 203076 570148 203082 570212
rect 220670 570148 220676 570212
rect 220740 570210 220787 570212
rect 220740 570208 220832 570210
rect 220782 570152 220832 570208
rect 220740 570150 220832 570152
rect 220740 570148 220787 570150
rect 238702 570148 238708 570212
rect 238772 570210 238819 570212
rect 238772 570208 238864 570210
rect 238814 570152 238864 570208
rect 238772 570150 238864 570152
rect 238772 570148 238819 570150
rect 220721 570147 220787 570148
rect 238753 570147 238819 570148
rect 113633 569804 113699 569805
rect 118325 569804 118391 569805
rect 120717 569804 120783 569805
rect 113633 569800 113664 569804
rect 113728 569802 113734 569804
rect 113633 569744 113638 569800
rect 113633 569740 113664 569744
rect 113728 569742 113790 569802
rect 118325 569800 118336 569804
rect 118400 569802 118406 569804
rect 118325 569744 118330 569800
rect 113728 569740 113734 569742
rect 118325 569740 118336 569744
rect 118400 569742 118482 569802
rect 118400 569740 118406 569742
rect 120666 569740 120672 569804
rect 120736 569802 120783 569804
rect 120736 569800 120828 569802
rect 120778 569744 120828 569800
rect 120736 569742 120828 569744
rect 120736 569740 120783 569742
rect 113633 569739 113699 569740
rect 118325 569739 118391 569740
rect 120717 569739 120783 569740
rect 113782 569604 113788 569668
rect 113852 569666 113858 569668
rect 114461 569666 114527 569669
rect 117129 569668 117195 569669
rect 117129 569666 117168 569668
rect 113852 569664 114527 569666
rect 113852 569608 114466 569664
rect 114522 569608 114527 569664
rect 113852 569606 114527 569608
rect 117076 569664 117168 569666
rect 117076 569608 117134 569664
rect 117076 569606 117168 569608
rect 113852 569604 113858 569606
rect 114461 569603 114527 569606
rect 117129 569604 117168 569606
rect 117232 569604 117238 569668
rect 118454 569604 118460 569668
rect 118524 569666 118530 569668
rect 120073 569666 120139 569669
rect 217869 569668 217935 569669
rect 217818 569666 217824 569668
rect 118524 569664 120139 569666
rect 118524 569608 120078 569664
rect 120134 569608 120139 569664
rect 118524 569606 120139 569608
rect 217778 569606 217824 569666
rect 217888 569664 217935 569668
rect 217930 569608 217935 569664
rect 118524 569604 118530 569606
rect 117129 569603 117195 569604
rect 120073 569603 120139 569606
rect 217818 569604 217824 569606
rect 217888 569604 217935 569608
rect 217869 569603 217935 569604
rect 119429 569124 119495 569125
rect 120993 569124 121059 569125
rect 119429 569120 119476 569124
rect 119540 569122 119546 569124
rect 120942 569122 120948 569124
rect 119429 569064 119434 569120
rect 119429 569060 119476 569064
rect 119540 569062 119586 569122
rect 120902 569062 120948 569122
rect 121012 569120 121059 569124
rect 121054 569064 121059 569120
rect 119540 569060 119546 569062
rect 120942 569060 120948 569062
rect 121012 569060 121059 569064
rect 119429 569059 119495 569060
rect 120993 569059 121059 569060
rect 116710 568924 116716 568988
rect 116780 568986 116786 568988
rect 119245 568986 119311 568989
rect 116780 568984 119311 568986
rect 116780 568928 119250 568984
rect 119306 568928 119311 568984
rect 116780 568926 119311 568928
rect 116780 568924 116786 568926
rect 119245 568923 119311 568926
rect 122598 568788 122604 568852
rect 122668 568850 122674 568852
rect 122741 568850 122807 568853
rect 122668 568848 122807 568850
rect 122668 568792 122746 568848
rect 122802 568792 122807 568848
rect 583520 568836 584960 569076
rect 122668 568790 122807 568792
rect 122668 568788 122674 568790
rect 122741 568787 122807 568790
rect 114737 568716 114803 568717
rect 114686 568714 114692 568716
rect 114646 568654 114692 568714
rect 114756 568712 114803 568716
rect 114798 568656 114803 568712
rect 114686 568652 114692 568654
rect 114756 568652 114803 568656
rect 115054 568652 115060 568716
rect 115124 568714 115130 568716
rect 118049 568714 118115 568717
rect 115124 568712 118115 568714
rect 115124 568656 118054 568712
rect 118110 568656 118115 568712
rect 115124 568654 118115 568656
rect 115124 568652 115130 568654
rect 114737 568651 114803 568652
rect 118049 568651 118115 568654
rect 86534 568516 86540 568580
rect 86604 568578 86610 568580
rect 86769 568578 86835 568581
rect 86604 568576 86835 568578
rect 86604 568520 86774 568576
rect 86830 568520 86835 568576
rect 86604 568518 86835 568520
rect 86604 568516 86610 568518
rect 86769 568515 86835 568518
rect 93894 568516 93900 568580
rect 93964 568578 93970 568580
rect 95141 568578 95207 568581
rect 93964 568576 95207 568578
rect 93964 568520 95146 568576
rect 95202 568520 95207 568576
rect 93964 568518 95207 568520
rect 93964 568516 93970 568518
rect 95141 568515 95207 568518
rect 101438 568516 101444 568580
rect 101508 568578 101514 568580
rect 101949 568578 102015 568581
rect 101508 568576 102015 568578
rect 101508 568520 101954 568576
rect 102010 568520 102015 568576
rect 101508 568518 102015 568520
rect 101508 568516 101514 568518
rect 101949 568515 102015 568518
rect 102726 568516 102732 568580
rect 102796 568578 102802 568580
rect 102961 568578 103027 568581
rect 103145 568580 103211 568581
rect 104065 568580 104131 568581
rect 104801 568580 104867 568581
rect 102796 568576 103027 568578
rect 102796 568520 102966 568576
rect 103022 568520 103027 568576
rect 102796 568518 103027 568520
rect 102796 568516 102802 568518
rect 102961 568515 103027 568518
rect 103094 568516 103100 568580
rect 103164 568578 103211 568580
rect 104014 568578 104020 568580
rect 103164 568576 103256 568578
rect 103206 568520 103256 568576
rect 103164 568518 103256 568520
rect 103974 568518 104020 568578
rect 104084 568576 104131 568580
rect 104126 568520 104131 568576
rect 103164 568516 103211 568518
rect 104014 568516 104020 568518
rect 104084 568516 104131 568520
rect 104750 568516 104756 568580
rect 104820 568578 104867 568580
rect 105261 568580 105327 568581
rect 104820 568576 104912 568578
rect 104862 568520 104912 568576
rect 104820 568518 104912 568520
rect 105261 568576 105308 568580
rect 105372 568578 105378 568580
rect 105261 568520 105266 568576
rect 104820 568516 104867 568518
rect 103145 568515 103211 568516
rect 104065 568515 104131 568516
rect 104801 568515 104867 568516
rect 105261 568516 105308 568520
rect 105372 568518 105418 568578
rect 105372 568516 105378 568518
rect 105854 568516 105860 568580
rect 105924 568578 105930 568580
rect 106181 568578 106247 568581
rect 106641 568580 106707 568581
rect 106590 568578 106596 568580
rect 105924 568576 106247 568578
rect 105924 568520 106186 568576
rect 106242 568520 106247 568576
rect 105924 568518 106247 568520
rect 106550 568518 106596 568578
rect 106660 568576 106707 568580
rect 106702 568520 106707 568576
rect 105924 568516 105930 568518
rect 105261 568515 105327 568516
rect 106181 568515 106247 568518
rect 106590 568516 106596 568518
rect 106660 568516 106707 568520
rect 106774 568516 106780 568580
rect 106844 568578 106850 568580
rect 107561 568578 107627 568581
rect 107745 568580 107811 568581
rect 106844 568576 107627 568578
rect 106844 568520 107566 568576
rect 107622 568520 107627 568576
rect 106844 568518 107627 568520
rect 106844 568516 106850 568518
rect 106641 568515 106707 568516
rect 107561 568515 107627 568518
rect 107694 568516 107700 568580
rect 107764 568578 107811 568580
rect 107764 568576 107856 568578
rect 107806 568520 107856 568576
rect 107764 568518 107856 568520
rect 107764 568516 107811 568518
rect 108614 568516 108620 568580
rect 108684 568578 108690 568580
rect 108941 568578 109007 568581
rect 108684 568576 109007 568578
rect 108684 568520 108946 568576
rect 109002 568520 109007 568576
rect 108684 568518 109007 568520
rect 108684 568516 108690 568518
rect 107745 568515 107811 568516
rect 108941 568515 109007 568518
rect 109718 568516 109724 568580
rect 109788 568578 109794 568580
rect 110321 568578 110387 568581
rect 109788 568576 110387 568578
rect 109788 568520 110326 568576
rect 110382 568520 110387 568576
rect 109788 568518 110387 568520
rect 109788 568516 109794 568518
rect 110321 568515 110387 568518
rect 110689 568578 110755 568581
rect 110822 568578 110828 568580
rect 110689 568576 110828 568578
rect 110689 568520 110694 568576
rect 110750 568520 110828 568576
rect 110689 568518 110828 568520
rect 110689 568515 110755 568518
rect 110822 568516 110828 568518
rect 110892 568516 110898 568580
rect 111558 568516 111564 568580
rect 111628 568578 111634 568580
rect 111701 568578 111767 568581
rect 115841 568580 115907 568581
rect 115790 568578 115796 568580
rect 111628 568576 111767 568578
rect 111628 568520 111706 568576
rect 111762 568520 111767 568576
rect 111628 568518 111767 568520
rect 115750 568518 115796 568578
rect 115860 568576 115907 568580
rect 115902 568520 115907 568576
rect 111628 568516 111634 568518
rect 111701 568515 111767 568518
rect 115790 568516 115796 568518
rect 115860 568516 115907 568520
rect 126462 568516 126468 568580
rect 126532 568578 126538 568580
rect 126605 568578 126671 568581
rect 126532 568576 126671 568578
rect 126532 568520 126610 568576
rect 126666 568520 126671 568576
rect 126532 568518 126671 568520
rect 126532 568516 126538 568518
rect 115841 568515 115907 568516
rect 126605 568515 126671 568518
rect 128445 568580 128511 568581
rect 128445 568576 128492 568580
rect 128556 568578 128562 568580
rect 195973 568578 196039 568581
rect 196198 568578 196204 568580
rect 128445 568520 128450 568576
rect 128445 568516 128492 568520
rect 128556 568518 128602 568578
rect 195973 568576 196204 568578
rect 195973 568520 195978 568576
rect 196034 568520 196204 568576
rect 195973 568518 196204 568520
rect 128556 568516 128562 568518
rect 128445 568515 128511 568516
rect 195973 568515 196039 568518
rect 196198 568516 196204 568518
rect 196268 568516 196274 568580
rect 197445 568578 197511 568581
rect 202229 568580 202295 568581
rect 197670 568578 197676 568580
rect 197445 568576 197676 568578
rect 197445 568520 197450 568576
rect 197506 568520 197676 568576
rect 197445 568518 197676 568520
rect 197445 568515 197511 568518
rect 197670 568516 197676 568518
rect 197740 568516 197746 568580
rect 202229 568576 202276 568580
rect 202340 568578 202346 568580
rect 202229 568520 202234 568576
rect 202229 568516 202276 568520
rect 202340 568518 202386 568578
rect 202340 568516 202346 568518
rect 203926 568516 203932 568580
rect 203996 568578 204002 568580
rect 204161 568578 204227 568581
rect 203996 568576 204227 568578
rect 203996 568520 204166 568576
rect 204222 568520 204227 568576
rect 203996 568518 204227 568520
rect 203996 568516 204002 568518
rect 202229 568515 202295 568516
rect 204161 568515 204227 568518
rect 204805 568580 204871 568581
rect 204805 568576 204852 568580
rect 204916 568578 204922 568580
rect 204805 568520 204810 568576
rect 204805 568516 204852 568520
rect 204916 568518 204962 568578
rect 204916 568516 204922 568518
rect 205398 568516 205404 568580
rect 205468 568578 205474 568580
rect 205541 568578 205607 568581
rect 205468 568576 205607 568578
rect 205468 568520 205546 568576
rect 205602 568520 205607 568576
rect 205468 568518 205607 568520
rect 205468 568516 205474 568518
rect 204805 568515 204871 568516
rect 205541 568515 205607 568518
rect 207013 568580 207079 568581
rect 207013 568576 207060 568580
rect 207124 568578 207130 568580
rect 207013 568520 207018 568576
rect 207013 568516 207060 568520
rect 207124 568518 207170 568578
rect 207124 568516 207130 568518
rect 209446 568516 209452 568580
rect 209516 568578 209522 568580
rect 209589 568578 209655 568581
rect 211889 568580 211955 568581
rect 211838 568578 211844 568580
rect 209516 568576 209655 568578
rect 209516 568520 209594 568576
rect 209650 568520 209655 568576
rect 209516 568518 209655 568520
rect 211798 568518 211844 568578
rect 211908 568576 211955 568580
rect 211950 568520 211955 568576
rect 209516 568516 209522 568518
rect 207013 568515 207079 568516
rect 209589 568515 209655 568518
rect 211838 568516 211844 568518
rect 211908 568516 211955 568520
rect 211889 568515 211955 568516
rect 213085 568580 213151 568581
rect 214097 568580 214163 568581
rect 215569 568580 215635 568581
rect 213085 568576 213132 568580
rect 213196 568578 213202 568580
rect 214046 568578 214052 568580
rect 213085 568520 213090 568576
rect 213085 568516 213132 568520
rect 213196 568518 213242 568578
rect 214006 568518 214052 568578
rect 214116 568576 214163 568580
rect 215518 568578 215524 568580
rect 214158 568520 214163 568576
rect 213196 568516 213202 568518
rect 214046 568516 214052 568518
rect 214116 568516 214163 568520
rect 215478 568518 215524 568578
rect 215588 568576 215635 568580
rect 215630 568520 215635 568576
rect 215518 568516 215524 568518
rect 215588 568516 215635 568520
rect 216622 568516 216628 568580
rect 216692 568578 216698 568580
rect 217133 568578 217199 568581
rect 216692 568576 217199 568578
rect 216692 568520 217138 568576
rect 217194 568520 217199 568576
rect 216692 568518 217199 568520
rect 216692 568516 216698 568518
rect 213085 568515 213151 568516
rect 214097 568515 214163 568516
rect 215569 568515 215635 568516
rect 217133 568515 217199 568518
rect 218830 568516 218836 568580
rect 218900 568578 218906 568580
rect 218973 568578 219039 568581
rect 221457 568580 221523 568581
rect 222377 568580 222443 568581
rect 223665 568580 223731 568581
rect 225873 568580 225939 568581
rect 226241 568580 226307 568581
rect 227161 568580 227227 568581
rect 221406 568578 221412 568580
rect 218900 568576 219039 568578
rect 218900 568520 218978 568576
rect 219034 568520 219039 568576
rect 218900 568518 219039 568520
rect 221366 568518 221412 568578
rect 221476 568576 221523 568580
rect 222326 568578 222332 568580
rect 221518 568520 221523 568576
rect 218900 568516 218906 568518
rect 218973 568515 219039 568518
rect 221406 568516 221412 568518
rect 221476 568516 221523 568520
rect 222286 568518 222332 568578
rect 222396 568576 222443 568580
rect 223614 568578 223620 568580
rect 222438 568520 222443 568576
rect 222326 568516 222332 568518
rect 222396 568516 222443 568520
rect 223574 568518 223620 568578
rect 223684 568576 223731 568580
rect 225822 568578 225828 568580
rect 223726 568520 223731 568576
rect 223614 568516 223620 568518
rect 223684 568516 223731 568520
rect 225782 568518 225828 568578
rect 225892 568576 225939 568580
rect 225934 568520 225939 568576
rect 225822 568516 225828 568518
rect 225892 568516 225939 568520
rect 226190 568516 226196 568580
rect 226260 568578 226307 568580
rect 227110 568578 227116 568580
rect 226260 568576 226352 568578
rect 226302 568520 226352 568576
rect 226260 568518 226352 568520
rect 227070 568518 227116 568578
rect 227180 568576 227227 568580
rect 227222 568520 227227 568576
rect 226260 568516 226307 568518
rect 227110 568516 227116 568518
rect 227180 568516 227227 568520
rect 227294 568516 227300 568580
rect 227364 568578 227370 568580
rect 227621 568578 227687 568581
rect 227364 568576 227687 568578
rect 227364 568520 227626 568576
rect 227682 568520 227687 568576
rect 227364 568518 227687 568520
rect 227364 568516 227370 568518
rect 221457 568515 221523 568516
rect 222377 568515 222443 568516
rect 223665 568515 223731 568516
rect 225873 568515 225939 568516
rect 226241 568515 226307 568516
rect 227161 568515 227227 568516
rect 227621 568515 227687 568518
rect 228357 568580 228423 568581
rect 228357 568576 228404 568580
rect 228468 568578 228474 568580
rect 228357 568520 228362 568576
rect 228357 568516 228404 568520
rect 228468 568518 228514 568578
rect 228468 568516 228474 568518
rect 228766 568516 228772 568580
rect 228836 568578 228842 568580
rect 229001 568578 229067 568581
rect 229369 568580 229435 568581
rect 229318 568578 229324 568580
rect 228836 568576 229067 568578
rect 228836 568520 229006 568576
rect 229062 568520 229067 568576
rect 228836 568518 229067 568520
rect 229278 568518 229324 568578
rect 229388 568576 229435 568580
rect 229430 568520 229435 568576
rect 228836 568516 228842 568518
rect 228357 568515 228423 568516
rect 229001 568515 229067 568518
rect 229318 568516 229324 568518
rect 229388 568516 229435 568520
rect 230238 568516 230244 568580
rect 230308 568578 230314 568580
rect 230381 568578 230447 568581
rect 230308 568576 230447 568578
rect 230308 568520 230386 568576
rect 230442 568520 230447 568576
rect 230308 568518 230447 568520
rect 230308 568516 230314 568518
rect 229369 568515 229435 568516
rect 230381 568515 230447 568518
rect 230790 568516 230796 568580
rect 230860 568578 230866 568580
rect 231761 568578 231827 568581
rect 233049 568580 233115 568581
rect 234521 568580 234587 568581
rect 230860 568576 231827 568578
rect 230860 568520 231766 568576
rect 231822 568520 231827 568576
rect 230860 568518 231827 568520
rect 230860 568516 230866 568518
rect 231761 568515 231827 568518
rect 232998 568516 233004 568580
rect 233068 568578 233115 568580
rect 233068 568576 233160 568578
rect 233110 568520 233160 568576
rect 233068 568518 233160 568520
rect 233068 568516 233115 568518
rect 234470 568516 234476 568580
rect 234540 568578 234587 568580
rect 234540 568576 234632 568578
rect 234582 568520 234632 568576
rect 234540 568518 234632 568520
rect 234540 568516 234587 568518
rect 235758 568516 235764 568580
rect 235828 568578 235834 568580
rect 235901 568578 235967 568581
rect 237281 568580 237347 568581
rect 235828 568576 235967 568578
rect 235828 568520 235906 568576
rect 235962 568520 235967 568576
rect 235828 568518 235967 568520
rect 235828 568516 235834 568518
rect 233049 568515 233115 568516
rect 234521 568515 234587 568516
rect 235901 568515 235967 568518
rect 237230 568516 237236 568580
rect 237300 568578 237347 568580
rect 237300 568576 237392 568578
rect 237342 568520 237392 568576
rect 237300 568518 237392 568520
rect 237300 568516 237347 568518
rect 238150 568516 238156 568580
rect 238220 568578 238226 568580
rect 238661 568578 238727 568581
rect 238220 568576 238727 568578
rect 238220 568520 238666 568576
rect 238722 568520 238727 568576
rect 238220 568518 238727 568520
rect 238220 568516 238226 568518
rect 237281 568515 237347 568516
rect 238661 568515 238727 568518
rect 239622 568516 239628 568580
rect 239692 568578 239698 568580
rect 240041 568578 240107 568581
rect 239692 568576 240107 568578
rect 239692 568520 240046 568576
rect 240102 568520 240107 568576
rect 239692 568518 240107 568520
rect 239692 568516 239698 568518
rect 240041 568515 240107 568518
rect 95141 568444 95207 568445
rect 109861 568444 109927 568445
rect 194409 568444 194475 568445
rect 95141 568442 95188 568444
rect 95096 568440 95188 568442
rect 95096 568384 95146 568440
rect 95096 568382 95188 568384
rect 95141 568380 95188 568382
rect 95252 568380 95258 568444
rect 109861 568440 109908 568444
rect 109972 568442 109978 568444
rect 194358 568442 194364 568444
rect 109861 568384 109866 568440
rect 109861 568380 109908 568384
rect 109972 568382 110018 568442
rect 194318 568382 194364 568442
rect 194428 568440 194475 568444
rect 194470 568384 194475 568440
rect 109972 568380 109978 568382
rect 194358 568380 194364 568382
rect 194428 568380 194475 568384
rect 95141 568379 95207 568380
rect 109861 568379 109927 568380
rect 194409 568379 194475 568380
rect 203701 568444 203767 568445
rect 220077 568444 220143 568445
rect 203701 568440 203748 568444
rect 203812 568442 203818 568444
rect 203701 568384 203706 568440
rect 203701 568380 203748 568384
rect 203812 568382 203858 568442
rect 220077 568440 220124 568444
rect 220188 568442 220194 568444
rect 220077 568384 220082 568440
rect 203812 568380 203818 568382
rect 220077 568380 220124 568384
rect 220188 568382 220234 568442
rect 220188 568380 220194 568382
rect 225638 568380 225644 568444
rect 225708 568442 225714 568444
rect 226149 568442 226215 568445
rect 225708 568440 226215 568442
rect 225708 568384 226154 568440
rect 226210 568384 226215 568440
rect 225708 568382 226215 568384
rect 225708 568380 225714 568382
rect 203701 568379 203767 568380
rect 220077 568379 220143 568380
rect 226149 568379 226215 568382
rect 232630 568380 232636 568444
rect 232700 568442 232706 568444
rect 233141 568442 233207 568445
rect 234613 568444 234679 568445
rect 234613 568442 234660 568444
rect 232700 568440 233207 568442
rect 232700 568384 233146 568440
rect 233202 568384 233207 568440
rect 232700 568382 233207 568384
rect 234568 568440 234660 568442
rect 234568 568384 234618 568440
rect 234568 568382 234660 568384
rect 232700 568380 232706 568382
rect 233141 568379 233207 568382
rect 234613 568380 234660 568382
rect 234724 568380 234730 568444
rect 234613 568379 234679 568380
rect 92606 568244 92612 568308
rect 92676 568306 92682 568308
rect 93761 568306 93827 568309
rect 92676 568304 93827 568306
rect 92676 568248 93766 568304
rect 93822 568248 93827 568304
rect 92676 568246 93827 568248
rect 92676 568244 92682 568246
rect 93761 568243 93827 568246
rect 96102 568244 96108 568308
rect 96172 568306 96178 568308
rect 96521 568306 96587 568309
rect 96172 568304 96587 568306
rect 96172 568248 96526 568304
rect 96582 568248 96587 568304
rect 96172 568246 96587 568248
rect 96172 568244 96178 568246
rect 96521 568243 96587 568246
rect 97390 568244 97396 568308
rect 97460 568306 97466 568308
rect 97901 568306 97967 568309
rect 97460 568304 97967 568306
rect 97460 568248 97906 568304
rect 97962 568248 97967 568304
rect 97460 568246 97967 568248
rect 97460 568244 97466 568246
rect 97901 568243 97967 568246
rect 99598 568244 99604 568308
rect 99668 568306 99674 568308
rect 100661 568306 100727 568309
rect 99668 568304 100727 568306
rect 99668 568248 100666 568304
rect 100722 568248 100727 568304
rect 99668 568246 100727 568248
rect 99668 568244 99674 568246
rect 100661 568243 100727 568246
rect 100886 568244 100892 568308
rect 100956 568306 100962 568308
rect 102041 568306 102107 568309
rect 100956 568304 102107 568306
rect 100956 568248 102046 568304
rect 102102 568248 102107 568304
rect 100956 568246 102107 568248
rect 100956 568244 100962 568246
rect 102041 568243 102107 568246
rect 123702 568244 123708 568308
rect 123772 568306 123778 568308
rect 124121 568306 124187 568309
rect 124305 568308 124371 568309
rect 123772 568304 124187 568306
rect 123772 568248 124126 568304
rect 124182 568248 124187 568304
rect 123772 568246 124187 568248
rect 123772 568244 123778 568246
rect 124121 568243 124187 568246
rect 124254 568244 124260 568308
rect 124324 568306 124371 568308
rect 124324 568304 124416 568306
rect 124366 568248 124416 568304
rect 124324 568246 124416 568248
rect 124324 568244 124371 568246
rect 125358 568244 125364 568308
rect 125428 568306 125434 568308
rect 125501 568306 125567 568309
rect 125428 568304 125567 568306
rect 125428 568248 125506 568304
rect 125562 568248 125567 568304
rect 125428 568246 125567 568248
rect 125428 568244 125434 568246
rect 124305 568243 124371 568244
rect 125501 568243 125567 568246
rect 129590 568244 129596 568308
rect 129660 568306 129666 568308
rect 145557 568306 145623 568309
rect 224769 568308 224835 568309
rect 129660 568304 145623 568306
rect 129660 568248 145562 568304
rect 145618 568248 145623 568304
rect 129660 568246 145623 568248
rect 129660 568244 129666 568246
rect 145557 568243 145623 568246
rect 224718 568244 224724 568308
rect 224788 568306 224835 568308
rect 233233 568306 233299 568309
rect 237373 568308 237439 568309
rect 233550 568306 233556 568308
rect 224788 568304 224880 568306
rect 224830 568248 224880 568304
rect 224788 568246 224880 568248
rect 233233 568304 233556 568306
rect 233233 568248 233238 568304
rect 233294 568248 233556 568304
rect 233233 568246 233556 568248
rect 224788 568244 224835 568246
rect 224769 568243 224835 568244
rect 233233 568243 233299 568246
rect 233550 568244 233556 568246
rect 233620 568244 233626 568308
rect 237373 568306 237420 568308
rect 237328 568304 237420 568306
rect 237328 568248 237378 568304
rect 237328 568246 237420 568248
rect 237373 568244 237420 568246
rect 237484 568244 237490 568308
rect 237373 568243 237439 568244
rect 75821 568170 75887 568173
rect 200246 568170 200252 568172
rect 75821 568168 200252 568170
rect 75821 568112 75826 568168
rect 75882 568112 200252 568168
rect 75821 568110 200252 568112
rect 75821 568107 75887 568110
rect 200246 568108 200252 568110
rect 200316 568108 200322 568172
rect 230473 568170 230539 568173
rect 230606 568170 230612 568172
rect 230473 568168 230612 568170
rect 230473 568112 230478 568168
rect 230534 568112 230612 568168
rect 230473 568110 230612 568112
rect 230473 568107 230539 568110
rect 230606 568108 230612 568110
rect 230676 568108 230682 568172
rect 231945 568170 232011 568173
rect 232814 568170 232820 568172
rect 231945 568168 232820 568170
rect 231945 568112 231950 568168
rect 232006 568112 232820 568168
rect 231945 568110 232820 568112
rect 231945 568107 232011 568110
rect 232814 568108 232820 568110
rect 232884 568108 232890 568172
rect 235993 568170 236059 568173
rect 236126 568170 236132 568172
rect 235993 568168 236132 568170
rect 235993 568112 235998 568168
rect 236054 568112 236132 568168
rect 235993 568110 236132 568112
rect 235993 568107 236059 568110
rect 236126 568108 236132 568110
rect 236196 568108 236202 568172
rect 77201 568034 77267 568037
rect 231853 568036 231919 568037
rect 201534 568034 201540 568036
rect 77201 568032 201540 568034
rect 77201 567976 77206 568032
rect 77262 567976 201540 568032
rect 77201 567974 201540 567976
rect 77201 567971 77267 567974
rect 201534 567972 201540 567974
rect 201604 567972 201610 568036
rect 231853 568034 231900 568036
rect 231808 568032 231900 568034
rect 231808 567976 231858 568032
rect 231808 567974 231900 567976
rect 231853 567972 231900 567974
rect 231964 567972 231970 568036
rect 231853 567971 231919 567972
rect 73061 567898 73127 567901
rect 199510 567898 199516 567900
rect 73061 567896 199516 567898
rect 73061 567840 73066 567896
rect 73122 567840 199516 567896
rect 73061 567838 199516 567840
rect 73061 567835 73127 567838
rect 199510 567836 199516 567838
rect 199580 567836 199586 567900
rect 91093 567762 91159 567765
rect 91502 567762 91508 567764
rect 91093 567760 91508 567762
rect 91093 567704 91098 567760
rect 91154 567704 91508 567760
rect 91093 567702 91508 567704
rect 91093 567699 91159 567702
rect 91502 567700 91508 567702
rect 91572 567700 91578 567764
rect 97758 567700 97764 567764
rect 97828 567762 97834 567764
rect 97901 567762 97967 567765
rect 97828 567760 97967 567762
rect 97828 567704 97906 567760
rect 97962 567704 97967 567760
rect 97828 567702 97967 567704
rect 97828 567700 97834 567702
rect 97901 567699 97967 567702
rect 100334 567700 100340 567764
rect 100404 567762 100410 567764
rect 100661 567762 100727 567765
rect 110321 567764 110387 567765
rect 100404 567760 100727 567762
rect 100404 567704 100666 567760
rect 100722 567704 100727 567760
rect 100404 567702 100727 567704
rect 100404 567700 100410 567702
rect 100661 567699 100727 567702
rect 110270 567700 110276 567764
rect 110340 567762 110387 567764
rect 124857 567762 124923 567765
rect 124990 567762 124996 567764
rect 110340 567760 110432 567762
rect 110382 567704 110432 567760
rect 110340 567702 110432 567704
rect 124857 567760 124996 567762
rect 124857 567704 124862 567760
rect 124918 567704 124996 567760
rect 124857 567702 124996 567704
rect 110340 567700 110387 567702
rect 110321 567699 110387 567700
rect 124857 567699 124923 567702
rect 124990 567700 124996 567702
rect 125060 567700 125066 567764
rect 83406 567564 83412 567628
rect 83476 567626 83482 567628
rect 194409 567626 194475 567629
rect 83476 567624 194475 567626
rect 83476 567568 194414 567624
rect 194470 567568 194475 567624
rect 83476 567566 194475 567568
rect 83476 567564 83482 567566
rect 194409 567563 194475 567566
rect 88333 567490 88399 567493
rect 88558 567490 88564 567492
rect 88333 567488 88564 567490
rect -960 567204 480 567444
rect 88333 567432 88338 567488
rect 88394 567432 88564 567488
rect 88333 567430 88564 567432
rect 88333 567427 88399 567430
rect 88558 567428 88564 567430
rect 88628 567428 88634 567492
rect 86953 567354 87019 567357
rect 89989 567356 90055 567357
rect 87454 567354 87460 567356
rect 86953 567352 87460 567354
rect 86953 567296 86958 567352
rect 87014 567296 87460 567352
rect 86953 567294 87460 567296
rect 86953 567291 87019 567294
rect 87454 567292 87460 567294
rect 87524 567292 87530 567356
rect 89989 567354 90036 567356
rect 89944 567352 90036 567354
rect 89944 567296 89994 567352
rect 89944 567294 90036 567296
rect 89989 567292 90036 567294
rect 90100 567292 90106 567356
rect 120625 567354 120691 567357
rect 121494 567354 121500 567356
rect 120625 567352 121500 567354
rect 120625 567296 120630 567352
rect 120686 567296 121500 567352
rect 120625 567294 121500 567296
rect 89989 567291 90055 567292
rect 120625 567291 120691 567294
rect 121494 567292 121500 567294
rect 121564 567292 121570 567356
rect 124254 567292 124260 567356
rect 124324 567354 124330 567356
rect 125041 567354 125107 567357
rect 124324 567352 125107 567354
rect 124324 567296 125046 567352
rect 125102 567296 125107 567352
rect 124324 567294 125107 567296
rect 124324 567292 124330 567294
rect 125041 567291 125107 567294
rect 208342 567292 208348 567356
rect 208412 567354 208418 567356
rect 209037 567354 209103 567357
rect 208412 567352 209103 567354
rect 208412 567296 209042 567352
rect 209098 567296 209103 567352
rect 208412 567294 209103 567296
rect 208412 567292 208418 567294
rect 209037 567291 209103 567294
rect 210366 567292 210372 567356
rect 210436 567354 210442 567356
rect 211061 567354 211127 567357
rect 210436 567352 211127 567354
rect 210436 567296 211066 567352
rect 211122 567296 211127 567352
rect 210436 567294 211127 567296
rect 210436 567292 210442 567294
rect 211061 567291 211127 567294
rect 217542 567292 217548 567356
rect 217612 567354 217618 567356
rect 217961 567354 218027 567357
rect 217612 567352 218027 567354
rect 217612 567296 217966 567352
rect 218022 567296 218027 567352
rect 217612 567294 218027 567296
rect 217612 567292 217618 567294
rect 217961 567291 218027 567294
rect 93342 567156 93348 567220
rect 93412 567218 93418 567220
rect 93669 567218 93735 567221
rect 93412 567216 93735 567218
rect 93412 567160 93674 567216
rect 93730 567160 93735 567216
rect 93412 567158 93735 567160
rect 93412 567156 93418 567158
rect 93669 567155 93735 567158
rect 94262 567156 94268 567220
rect 94332 567218 94338 567220
rect 95049 567218 95115 567221
rect 94332 567216 95115 567218
rect 94332 567160 95054 567216
rect 95110 567160 95115 567216
rect 94332 567158 95115 567160
rect 94332 567156 94338 567158
rect 95049 567155 95115 567158
rect 96286 567156 96292 567220
rect 96356 567218 96362 567220
rect 96429 567218 96495 567221
rect 96356 567216 96495 567218
rect 96356 567160 96434 567216
rect 96490 567160 96495 567216
rect 96356 567158 96495 567160
rect 96356 567156 96362 567158
rect 96429 567155 96495 567158
rect 98862 567156 98868 567220
rect 98932 567218 98938 567220
rect 99189 567218 99255 567221
rect 98932 567216 99255 567218
rect 98932 567160 99194 567216
rect 99250 567160 99255 567216
rect 98932 567158 99255 567160
rect 98932 567156 98938 567158
rect 99189 567155 99255 567158
rect 122966 567156 122972 567220
rect 123036 567218 123042 567220
rect 123477 567218 123543 567221
rect 123036 567216 123543 567218
rect 123036 567160 123482 567216
rect 123538 567160 123543 567216
rect 123036 567158 123543 567160
rect 123036 567156 123042 567158
rect 123477 567155 123543 567158
rect 124806 567156 124812 567220
rect 124876 567218 124882 567220
rect 125317 567218 125383 567221
rect 124876 567216 125383 567218
rect 124876 567160 125322 567216
rect 125378 567160 125383 567216
rect 124876 567158 125383 567160
rect 124876 567156 124882 567158
rect 125317 567155 125383 567158
rect 126646 567156 126652 567220
rect 126716 567218 126722 567220
rect 126881 567218 126947 567221
rect 126716 567216 126947 567218
rect 126716 567160 126886 567216
rect 126942 567160 126947 567216
rect 126716 567158 126947 567160
rect 126716 567156 126722 567158
rect 126881 567155 126947 567158
rect 127617 567218 127683 567221
rect 128169 567220 128235 567221
rect 127750 567218 127756 567220
rect 127617 567216 127756 567218
rect 127617 567160 127622 567216
rect 127678 567160 127756 567216
rect 127617 567158 127756 567160
rect 127617 567155 127683 567158
rect 127750 567156 127756 567158
rect 127820 567156 127826 567220
rect 128118 567156 128124 567220
rect 128188 567218 128235 567220
rect 128188 567216 128280 567218
rect 128230 567160 128280 567216
rect 128188 567158 128280 567160
rect 128188 567156 128235 567158
rect 205766 567156 205772 567220
rect 205836 567218 205842 567220
rect 206277 567218 206343 567221
rect 206921 567220 206987 567221
rect 205836 567216 206343 567218
rect 205836 567160 206282 567216
rect 206338 567160 206343 567216
rect 205836 567158 206343 567160
rect 205836 567156 205842 567158
rect 128169 567155 128235 567156
rect 206277 567155 206343 567158
rect 206870 567156 206876 567220
rect 206940 567218 206987 567220
rect 206940 567216 207032 567218
rect 206982 567160 207032 567216
rect 206940 567158 207032 567160
rect 206940 567156 206987 567158
rect 207974 567156 207980 567220
rect 208044 567218 208050 567220
rect 208301 567218 208367 567221
rect 208044 567216 208367 567218
rect 208044 567160 208306 567216
rect 208362 567160 208367 567216
rect 208044 567158 208367 567160
rect 208044 567156 208050 567158
rect 206921 567155 206987 567156
rect 208301 567155 208367 567158
rect 209262 567156 209268 567220
rect 209332 567218 209338 567220
rect 209681 567218 209747 567221
rect 209332 567216 209747 567218
rect 209332 567160 209686 567216
rect 209742 567160 209747 567216
rect 209332 567158 209747 567160
rect 209332 567156 209338 567158
rect 209681 567155 209747 567158
rect 210417 567218 210483 567221
rect 210969 567220 211035 567221
rect 212441 567220 212507 567221
rect 210550 567218 210556 567220
rect 210417 567216 210556 567218
rect 210417 567160 210422 567216
rect 210478 567160 210556 567216
rect 210417 567158 210556 567160
rect 210417 567155 210483 567158
rect 210550 567156 210556 567158
rect 210620 567156 210626 567220
rect 210918 567156 210924 567220
rect 210988 567218 211035 567220
rect 210988 567216 211080 567218
rect 211030 567160 211080 567216
rect 210988 567158 211080 567160
rect 210988 567156 211035 567158
rect 212390 567156 212396 567220
rect 212460 567218 212507 567220
rect 212460 567216 212552 567218
rect 212502 567160 212552 567216
rect 212460 567158 212552 567160
rect 212460 567156 212507 567158
rect 213494 567156 213500 567220
rect 213564 567218 213570 567220
rect 213821 567218 213887 567221
rect 213564 567216 213887 567218
rect 213564 567160 213826 567216
rect 213882 567160 213887 567216
rect 213564 567158 213887 567160
rect 213564 567156 213570 567158
rect 210969 567155 211035 567156
rect 212441 567155 212507 567156
rect 213821 567155 213887 567158
rect 214782 567156 214788 567220
rect 214852 567218 214858 567220
rect 215201 567218 215267 567221
rect 214852 567216 215267 567218
rect 214852 567160 215206 567216
rect 215262 567160 215267 567216
rect 214852 567158 215267 567160
rect 214852 567156 214858 567158
rect 215201 567155 215267 567158
rect 216254 567156 216260 567220
rect 216324 567218 216330 567220
rect 216581 567218 216647 567221
rect 217869 567220 217935 567221
rect 217869 567218 217916 567220
rect 216324 567216 216647 567218
rect 216324 567160 216586 567216
rect 216642 567160 216647 567216
rect 216324 567158 216647 567160
rect 217824 567216 217916 567218
rect 217824 567160 217874 567216
rect 217824 567158 217916 567160
rect 216324 567156 216330 567158
rect 216581 567155 216647 567158
rect 217869 567156 217916 567158
rect 217980 567156 217986 567220
rect 219198 567156 219204 567220
rect 219268 567218 219274 567220
rect 219341 567218 219407 567221
rect 219268 567216 219407 567218
rect 219268 567160 219346 567216
rect 219402 567160 219407 567216
rect 219268 567158 219407 567160
rect 219268 567156 219274 567158
rect 217869 567155 217935 567156
rect 219341 567155 219407 567158
rect 221958 567156 221964 567220
rect 222028 567218 222034 567220
rect 222101 567218 222167 567221
rect 222028 567216 222167 567218
rect 222028 567160 222106 567216
rect 222162 567160 222167 567216
rect 222028 567158 222167 567160
rect 222028 567156 222034 567158
rect 222101 567155 222167 567158
rect 223246 567156 223252 567220
rect 223316 567218 223322 567220
rect 223481 567218 223547 567221
rect 223316 567216 223547 567218
rect 223316 567160 223486 567216
rect 223542 567160 223547 567216
rect 223316 567158 223547 567160
rect 223316 567156 223322 567158
rect 223481 567155 223547 567158
rect 223798 567156 223804 567220
rect 223868 567218 223874 567220
rect 224861 567218 224927 567221
rect 223868 567216 224927 567218
rect 223868 567160 224866 567216
rect 224922 567160 224927 567216
rect 223868 567158 224927 567160
rect 223868 567156 223874 567158
rect 224861 567155 224927 567158
rect 117262 566476 117268 566540
rect 117332 566538 117338 566540
rect 118509 566538 118575 566541
rect 117332 566536 118575 566538
rect 117332 566480 118514 566536
rect 118570 566480 118575 566536
rect 117332 566478 118575 566480
rect 117332 566476 117338 566478
rect 118509 566475 118575 566478
rect 121494 566068 121500 566132
rect 121564 566130 121570 566132
rect 122097 566130 122163 566133
rect 121564 566128 122163 566130
rect 121564 566072 122102 566128
rect 122158 566072 122163 566128
rect 121564 566070 122163 566072
rect 121564 566068 121570 566070
rect 122097 566067 122163 566070
rect 583520 557140 584960 557380
rect -960 552924 480 553164
rect 583520 545444 584960 545684
rect -960 538508 480 538748
rect 583520 533748 584960 533988
rect -960 524092 480 524332
rect 152457 524242 152523 524245
rect 204345 524242 204411 524245
rect 152457 524240 204411 524242
rect 152457 524184 152462 524240
rect 152518 524184 204350 524240
rect 204406 524184 204411 524240
rect 152457 524182 204411 524184
rect 152457 524179 152523 524182
rect 204345 524179 204411 524182
rect 145557 524106 145623 524109
rect 210049 524106 210115 524109
rect 145557 524104 210115 524106
rect 145557 524048 145562 524104
rect 145618 524048 210054 524104
rect 210110 524048 210115 524104
rect 145557 524046 210115 524048
rect 145557 524043 145623 524046
rect 210049 524043 210115 524046
rect 125317 523970 125383 523973
rect 202413 523970 202479 523973
rect 125317 523968 202479 523970
rect 125317 523912 125322 523968
rect 125378 523912 202418 523968
rect 202474 523912 202479 523968
rect 125317 523910 202479 523912
rect 125317 523907 125383 523910
rect 202413 523907 202479 523910
rect 126881 523834 126947 523837
rect 206185 523834 206251 523837
rect 126881 523832 206251 523834
rect 126881 523776 126886 523832
rect 126942 523776 206190 523832
rect 206246 523776 206251 523832
rect 126881 523774 206251 523776
rect 126881 523771 126947 523774
rect 206185 523771 206251 523774
rect 70945 523698 71011 523701
rect 197445 523698 197511 523701
rect 70945 523696 197511 523698
rect 70945 523640 70950 523696
rect 71006 523640 197450 523696
rect 197506 523640 197511 523696
rect 70945 523638 197511 523640
rect 70945 523635 71011 523638
rect 197445 523635 197511 523638
rect 583520 521916 584960 522156
rect 273989 520978 274055 520981
rect 271860 520976 274055 520978
rect 271860 520920 273994 520976
rect 274050 520920 274055 520976
rect 271860 520918 274055 520920
rect 273989 520915 274055 520918
rect 274265 519074 274331 519077
rect 271860 519072 274331 519074
rect 271860 519016 274270 519072
rect 274326 519016 274331 519072
rect 271860 519014 274331 519016
rect 274265 519011 274331 519014
rect 337745 517442 337811 517445
rect 337745 517440 340285 517442
rect 337745 517384 337750 517440
rect 337806 517384 340285 517440
rect 337745 517382 340285 517384
rect 337745 517379 337811 517382
rect 340225 517276 340285 517382
rect 274081 517170 274147 517173
rect 271860 517168 274147 517170
rect 271860 517112 274086 517168
rect 274142 517112 274147 517168
rect 271860 517110 274147 517112
rect 274081 517107 274147 517110
rect 320173 516764 320239 516765
rect 320173 516762 320220 516764
rect 320128 516760 320220 516762
rect 320128 516704 320178 516760
rect 320128 516702 320220 516704
rect 320173 516700 320220 516702
rect 320284 516700 320290 516764
rect 398833 516762 398899 516765
rect 398833 516760 399832 516762
rect 398833 516704 398838 516760
rect 398894 516704 399832 516760
rect 398833 516702 399832 516704
rect 320173 516699 320239 516700
rect 398833 516699 398899 516702
rect 400213 516626 400279 516629
rect 401593 516626 401659 516629
rect 400213 516624 400936 516626
rect 400213 516568 400218 516624
rect 400274 516568 400936 516624
rect 400213 516566 400936 516568
rect 401593 516624 402631 516626
rect 401593 516568 401598 516624
rect 401654 516568 402631 516624
rect 401593 516566 402631 516568
rect 400213 516563 400279 516566
rect 401593 516563 401659 516566
rect 273846 516428 273852 516492
rect 273916 516490 273922 516492
rect 338389 516490 338455 516493
rect 273916 516488 338455 516490
rect 273916 516432 338394 516488
rect 338450 516432 338455 516488
rect 273916 516430 338455 516432
rect 273916 516428 273922 516430
rect 338389 516427 338455 516430
rect 340873 516490 340939 516493
rect 403341 516490 403407 516493
rect 404353 516490 404419 516493
rect 406009 516490 406075 516493
rect 340873 516488 398084 516490
rect 340873 516432 340878 516488
rect 340934 516432 398084 516488
rect 340873 516430 398084 516432
rect 403341 516488 403788 516490
rect 403341 516432 403346 516488
rect 403402 516432 403788 516488
rect 403341 516430 403788 516432
rect 404353 516488 405444 516490
rect 404353 516432 404358 516488
rect 404414 516432 405444 516488
rect 404353 516430 405444 516432
rect 406009 516488 406587 516490
rect 406009 516432 406014 516488
rect 406070 516432 406587 516488
rect 406009 516430 406587 516432
rect 340873 516427 340939 516430
rect 403341 516427 403407 516430
rect 404353 516427 404419 516430
rect 406009 516427 406075 516430
rect 273621 515266 273687 515269
rect 271860 515264 273687 515266
rect 271860 515208 273626 515264
rect 273682 515208 273687 515264
rect 271860 515206 273687 515208
rect 273621 515203 273687 515206
rect 274173 513362 274239 513365
rect 271860 513360 274239 513362
rect 271860 513304 274178 513360
rect 274234 513304 274239 513360
rect 271860 513302 274239 513304
rect 274173 513299 274239 513302
rect 320173 512140 320239 512141
rect 320173 512138 320220 512140
rect 320128 512136 320220 512138
rect 320128 512080 320178 512136
rect 320128 512078 320220 512080
rect 320173 512076 320220 512078
rect 320284 512076 320290 512140
rect 320173 512075 320239 512076
rect 273529 511458 273595 511461
rect 271860 511456 273595 511458
rect 271860 511400 273534 511456
rect 273590 511400 273595 511456
rect 271860 511398 273595 511400
rect 273529 511395 273595 511398
rect 583520 510220 584960 510460
rect -960 509812 480 510052
rect 274265 509554 274331 509557
rect 271860 509552 274331 509554
rect 271860 509496 274270 509552
rect 274326 509496 274331 509552
rect 271860 509494 274331 509496
rect 274265 509491 274331 509494
rect 316677 509146 316743 509149
rect 320030 509146 320036 509148
rect 316677 509144 320036 509146
rect 316677 509088 316682 509144
rect 316738 509088 320036 509144
rect 316677 509086 320036 509088
rect 316677 509083 316743 509086
rect 320030 509084 320036 509086
rect 320100 509084 320106 509148
rect 319437 507922 319503 507925
rect 320030 507922 320036 507924
rect 319437 507920 320036 507922
rect 319437 507864 319442 507920
rect 319498 507864 320036 507920
rect 319437 507862 320036 507864
rect 319437 507859 319503 507862
rect 320030 507860 320036 507862
rect 320100 507860 320106 507924
rect 273713 507650 273779 507653
rect 271860 507648 273779 507650
rect 271860 507592 273718 507648
rect 273774 507592 273779 507648
rect 271860 507590 273779 507592
rect 273713 507587 273779 507590
rect 320357 507516 320423 507517
rect 320357 507514 320404 507516
rect 320312 507512 320404 507514
rect 320312 507456 320362 507512
rect 320312 507454 320404 507456
rect 320357 507452 320404 507454
rect 320468 507452 320474 507516
rect 320357 507451 320423 507452
rect 319805 506292 319871 506293
rect 320173 506292 320239 506293
rect 319805 506290 319852 506292
rect 319760 506288 319852 506290
rect 319760 506232 319810 506288
rect 319760 506230 319852 506232
rect 319805 506228 319852 506230
rect 319916 506228 319922 506292
rect 320173 506290 320220 506292
rect 320128 506288 320220 506290
rect 320128 506232 320178 506288
rect 320128 506230 320220 506232
rect 320173 506228 320220 506230
rect 320284 506228 320290 506292
rect 319805 506227 319871 506228
rect 320173 506227 320239 506228
rect 273529 505746 273595 505749
rect 271860 505744 273595 505746
rect 271860 505688 273534 505744
rect 273590 505688 273595 505744
rect 271860 505686 273595 505688
rect 273529 505683 273595 505686
rect 320725 504796 320791 504797
rect 320725 504794 320772 504796
rect 320680 504792 320772 504794
rect 320680 504736 320730 504792
rect 320680 504734 320772 504736
rect 320725 504732 320772 504734
rect 320836 504732 320842 504796
rect 320725 504731 320791 504732
rect 273529 503842 273595 503845
rect 271860 503840 273595 503842
rect 271860 503784 273534 503840
rect 273590 503784 273595 503840
rect 271860 503782 273595 503784
rect 273529 503779 273595 503782
rect 276606 503780 276612 503844
rect 276676 503842 276682 503844
rect 319846 503842 319852 503844
rect 276676 503782 319852 503842
rect 276676 503780 276682 503782
rect 319846 503780 319852 503782
rect 319916 503780 319922 503844
rect 320541 503708 320607 503709
rect 320541 503706 320588 503708
rect 320496 503704 320588 503706
rect 320496 503648 320546 503704
rect 320496 503646 320588 503648
rect 320541 503644 320588 503646
rect 320652 503644 320658 503708
rect 320541 503643 320607 503644
rect 320173 503164 320239 503165
rect 320173 503162 320220 503164
rect 320128 503160 320220 503162
rect 320128 503104 320178 503160
rect 320128 503102 320220 503104
rect 320173 503100 320220 503102
rect 320284 503100 320290 503164
rect 320173 503099 320239 503100
rect 320357 502484 320423 502485
rect 320357 502482 320404 502484
rect 320312 502480 320404 502482
rect 320312 502424 320362 502480
rect 320312 502422 320404 502424
rect 320357 502420 320404 502422
rect 320468 502420 320474 502484
rect 320357 502419 320423 502420
rect 273621 501938 273687 501941
rect 271860 501936 273687 501938
rect 271860 501880 273626 501936
rect 273682 501880 273687 501936
rect 271860 501878 273687 501880
rect 273621 501875 273687 501878
rect 320817 501396 320883 501397
rect 320766 501332 320772 501396
rect 320836 501394 320883 501396
rect 320836 501392 320928 501394
rect 320878 501336 320928 501392
rect 320836 501334 320928 501336
rect 320836 501332 320883 501334
rect 320817 501331 320883 501332
rect 319805 500988 319871 500989
rect 319805 500986 319852 500988
rect 319760 500984 319852 500986
rect 319760 500928 319810 500984
rect 319760 500926 319852 500928
rect 319805 500924 319852 500926
rect 319916 500924 319922 500988
rect 319805 500923 319871 500924
rect 319989 500852 320055 500853
rect 319989 500850 320036 500852
rect 319944 500848 320036 500850
rect 319944 500792 319994 500848
rect 319944 500790 320036 500792
rect 319989 500788 320036 500790
rect 320100 500788 320106 500852
rect 319989 500787 320055 500788
rect 320633 500172 320699 500173
rect 320582 500108 320588 500172
rect 320652 500170 320699 500172
rect 320652 500168 320744 500170
rect 320694 500112 320744 500168
rect 320652 500110 320744 500112
rect 320652 500108 320699 500110
rect 320633 500107 320699 500108
rect 273713 500034 273779 500037
rect 271860 500032 273779 500034
rect 271860 499976 273718 500032
rect 273774 499976 273779 500032
rect 271860 499974 273779 499976
rect 273713 499971 273779 499974
rect 320265 499628 320331 499629
rect 320214 499564 320220 499628
rect 320284 499626 320331 499628
rect 320284 499624 320376 499626
rect 320326 499568 320376 499624
rect 320284 499566 320376 499568
rect 320284 499564 320331 499566
rect 320265 499563 320331 499564
rect 320725 498948 320791 498949
rect 320725 498946 320772 498948
rect 320680 498944 320772 498946
rect 320680 498888 320730 498944
rect 320680 498886 320772 498888
rect 320725 498884 320772 498886
rect 320836 498884 320842 498948
rect 320725 498883 320791 498884
rect 583520 498524 584960 498764
rect 273713 498130 273779 498133
rect 271860 498128 273779 498130
rect 271860 498072 273718 498128
rect 273774 498072 273779 498128
rect 271860 498070 273779 498072
rect 273713 498067 273779 498070
rect 319805 497996 319871 497997
rect 319805 497994 319852 497996
rect 319760 497992 319852 497994
rect 319760 497936 319810 497992
rect 319760 497934 319852 497936
rect 319805 497932 319852 497934
rect 319916 497932 319922 497996
rect 319805 497931 319871 497932
rect 320265 497860 320331 497861
rect 320214 497796 320220 497860
rect 320284 497858 320331 497860
rect 320284 497856 320376 497858
rect 320326 497800 320376 497856
rect 320284 497798 320376 497800
rect 320284 497796 320331 497798
rect 320265 497795 320331 497796
rect 320173 497316 320239 497317
rect 320173 497314 320220 497316
rect 320128 497312 320220 497314
rect 320128 497256 320178 497312
rect 320128 497254 320220 497256
rect 320173 497252 320220 497254
rect 320284 497252 320290 497316
rect 320173 497251 320239 497252
rect 320449 496636 320515 496637
rect 320398 496572 320404 496636
rect 320468 496634 320515 496636
rect 320468 496632 320560 496634
rect 320510 496576 320560 496632
rect 320468 496574 320560 496576
rect 320468 496572 320515 496574
rect 320449 496571 320515 496572
rect 273713 496226 273779 496229
rect 271860 496224 273779 496226
rect 271860 496168 273718 496224
rect 273774 496168 273779 496224
rect 271860 496166 273779 496168
rect 273713 496163 273779 496166
rect -960 495396 480 495636
rect 320817 495548 320883 495549
rect 320766 495546 320772 495548
rect 320726 495486 320772 495546
rect 320836 495544 320883 495548
rect 320878 495488 320883 495544
rect 320766 495484 320772 495486
rect 320836 495484 320883 495488
rect 320817 495483 320883 495484
rect 319805 495276 319871 495277
rect 319805 495274 319852 495276
rect 319760 495272 319852 495274
rect 319760 495216 319810 495272
rect 319760 495214 319852 495216
rect 319805 495212 319852 495214
rect 319916 495212 319922 495276
rect 319805 495211 319871 495212
rect 320173 495004 320239 495005
rect 320173 495002 320220 495004
rect 320128 495000 320220 495002
rect 320128 494944 320178 495000
rect 320128 494942 320220 494944
rect 320173 494940 320220 494942
rect 320284 494940 320290 495004
rect 320173 494939 320239 494940
rect 320541 494596 320607 494597
rect 320541 494592 320588 494596
rect 320652 494594 320658 494596
rect 320541 494536 320546 494592
rect 320541 494532 320588 494536
rect 320652 494534 320698 494594
rect 320652 494532 320658 494534
rect 320541 494531 320607 494532
rect 273621 494322 273687 494325
rect 271860 494320 273687 494322
rect 271860 494264 273626 494320
rect 273682 494264 273687 494320
rect 271860 494262 273687 494264
rect 273621 494259 273687 494262
rect 319805 493780 319871 493781
rect 319805 493778 319852 493780
rect 319760 493776 319852 493778
rect 319760 493720 319810 493776
rect 319760 493718 319852 493720
rect 319805 493716 319852 493718
rect 319916 493716 319922 493780
rect 319805 493715 319871 493716
rect 320357 493508 320423 493509
rect 320357 493504 320404 493508
rect 320468 493506 320474 493508
rect 320357 493448 320362 493504
rect 320357 493444 320404 493448
rect 320468 493446 320514 493506
rect 320468 493444 320474 493446
rect 320357 493443 320423 493444
rect 319989 492692 320055 492693
rect 319989 492690 320036 492692
rect 319944 492688 320036 492690
rect 319944 492632 319994 492688
rect 319944 492630 320036 492632
rect 319989 492628 320036 492630
rect 320100 492628 320106 492692
rect 319989 492627 320055 492628
rect 273621 492418 273687 492421
rect 271860 492416 273687 492418
rect 271860 492360 273626 492416
rect 273682 492360 273687 492416
rect 271860 492358 273687 492360
rect 273621 492355 273687 492358
rect 320633 492284 320699 492285
rect 320582 492282 320588 492284
rect 320542 492222 320588 492282
rect 320652 492280 320699 492284
rect 320694 492224 320699 492280
rect 320582 492220 320588 492222
rect 320652 492220 320699 492224
rect 320633 492219 320699 492220
rect 319805 491196 319871 491197
rect 319805 491194 319852 491196
rect 319760 491192 319852 491194
rect 319760 491136 319810 491192
rect 319760 491134 319852 491136
rect 319805 491132 319852 491134
rect 319916 491132 319922 491196
rect 319805 491131 319871 491132
rect 320633 490924 320699 490925
rect 320582 490922 320588 490924
rect 320542 490862 320588 490922
rect 320652 490920 320699 490924
rect 320694 490864 320699 490920
rect 320582 490860 320588 490862
rect 320652 490860 320699 490864
rect 320633 490859 320699 490860
rect 273437 490514 273503 490517
rect 271860 490512 273503 490514
rect 271860 490456 273442 490512
rect 273498 490456 273503 490512
rect 271860 490454 273503 490456
rect 273437 490451 273503 490454
rect 320173 490380 320239 490381
rect 320173 490378 320220 490380
rect 320128 490376 320220 490378
rect 320128 490320 320178 490376
rect 320128 490318 320220 490320
rect 320173 490316 320220 490318
rect 320284 490316 320290 490380
rect 320173 490315 320239 490316
rect 320081 489834 320147 489837
rect 320214 489834 320220 489836
rect 320081 489832 320220 489834
rect 320081 489776 320086 489832
rect 320142 489776 320220 489832
rect 320081 489774 320220 489776
rect 320081 489771 320147 489774
rect 320214 489772 320220 489774
rect 320284 489772 320290 489836
rect 273621 488610 273687 488613
rect 271860 488608 273687 488610
rect 271860 488552 273626 488608
rect 273682 488552 273687 488608
rect 271860 488550 273687 488552
rect 273621 488547 273687 488550
rect 320265 488474 320331 488477
rect 320725 488476 320791 488477
rect 320725 488474 320772 488476
rect 320265 488472 320772 488474
rect 320836 488474 320842 488476
rect 320265 488416 320270 488472
rect 320326 488416 320730 488472
rect 320265 488414 320772 488416
rect 320265 488411 320331 488414
rect 320725 488412 320772 488414
rect 320836 488414 320882 488474
rect 320836 488412 320842 488414
rect 320725 488411 320791 488412
rect 319805 487932 319871 487933
rect 320173 487932 320239 487933
rect 319805 487930 319852 487932
rect 319760 487928 319852 487930
rect 319760 487872 319810 487928
rect 319760 487870 319852 487872
rect 319805 487868 319852 487870
rect 319916 487868 319922 487932
rect 320173 487930 320220 487932
rect 320128 487928 320220 487930
rect 320128 487872 320178 487928
rect 320128 487870 320220 487872
rect 320173 487868 320220 487870
rect 320284 487868 320290 487932
rect 319805 487867 319871 487868
rect 320173 487867 320239 487868
rect 320265 487388 320331 487389
rect 320214 487386 320220 487388
rect 320174 487326 320220 487386
rect 320284 487386 320331 487388
rect 320449 487386 320515 487389
rect 320284 487384 320515 487386
rect 320326 487328 320454 487384
rect 320510 487328 320515 487384
rect 320214 487324 320220 487326
rect 320284 487326 320515 487328
rect 320284 487324 320331 487326
rect 320265 487323 320331 487324
rect 320449 487323 320515 487326
rect 273529 486706 273595 486709
rect 271860 486704 273595 486706
rect 271860 486648 273534 486704
rect 273590 486648 273595 486704
rect 271860 486646 273595 486648
rect 273529 486643 273595 486646
rect 319713 486706 319779 486709
rect 319846 486706 319852 486708
rect 319713 486704 319852 486706
rect 319713 486648 319718 486704
rect 319774 486648 319852 486704
rect 319713 486646 319852 486648
rect 319713 486643 319779 486646
rect 319846 486644 319852 486646
rect 319916 486644 319922 486708
rect 583520 486692 584960 486932
rect 320449 486164 320515 486165
rect 320398 486162 320404 486164
rect 320358 486102 320404 486162
rect 320468 486160 320515 486164
rect 320510 486104 320515 486160
rect 320398 486100 320404 486102
rect 320468 486100 320515 486104
rect 320449 486099 320515 486100
rect 319805 485620 319871 485621
rect 319805 485618 319852 485620
rect 319760 485616 319852 485618
rect 319760 485560 319810 485616
rect 319760 485558 319852 485560
rect 319805 485556 319852 485558
rect 319916 485556 319922 485620
rect 319805 485555 319871 485556
rect 320541 484940 320607 484941
rect 320541 484936 320588 484940
rect 320652 484938 320658 484940
rect 320541 484880 320546 484936
rect 320541 484876 320588 484880
rect 320652 484878 320698 484938
rect 320652 484876 320658 484878
rect 320541 484875 320607 484876
rect 273621 484802 273687 484805
rect 271860 484800 273687 484802
rect 271860 484744 273626 484800
rect 273682 484744 273687 484800
rect 271860 484742 273687 484744
rect 273621 484739 273687 484742
rect 320173 484532 320239 484533
rect 320173 484530 320220 484532
rect 320128 484528 320220 484530
rect 320128 484472 320178 484528
rect 320128 484470 320220 484472
rect 320173 484468 320220 484470
rect 320284 484468 320290 484532
rect 320173 484467 320239 484468
rect 320357 484124 320423 484125
rect 320357 484120 320404 484124
rect 320468 484122 320474 484124
rect 320357 484064 320362 484120
rect 320357 484060 320404 484064
rect 320468 484062 320514 484122
rect 320468 484060 320474 484062
rect 320357 484059 320423 484060
rect 319805 483036 319871 483037
rect 319805 483034 319852 483036
rect 319760 483032 319852 483034
rect 319760 482976 319810 483032
rect 319760 482974 319852 482976
rect 319805 482972 319852 482974
rect 319916 482972 319922 483036
rect 319805 482971 319871 482972
rect 273621 482898 273687 482901
rect 271860 482896 273687 482898
rect 271860 482840 273626 482896
rect 273682 482840 273687 482896
rect 271860 482838 273687 482840
rect 273621 482835 273687 482838
rect 320725 482762 320791 482765
rect 320725 482760 320834 482762
rect 320725 482704 320730 482760
rect 320786 482704 320834 482760
rect 320725 482699 320834 482704
rect 320633 482628 320699 482629
rect 320582 482626 320588 482628
rect 320542 482566 320588 482626
rect 320652 482624 320699 482628
rect 320694 482568 320699 482624
rect 320582 482564 320588 482566
rect 320652 482564 320699 482568
rect 320633 482563 320699 482564
rect 320633 482354 320699 482357
rect 320774 482354 320834 482699
rect 320633 482352 320834 482354
rect 320633 482296 320638 482352
rect 320694 482296 320834 482352
rect 320633 482294 320834 482296
rect 320633 482291 320699 482294
rect 320173 482084 320239 482085
rect 320173 482082 320220 482084
rect 320128 482080 320220 482082
rect 320128 482024 320178 482080
rect 320128 482022 320220 482024
rect 320173 482020 320220 482022
rect 320284 482020 320290 482084
rect 320173 482019 320239 482020
rect 320449 481540 320515 481541
rect 320398 481538 320404 481540
rect 320358 481478 320404 481538
rect 320468 481536 320515 481540
rect 320510 481480 320515 481536
rect 320398 481476 320404 481478
rect 320468 481476 320515 481480
rect 320449 481475 320515 481476
rect -960 480980 480 481220
rect 273621 480994 273687 480997
rect 271860 480992 273687 480994
rect 271860 480936 273626 480992
rect 273682 480936 273687 480992
rect 271860 480934 273687 480936
rect 273621 480931 273687 480934
rect 320541 480316 320607 480317
rect 320541 480312 320588 480316
rect 320652 480314 320658 480316
rect 320541 480256 320546 480312
rect 320541 480252 320588 480256
rect 320652 480254 320698 480314
rect 320652 480252 320658 480254
rect 320541 480251 320607 480252
rect 319805 479772 319871 479773
rect 320173 479772 320239 479773
rect 319805 479770 319852 479772
rect 319760 479768 319852 479770
rect 319760 479712 319810 479768
rect 319760 479710 319852 479712
rect 319805 479708 319852 479710
rect 319916 479708 319922 479772
rect 320173 479770 320220 479772
rect 320128 479768 320220 479770
rect 320128 479712 320178 479768
rect 320128 479710 320220 479712
rect 320173 479708 320220 479710
rect 320284 479708 320290 479772
rect 319805 479707 319871 479708
rect 320173 479707 320239 479708
rect 273621 479090 273687 479093
rect 320633 479092 320699 479093
rect 320582 479090 320588 479092
rect 271860 479088 273687 479090
rect 271860 479032 273626 479088
rect 273682 479032 273687 479088
rect 271860 479030 273687 479032
rect 320542 479030 320588 479090
rect 320652 479088 320699 479092
rect 320694 479032 320699 479088
rect 273621 479027 273687 479030
rect 320582 479028 320588 479030
rect 320652 479028 320699 479032
rect 320633 479027 320699 479028
rect 320633 478004 320699 478005
rect 320582 477940 320588 478004
rect 320652 478002 320699 478004
rect 320652 478000 320744 478002
rect 320694 477944 320744 478000
rect 320652 477942 320744 477944
rect 320652 477940 320699 477942
rect 320633 477939 320699 477940
rect 273621 477186 273687 477189
rect 271860 477184 273687 477186
rect 271860 477128 273626 477184
rect 273682 477128 273687 477184
rect 271860 477126 273687 477128
rect 273621 477123 273687 477126
rect 320173 476780 320239 476781
rect 320357 476780 320423 476781
rect 320173 476778 320220 476780
rect 320128 476776 320220 476778
rect 320128 476720 320178 476776
rect 320128 476718 320220 476720
rect 320173 476716 320220 476718
rect 320284 476716 320290 476780
rect 320357 476776 320404 476780
rect 320468 476778 320474 476780
rect 320357 476720 320362 476776
rect 320357 476716 320404 476720
rect 320468 476718 320514 476778
rect 320468 476716 320474 476718
rect 320173 476715 320239 476716
rect 320357 476715 320423 476716
rect 320449 475962 320515 475965
rect 320725 475962 320791 475965
rect 320449 475960 320791 475962
rect 320449 475904 320454 475960
rect 320510 475904 320730 475960
rect 320786 475904 320791 475960
rect 320449 475902 320791 475904
rect 320449 475899 320515 475902
rect 320725 475899 320791 475902
rect 319846 475764 319852 475828
rect 319916 475826 319922 475828
rect 320633 475826 320699 475829
rect 320817 475828 320883 475829
rect 319916 475824 320699 475826
rect 319916 475768 320638 475824
rect 320694 475768 320699 475824
rect 319916 475766 320699 475768
rect 319916 475764 319922 475766
rect 320633 475763 320699 475766
rect 320766 475764 320772 475828
rect 320836 475826 320883 475828
rect 320836 475824 320928 475826
rect 320878 475768 320928 475824
rect 320836 475766 320928 475768
rect 320836 475764 320883 475766
rect 320817 475763 320883 475764
rect 320582 475628 320588 475692
rect 320652 475690 320658 475692
rect 320652 475630 320834 475690
rect 320652 475628 320658 475630
rect 320774 475557 320834 475630
rect 320774 475552 320883 475557
rect 320774 475496 320822 475552
rect 320878 475496 320883 475552
rect 320774 475494 320883 475496
rect 320817 475491 320883 475494
rect 273621 475282 273687 475285
rect 271860 475280 273687 475282
rect 271860 475224 273626 475280
rect 273682 475224 273687 475280
rect 271860 475222 273687 475224
rect 273621 475219 273687 475222
rect 583520 474996 584960 475236
rect 320173 474468 320239 474469
rect 320725 474468 320791 474469
rect 320173 474466 320220 474468
rect 320128 474464 320220 474466
rect 320128 474408 320178 474464
rect 320128 474406 320220 474408
rect 320173 474404 320220 474406
rect 320284 474404 320290 474468
rect 320725 474464 320772 474468
rect 320836 474466 320842 474468
rect 320725 474408 320730 474464
rect 320725 474404 320772 474408
rect 320836 474406 320882 474466
rect 320836 474404 320842 474406
rect 320173 474403 320239 474404
rect 320725 474403 320791 474404
rect 273621 473378 273687 473381
rect 271860 473376 273687 473378
rect 271860 473320 273626 473376
rect 273682 473320 273687 473376
rect 271860 473318 273687 473320
rect 273621 473315 273687 473318
rect 320265 473378 320331 473381
rect 320265 473376 320650 473378
rect 320265 473320 320270 473376
rect 320326 473320 320650 473376
rect 320265 473318 320650 473320
rect 320265 473315 320331 473318
rect 320590 473245 320650 473318
rect 320265 473244 320331 473245
rect 320214 473180 320220 473244
rect 320284 473242 320331 473244
rect 320541 473244 320650 473245
rect 320284 473240 320376 473242
rect 320326 473184 320376 473240
rect 320284 473182 320376 473184
rect 320541 473240 320588 473244
rect 320652 473242 320658 473244
rect 320541 473184 320546 473240
rect 320284 473180 320331 473182
rect 320265 473179 320331 473180
rect 320541 473180 320588 473184
rect 320652 473182 320698 473242
rect 320652 473180 320658 473182
rect 320541 473179 320607 473180
rect 320214 472228 320220 472292
rect 320284 472290 320290 472292
rect 320357 472290 320423 472293
rect 320284 472288 320423 472290
rect 320284 472232 320362 472288
rect 320418 472232 320423 472288
rect 320284 472230 320423 472232
rect 320284 472228 320290 472230
rect 320357 472227 320423 472230
rect 320357 472156 320423 472157
rect 320357 472154 320404 472156
rect 320312 472152 320404 472154
rect 320312 472096 320362 472152
rect 320312 472094 320404 472096
rect 320357 472092 320404 472094
rect 320468 472092 320474 472156
rect 320357 472091 320423 472092
rect 273529 471474 273595 471477
rect 271860 471472 273595 471474
rect 271860 471416 273534 471472
rect 273590 471416 273595 471472
rect 271860 471414 273595 471416
rect 273529 471411 273595 471414
rect 320173 471066 320239 471069
rect 320449 471066 320515 471069
rect 320582 471066 320588 471068
rect 320173 471064 320588 471066
rect 320173 471008 320178 471064
rect 320234 471008 320454 471064
rect 320510 471008 320588 471064
rect 320173 471006 320588 471008
rect 320173 471003 320239 471006
rect 320449 471003 320515 471006
rect 320582 471004 320588 471006
rect 320652 471004 320658 471068
rect 320449 470932 320515 470933
rect 320398 470868 320404 470932
rect 320468 470930 320515 470932
rect 320468 470928 320560 470930
rect 320510 470872 320560 470928
rect 320468 470870 320560 470872
rect 320468 470868 320515 470870
rect 320449 470867 320515 470868
rect 320265 470114 320331 470117
rect 320398 470114 320404 470116
rect 320265 470112 320404 470114
rect 320265 470056 320270 470112
rect 320326 470056 320404 470112
rect 320265 470054 320404 470056
rect 320265 470051 320331 470054
rect 320398 470052 320404 470054
rect 320468 470052 320474 470116
rect 320265 469844 320331 469845
rect 320214 469780 320220 469844
rect 320284 469842 320331 469844
rect 320284 469840 320376 469842
rect 320326 469784 320376 469840
rect 320284 469782 320376 469784
rect 320284 469780 320331 469782
rect 320265 469779 320331 469780
rect 273529 469570 273595 469573
rect 271860 469568 273595 469570
rect 271860 469512 273534 469568
rect 273590 469512 273595 469568
rect 271860 469510 273595 469512
rect 273529 469507 273595 469510
rect 319846 469100 319852 469164
rect 319916 469162 319922 469164
rect 320357 469162 320423 469165
rect 319916 469160 320423 469162
rect 319916 469104 320362 469160
rect 320418 469104 320423 469160
rect 319916 469102 320423 469104
rect 319916 469100 319922 469102
rect 320357 469099 320423 469102
rect 320633 468892 320699 468893
rect 320582 468890 320588 468892
rect 320542 468830 320588 468890
rect 320652 468888 320699 468892
rect 320694 468832 320699 468888
rect 320582 468828 320588 468830
rect 320652 468828 320699 468832
rect 320633 468827 320699 468828
rect 320173 468620 320239 468621
rect 320173 468618 320220 468620
rect 320128 468616 320220 468618
rect 320128 468560 320178 468616
rect 320128 468558 320220 468560
rect 320173 468556 320220 468558
rect 320284 468556 320290 468620
rect 320173 468555 320239 468556
rect 273529 467666 273595 467669
rect 271860 467664 273595 467666
rect 271860 467608 273534 467664
rect 273590 467608 273595 467664
rect 271860 467606 273595 467608
rect 273529 467603 273595 467606
rect 320398 467604 320404 467668
rect 320468 467666 320474 467668
rect 320633 467666 320699 467669
rect 320468 467664 320699 467666
rect 320468 467608 320638 467664
rect 320694 467608 320699 467664
rect 320468 467606 320699 467608
rect 320468 467604 320474 467606
rect 320633 467603 320699 467606
rect -960 466700 480 466940
rect 273529 465762 273595 465765
rect 271860 465760 273595 465762
rect 271860 465704 273534 465760
rect 273590 465704 273595 465760
rect 271860 465702 273595 465704
rect 273529 465699 273595 465702
rect 320173 465220 320239 465221
rect 320173 465218 320220 465220
rect 320128 465216 320220 465218
rect 320128 465160 320178 465216
rect 320128 465158 320220 465160
rect 320173 465156 320220 465158
rect 320284 465156 320290 465220
rect 320398 465156 320404 465220
rect 320468 465156 320474 465220
rect 320173 465155 320239 465156
rect 320173 464946 320239 464949
rect 320406 464946 320466 465156
rect 320173 464944 320466 464946
rect 320173 464888 320178 464944
rect 320234 464888 320466 464944
rect 320173 464886 320466 464888
rect 320173 464883 320239 464886
rect 273253 463858 273319 463861
rect 271860 463856 273319 463858
rect 271860 463800 273258 463856
rect 273314 463800 273319 463856
rect 271860 463798 273319 463800
rect 273253 463795 273319 463798
rect 583520 463300 584960 463540
rect 273253 461954 273319 461957
rect 271860 461952 273319 461954
rect 271860 461896 273258 461952
rect 273314 461896 273319 461952
rect 271860 461894 273319 461896
rect 273253 461891 273319 461894
rect 273253 460050 273319 460053
rect 271860 460048 273319 460050
rect 271860 459992 273258 460048
rect 273314 459992 273319 460048
rect 271860 459990 273319 459992
rect 273253 459987 273319 459990
rect 273253 458146 273319 458149
rect 271860 458144 273319 458146
rect 271860 458088 273258 458144
rect 273314 458088 273319 458144
rect 271860 458086 273319 458088
rect 273253 458083 273319 458086
rect 273253 456242 273319 456245
rect 271860 456240 273319 456242
rect 271860 456184 273258 456240
rect 273314 456184 273319 456240
rect 271860 456182 273319 456184
rect 273253 456179 273319 456182
rect 273253 454338 273319 454341
rect 271860 454336 273319 454338
rect 271860 454280 273258 454336
rect 273314 454280 273319 454336
rect 271860 454278 273319 454280
rect 273253 454275 273319 454278
rect -960 452284 480 452524
rect 273253 452434 273319 452437
rect 271860 452432 273319 452434
rect 271860 452376 273258 452432
rect 273314 452376 273319 452432
rect 271860 452374 273319 452376
rect 273253 452371 273319 452374
rect 583520 451604 584960 451844
rect 273345 450530 273411 450533
rect 271860 450528 273411 450530
rect 271860 450472 273350 450528
rect 273406 450472 273411 450528
rect 271860 450470 273411 450472
rect 273345 450467 273411 450470
rect 273437 448626 273503 448629
rect 271860 448624 273503 448626
rect 271860 448568 273442 448624
rect 273498 448568 273503 448624
rect 271860 448566 273503 448568
rect 273437 448563 273503 448566
rect 273437 446722 273503 446725
rect 271860 446720 273503 446722
rect 271860 446664 273442 446720
rect 273498 446664 273503 446720
rect 271860 446662 273503 446664
rect 273437 446659 273503 446662
rect 273437 444818 273503 444821
rect 271860 444816 273503 444818
rect 271860 444760 273442 444816
rect 273498 444760 273503 444816
rect 271860 444758 273503 444760
rect 273437 444755 273503 444758
rect 273437 442914 273503 442917
rect 271860 442912 273503 442914
rect 271860 442856 273442 442912
rect 273498 442856 273503 442912
rect 271860 442854 273503 442856
rect 273437 442851 273503 442854
rect 320449 442370 320515 442373
rect 320725 442370 320791 442373
rect 320449 442368 320791 442370
rect 320449 442312 320454 442368
rect 320510 442312 320730 442368
rect 320786 442312 320791 442368
rect 320449 442310 320791 442312
rect 320449 442307 320515 442310
rect 320725 442307 320791 442310
rect 273437 441010 273503 441013
rect 271860 441008 273503 441010
rect 271860 440952 273442 441008
rect 273498 440952 273503 441008
rect 271860 440950 273503 440952
rect 273437 440947 273503 440950
rect 583520 439772 584960 440012
rect 273437 439106 273503 439109
rect 271860 439104 273503 439106
rect 271860 439048 273442 439104
rect 273498 439048 273503 439104
rect 271860 439046 273503 439048
rect 273437 439043 273503 439046
rect -960 437868 480 438108
rect 274633 437202 274699 437205
rect 271860 437200 274699 437202
rect 271860 437144 274638 437200
rect 274694 437144 274699 437200
rect 271860 437142 274699 437144
rect 274633 437139 274699 437142
rect 274725 435298 274791 435301
rect 271860 435296 274791 435298
rect 271860 435240 274730 435296
rect 274786 435240 274791 435296
rect 271860 435238 274791 435240
rect 274725 435235 274791 435238
rect 273253 433394 273319 433397
rect 271860 433392 273319 433394
rect 271860 433336 273258 433392
rect 273314 433336 273319 433392
rect 271860 433334 273319 433336
rect 273253 433331 273319 433334
rect 273253 431490 273319 431493
rect 271860 431488 273319 431490
rect 271860 431432 273258 431488
rect 273314 431432 273319 431488
rect 271860 431430 273319 431432
rect 273253 431427 273319 431430
rect 273253 429586 273319 429589
rect 271860 429584 273319 429586
rect 271860 429528 273258 429584
rect 273314 429528 273319 429584
rect 271860 429526 273319 429528
rect 273253 429523 273319 429526
rect 583520 428076 584960 428316
rect 273253 427682 273319 427685
rect 271860 427680 273319 427682
rect 271860 427624 273258 427680
rect 273314 427624 273319 427680
rect 271860 427622 273319 427624
rect 273253 427619 273319 427622
rect 273253 425778 273319 425781
rect 271860 425776 273319 425778
rect 271860 425720 273258 425776
rect 273314 425720 273319 425776
rect 271860 425718 273319 425720
rect 273253 425715 273319 425718
rect 273437 423874 273503 423877
rect 271860 423872 273503 423874
rect -960 423588 480 423828
rect 271860 423816 273442 423872
rect 273498 423816 273503 423872
rect 271860 423814 273503 423816
rect 273437 423811 273503 423814
rect 273437 421970 273503 421973
rect 271860 421968 273503 421970
rect 271860 421912 273442 421968
rect 273498 421912 273503 421968
rect 271860 421910 273503 421912
rect 273437 421907 273503 421910
rect 273437 420066 273503 420069
rect 271860 420064 273503 420066
rect 271860 420008 273442 420064
rect 273498 420008 273503 420064
rect 271860 420006 273503 420008
rect 273437 420003 273503 420006
rect 273437 418162 273503 418165
rect 271860 418160 273503 418162
rect 271860 418104 273442 418160
rect 273498 418104 273503 418160
rect 271860 418102 273503 418104
rect 273437 418099 273503 418102
rect 583520 416380 584960 416620
rect 273437 416258 273503 416261
rect 271860 416256 273503 416258
rect 271860 416200 273442 416256
rect 273498 416200 273503 416256
rect 271860 416198 273503 416200
rect 273437 416195 273503 416198
rect 273437 414354 273503 414357
rect 271860 414352 273503 414354
rect 271860 414296 273442 414352
rect 273498 414296 273503 414352
rect 271860 414294 273503 414296
rect 273437 414291 273503 414294
rect 273437 412450 273503 412453
rect 271860 412448 273503 412450
rect 271860 412392 273442 412448
rect 273498 412392 273503 412448
rect 271860 412390 273503 412392
rect 273437 412387 273503 412390
rect 273437 410546 273503 410549
rect 271860 410544 273503 410546
rect 271860 410488 273442 410544
rect 273498 410488 273503 410544
rect 271860 410486 273503 410488
rect 273437 410483 273503 410486
rect -960 409172 480 409412
rect 273437 408642 273503 408645
rect 271860 408640 273503 408642
rect 271860 408584 273442 408640
rect 273498 408584 273503 408640
rect 271860 408582 273503 408584
rect 273437 408579 273503 408582
rect 273437 406738 273503 406741
rect 271860 406736 273503 406738
rect 271860 406680 273442 406736
rect 273498 406680 273503 406736
rect 271860 406678 273503 406680
rect 273437 406675 273503 406678
rect 276606 404834 276612 404836
rect 271860 404774 276612 404834
rect 276606 404772 276612 404774
rect 276676 404772 276682 404836
rect 583520 404684 584960 404924
rect 273437 402930 273503 402933
rect 271860 402928 273503 402930
rect 271860 402872 273442 402928
rect 273498 402872 273503 402928
rect 271860 402870 273503 402872
rect 273437 402867 273503 402870
rect 273437 401026 273503 401029
rect 271860 401024 273503 401026
rect 271860 400968 273442 401024
rect 273498 400968 273503 401024
rect 271860 400966 273503 400968
rect 273437 400963 273503 400966
rect 273437 399122 273503 399125
rect 271860 399120 273503 399122
rect 271860 399064 273442 399120
rect 273498 399064 273503 399120
rect 271860 399062 273503 399064
rect 273437 399059 273503 399062
rect 273437 397218 273503 397221
rect 271860 397216 273503 397218
rect 271860 397160 273442 397216
rect 273498 397160 273503 397216
rect 271860 397158 273503 397160
rect 273437 397155 273503 397158
rect 338665 396810 338731 396813
rect 397453 396810 397519 396813
rect 338665 396808 340255 396810
rect 338665 396752 338670 396808
rect 338726 396752 340255 396808
rect 338665 396750 340255 396752
rect 397453 396808 398084 396810
rect 397453 396752 397458 396808
rect 397514 396752 398084 396808
rect 397453 396750 398084 396752
rect 338665 396747 338731 396750
rect 397453 396747 397519 396750
rect 398833 396674 398899 396677
rect 400213 396674 400279 396677
rect 398833 396672 399832 396674
rect 398833 396616 398838 396672
rect 398894 396616 399832 396672
rect 398833 396614 399832 396616
rect 400213 396672 400936 396674
rect 400213 396616 400218 396672
rect 400274 396616 400936 396672
rect 400213 396614 400936 396616
rect 398833 396611 398899 396614
rect 400213 396611 400279 396614
rect 401593 396538 401659 396541
rect 403341 396538 403407 396541
rect 404353 396538 404419 396541
rect 406009 396538 406075 396541
rect 401593 396536 402631 396538
rect 401593 396480 401598 396536
rect 401654 396480 402631 396536
rect 401593 396478 402631 396480
rect 403341 396536 403788 396538
rect 403341 396480 403346 396536
rect 403402 396480 403788 396536
rect 403341 396478 403788 396480
rect 404353 396536 405444 396538
rect 404353 396480 404358 396536
rect 404414 396480 405444 396536
rect 404353 396478 405444 396480
rect 406009 396536 406587 396538
rect 406009 396480 406014 396536
rect 406070 396480 406587 396536
rect 406009 396478 406587 396480
rect 401593 396475 401659 396478
rect 403341 396475 403407 396478
rect 404353 396475 404419 396478
rect 406009 396475 406075 396478
rect 279918 396068 279924 396132
rect 279988 396130 279994 396132
rect 280061 396130 280127 396133
rect 279988 396128 280127 396130
rect 279988 396072 280066 396128
rect 280122 396072 280127 396128
rect 279988 396070 280127 396072
rect 279988 396068 279994 396070
rect 280061 396067 280127 396070
rect 273437 395314 273503 395317
rect 271860 395312 273503 395314
rect 271860 395256 273442 395312
rect 273498 395256 273503 395312
rect 271860 395254 273503 395256
rect 273437 395251 273503 395254
rect -960 394892 480 395132
rect 273437 393410 273503 393413
rect 271860 393408 273503 393410
rect 271860 393352 273442 393408
rect 273498 393352 273503 393408
rect 271860 393350 273503 393352
rect 273437 393347 273503 393350
rect 583520 392852 584960 393092
rect 320173 392052 320239 392053
rect 320173 392050 320220 392052
rect 320128 392048 320220 392050
rect 320128 391992 320178 392048
rect 320128 391990 320220 391992
rect 320173 391988 320220 391990
rect 320284 391988 320290 392052
rect 320173 391987 320239 391988
rect 273437 391506 273503 391509
rect 271860 391504 273503 391506
rect 271860 391448 273442 391504
rect 273498 391448 273503 391504
rect 271860 391446 273503 391448
rect 273437 391443 273503 391446
rect 320265 389876 320331 389877
rect 320214 389812 320220 389876
rect 320284 389874 320331 389876
rect 320284 389872 320376 389874
rect 320326 389816 320376 389872
rect 320284 389814 320376 389816
rect 320284 389812 320331 389814
rect 320265 389811 320331 389812
rect 273529 389602 273595 389605
rect 271860 389600 273595 389602
rect 271860 389544 273534 389600
rect 273590 389544 273595 389600
rect 271860 389542 273595 389544
rect 273529 389539 273595 389542
rect 320081 389058 320147 389061
rect 320214 389058 320220 389060
rect 320081 389056 320220 389058
rect 320081 389000 320086 389056
rect 320142 389000 320220 389056
rect 320081 388998 320220 389000
rect 320081 388995 320147 388998
rect 320214 388996 320220 388998
rect 320284 388996 320290 389060
rect 273621 387698 273687 387701
rect 271860 387696 273687 387698
rect 271860 387640 273626 387696
rect 273682 387640 273687 387696
rect 271860 387638 273687 387640
rect 273621 387635 273687 387638
rect 320265 387564 320331 387565
rect 320214 387500 320220 387564
rect 320284 387562 320331 387564
rect 320284 387560 320376 387562
rect 320326 387504 320376 387560
rect 320284 387502 320376 387504
rect 320284 387500 320331 387502
rect 320265 387499 320331 387500
rect 319846 386412 319852 386476
rect 319916 386474 319922 386476
rect 320357 386474 320423 386477
rect 319916 386472 320423 386474
rect 319916 386416 320362 386472
rect 320418 386416 320423 386472
rect 319916 386414 320423 386416
rect 319916 386412 319922 386414
rect 320357 386411 320423 386414
rect 320173 386340 320239 386341
rect 320173 386338 320220 386340
rect 320128 386336 320220 386338
rect 320128 386280 320178 386336
rect 320128 386278 320220 386280
rect 320173 386276 320220 386278
rect 320284 386276 320290 386340
rect 320173 386275 320239 386276
rect 273529 385794 273595 385797
rect 271860 385792 273595 385794
rect 271860 385736 273534 385792
rect 273590 385736 273595 385792
rect 271860 385734 273595 385736
rect 273529 385731 273595 385734
rect 320633 384844 320699 384845
rect 320582 384780 320588 384844
rect 320652 384842 320699 384844
rect 320652 384840 320744 384842
rect 320694 384784 320744 384840
rect 320652 384782 320744 384784
rect 320652 384780 320699 384782
rect 320633 384779 320699 384780
rect 274633 383890 274699 383893
rect 271860 383888 274699 383890
rect 271860 383832 274638 383888
rect 274694 383832 274699 383888
rect 271860 383830 274699 383832
rect 274633 383827 274699 383830
rect 319846 383692 319852 383756
rect 319916 383754 319922 383756
rect 320173 383754 320239 383757
rect 319916 383752 320239 383754
rect 319916 383696 320178 383752
rect 320234 383696 320239 383752
rect 319916 383694 320239 383696
rect 319916 383692 319922 383694
rect 320173 383691 320239 383694
rect 320725 383620 320791 383621
rect 320725 383618 320772 383620
rect 320680 383616 320772 383618
rect 320680 383560 320730 383616
rect 320680 383558 320772 383560
rect 320725 383556 320772 383558
rect 320836 383556 320842 383620
rect 320725 383555 320791 383556
rect 320265 383212 320331 383213
rect 320214 383148 320220 383212
rect 320284 383210 320331 383212
rect 320284 383208 320376 383210
rect 320326 383152 320376 383208
rect 320284 383150 320376 383152
rect 320284 383148 320331 383150
rect 320265 383147 320331 383148
rect 320817 382532 320883 382533
rect 320766 382468 320772 382532
rect 320836 382530 320883 382532
rect 320836 382528 320928 382530
rect 320878 382472 320928 382528
rect 320836 382470 320928 382472
rect 320836 382468 320883 382470
rect 320817 382467 320883 382468
rect 273529 381986 273595 381989
rect 271860 381984 273595 381986
rect 271860 381928 273534 381984
rect 273590 381928 273595 381984
rect 271860 381926 273595 381928
rect 273529 381923 273595 381926
rect 320633 381308 320699 381309
rect 320582 381244 320588 381308
rect 320652 381306 320699 381308
rect 320652 381304 320744 381306
rect 320694 381248 320744 381304
rect 320652 381246 320744 381248
rect 320652 381244 320699 381246
rect 320633 381243 320699 381244
rect 583520 381156 584960 381396
rect 320357 380900 320423 380901
rect 320357 380898 320404 380900
rect 320312 380896 320404 380898
rect 320312 380840 320362 380896
rect 320312 380838 320404 380840
rect 320357 380836 320404 380838
rect 320468 380836 320474 380900
rect 320357 380835 320423 380836
rect -960 380476 480 380716
rect 273621 380354 273687 380357
rect 271646 380352 273687 380354
rect 271646 380296 273626 380352
rect 273682 380296 273687 380352
rect 271646 380294 273687 380296
rect 271646 380052 271706 380294
rect 273621 380291 273687 380294
rect 320817 380220 320883 380221
rect 320766 380156 320772 380220
rect 320836 380218 320883 380220
rect 320836 380216 320928 380218
rect 320878 380160 320928 380216
rect 320836 380158 320928 380160
rect 320836 380156 320883 380158
rect 320817 380155 320883 380156
rect 320265 379676 320331 379677
rect 320214 379612 320220 379676
rect 320284 379674 320331 379676
rect 320284 379672 320376 379674
rect 320326 379616 320376 379672
rect 320284 379614 320376 379616
rect 320284 379612 320331 379614
rect 320265 379611 320331 379612
rect 319846 379476 319852 379540
rect 319916 379538 319922 379540
rect 320173 379538 320239 379541
rect 319916 379536 320239 379538
rect 319916 379480 320178 379536
rect 320234 379480 320239 379536
rect 319916 379478 320239 379480
rect 319916 379476 319922 379478
rect 320173 379475 320239 379478
rect 320449 378996 320515 378997
rect 320398 378994 320404 378996
rect 320358 378934 320404 378994
rect 320468 378992 320515 378996
rect 320510 378936 320515 378992
rect 320398 378932 320404 378934
rect 320468 378932 320515 378936
rect 320449 378931 320515 378932
rect 320541 378452 320607 378453
rect 320541 378450 320588 378452
rect 320496 378448 320588 378450
rect 320496 378392 320546 378448
rect 320496 378390 320588 378392
rect 320541 378388 320588 378390
rect 320652 378388 320658 378452
rect 320541 378387 320607 378388
rect 274449 378178 274515 378181
rect 271860 378176 274515 378178
rect 271860 378120 274454 378176
rect 274510 378120 274515 378176
rect 271860 378118 274515 378120
rect 274449 378115 274515 378118
rect 320173 377770 320239 377773
rect 320817 377772 320883 377773
rect 320766 377770 320772 377772
rect 320173 377768 320772 377770
rect 320836 377768 320883 377772
rect 320173 377712 320178 377768
rect 320234 377712 320772 377768
rect 320878 377712 320883 377768
rect 320173 377710 320772 377712
rect 320173 377707 320239 377710
rect 320766 377708 320772 377710
rect 320836 377708 320883 377712
rect 320817 377707 320883 377708
rect 320173 376818 320239 376821
rect 320725 376818 320791 376821
rect 320173 376816 320791 376818
rect 320173 376760 320178 376816
rect 320234 376760 320730 376816
rect 320786 376760 320791 376816
rect 320173 376758 320791 376760
rect 320173 376755 320239 376758
rect 320725 376755 320791 376758
rect 320030 376620 320036 376684
rect 320100 376682 320106 376684
rect 320357 376682 320423 376685
rect 320100 376680 320423 376682
rect 320100 376624 320362 376680
rect 320418 376624 320423 376680
rect 320100 376622 320423 376624
rect 320100 376620 320106 376622
rect 320357 376619 320423 376622
rect 274449 376274 274515 376277
rect 271860 376272 274515 376274
rect 271860 376216 274454 376272
rect 274510 376216 274515 376272
rect 271860 376214 274515 376216
rect 274449 376211 274515 376214
rect 320265 376140 320331 376141
rect 320214 376076 320220 376140
rect 320284 376138 320331 376140
rect 320284 376136 320376 376138
rect 320326 376080 320376 376136
rect 320284 376078 320376 376080
rect 320284 376076 320331 376078
rect 320265 376075 320331 376076
rect 320173 375460 320239 375461
rect 320173 375456 320220 375460
rect 320284 375458 320290 375460
rect 320173 375400 320178 375456
rect 320173 375396 320220 375400
rect 320284 375398 320330 375458
rect 320284 375396 320290 375398
rect 320173 375395 320239 375396
rect 319805 375188 319871 375189
rect 319805 375186 319852 375188
rect 319760 375184 319852 375186
rect 319760 375128 319810 375184
rect 319760 375126 319852 375128
rect 319805 375124 319852 375126
rect 319916 375124 319922 375188
rect 319805 375123 319871 375124
rect 274449 374370 274515 374373
rect 271860 374368 274515 374370
rect 271860 374312 274454 374368
rect 274510 374312 274515 374368
rect 271860 374310 274515 374312
rect 274449 374307 274515 374310
rect 320541 374372 320607 374373
rect 320541 374368 320588 374372
rect 320652 374370 320658 374372
rect 320541 374312 320546 374368
rect 320541 374308 320588 374312
rect 320652 374310 320698 374370
rect 320652 374308 320658 374310
rect 320541 374307 320607 374308
rect 319989 373828 320055 373829
rect 319989 373826 320036 373828
rect 319944 373824 320036 373826
rect 319944 373768 319994 373824
rect 319944 373766 320036 373768
rect 319989 373764 320036 373766
rect 320100 373764 320106 373828
rect 319989 373763 320055 373764
rect 320081 373148 320147 373149
rect 320030 373146 320036 373148
rect 319990 373086 320036 373146
rect 320100 373144 320147 373148
rect 320142 373088 320147 373144
rect 320030 373084 320036 373086
rect 320100 373084 320147 373088
rect 320081 373083 320147 373084
rect 319846 372676 319852 372740
rect 319916 372738 319922 372740
rect 320173 372738 320239 372741
rect 319916 372736 320239 372738
rect 319916 372680 320178 372736
rect 320234 372680 320239 372736
rect 319916 372678 320239 372680
rect 319916 372676 319922 372678
rect 320173 372675 320239 372678
rect 320357 372604 320423 372605
rect 320357 372602 320404 372604
rect 320312 372600 320404 372602
rect 320312 372544 320362 372600
rect 320312 372542 320404 372544
rect 320357 372540 320404 372542
rect 320468 372540 320474 372604
rect 320357 372539 320423 372540
rect 274449 372466 274515 372469
rect 271860 372464 274515 372466
rect 271860 372408 274454 372464
rect 274510 372408 274515 372464
rect 271860 372406 274515 372408
rect 274449 372403 274515 372406
rect 320633 372332 320699 372333
rect 320582 372330 320588 372332
rect 320542 372270 320588 372330
rect 320652 372328 320699 372332
rect 320694 372272 320699 372328
rect 320582 372268 320588 372270
rect 320652 372268 320699 372272
rect 320633 372267 320699 372268
rect 320265 371516 320331 371517
rect 320214 371452 320220 371516
rect 320284 371514 320331 371516
rect 320284 371512 320376 371514
rect 320326 371456 320376 371512
rect 320284 371454 320376 371456
rect 320284 371452 320331 371454
rect 320265 371451 320331 371452
rect 320817 371244 320883 371245
rect 320766 371242 320772 371244
rect 320726 371182 320772 371242
rect 320836 371240 320883 371244
rect 320878 371184 320883 371240
rect 320766 371180 320772 371182
rect 320836 371180 320883 371184
rect 320817 371179 320883 371180
rect 274449 370562 274515 370565
rect 271860 370560 274515 370562
rect 271860 370504 274454 370560
rect 274510 370504 274515 370560
rect 271860 370502 274515 370504
rect 274449 370499 274515 370502
rect 320449 369748 320515 369749
rect 320398 369746 320404 369748
rect 320358 369686 320404 369746
rect 320468 369744 320515 369748
rect 320510 369688 320515 369744
rect 320398 369684 320404 369686
rect 320468 369684 320515 369688
rect 320406 369683 320515 369684
rect 320406 369474 320466 369683
rect 320725 369474 320791 369477
rect 320406 369472 320791 369474
rect 320406 369416 320730 369472
rect 320786 369416 320791 369472
rect 583520 369460 584960 369700
rect 320406 369414 320791 369416
rect 320725 369411 320791 369414
rect 320357 369204 320423 369205
rect 320357 369202 320404 369204
rect 320312 369200 320404 369202
rect 320312 369144 320362 369200
rect 320312 369142 320404 369144
rect 320357 369140 320404 369142
rect 320468 369140 320474 369204
rect 320357 369139 320423 369140
rect 273621 368658 273687 368661
rect 271860 368656 273687 368658
rect 271860 368600 273626 368656
rect 273682 368600 273687 368656
rect 271860 368598 273687 368600
rect 273621 368595 273687 368598
rect 319846 368460 319852 368524
rect 319916 368522 319922 368524
rect 320173 368522 320239 368525
rect 320817 368524 320883 368525
rect 320766 368522 320772 368524
rect 319916 368520 320239 368522
rect 319916 368464 320178 368520
rect 320234 368464 320239 368520
rect 319916 368462 320239 368464
rect 320726 368462 320772 368522
rect 320836 368520 320883 368524
rect 320878 368464 320883 368520
rect 319916 368460 319922 368462
rect 320173 368459 320239 368462
rect 320766 368460 320772 368462
rect 320836 368460 320883 368464
rect 320817 368459 320883 368460
rect 320265 367980 320331 367981
rect 320214 367916 320220 367980
rect 320284 367978 320331 367980
rect 320284 367976 320376 367978
rect 320326 367920 320376 367976
rect 320284 367918 320376 367920
rect 320284 367916 320331 367918
rect 320265 367915 320331 367916
rect 320817 367300 320883 367301
rect 319662 367236 319668 367300
rect 319732 367298 319738 367300
rect 320766 367298 320772 367300
rect 319732 367238 320772 367298
rect 320836 367296 320883 367300
rect 320878 367240 320883 367296
rect 319732 367236 319738 367238
rect 320766 367236 320772 367238
rect 320836 367236 320883 367240
rect 320817 367235 320883 367236
rect 274541 366754 274607 366757
rect 271860 366752 274607 366754
rect 271860 366696 274546 366752
rect 274602 366696 274607 366752
rect 271860 366694 274607 366696
rect 274541 366691 274607 366694
rect -960 366060 480 366300
rect 320633 366212 320699 366213
rect 320582 366210 320588 366212
rect 320542 366150 320588 366210
rect 320652 366208 320699 366212
rect 320694 366152 320699 366208
rect 320582 366148 320588 366150
rect 320652 366148 320699 366152
rect 320633 366147 320699 366148
rect 319805 365666 319871 365669
rect 320030 365666 320036 365668
rect 319805 365664 320036 365666
rect 319805 365608 319810 365664
rect 319866 365608 320036 365664
rect 319805 365606 320036 365608
rect 319805 365603 319871 365606
rect 320030 365604 320036 365606
rect 320100 365604 320106 365668
rect 320173 364988 320239 364989
rect 320173 364984 320220 364988
rect 320284 364986 320290 364988
rect 320633 364986 320699 364989
rect 320284 364984 320699 364986
rect 320173 364928 320178 364984
rect 320284 364928 320638 364984
rect 320694 364928 320699 364984
rect 320173 364924 320220 364928
rect 320284 364926 320699 364928
rect 320284 364924 320290 364926
rect 320173 364923 320239 364924
rect 320633 364923 320699 364926
rect 273805 364850 273871 364853
rect 271860 364848 273871 364850
rect 271860 364792 273810 364848
rect 273866 364792 273871 364848
rect 271860 364790 273871 364792
rect 273805 364787 273871 364790
rect 320449 364444 320515 364445
rect 320398 364380 320404 364444
rect 320468 364442 320515 364444
rect 320468 364440 320560 364442
rect 320510 364384 320560 364440
rect 320468 364382 320560 364384
rect 320468 364380 320515 364382
rect 320449 364379 320515 364380
rect 319989 363764 320055 363765
rect 319989 363760 320036 363764
rect 320100 363762 320106 363764
rect 319989 363704 319994 363760
rect 319989 363700 320036 363704
rect 320100 363702 320146 363762
rect 320100 363700 320106 363702
rect 319989 363699 320055 363700
rect 318793 363490 318859 363493
rect 319478 363490 319484 363492
rect 318793 363488 319484 363490
rect 318793 363432 318798 363488
rect 318854 363432 319484 363488
rect 318793 363430 319484 363432
rect 318793 363427 318859 363430
rect 319478 363428 319484 363430
rect 319548 363428 319554 363492
rect 274357 362946 274423 362949
rect 271860 362944 274423 362946
rect 271860 362888 274362 362944
rect 274418 362888 274423 362944
rect 271860 362886 274423 362888
rect 274357 362883 274423 362886
rect 320081 362676 320147 362677
rect 320030 362674 320036 362676
rect 319990 362614 320036 362674
rect 320100 362672 320147 362676
rect 320142 362616 320147 362672
rect 320030 362612 320036 362614
rect 320100 362612 320147 362616
rect 320081 362611 320147 362612
rect 320357 362132 320423 362133
rect 320357 362130 320404 362132
rect 320312 362128 320404 362130
rect 320312 362072 320362 362128
rect 320312 362070 320404 362072
rect 320357 362068 320404 362070
rect 320468 362068 320474 362132
rect 320357 362067 320423 362068
rect 319805 361452 319871 361453
rect 320173 361452 320239 361453
rect 319805 361450 319852 361452
rect 319760 361448 319852 361450
rect 319760 361392 319810 361448
rect 319760 361390 319852 361392
rect 319805 361388 319852 361390
rect 319916 361388 319922 361452
rect 320173 361448 320220 361452
rect 320284 361450 320290 361452
rect 320173 361392 320178 361448
rect 320173 361388 320220 361392
rect 320284 361390 320330 361450
rect 320284 361388 320290 361390
rect 319805 361387 319871 361388
rect 320173 361387 320239 361388
rect 273529 361042 273595 361045
rect 320265 361044 320331 361045
rect 271860 361040 273595 361042
rect 271860 360984 273534 361040
rect 273590 360984 273595 361040
rect 271860 360982 273595 360984
rect 273529 360979 273595 360982
rect 320214 360980 320220 361044
rect 320284 361042 320331 361044
rect 320284 361040 320376 361042
rect 320326 360984 320376 361040
rect 320284 360982 320376 360984
rect 320284 360980 320331 360982
rect 320265 360979 320331 360980
rect 320265 360364 320331 360365
rect 320214 360362 320220 360364
rect 320174 360302 320220 360362
rect 320284 360360 320331 360364
rect 320326 360304 320331 360360
rect 320214 360300 320220 360302
rect 320284 360300 320331 360304
rect 320265 360299 320331 360300
rect 320449 359820 320515 359821
rect 320398 359818 320404 359820
rect 320358 359758 320404 359818
rect 320468 359818 320515 359820
rect 320725 359818 320791 359821
rect 320468 359816 320791 359818
rect 320510 359760 320730 359816
rect 320786 359760 320791 359816
rect 320398 359756 320404 359758
rect 320468 359758 320791 359760
rect 320468 359756 320515 359758
rect 320449 359755 320515 359756
rect 320725 359755 320791 359758
rect 273805 359138 273871 359141
rect 271860 359136 273871 359138
rect 271860 359080 273810 359136
rect 273866 359080 273871 359136
rect 271860 359078 273871 359080
rect 273805 359075 273871 359078
rect 320357 358596 320423 358597
rect 320357 358594 320404 358596
rect 320312 358592 320404 358594
rect 320312 358536 320362 358592
rect 320312 358534 320404 358536
rect 320357 358532 320404 358534
rect 320468 358532 320474 358596
rect 320357 358531 320423 358532
rect 320265 357916 320331 357917
rect 320214 357914 320220 357916
rect 320174 357854 320220 357914
rect 320284 357912 320331 357916
rect 320326 357856 320331 357912
rect 320214 357852 320220 357854
rect 320284 357852 320331 357856
rect 320265 357851 320331 357852
rect 583520 357764 584960 358004
rect 273846 357234 273852 357236
rect 271860 357174 273852 357234
rect 273846 357172 273852 357174
rect 273916 357172 273922 357236
rect 320541 357100 320607 357101
rect 320541 357098 320588 357100
rect 320496 357096 320588 357098
rect 320496 357040 320546 357096
rect 320496 357038 320588 357040
rect 320541 357036 320588 357038
rect 320652 357036 320658 357100
rect 320541 357035 320607 357036
rect 320173 356828 320239 356829
rect 320173 356826 320220 356828
rect 320128 356824 320220 356826
rect 320128 356768 320178 356824
rect 320128 356766 320220 356768
rect 320173 356764 320220 356766
rect 320284 356764 320290 356828
rect 320173 356763 320239 356764
rect 320633 356012 320699 356013
rect 320582 355948 320588 356012
rect 320652 356010 320699 356012
rect 320652 356008 320744 356010
rect 320694 355952 320744 356008
rect 320652 355950 320744 355952
rect 320652 355948 320699 355950
rect 320633 355947 320699 355948
rect 320173 355604 320239 355605
rect 320173 355602 320220 355604
rect 320128 355600 320220 355602
rect 320128 355544 320178 355600
rect 320128 355542 320220 355544
rect 320173 355540 320220 355542
rect 320284 355540 320290 355604
rect 320173 355539 320239 355540
rect 274357 355330 274423 355333
rect 271860 355328 274423 355330
rect 271860 355272 274362 355328
rect 274418 355272 274423 355328
rect 271860 355270 274423 355272
rect 274357 355267 274423 355270
rect 320817 354652 320883 354653
rect 320766 354650 320772 354652
rect 320726 354590 320772 354650
rect 320836 354648 320883 354652
rect 320878 354592 320883 354648
rect 320766 354588 320772 354590
rect 320836 354588 320883 354592
rect 320817 354587 320883 354588
rect 320173 354516 320239 354517
rect 320173 354514 320220 354516
rect 320128 354512 320220 354514
rect 320128 354456 320178 354512
rect 320128 354454 320220 354456
rect 320173 354452 320220 354454
rect 320284 354452 320290 354516
rect 320173 354451 320239 354452
rect 273805 353426 273871 353429
rect 271860 353424 273871 353426
rect 271860 353368 273810 353424
rect 273866 353368 273871 353424
rect 271860 353366 273871 353368
rect 273805 353363 273871 353366
rect 319846 353364 319852 353428
rect 319916 353426 319922 353428
rect 320265 353426 320331 353429
rect 319916 353424 320331 353426
rect 319916 353368 320270 353424
rect 320326 353368 320331 353424
rect 319916 353366 320331 353368
rect 319916 353364 319922 353366
rect 320265 353363 320331 353366
rect 320265 353292 320331 353293
rect 320817 353292 320883 353293
rect 320214 353228 320220 353292
rect 320284 353290 320331 353292
rect 320766 353290 320772 353292
rect 320284 353288 320376 353290
rect 320326 353232 320376 353288
rect 320284 353230 320376 353232
rect 320726 353230 320772 353290
rect 320836 353288 320883 353292
rect 320878 353232 320883 353288
rect 320284 353228 320331 353230
rect 320766 353228 320772 353230
rect 320836 353228 320883 353232
rect 320265 353227 320331 353228
rect 320817 353227 320883 353228
rect 320173 352612 320239 352613
rect 320173 352610 320220 352612
rect 320128 352608 320220 352610
rect 320128 352552 320178 352608
rect 320128 352550 320220 352552
rect 320173 352548 320220 352550
rect 320284 352548 320290 352612
rect 320173 352547 320239 352548
rect 320357 352476 320423 352477
rect 320357 352474 320404 352476
rect 320312 352472 320404 352474
rect 320312 352416 320362 352472
rect 320312 352414 320404 352416
rect 320357 352412 320404 352414
rect 320468 352412 320474 352476
rect 320357 352411 320423 352412
rect -960 351780 480 352020
rect 274541 351522 274607 351525
rect 271860 351520 274607 351522
rect 271860 351464 274546 351520
rect 274602 351464 274607 351520
rect 271860 351462 274607 351464
rect 274541 351459 274607 351462
rect 320633 351252 320699 351253
rect 320582 351188 320588 351252
rect 320652 351250 320699 351252
rect 320652 351248 320744 351250
rect 320694 351192 320744 351248
rect 320652 351190 320744 351192
rect 320652 351188 320699 351190
rect 320633 351187 320699 351188
rect 320357 350980 320423 350981
rect 320357 350978 320404 350980
rect 320312 350976 320404 350978
rect 320312 350920 320362 350976
rect 320312 350918 320404 350920
rect 320357 350916 320404 350918
rect 320468 350916 320474 350980
rect 320357 350915 320423 350916
rect 320725 350164 320791 350165
rect 320725 350160 320772 350164
rect 320836 350162 320842 350164
rect 320725 350104 320730 350160
rect 320725 350100 320772 350104
rect 320836 350102 320882 350162
rect 320836 350100 320842 350102
rect 320725 350099 320791 350100
rect 320173 349756 320239 349757
rect 320173 349754 320220 349756
rect 320128 349752 320220 349754
rect 320128 349696 320178 349752
rect 320128 349694 320220 349696
rect 320173 349692 320220 349694
rect 320284 349692 320290 349756
rect 320173 349691 320239 349692
rect 273529 349618 273595 349621
rect 271860 349616 273595 349618
rect 271860 349560 273534 349616
rect 273590 349560 273595 349616
rect 271860 349558 273595 349560
rect 273529 349555 273595 349558
rect 320173 348668 320239 348669
rect 320173 348666 320220 348668
rect 320128 348664 320220 348666
rect 320128 348608 320178 348664
rect 320128 348606 320220 348608
rect 320173 348604 320220 348606
rect 320284 348604 320290 348668
rect 320173 348603 320239 348604
rect 273529 347714 273595 347717
rect 271860 347712 273595 347714
rect 271860 347656 273534 347712
rect 273590 347656 273595 347712
rect 271860 347654 273595 347656
rect 273529 347651 273595 347654
rect 320173 346356 320239 346357
rect 320173 346354 320220 346356
rect 320128 346352 320220 346354
rect 320128 346296 320178 346352
rect 320128 346294 320220 346296
rect 320173 346292 320220 346294
rect 320284 346292 320290 346356
rect 320173 346291 320239 346292
rect 583520 345932 584960 346172
rect 273529 345810 273595 345813
rect 271860 345808 273595 345810
rect 271860 345752 273534 345808
rect 273590 345752 273595 345808
rect 271860 345750 273595 345752
rect 273529 345747 273595 345750
rect 273621 343906 273687 343909
rect 271860 343904 273687 343906
rect 271860 343848 273626 343904
rect 273682 343848 273687 343904
rect 271860 343846 273687 343848
rect 273621 343843 273687 343846
rect 273529 342002 273595 342005
rect 271860 342000 273595 342002
rect 271860 341944 273534 342000
rect 273590 341944 273595 342000
rect 271860 341942 273595 341944
rect 273529 341939 273595 341942
rect 273529 340098 273595 340101
rect 271860 340096 273595 340098
rect 271860 340040 273534 340096
rect 273590 340040 273595 340096
rect 271860 340038 273595 340040
rect 273529 340035 273595 340038
rect 273897 338194 273963 338197
rect 271860 338192 273963 338194
rect 271860 338136 273902 338192
rect 273958 338136 273963 338192
rect 271860 338134 273963 338136
rect 273897 338131 273963 338134
rect -960 337364 480 337604
rect 273253 336290 273319 336293
rect 271860 336288 273319 336290
rect 271860 336232 273258 336288
rect 273314 336232 273319 336288
rect 271860 336230 273319 336232
rect 273253 336227 273319 336230
rect 273805 334386 273871 334389
rect 271860 334384 273871 334386
rect 271860 334328 273810 334384
rect 273866 334328 273871 334384
rect 271860 334326 273871 334328
rect 273805 334323 273871 334326
rect 583520 334236 584960 334476
rect 274265 332482 274331 332485
rect 271860 332480 274331 332482
rect 271860 332424 274270 332480
rect 274326 332424 274331 332480
rect 271860 332422 274331 332424
rect 274265 332419 274331 332422
rect 273345 330578 273411 330581
rect 271860 330576 273411 330578
rect 271860 330520 273350 330576
rect 273406 330520 273411 330576
rect 271860 330518 273411 330520
rect 273345 330515 273411 330518
rect 273989 328674 274055 328677
rect 271860 328672 274055 328674
rect 271860 328616 273994 328672
rect 274050 328616 274055 328672
rect 271860 328614 274055 328616
rect 273989 328611 274055 328614
rect 273529 326770 273595 326773
rect 271860 326768 273595 326770
rect 271860 326712 273534 326768
rect 273590 326712 273595 326768
rect 271860 326710 273595 326712
rect 273529 326707 273595 326710
rect 273437 324866 273503 324869
rect 271860 324864 273503 324866
rect 271860 324808 273442 324864
rect 273498 324808 273503 324864
rect 271860 324806 273503 324808
rect 273437 324803 273503 324806
rect -960 322948 480 323188
rect 273529 322962 273595 322965
rect 271860 322960 273595 322962
rect 271860 322904 273534 322960
rect 273590 322904 273595 322960
rect 271860 322902 273595 322904
rect 273529 322899 273595 322902
rect 583520 322540 584960 322780
rect 273437 321058 273503 321061
rect 271860 321056 273503 321058
rect 271860 321000 273442 321056
rect 273498 321000 273503 321056
rect 271860 320998 273503 321000
rect 273437 320995 273503 320998
rect 70158 320588 70164 320652
rect 70228 320650 70234 320652
rect 70301 320650 70367 320653
rect 70228 320648 70367 320650
rect 70228 320592 70306 320648
rect 70362 320592 70367 320648
rect 70228 320590 70367 320592
rect 70228 320588 70234 320590
rect 70301 320587 70367 320590
rect 69013 318746 69079 318749
rect 70209 318746 70275 318749
rect 69013 318744 70275 318746
rect 69013 318688 69018 318744
rect 69074 318688 70214 318744
rect 70270 318688 70275 318744
rect 69013 318686 70275 318688
rect 69013 318683 69079 318686
rect 70209 318683 70275 318686
rect 164233 318746 164299 318749
rect 166993 318746 167059 318749
rect 164233 318744 167059 318746
rect 164233 318688 164238 318744
rect 164294 318688 166998 318744
rect 167054 318688 167059 318744
rect 164233 318686 167059 318688
rect 164233 318683 164299 318686
rect 166993 318683 167059 318686
rect 23381 318610 23447 318613
rect 78029 318610 78095 318613
rect 23381 318608 78095 318610
rect 23381 318552 23386 318608
rect 23442 318552 78034 318608
rect 78090 318552 78095 318608
rect 23381 318550 78095 318552
rect 23381 318547 23447 318550
rect 78029 318547 78095 318550
rect 229737 318610 229803 318613
rect 237189 318610 237255 318613
rect 374637 318610 374703 318613
rect 229737 318608 237114 318610
rect 229737 318552 229742 318608
rect 229798 318552 237114 318608
rect 229737 318550 237114 318552
rect 229737 318547 229803 318550
rect 17861 318474 17927 318477
rect 75913 318474 75979 318477
rect 17861 318472 75979 318474
rect 17861 318416 17866 318472
rect 17922 318416 75918 318472
rect 75974 318416 75979 318472
rect 17861 318414 75979 318416
rect 237054 318474 237114 318550
rect 237189 318608 374703 318610
rect 237189 318552 237194 318608
rect 237250 318552 374642 318608
rect 374698 318552 374703 318608
rect 237189 318550 374703 318552
rect 237189 318547 237255 318550
rect 374637 318547 374703 318550
rect 367737 318474 367803 318477
rect 237054 318472 367803 318474
rect 237054 318416 367742 318472
rect 367798 318416 367803 318472
rect 237054 318414 367803 318416
rect 17861 318411 17927 318414
rect 75913 318411 75979 318414
rect 367737 318411 367803 318414
rect 16481 318338 16547 318341
rect 75545 318338 75611 318341
rect 16481 318336 75611 318338
rect 16481 318280 16486 318336
rect 16542 318280 75550 318336
rect 75606 318280 75611 318336
rect 16481 318278 75611 318280
rect 16481 318275 16547 318278
rect 75545 318275 75611 318278
rect 234705 318338 234771 318341
rect 373257 318338 373323 318341
rect 234705 318336 373323 318338
rect 234705 318280 234710 318336
rect 234766 318280 373262 318336
rect 373318 318280 373323 318336
rect 234705 318278 373323 318280
rect 234705 318275 234771 318278
rect 373257 318275 373323 318278
rect 15101 318202 15167 318205
rect 75085 318202 75151 318205
rect 15101 318200 75151 318202
rect 15101 318144 15106 318200
rect 15162 318144 75090 318200
rect 75146 318144 75151 318200
rect 15101 318142 75151 318144
rect 15101 318139 15167 318142
rect 75085 318139 75151 318142
rect 147397 318202 147463 318205
rect 147857 318202 147923 318205
rect 147397 318200 147923 318202
rect 147397 318144 147402 318200
rect 147458 318144 147862 318200
rect 147918 318144 147923 318200
rect 147397 318142 147923 318144
rect 147397 318139 147463 318142
rect 147857 318139 147923 318142
rect 227253 318202 227319 318205
rect 364977 318202 365043 318205
rect 227253 318200 365043 318202
rect 227253 318144 227258 318200
rect 227314 318144 364982 318200
rect 365038 318144 365043 318200
rect 227253 318142 365043 318144
rect 227253 318139 227319 318142
rect 364977 318139 365043 318142
rect 13721 318066 13787 318069
rect 74717 318066 74783 318069
rect 13721 318064 74783 318066
rect 13721 318008 13726 318064
rect 13782 318008 74722 318064
rect 74778 318008 74783 318064
rect 13721 318006 74783 318008
rect 13721 318003 13787 318006
rect 74717 318003 74783 318006
rect 143165 318066 143231 318069
rect 163497 318066 163563 318069
rect 143165 318064 163563 318066
rect 143165 318008 143170 318064
rect 143226 318008 163502 318064
rect 163558 318008 163563 318064
rect 143165 318006 163563 318008
rect 143165 318003 143231 318006
rect 163497 318003 163563 318006
rect 232221 318066 232287 318069
rect 371877 318066 371943 318069
rect 232221 318064 371943 318066
rect 232221 318008 232226 318064
rect 232282 318008 371882 318064
rect 371938 318008 371943 318064
rect 232221 318006 371943 318008
rect 232221 318003 232287 318006
rect 371877 318003 371943 318006
rect 265341 314666 265407 314669
rect 265801 314666 265867 314669
rect 265341 314664 265867 314666
rect 265341 314608 265346 314664
rect 265402 314608 265806 314664
rect 265862 314608 265867 314664
rect 265341 314606 265867 314608
rect 265341 314603 265407 314606
rect 265801 314603 265867 314606
rect 583520 310708 584960 310948
rect 252921 309226 252987 309229
rect 252694 309224 252987 309226
rect 252694 309168 252926 309224
rect 252982 309168 252987 309224
rect 252694 309166 252987 309168
rect 252694 309093 252754 309166
rect 252921 309163 252987 309166
rect 252694 309088 252803 309093
rect 252694 309032 252742 309088
rect 252798 309032 252803 309088
rect 252694 309030 252803 309032
rect 252737 309027 252803 309030
rect -960 308668 480 308908
rect 90449 307866 90515 307869
rect 90222 307864 90515 307866
rect 90222 307808 90454 307864
rect 90510 307808 90515 307864
rect 90222 307806 90515 307808
rect 90222 307733 90282 307806
rect 90449 307803 90515 307806
rect 90173 307728 90282 307733
rect 90173 307672 90178 307728
rect 90234 307672 90282 307728
rect 90173 307670 90282 307672
rect 90173 307667 90239 307670
rect 583520 299012 584960 299252
rect 105169 298074 105235 298077
rect 105353 298074 105419 298077
rect 105169 298072 105419 298074
rect 105169 298016 105174 298072
rect 105230 298016 105358 298072
rect 105414 298016 105419 298072
rect 105169 298014 105419 298016
rect 105169 298011 105235 298014
rect 105353 298011 105419 298014
rect 89989 296714 90055 296717
rect 90265 296714 90331 296717
rect 89989 296712 90331 296714
rect 89989 296656 89994 296712
rect 90050 296656 90270 296712
rect 90326 296656 90331 296712
rect 89989 296654 90331 296656
rect 89989 296651 90055 296654
rect 90265 296651 90331 296654
rect 233969 296714 234035 296717
rect 234245 296714 234311 296717
rect 233969 296712 234311 296714
rect 233969 296656 233974 296712
rect 234030 296656 234250 296712
rect 234306 296656 234311 296712
rect 233969 296654 234311 296656
rect 233969 296651 234035 296654
rect 234245 296651 234311 296654
rect -960 294252 480 294492
rect 263685 293994 263751 293997
rect 264697 293994 264763 293997
rect 263685 293992 264763 293994
rect 263685 293936 263690 293992
rect 263746 293936 264702 293992
rect 264758 293936 264763 293992
rect 263685 293934 264763 293936
rect 263685 293931 263751 293934
rect 264697 293931 264763 293934
rect 583520 287316 584960 287556
rect 72325 287058 72391 287061
rect 72509 287058 72575 287061
rect 72325 287056 72575 287058
rect 72325 287000 72330 287056
rect 72386 287000 72514 287056
rect 72570 287000 72575 287056
rect 72325 286998 72575 287000
rect 72325 286995 72391 286998
rect 72509 286995 72575 286998
rect 81617 287058 81683 287061
rect 81801 287058 81867 287061
rect 81617 287056 81867 287058
rect 81617 287000 81622 287056
rect 81678 287000 81806 287056
rect 81862 287000 81867 287056
rect 81617 286998 81867 287000
rect 81617 286995 81683 286998
rect 81801 286995 81867 286998
rect 94129 287058 94195 287061
rect 94313 287058 94379 287061
rect 94129 287056 94379 287058
rect 94129 287000 94134 287056
rect 94190 287000 94318 287056
rect 94374 287000 94379 287056
rect 94129 286998 94379 287000
rect 94129 286995 94195 286998
rect 94313 286995 94379 286998
rect -960 279972 480 280212
rect 193673 278762 193739 278765
rect 193857 278762 193923 278765
rect 255221 278762 255287 278765
rect 193673 278760 193923 278762
rect 193673 278704 193678 278760
rect 193734 278704 193862 278760
rect 193918 278704 193923 278760
rect 193673 278702 193923 278704
rect 193673 278699 193739 278702
rect 193857 278699 193923 278702
rect 255086 278760 255287 278762
rect 255086 278704 255226 278760
rect 255282 278704 255287 278760
rect 255086 278702 255287 278704
rect 255086 278626 255146 278702
rect 255221 278699 255287 278702
rect 255313 278626 255379 278629
rect 255086 278624 255379 278626
rect 255086 278568 255318 278624
rect 255374 278568 255379 278624
rect 255086 278566 255379 278568
rect 255313 278563 255379 278566
rect 72325 277402 72391 277405
rect 72601 277402 72667 277405
rect 72325 277400 72667 277402
rect 72325 277344 72330 277400
rect 72386 277344 72606 277400
rect 72662 277344 72667 277400
rect 72325 277342 72667 277344
rect 72325 277339 72391 277342
rect 72601 277339 72667 277342
rect 73429 277402 73495 277405
rect 73613 277402 73679 277405
rect 73429 277400 73679 277402
rect 73429 277344 73434 277400
rect 73490 277344 73618 277400
rect 73674 277344 73679 277400
rect 73429 277342 73679 277344
rect 73429 277339 73495 277342
rect 73613 277339 73679 277342
rect 583520 275620 584960 275860
rect 264513 274682 264579 274685
rect 264697 274682 264763 274685
rect 264513 274680 264763 274682
rect 264513 274624 264518 274680
rect 264574 274624 264702 274680
rect 264758 274624 264763 274680
rect 264513 274622 264763 274624
rect 264513 274619 264579 274622
rect 264697 274619 264763 274622
rect 78673 267746 78739 267749
rect 78949 267746 79015 267749
rect 78673 267744 79015 267746
rect 78673 267688 78678 267744
rect 78734 267688 78954 267744
rect 79010 267688 79015 267744
rect 78673 267686 79015 267688
rect 78673 267683 78739 267686
rect 78949 267683 79015 267686
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 193673 259450 193739 259453
rect 193857 259450 193923 259453
rect 193673 259448 193923 259450
rect 193673 259392 193678 259448
rect 193734 259392 193862 259448
rect 193918 259392 193923 259448
rect 193673 259390 193923 259392
rect 193673 259387 193739 259390
rect 193857 259387 193923 259390
rect 246941 259450 247007 259453
rect 247125 259450 247191 259453
rect 246941 259448 247191 259450
rect 246941 259392 246946 259448
rect 247002 259392 247130 259448
rect 247186 259392 247191 259448
rect 246941 259390 247191 259392
rect 246941 259387 247007 259390
rect 247125 259387 247191 259390
rect 81709 258090 81775 258093
rect 81893 258090 81959 258093
rect 81709 258088 81959 258090
rect 81709 258032 81714 258088
rect 81770 258032 81898 258088
rect 81954 258032 81959 258088
rect 81709 258030 81959 258032
rect 81709 258027 81775 258030
rect 81893 258027 81959 258030
rect 583520 252092 584960 252332
rect -960 251140 480 251380
rect 242341 249794 242407 249797
rect 242525 249794 242591 249797
rect 242341 249792 242591 249794
rect 242341 249736 242346 249792
rect 242402 249736 242530 249792
rect 242586 249736 242591 249792
rect 242341 249734 242591 249736
rect 242341 249731 242407 249734
rect 242525 249731 242591 249734
rect 77477 248434 77543 248437
rect 77845 248434 77911 248437
rect 77477 248432 77911 248434
rect 77477 248376 77482 248432
rect 77538 248376 77850 248432
rect 77906 248376 77911 248432
rect 77477 248374 77911 248376
rect 77477 248371 77543 248374
rect 77845 248371 77911 248374
rect 193857 241770 193923 241773
rect 193857 241768 194058 241770
rect 193857 241712 193862 241768
rect 193918 241712 194058 241768
rect 193857 241710 194058 241712
rect 193857 241707 193923 241710
rect 193857 241634 193923 241637
rect 193998 241634 194058 241710
rect 193857 241632 194058 241634
rect 193857 241576 193862 241632
rect 193918 241576 194058 241632
rect 193857 241574 194058 241576
rect 193857 241571 193923 241574
rect 106641 241500 106707 241501
rect 106590 241498 106596 241500
rect 106550 241438 106596 241498
rect 106660 241496 106707 241500
rect 106702 241440 106707 241496
rect 106590 241436 106596 241438
rect 106660 241436 106707 241440
rect 106641 241435 106707 241436
rect 151077 241498 151143 241501
rect 151077 241496 151186 241498
rect 151077 241440 151082 241496
rect 151138 241440 151186 241496
rect 151077 241435 151186 241440
rect 150985 241362 151051 241365
rect 151126 241362 151186 241435
rect 150985 241360 151186 241362
rect 150985 241304 150990 241360
rect 151046 241304 151186 241360
rect 150985 241302 151186 241304
rect 150985 241299 151051 241302
rect 583520 240396 584960 240636
rect 89989 240138 90055 240141
rect 90173 240138 90239 240141
rect 89989 240136 90239 240138
rect 89989 240080 89994 240136
rect 90050 240080 90178 240136
rect 90234 240080 90239 240136
rect 89989 240078 90239 240080
rect 89989 240075 90055 240078
rect 90173 240075 90239 240078
rect 193673 240138 193739 240141
rect 193857 240138 193923 240141
rect 193673 240136 193923 240138
rect 193673 240080 193678 240136
rect 193734 240080 193862 240136
rect 193918 240080 193923 240136
rect 193673 240078 193923 240080
rect 193673 240075 193739 240078
rect 193857 240075 193923 240078
rect 246941 240138 247007 240141
rect 247125 240138 247191 240141
rect 246941 240136 247191 240138
rect 246941 240080 246946 240136
rect 247002 240080 247130 240136
rect 247186 240080 247191 240136
rect 246941 240078 247191 240080
rect 246941 240075 247007 240078
rect 247125 240075 247191 240078
rect 250805 240138 250871 240141
rect 250989 240138 251055 240141
rect 250805 240136 251055 240138
rect 250805 240080 250810 240136
rect 250866 240080 250994 240136
rect 251050 240080 251055 240136
rect 250805 240078 251055 240080
rect 250805 240075 250871 240078
rect 250989 240075 251055 240078
rect 252093 240138 252159 240141
rect 252277 240138 252343 240141
rect 252093 240136 252343 240138
rect 252093 240080 252098 240136
rect 252154 240080 252282 240136
rect 252338 240080 252343 240136
rect 252093 240078 252343 240080
rect 252093 240075 252159 240078
rect 252277 240075 252343 240078
rect 259085 240138 259151 240141
rect 259269 240138 259335 240141
rect 259085 240136 259335 240138
rect 259085 240080 259090 240136
rect 259146 240080 259274 240136
rect 259330 240080 259335 240136
rect 259085 240078 259335 240080
rect 259085 240075 259151 240078
rect 259269 240075 259335 240078
rect -960 236860 480 237100
rect 106549 235380 106615 235381
rect 106549 235378 106596 235380
rect 106504 235376 106596 235378
rect 106504 235320 106554 235376
rect 106504 235318 106596 235320
rect 106549 235316 106596 235318
rect 106660 235316 106666 235380
rect 106549 235315 106615 235316
rect 73429 231842 73495 231845
rect 73705 231842 73771 231845
rect 73429 231840 73771 231842
rect 73429 231784 73434 231840
rect 73490 231784 73710 231840
rect 73766 231784 73771 231840
rect 73429 231782 73771 231784
rect 73429 231779 73495 231782
rect 73705 231779 73771 231782
rect 324865 231842 324931 231845
rect 325049 231842 325115 231845
rect 324865 231840 325115 231842
rect 324865 231784 324870 231840
rect 324926 231784 325054 231840
rect 325110 231784 325115 231840
rect 324865 231782 325115 231784
rect 324865 231779 324931 231782
rect 325049 231779 325115 231782
rect 90633 230482 90699 230485
rect 90817 230482 90883 230485
rect 90633 230480 90883 230482
rect 90633 230424 90638 230480
rect 90694 230424 90822 230480
rect 90878 230424 90883 230480
rect 90633 230422 90883 230424
rect 90633 230419 90699 230422
rect 90817 230419 90883 230422
rect 242341 230482 242407 230485
rect 242525 230482 242591 230485
rect 242341 230480 242591 230482
rect 242341 230424 242346 230480
rect 242402 230424 242530 230480
rect 242586 230424 242591 230480
rect 242341 230422 242591 230424
rect 242341 230419 242407 230422
rect 242525 230419 242591 230422
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 81709 222186 81775 222189
rect 94037 222186 94103 222189
rect 94313 222186 94379 222189
rect 81709 222184 81818 222186
rect 81709 222128 81714 222184
rect 81770 222128 81818 222184
rect 81709 222123 81818 222128
rect 94037 222184 94379 222186
rect 94037 222128 94042 222184
rect 94098 222128 94318 222184
rect 94374 222128 94379 222184
rect 94037 222126 94379 222128
rect 94037 222123 94103 222126
rect 94313 222123 94379 222126
rect 151077 222186 151143 222189
rect 151077 222184 151186 222186
rect 151077 222128 151082 222184
rect 151138 222128 151186 222184
rect 151077 222123 151186 222128
rect 81758 222053 81818 222123
rect 81758 222048 81867 222053
rect 81758 221992 81806 222048
rect 81862 221992 81867 222048
rect 81758 221990 81867 221992
rect 81801 221987 81867 221990
rect 150985 222050 151051 222053
rect 151126 222050 151186 222123
rect 150985 222048 151186 222050
rect 150985 221992 150990 222048
rect 151046 221992 151186 222048
rect 150985 221990 151186 221992
rect 150985 221987 151051 221990
rect 193673 220826 193739 220829
rect 193857 220826 193923 220829
rect 193673 220824 193923 220826
rect 193673 220768 193678 220824
rect 193734 220768 193862 220824
rect 193918 220768 193923 220824
rect 193673 220766 193923 220768
rect 193673 220763 193739 220766
rect 193857 220763 193923 220766
rect 246941 220826 247007 220829
rect 247125 220826 247191 220829
rect 246941 220824 247191 220826
rect 246941 220768 246946 220824
rect 247002 220768 247130 220824
rect 247186 220768 247191 220824
rect 246941 220766 247191 220768
rect 246941 220763 247007 220766
rect 247125 220763 247191 220766
rect 250805 220826 250871 220829
rect 250989 220826 251055 220829
rect 250805 220824 251055 220826
rect 250805 220768 250810 220824
rect 250866 220768 250994 220824
rect 251050 220768 251055 220824
rect 250805 220766 251055 220768
rect 250805 220763 250871 220766
rect 250989 220763 251055 220766
rect 252093 220826 252159 220829
rect 252277 220826 252343 220829
rect 252093 220824 252343 220826
rect 252093 220768 252098 220824
rect 252154 220768 252282 220824
rect 252338 220768 252343 220824
rect 252093 220766 252343 220768
rect 252093 220763 252159 220766
rect 252277 220763 252343 220766
rect 259085 220826 259151 220829
rect 259269 220826 259335 220829
rect 259085 220824 259335 220826
rect 259085 220768 259090 220824
rect 259146 220768 259274 220824
rect 259330 220768 259335 220824
rect 259085 220766 259335 220768
rect 259085 220763 259151 220766
rect 259269 220763 259335 220766
rect 255313 219466 255379 219469
rect 255497 219466 255563 219469
rect 255313 219464 255563 219466
rect 255313 219408 255318 219464
rect 255374 219408 255502 219464
rect 255558 219408 255563 219464
rect 255313 219406 255563 219408
rect 255313 219403 255379 219406
rect 255497 219403 255563 219406
rect 233785 217970 233851 217973
rect 234061 217970 234127 217973
rect 233785 217968 234127 217970
rect 233785 217912 233790 217968
rect 233846 217912 234066 217968
rect 234122 217912 234127 217968
rect 233785 217910 234127 217912
rect 233785 217907 233851 217910
rect 234061 217907 234127 217910
rect 583520 216868 584960 217108
rect 73429 212530 73495 212533
rect 73705 212530 73771 212533
rect 73429 212528 73771 212530
rect 73429 212472 73434 212528
rect 73490 212472 73710 212528
rect 73766 212472 73771 212528
rect 73429 212470 73771 212472
rect 73429 212467 73495 212470
rect 73705 212467 73771 212470
rect 92749 212530 92815 212533
rect 92933 212530 92999 212533
rect 92749 212528 92999 212530
rect 92749 212472 92754 212528
rect 92810 212472 92938 212528
rect 92994 212472 92999 212528
rect 92749 212470 92999 212472
rect 92749 212467 92815 212470
rect 92933 212467 92999 212470
rect 324865 212530 324931 212533
rect 325049 212530 325115 212533
rect 324865 212528 325115 212530
rect 324865 212472 324870 212528
rect 324926 212472 325054 212528
rect 325110 212472 325115 212528
rect 324865 212470 325115 212472
rect 324865 212467 324931 212470
rect 325049 212467 325115 212470
rect 193673 211170 193739 211173
rect 193857 211170 193923 211173
rect 193673 211168 193923 211170
rect 193673 211112 193678 211168
rect 193734 211112 193862 211168
rect 193918 211112 193923 211168
rect 193673 211110 193923 211112
rect 193673 211107 193739 211110
rect 193857 211107 193923 211110
rect 246941 211170 247007 211173
rect 247125 211170 247191 211173
rect 246941 211168 247191 211170
rect 246941 211112 246946 211168
rect 247002 211112 247130 211168
rect 247186 211112 247191 211168
rect 246941 211110 247191 211112
rect 246941 211107 247007 211110
rect 247125 211107 247191 211110
rect 250805 211170 250871 211173
rect 250989 211170 251055 211173
rect 250805 211168 251055 211170
rect 250805 211112 250810 211168
rect 250866 211112 250994 211168
rect 251050 211112 251055 211168
rect 250805 211110 251055 211112
rect 250805 211107 250871 211110
rect 250989 211107 251055 211110
rect 252093 211170 252159 211173
rect 252277 211170 252343 211173
rect 252093 211168 252343 211170
rect 252093 211112 252098 211168
rect 252154 211112 252282 211168
rect 252338 211112 252343 211168
rect 252093 211110 252343 211112
rect 252093 211107 252159 211110
rect 252277 211107 252343 211110
rect 259085 211170 259151 211173
rect 259269 211170 259335 211173
rect 259085 211168 259335 211170
rect 259085 211112 259090 211168
rect 259146 211112 259274 211168
rect 259330 211112 259335 211168
rect 259085 211110 259335 211112
rect 259085 211107 259151 211110
rect 259269 211107 259335 211110
rect -960 208028 480 208268
rect 583520 205172 584960 205412
rect 77477 202876 77543 202877
rect 77477 202874 77524 202876
rect 77432 202872 77524 202874
rect 77432 202816 77482 202872
rect 77432 202814 77524 202816
rect 77477 202812 77524 202814
rect 77588 202812 77594 202876
rect 78765 202874 78831 202877
rect 78630 202872 78831 202874
rect 78630 202816 78770 202872
rect 78826 202816 78831 202872
rect 78630 202814 78831 202816
rect 77477 202811 77543 202812
rect 78630 202738 78690 202814
rect 78765 202811 78831 202814
rect 151077 202874 151143 202877
rect 151077 202872 151186 202874
rect 151077 202816 151082 202872
rect 151138 202816 151186 202872
rect 151077 202811 151186 202816
rect 78857 202738 78923 202741
rect 78630 202736 78923 202738
rect 78630 202680 78862 202736
rect 78918 202680 78923 202736
rect 78630 202678 78923 202680
rect 78857 202675 78923 202678
rect 150985 202738 151051 202741
rect 151126 202738 151186 202811
rect 150985 202736 151186 202738
rect 150985 202680 150990 202736
rect 151046 202680 151186 202736
rect 150985 202678 151186 202680
rect 150985 202675 151051 202678
rect 242341 201514 242407 201517
rect 242525 201514 242591 201517
rect 242341 201512 242591 201514
rect 242341 201456 242346 201512
rect 242402 201456 242530 201512
rect 242586 201456 242591 201512
rect 242341 201454 242591 201456
rect 242341 201451 242407 201454
rect 242525 201451 242591 201454
rect 77569 195804 77635 195805
rect 77518 195802 77524 195804
rect 77478 195742 77524 195802
rect 77588 195800 77635 195804
rect 77630 195744 77635 195800
rect 77518 195740 77524 195742
rect 77588 195740 77635 195744
rect 77569 195739 77635 195740
rect -960 193748 480 193988
rect 583520 193476 584960 193716
rect 89989 193218 90055 193221
rect 90173 193218 90239 193221
rect 89989 193216 90239 193218
rect 89989 193160 89994 193216
rect 90050 193160 90178 193216
rect 90234 193160 90239 193216
rect 89989 193158 90239 193160
rect 89989 193155 90055 193158
rect 90173 193155 90239 193158
rect 106641 193218 106707 193221
rect 106825 193218 106891 193221
rect 106641 193216 106891 193218
rect 106641 193160 106646 193216
rect 106702 193160 106830 193216
rect 106886 193160 106891 193216
rect 106641 193158 106891 193160
rect 106641 193155 106707 193158
rect 106825 193155 106891 193158
rect 324865 193218 324931 193221
rect 325049 193218 325115 193221
rect 324865 193216 325115 193218
rect 324865 193160 324870 193216
rect 324926 193160 325054 193216
rect 325110 193160 325115 193216
rect 324865 193158 325115 193160
rect 324865 193155 324931 193158
rect 325049 193155 325115 193158
rect 193673 191858 193739 191861
rect 193857 191858 193923 191861
rect 193673 191856 193923 191858
rect 193673 191800 193678 191856
rect 193734 191800 193862 191856
rect 193918 191800 193923 191856
rect 193673 191798 193923 191800
rect 193673 191795 193739 191798
rect 193857 191795 193923 191798
rect 246941 191858 247007 191861
rect 247125 191858 247191 191861
rect 246941 191856 247191 191858
rect 246941 191800 246946 191856
rect 247002 191800 247130 191856
rect 247186 191800 247191 191856
rect 246941 191798 247191 191800
rect 246941 191795 247007 191798
rect 247125 191795 247191 191798
rect 81709 183562 81775 183565
rect 81893 183562 81959 183565
rect 81709 183560 81959 183562
rect 81709 183504 81714 183560
rect 81770 183504 81898 183560
rect 81954 183504 81959 183560
rect 81709 183502 81959 183504
rect 81709 183499 81775 183502
rect 81893 183499 81959 183502
rect 151077 183562 151143 183565
rect 211705 183562 211771 183565
rect 211889 183562 211955 183565
rect 151077 183560 151186 183562
rect 151077 183504 151082 183560
rect 151138 183504 151186 183560
rect 151077 183499 151186 183504
rect 211705 183560 211955 183562
rect 211705 183504 211710 183560
rect 211766 183504 211894 183560
rect 211950 183504 211955 183560
rect 211705 183502 211955 183504
rect 211705 183499 211771 183502
rect 211889 183499 211955 183502
rect 227161 183562 227227 183565
rect 227345 183562 227411 183565
rect 227161 183560 227411 183562
rect 227161 183504 227166 183560
rect 227222 183504 227350 183560
rect 227406 183504 227411 183560
rect 227161 183502 227411 183504
rect 227161 183499 227227 183502
rect 227345 183499 227411 183502
rect 150985 183426 151051 183429
rect 151126 183426 151186 183499
rect 150985 183424 151186 183426
rect 150985 183368 150990 183424
rect 151046 183368 151186 183424
rect 150985 183366 151186 183368
rect 150985 183363 151051 183366
rect 72049 182202 72115 182205
rect 72325 182202 72391 182205
rect 72049 182200 72391 182202
rect 72049 182144 72054 182200
rect 72110 182144 72330 182200
rect 72386 182144 72391 182200
rect 72049 182142 72391 182144
rect 72049 182139 72115 182142
rect 72325 182139 72391 182142
rect 73337 182202 73403 182205
rect 73613 182202 73679 182205
rect 73337 182200 73679 182202
rect 73337 182144 73342 182200
rect 73398 182144 73618 182200
rect 73674 182144 73679 182200
rect 73337 182142 73679 182144
rect 73337 182139 73403 182142
rect 73613 182139 73679 182142
rect 242341 182202 242407 182205
rect 242525 182202 242591 182205
rect 242341 182200 242591 182202
rect 242341 182144 242346 182200
rect 242402 182144 242530 182200
rect 242586 182144 242591 182200
rect 242341 182142 242591 182144
rect 242341 182139 242407 182142
rect 242525 182139 242591 182142
rect 583520 181780 584960 182020
rect 235533 180842 235599 180845
rect 235717 180842 235783 180845
rect 235533 180840 235783 180842
rect 235533 180784 235538 180840
rect 235594 180784 235722 180840
rect 235778 180784 235783 180840
rect 235533 180782 235783 180784
rect 235533 180779 235599 180782
rect 235717 180779 235783 180782
rect 260281 180842 260347 180845
rect 260465 180842 260531 180845
rect 260281 180840 260531 180842
rect 260281 180784 260286 180840
rect 260342 180784 260470 180840
rect 260526 180784 260531 180840
rect 260281 180782 260531 180784
rect 260281 180779 260347 180782
rect 260465 180779 260531 180782
rect 267089 180842 267155 180845
rect 267273 180842 267339 180845
rect 267089 180840 267339 180842
rect 267089 180784 267094 180840
rect 267150 180784 267278 180840
rect 267334 180784 267339 180840
rect 267089 180782 267339 180784
rect 267089 180779 267155 180782
rect 267273 180779 267339 180782
rect -960 179332 480 179572
rect 106457 173906 106523 173909
rect 106733 173906 106799 173909
rect 106457 173904 106799 173906
rect 106457 173848 106462 173904
rect 106518 173848 106738 173904
rect 106794 173848 106799 173904
rect 106457 173846 106799 173848
rect 106457 173843 106523 173846
rect 106733 173843 106799 173846
rect 234153 173906 234219 173909
rect 234337 173906 234403 173909
rect 234153 173904 234403 173906
rect 234153 173848 234158 173904
rect 234214 173848 234342 173904
rect 234398 173848 234403 173904
rect 234153 173846 234403 173848
rect 234153 173843 234219 173846
rect 234337 173843 234403 173846
rect 324865 173906 324931 173909
rect 325049 173906 325115 173909
rect 324865 173904 325115 173906
rect 324865 173848 324870 173904
rect 324926 173848 325054 173904
rect 325110 173848 325115 173904
rect 324865 173846 325115 173848
rect 324865 173843 324931 173846
rect 325049 173843 325115 173846
rect 193673 172546 193739 172549
rect 193857 172546 193923 172549
rect 193673 172544 193923 172546
rect 193673 172488 193678 172544
rect 193734 172488 193862 172544
rect 193918 172488 193923 172544
rect 193673 172486 193923 172488
rect 193673 172483 193739 172486
rect 193857 172483 193923 172486
rect 246941 172546 247007 172549
rect 247125 172546 247191 172549
rect 246941 172544 247191 172546
rect 246941 172488 246946 172544
rect 247002 172488 247130 172544
rect 247186 172488 247191 172544
rect 246941 172486 247191 172488
rect 246941 172483 247007 172486
rect 247125 172483 247191 172486
rect 250805 172546 250871 172549
rect 250989 172546 251055 172549
rect 250805 172544 251055 172546
rect 250805 172488 250810 172544
rect 250866 172488 250994 172544
rect 251050 172488 251055 172544
rect 250805 172486 251055 172488
rect 250805 172483 250871 172486
rect 250989 172483 251055 172486
rect 252093 172546 252159 172549
rect 252277 172546 252343 172549
rect 252093 172544 252343 172546
rect 252093 172488 252098 172544
rect 252154 172488 252282 172544
rect 252338 172488 252343 172544
rect 252093 172486 252343 172488
rect 252093 172483 252159 172486
rect 252277 172483 252343 172486
rect 259085 172546 259151 172549
rect 259269 172546 259335 172549
rect 259085 172544 259335 172546
rect 259085 172488 259090 172544
rect 259146 172488 259274 172544
rect 259330 172488 259335 172544
rect 259085 172486 259335 172488
rect 259085 172483 259151 172486
rect 259269 172483 259335 172486
rect 583520 169948 584960 170188
rect -960 164916 480 165156
rect 104893 164250 104959 164253
rect 105077 164250 105143 164253
rect 104893 164248 105143 164250
rect 104893 164192 104898 164248
rect 104954 164192 105082 164248
rect 105138 164192 105143 164248
rect 104893 164190 105143 164192
rect 104893 164187 104959 164190
rect 105077 164187 105143 164190
rect 106457 164250 106523 164253
rect 106641 164250 106707 164253
rect 106457 164248 106707 164250
rect 106457 164192 106462 164248
rect 106518 164192 106646 164248
rect 106702 164192 106707 164248
rect 106457 164190 106707 164192
rect 106457 164187 106523 164190
rect 106641 164187 106707 164190
rect 73337 162890 73403 162893
rect 73613 162890 73679 162893
rect 91185 162890 91251 162893
rect 73337 162888 73679 162890
rect 73337 162832 73342 162888
rect 73398 162832 73618 162888
rect 73674 162832 73679 162888
rect 73337 162830 73679 162832
rect 73337 162827 73403 162830
rect 73613 162827 73679 162830
rect 91142 162888 91251 162890
rect 91142 162832 91190 162888
rect 91246 162832 91251 162888
rect 91142 162827 91251 162832
rect 94129 162890 94195 162893
rect 94313 162890 94379 162893
rect 94129 162888 94379 162890
rect 94129 162832 94134 162888
rect 94190 162832 94318 162888
rect 94374 162832 94379 162888
rect 94129 162830 94379 162832
rect 94129 162827 94195 162830
rect 94313 162827 94379 162830
rect 91142 162621 91202 162827
rect 91093 162616 91202 162621
rect 91093 162560 91098 162616
rect 91154 162560 91202 162616
rect 91093 162558 91202 162560
rect 91093 162555 91159 162558
rect 583520 158252 584960 158492
rect 204805 154730 204871 154733
rect 204805 154728 204914 154730
rect 204805 154672 204810 154728
rect 204866 154672 204914 154728
rect 204805 154667 204914 154672
rect 204854 154597 204914 154667
rect 204854 154592 204963 154597
rect 204854 154536 204902 154592
rect 204958 154536 204963 154592
rect 204854 154534 204963 154536
rect 204897 154531 204963 154534
rect 235533 154594 235599 154597
rect 235717 154594 235783 154597
rect 235533 154592 235783 154594
rect 235533 154536 235538 154592
rect 235594 154536 235722 154592
rect 235778 154536 235783 154592
rect 235533 154534 235783 154536
rect 235533 154531 235599 154534
rect 235717 154531 235783 154534
rect 91093 153234 91159 153237
rect 90958 153232 91159 153234
rect 90958 153176 91098 153232
rect 91154 153176 91159 153232
rect 90958 153174 91159 153176
rect 90958 153098 91018 153174
rect 91093 153171 91159 153174
rect 250805 153234 250871 153237
rect 250989 153234 251055 153237
rect 250805 153232 251055 153234
rect 250805 153176 250810 153232
rect 250866 153176 250994 153232
rect 251050 153176 251055 153232
rect 250805 153174 251055 153176
rect 250805 153171 250871 153174
rect 250989 153171 251055 153174
rect 252093 153234 252159 153237
rect 252277 153234 252343 153237
rect 252093 153232 252343 153234
rect 252093 153176 252098 153232
rect 252154 153176 252282 153232
rect 252338 153176 252343 153232
rect 252093 153174 252343 153176
rect 252093 153171 252159 153174
rect 252277 153171 252343 153174
rect 255221 153234 255287 153237
rect 255405 153234 255471 153237
rect 255221 153232 255471 153234
rect 255221 153176 255226 153232
rect 255282 153176 255410 153232
rect 255466 153176 255471 153232
rect 255221 153174 255471 153176
rect 255221 153171 255287 153174
rect 255405 153171 255471 153174
rect 259085 153234 259151 153237
rect 259269 153234 259335 153237
rect 259085 153232 259335 153234
rect 259085 153176 259090 153232
rect 259146 153176 259274 153232
rect 259330 153176 259335 153232
rect 259085 153174 259335 153176
rect 259085 153171 259151 153174
rect 259269 153171 259335 153174
rect 91185 153098 91251 153101
rect 90958 153096 91251 153098
rect 90958 153040 91190 153096
rect 91246 153040 91251 153096
rect 90958 153038 91251 153040
rect 91185 153035 91251 153038
rect -960 150636 480 150876
rect 583520 146556 584960 146796
rect 324957 144938 325023 144941
rect 325233 144938 325299 144941
rect 324957 144936 325299 144938
rect 324957 144880 324962 144936
rect 325018 144880 325238 144936
rect 325294 144880 325299 144936
rect 324957 144878 325299 144880
rect 324957 144875 325023 144878
rect 325233 144875 325299 144878
rect 255221 143444 255287 143445
rect 255221 143442 255268 143444
rect 255176 143440 255268 143442
rect 255176 143384 255226 143440
rect 255176 143382 255268 143384
rect 255221 143380 255268 143382
rect 255332 143380 255338 143444
rect 255221 143379 255287 143380
rect -960 136220 480 136460
rect 89989 135418 90055 135421
rect 92749 135418 92815 135421
rect 204805 135418 204871 135421
rect 89989 135416 90098 135418
rect 89989 135360 89994 135416
rect 90050 135360 90098 135416
rect 89989 135355 90098 135360
rect 92749 135416 92858 135418
rect 92749 135360 92754 135416
rect 92810 135360 92858 135416
rect 92749 135355 92858 135360
rect 204805 135416 204914 135418
rect 204805 135360 204810 135416
rect 204866 135360 204914 135416
rect 204805 135355 204914 135360
rect 90038 135285 90098 135355
rect 92798 135285 92858 135355
rect 70761 135282 70827 135285
rect 70945 135282 71011 135285
rect 70761 135280 71011 135282
rect 70761 135224 70766 135280
rect 70822 135224 70950 135280
rect 71006 135224 71011 135280
rect 70761 135222 71011 135224
rect 70761 135219 70827 135222
rect 70945 135219 71011 135222
rect 89989 135280 90098 135285
rect 89989 135224 89994 135280
rect 90050 135224 90098 135280
rect 89989 135222 90098 135224
rect 92749 135280 92858 135285
rect 92749 135224 92754 135280
rect 92810 135224 92858 135280
rect 92749 135222 92858 135224
rect 204854 135285 204914 135355
rect 204854 135280 204963 135285
rect 204854 135224 204902 135280
rect 204958 135224 204963 135280
rect 204854 135222 204963 135224
rect 89989 135219 90055 135222
rect 92749 135219 92815 135222
rect 204897 135219 204963 135222
rect 583520 134724 584960 134964
rect 81893 133922 81959 133925
rect 82077 133922 82143 133925
rect 81893 133920 82143 133922
rect 81893 133864 81898 133920
rect 81954 133864 82082 133920
rect 82138 133864 82143 133920
rect 81893 133862 82143 133864
rect 81893 133859 81959 133862
rect 82077 133859 82143 133862
rect 94129 133922 94195 133925
rect 94313 133922 94379 133925
rect 94129 133920 94379 133922
rect 94129 133864 94134 133920
rect 94190 133864 94318 133920
rect 94374 133864 94379 133920
rect 94129 133862 94379 133864
rect 94129 133859 94195 133862
rect 94313 133859 94379 133862
rect 246941 133922 247007 133925
rect 247125 133922 247191 133925
rect 246941 133920 247191 133922
rect 246941 133864 246946 133920
rect 247002 133864 247130 133920
rect 247186 133864 247191 133920
rect 246941 133862 247191 133864
rect 246941 133859 247007 133862
rect 247125 133859 247191 133862
rect 248229 133922 248295 133925
rect 248413 133922 248479 133925
rect 248229 133920 248479 133922
rect 248229 133864 248234 133920
rect 248290 133864 248418 133920
rect 248474 133864 248479 133920
rect 248229 133862 248479 133864
rect 248229 133859 248295 133862
rect 248413 133859 248479 133862
rect 249425 133922 249491 133925
rect 249609 133922 249675 133925
rect 249425 133920 249675 133922
rect 249425 133864 249430 133920
rect 249486 133864 249614 133920
rect 249670 133864 249675 133920
rect 249425 133862 249675 133864
rect 249425 133859 249491 133862
rect 249609 133859 249675 133862
rect 250989 133922 251055 133925
rect 251173 133922 251239 133925
rect 250989 133920 251239 133922
rect 250989 133864 250994 133920
rect 251050 133864 251178 133920
rect 251234 133864 251239 133920
rect 250989 133862 251239 133864
rect 250989 133859 251055 133862
rect 251173 133859 251239 133862
rect 252093 133922 252159 133925
rect 252277 133922 252343 133925
rect 252093 133920 252343 133922
rect 252093 133864 252098 133920
rect 252154 133864 252282 133920
rect 252338 133864 252343 133920
rect 252093 133862 252343 133864
rect 252093 133859 252159 133862
rect 252277 133859 252343 133862
rect 255262 133860 255268 133924
rect 255332 133922 255338 133924
rect 255405 133922 255471 133925
rect 255332 133920 255471 133922
rect 255332 133864 255410 133920
rect 255466 133864 255471 133920
rect 255332 133862 255471 133864
rect 255332 133860 255338 133862
rect 255405 133859 255471 133862
rect 264789 133922 264855 133925
rect 264973 133922 265039 133925
rect 264789 133920 265039 133922
rect 264789 133864 264794 133920
rect 264850 133864 264978 133920
rect 265034 133864 265039 133920
rect 264789 133862 265039 133864
rect 264789 133859 264855 133862
rect 264973 133859 265039 133862
rect 77477 125626 77543 125629
rect 77661 125626 77727 125629
rect 77477 125624 77727 125626
rect 77477 125568 77482 125624
rect 77538 125568 77666 125624
rect 77722 125568 77727 125624
rect 77477 125566 77727 125568
rect 77477 125563 77543 125566
rect 77661 125563 77727 125566
rect 78765 125626 78831 125629
rect 78949 125626 79015 125629
rect 78765 125624 79015 125626
rect 78765 125568 78770 125624
rect 78826 125568 78954 125624
rect 79010 125568 79015 125624
rect 78765 125566 79015 125568
rect 78765 125563 78831 125566
rect 78949 125563 79015 125566
rect 81709 125626 81775 125629
rect 81893 125626 81959 125629
rect 81709 125624 81959 125626
rect 81709 125568 81714 125624
rect 81770 125568 81898 125624
rect 81954 125568 81959 125624
rect 81709 125566 81959 125568
rect 81709 125563 81775 125566
rect 81893 125563 81959 125566
rect 255221 125626 255287 125629
rect 255405 125626 255471 125629
rect 255221 125624 255471 125626
rect 255221 125568 255226 125624
rect 255282 125568 255410 125624
rect 255466 125568 255471 125624
rect 255221 125566 255471 125568
rect 255221 125563 255287 125566
rect 255405 125563 255471 125566
rect 259085 125626 259151 125629
rect 259269 125626 259335 125629
rect 259085 125624 259335 125626
rect 259085 125568 259090 125624
rect 259146 125568 259274 125624
rect 259330 125568 259335 125624
rect 259085 125566 259335 125568
rect 259085 125563 259151 125566
rect 259269 125563 259335 125566
rect 324957 125626 325023 125629
rect 325233 125626 325299 125629
rect 324957 125624 325299 125626
rect 324957 125568 324962 125624
rect 325018 125568 325238 125624
rect 325294 125568 325299 125624
rect 324957 125566 325299 125568
rect 324957 125563 325023 125566
rect 325233 125563 325299 125566
rect 583520 123028 584960 123268
rect -960 121940 480 122180
rect 89989 115970 90055 115973
rect 90173 115970 90239 115973
rect 89989 115968 90239 115970
rect 89989 115912 89994 115968
rect 90050 115912 90178 115968
rect 90234 115912 90239 115968
rect 89989 115910 90239 115912
rect 89989 115907 90055 115910
rect 90173 115907 90239 115910
rect 92749 115970 92815 115973
rect 92933 115970 92999 115973
rect 92749 115968 92999 115970
rect 92749 115912 92754 115968
rect 92810 115912 92938 115968
rect 92994 115912 92999 115968
rect 92749 115910 92999 115912
rect 92749 115907 92815 115910
rect 92933 115907 92999 115910
rect 91001 114610 91067 114613
rect 91185 114610 91251 114613
rect 91001 114608 91251 114610
rect 91001 114552 91006 114608
rect 91062 114552 91190 114608
rect 91246 114552 91251 114608
rect 91001 114550 91251 114552
rect 91001 114547 91067 114550
rect 91185 114547 91251 114550
rect 583520 111332 584960 111572
rect -960 107524 480 107764
rect 94129 106586 94195 106589
rect 93902 106584 94195 106586
rect 93902 106528 94134 106584
rect 94190 106528 94195 106584
rect 93902 106526 94195 106528
rect 93902 106314 93962 106526
rect 94129 106523 94195 106526
rect 94037 106314 94103 106317
rect 93902 106312 94103 106314
rect 93902 106256 94042 106312
rect 94098 106256 94103 106312
rect 93902 106254 94103 106256
rect 94037 106251 94103 106254
rect 259085 106314 259151 106317
rect 259269 106314 259335 106317
rect 259085 106312 259335 106314
rect 259085 106256 259090 106312
rect 259146 106256 259274 106312
rect 259330 106256 259335 106312
rect 259085 106254 259335 106256
rect 259085 106251 259151 106254
rect 259269 106251 259335 106254
rect 324957 106314 325023 106317
rect 325233 106314 325299 106317
rect 324957 106312 325299 106314
rect 324957 106256 324962 106312
rect 325018 106256 325238 106312
rect 325294 106256 325299 106312
rect 324957 106254 325299 106256
rect 324957 106251 325023 106254
rect 325233 106251 325299 106254
rect 583520 99636 584960 99876
rect 89989 96658 90055 96661
rect 90173 96658 90239 96661
rect 89989 96656 90239 96658
rect 89989 96600 89994 96656
rect 90050 96600 90178 96656
rect 90234 96600 90239 96656
rect 89989 96598 90239 96600
rect 89989 96595 90055 96598
rect 90173 96595 90239 96598
rect 92749 96658 92815 96661
rect 92933 96658 92999 96661
rect 92749 96656 92999 96658
rect 92749 96600 92754 96656
rect 92810 96600 92938 96656
rect 92994 96600 92999 96656
rect 92749 96598 92999 96600
rect 92749 96595 92815 96598
rect 92933 96595 92999 96598
rect -960 93108 480 93348
rect 583520 87804 584960 88044
rect 72233 87138 72299 87141
rect 77569 87138 77635 87141
rect 81801 87138 81867 87141
rect 72190 87136 72299 87138
rect 72190 87080 72238 87136
rect 72294 87080 72299 87136
rect 72190 87075 72299 87080
rect 77526 87136 77635 87138
rect 77526 87080 77574 87136
rect 77630 87080 77635 87136
rect 77526 87075 77635 87080
rect 81758 87136 81867 87138
rect 81758 87080 81806 87136
rect 81862 87080 81867 87136
rect 81758 87075 81867 87080
rect 94037 87138 94103 87141
rect 94037 87136 94146 87138
rect 94037 87080 94042 87136
rect 94098 87080 94146 87136
rect 94037 87075 94146 87080
rect 72190 87005 72250 87075
rect 77526 87005 77586 87075
rect 81758 87005 81818 87075
rect 94086 87005 94146 87075
rect 72141 87000 72250 87005
rect 72141 86944 72146 87000
rect 72202 86944 72250 87000
rect 72141 86942 72250 86944
rect 73429 87002 73495 87005
rect 73613 87002 73679 87005
rect 73429 87000 73679 87002
rect 73429 86944 73434 87000
rect 73490 86944 73618 87000
rect 73674 86944 73679 87000
rect 73429 86942 73679 86944
rect 72141 86939 72207 86942
rect 73429 86939 73495 86942
rect 73613 86939 73679 86942
rect 77477 87000 77586 87005
rect 77477 86944 77482 87000
rect 77538 86944 77586 87000
rect 77477 86942 77586 86944
rect 81709 87000 81818 87005
rect 81709 86944 81714 87000
rect 81770 86944 81818 87000
rect 81709 86942 81818 86944
rect 94037 87000 94146 87005
rect 94037 86944 94042 87000
rect 94098 86944 94146 87000
rect 94037 86942 94146 86944
rect 252093 87002 252159 87005
rect 252277 87002 252343 87005
rect 252093 87000 252343 87002
rect 252093 86944 252098 87000
rect 252154 86944 252282 87000
rect 252338 86944 252343 87000
rect 252093 86942 252343 86944
rect 77477 86939 77543 86942
rect 81709 86939 81775 86942
rect 94037 86939 94103 86942
rect 252093 86939 252159 86942
rect 252277 86939 252343 86942
rect 91001 85506 91067 85509
rect 91001 85504 91202 85506
rect 91001 85448 91006 85504
rect 91062 85448 91202 85504
rect 91001 85446 91202 85448
rect 91001 85443 91067 85446
rect 91142 85373 91202 85446
rect 91093 85368 91202 85373
rect 91093 85312 91098 85368
rect 91154 85312 91202 85368
rect 91093 85310 91202 85312
rect 91093 85307 91159 85310
rect -960 78828 480 79068
rect 70761 77346 70827 77349
rect 70945 77346 71011 77349
rect 70761 77344 71011 77346
rect 70761 77288 70766 77344
rect 70822 77288 70950 77344
rect 71006 77288 71011 77344
rect 70761 77286 71011 77288
rect 70761 77283 70827 77286
rect 70945 77283 71011 77286
rect 583520 76108 584960 76348
rect 81801 66330 81867 66333
rect 81574 66328 81867 66330
rect 81574 66272 81806 66328
rect 81862 66272 81867 66328
rect 81574 66270 81867 66272
rect 81574 66058 81634 66270
rect 81801 66267 81867 66270
rect 81801 66058 81867 66061
rect 81574 66056 81867 66058
rect 81574 66000 81806 66056
rect 81862 66000 81867 66056
rect 81574 65998 81867 66000
rect 81801 65995 81867 65998
rect -960 64412 480 64652
rect 583520 64412 584960 64652
rect 96981 60756 97047 60757
rect 96981 60752 97028 60756
rect 97092 60754 97098 60756
rect 96981 60696 96986 60752
rect 96981 60692 97028 60696
rect 97092 60694 97138 60754
rect 97092 60692 97098 60694
rect 96981 60691 97047 60692
rect 96981 56676 97047 56677
rect 96981 56672 97028 56676
rect 97092 56674 97098 56676
rect 96981 56616 96986 56672
rect 96981 56612 97028 56616
rect 97092 56614 97138 56674
rect 97092 56612 97098 56614
rect 96981 56611 97047 56612
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 243629 46882 243695 46885
rect 243813 46882 243879 46885
rect 243629 46880 243879 46882
rect 243629 46824 243634 46880
rect 243690 46824 243818 46880
rect 243874 46824 243879 46880
rect 243629 46822 243879 46824
rect 243629 46819 243695 46822
rect 243813 46819 243879 46822
rect 583520 40884 584960 41124
rect -960 35716 480 35956
rect 583520 29188 584960 29428
rect 227294 22068 227300 22132
rect 227364 22130 227370 22132
rect 227437 22130 227503 22133
rect 227364 22128 227503 22130
rect 227364 22072 227442 22128
rect 227498 22072 227503 22128
rect 227364 22070 227503 22072
rect 227364 22068 227370 22070
rect 227437 22067 227503 22070
rect -960 21300 480 21540
rect 227345 19412 227411 19413
rect 227294 19348 227300 19412
rect 227364 19410 227411 19412
rect 227364 19408 227456 19410
rect 227406 19352 227456 19408
rect 227364 19350 227456 19352
rect 227364 19348 227411 19350
rect 227345 19347 227411 19348
rect 583520 17492 584960 17732
rect 239857 15194 239923 15197
rect 256693 15194 256759 15197
rect 239857 15192 256759 15194
rect 239857 15136 239862 15192
rect 239918 15136 256698 15192
rect 256754 15136 256759 15192
rect 239857 15134 256759 15136
rect 239857 15131 239923 15134
rect 256693 15131 256759 15134
rect 264697 15192 264763 15197
rect 264697 15136 264702 15192
rect 264758 15136 264763 15192
rect 264697 15131 264763 15136
rect 266256 15132 266262 15196
rect 266326 15194 266332 15196
rect 489913 15194 489979 15197
rect 266326 15192 489979 15194
rect 266326 15136 489918 15192
rect 489974 15136 489979 15192
rect 266326 15134 489979 15136
rect 266326 15132 266332 15134
rect 489913 15131 489979 15134
rect 264700 15058 264760 15131
rect 265157 15058 265223 15061
rect 264700 15056 265223 15058
rect 264700 15000 265162 15056
rect 265218 15000 265223 15056
rect 264700 14998 265223 15000
rect 265157 14995 265223 14998
rect 268837 15058 268903 15061
rect 571333 15058 571399 15061
rect 268837 15056 571399 15058
rect 268837 15000 268842 15056
rect 268898 15000 571338 15056
rect 571394 15000 571399 15056
rect 268837 14998 571399 15000
rect 268837 14995 268903 14998
rect 571333 14995 571399 14998
rect 270309 14922 270375 14925
rect 574093 14922 574159 14925
rect 270309 14920 574159 14922
rect 270309 14864 270314 14920
rect 270370 14864 574098 14920
rect 574154 14864 574159 14920
rect 270309 14862 574159 14864
rect 270309 14859 270375 14862
rect 574093 14859 574159 14862
rect 256693 14786 256759 14789
rect 266256 14786 266262 14788
rect 256693 14784 266262 14786
rect 256693 14728 256698 14784
rect 256754 14728 266262 14784
rect 256693 14726 266262 14728
rect 256693 14723 256759 14726
rect 266256 14724 266262 14726
rect 266326 14724 266332 14788
rect 270217 14786 270283 14789
rect 576853 14786 576919 14789
rect 270217 14784 576919 14786
rect 270217 14728 270222 14784
rect 270278 14728 576858 14784
rect 576914 14728 576919 14784
rect 270217 14726 576919 14728
rect 270217 14723 270283 14726
rect 576853 14723 576919 14726
rect 271505 14650 271571 14653
rect 578233 14650 578299 14653
rect 271505 14648 578299 14650
rect 271505 14592 271510 14648
rect 271566 14592 578238 14648
rect 578294 14592 578299 14648
rect 271505 14590 578299 14592
rect 271505 14587 271571 14590
rect 578233 14587 578299 14590
rect 271597 14514 271663 14517
rect 580993 14514 581059 14517
rect 271597 14512 581059 14514
rect 271597 14456 271602 14512
rect 271658 14456 580998 14512
rect 581054 14456 581059 14512
rect 271597 14454 581059 14456
rect 271597 14451 271663 14454
rect 580993 14451 581059 14454
rect 262213 13834 262279 13837
rect 262397 13834 262463 13837
rect 262213 13832 262463 13834
rect 262213 13776 262218 13832
rect 262274 13776 262402 13832
rect 262458 13776 262463 13832
rect 262213 13774 262463 13776
rect 262213 13771 262279 13774
rect 262397 13771 262463 13774
rect 260557 13698 260623 13701
rect 549253 13698 549319 13701
rect 260557 13696 549319 13698
rect 260557 13640 260562 13696
rect 260618 13640 549258 13696
rect 549314 13640 549319 13696
rect 260557 13638 549319 13640
rect 260557 13635 260623 13638
rect 549253 13635 549319 13638
rect 261937 13562 262003 13565
rect 553393 13562 553459 13565
rect 261937 13560 553459 13562
rect 261937 13504 261942 13560
rect 261998 13504 553398 13560
rect 553454 13504 553459 13560
rect 261937 13502 553459 13504
rect 261937 13499 262003 13502
rect 553393 13499 553459 13502
rect 263225 13426 263291 13429
rect 556153 13426 556219 13429
rect 263225 13424 556219 13426
rect 263225 13368 263230 13424
rect 263286 13368 556158 13424
rect 556214 13368 556219 13424
rect 263225 13366 556219 13368
rect 263225 13363 263291 13366
rect 556153 13363 556219 13366
rect 265157 13290 265223 13293
rect 560293 13290 560359 13293
rect 265157 13288 560359 13290
rect 265157 13232 265162 13288
rect 265218 13232 560298 13288
rect 560354 13232 560359 13288
rect 265157 13230 560359 13232
rect 265157 13227 265223 13230
rect 560293 13227 560359 13230
rect 266077 13154 266143 13157
rect 563053 13154 563119 13157
rect 266077 13152 563119 13154
rect 266077 13096 266082 13152
rect 266138 13096 563058 13152
rect 563114 13096 563119 13152
rect 266077 13094 563119 13096
rect 266077 13091 266143 13094
rect 563053 13091 563119 13094
rect 267365 13018 267431 13021
rect 567193 13018 567259 13021
rect 267365 13016 567259 13018
rect 267365 12960 267370 13016
rect 267426 12960 567198 13016
rect 567254 12960 567259 13016
rect 267365 12958 567259 12960
rect 267365 12955 267431 12958
rect 567193 12955 567259 12958
rect 231485 12338 231551 12341
rect 462313 12338 462379 12341
rect 231485 12336 462379 12338
rect 231485 12280 231490 12336
rect 231546 12280 462318 12336
rect 462374 12280 462379 12336
rect 231485 12278 462379 12280
rect 231485 12275 231551 12278
rect 462313 12275 462379 12278
rect 231577 12202 231643 12205
rect 466453 12202 466519 12205
rect 231577 12200 466519 12202
rect 231577 12144 231582 12200
rect 231638 12144 466458 12200
rect 466514 12144 466519 12200
rect 231577 12142 466519 12144
rect 231577 12139 231643 12142
rect 466453 12139 466519 12142
rect 233049 12066 233115 12069
rect 469213 12066 469279 12069
rect 233049 12064 469279 12066
rect 233049 12008 233054 12064
rect 233110 12008 469218 12064
rect 469274 12008 469279 12064
rect 233049 12006 469279 12008
rect 233049 12003 233115 12006
rect 469213 12003 469279 12006
rect 234613 11930 234679 11933
rect 473353 11930 473419 11933
rect 234613 11928 473419 11930
rect 234613 11872 234618 11928
rect 234674 11872 473358 11928
rect 473414 11872 473419 11928
rect 234613 11870 473419 11872
rect 234613 11867 234679 11870
rect 473353 11867 473419 11870
rect 235809 11794 235875 11797
rect 477585 11794 477651 11797
rect 235809 11792 477651 11794
rect 235809 11736 235814 11792
rect 235870 11736 477590 11792
rect 477646 11736 477651 11792
rect 235809 11734 477651 11736
rect 235809 11731 235875 11734
rect 477585 11731 477651 11734
rect 237281 11658 237347 11661
rect 480253 11658 480319 11661
rect 237281 11656 480319 11658
rect 237281 11600 237286 11656
rect 237342 11600 480258 11656
rect 480314 11600 480319 11656
rect 237281 11598 480319 11600
rect 237281 11595 237347 11598
rect 480253 11595 480319 11598
rect 195697 10842 195763 10845
rect 362953 10842 363019 10845
rect 195697 10840 363019 10842
rect 195697 10784 195702 10840
rect 195758 10784 362958 10840
rect 363014 10784 363019 10840
rect 195697 10782 363019 10784
rect 195697 10779 195763 10782
rect 362953 10779 363019 10782
rect 197077 10706 197143 10709
rect 365713 10706 365779 10709
rect 197077 10704 365779 10706
rect 197077 10648 197082 10704
rect 197138 10648 365718 10704
rect 365774 10648 365779 10704
rect 197077 10646 365779 10648
rect 197077 10643 197143 10646
rect 365713 10643 365779 10646
rect 198549 10570 198615 10573
rect 369853 10570 369919 10573
rect 198549 10568 369919 10570
rect 198549 10512 198554 10568
rect 198610 10512 369858 10568
rect 369914 10512 369919 10568
rect 198549 10510 369919 10512
rect 198549 10507 198615 10510
rect 369853 10507 369919 10510
rect 199837 10434 199903 10437
rect 374085 10434 374151 10437
rect 199837 10432 374151 10434
rect 199837 10376 199842 10432
rect 199898 10376 374090 10432
rect 374146 10376 374151 10432
rect 199837 10374 374151 10376
rect 199837 10371 199903 10374
rect 374085 10371 374151 10374
rect 201309 10298 201375 10301
rect 376753 10298 376819 10301
rect 201309 10296 376819 10298
rect 201309 10240 201314 10296
rect 201370 10240 376758 10296
rect 376814 10240 376819 10296
rect 201309 10238 376819 10240
rect 201309 10235 201375 10238
rect 376753 10235 376819 10238
rect 246941 9890 247007 9893
rect 246806 9888 247007 9890
rect 246806 9832 246946 9888
rect 247002 9832 247007 9888
rect 246806 9830 247007 9832
rect 151077 9652 151143 9655
rect 150942 9650 151143 9652
rect 150942 9594 151082 9650
rect 151138 9594 151143 9650
rect 150942 9592 151143 9594
rect 150942 9482 151002 9592
rect 151077 9589 151143 9592
rect 153193 9482 153259 9485
rect 150942 9480 153259 9482
rect 150942 9424 153198 9480
rect 153254 9424 153259 9480
rect 150942 9422 153259 9424
rect 246806 9482 246866 9830
rect 246941 9827 247007 9830
rect 259177 9618 259243 9621
rect 545297 9618 545363 9621
rect 259177 9616 545363 9618
rect 259177 9560 259182 9616
rect 259238 9560 545302 9616
rect 545358 9560 545363 9616
rect 259177 9558 545363 9560
rect 259177 9555 259243 9558
rect 545297 9555 545363 9558
rect 249241 9482 249307 9485
rect 246806 9480 249307 9482
rect 246806 9424 249246 9480
rect 249302 9424 249307 9480
rect 246806 9422 249307 9424
rect 153193 9419 153259 9422
rect 249241 9419 249307 9422
rect 262397 9482 262463 9485
rect 552381 9482 552447 9485
rect 262397 9480 552447 9482
rect 262397 9424 262402 9480
rect 262458 9424 552386 9480
rect 552442 9424 552447 9480
rect 262397 9422 552447 9424
rect 262397 9419 262463 9422
rect 552381 9419 552447 9422
rect 263225 9346 263291 9349
rect 555969 9346 556035 9349
rect 263225 9344 556035 9346
rect 263225 9288 263230 9344
rect 263286 9288 555974 9344
rect 556030 9288 556035 9344
rect 263225 9286 556035 9288
rect 263225 9283 263291 9286
rect 555969 9283 556035 9286
rect 244089 9210 244155 9213
rect 249333 9210 249399 9213
rect 244089 9208 249399 9210
rect 244089 9152 244094 9208
rect 244150 9152 249338 9208
rect 249394 9152 249399 9208
rect 244089 9150 249399 9152
rect 244089 9147 244155 9150
rect 249333 9147 249399 9150
rect 264789 9210 264855 9213
rect 559557 9210 559623 9213
rect 264789 9208 559623 9210
rect 264789 9152 264794 9208
rect 264850 9152 559562 9208
rect 559618 9152 559623 9208
rect 264789 9150 559623 9152
rect 264789 9147 264855 9150
rect 559557 9147 559623 9150
rect 266169 9074 266235 9077
rect 563145 9074 563211 9077
rect 266169 9072 563211 9074
rect 266169 9016 266174 9072
rect 266230 9016 563150 9072
rect 563206 9016 563211 9072
rect 266169 9014 563211 9016
rect 266169 9011 266235 9014
rect 563145 9011 563211 9014
rect 268929 8938 268995 8941
rect 573817 8938 573883 8941
rect 268929 8936 573883 8938
rect 268929 8880 268934 8936
rect 268990 8880 573822 8936
rect 573878 8880 573883 8936
rect 268929 8878 573883 8880
rect 268929 8875 268995 8878
rect 573817 8875 573883 8878
rect 205633 8802 205699 8805
rect 215109 8802 215175 8805
rect 205633 8800 215175 8802
rect 205633 8744 205638 8800
rect 205694 8744 215114 8800
rect 215170 8744 215175 8800
rect 205633 8742 215175 8744
rect 205633 8739 205699 8742
rect 215109 8739 215175 8742
rect 224953 8802 225019 8805
rect 239581 8802 239647 8805
rect 224953 8800 239647 8802
rect 224953 8744 224958 8800
rect 225014 8744 239586 8800
rect 239642 8744 239647 8800
rect 224953 8742 239647 8744
rect 224953 8739 225019 8742
rect 239581 8739 239647 8742
rect 248137 8666 248203 8669
rect 249793 8666 249859 8669
rect 248137 8664 249859 8666
rect 248137 8608 248142 8664
rect 248198 8608 249798 8664
rect 249854 8608 249859 8664
rect 248137 8606 249859 8608
rect 248137 8603 248203 8606
rect 249793 8603 249859 8606
rect 234429 8394 234495 8397
rect 239765 8394 239831 8397
rect 234429 8392 239831 8394
rect 234429 8336 234434 8392
rect 234490 8336 239770 8392
rect 239826 8336 239831 8392
rect 234429 8334 239831 8336
rect 234429 8331 234495 8334
rect 239765 8331 239831 8334
rect 228909 8258 228975 8261
rect 458449 8258 458515 8261
rect 228909 8256 458515 8258
rect 228909 8200 228914 8256
rect 228970 8200 458454 8256
rect 458510 8200 458515 8256
rect 228909 8198 458515 8200
rect 228909 8195 228975 8198
rect 458449 8195 458515 8198
rect 230381 8122 230447 8125
rect 462037 8122 462103 8125
rect 230381 8120 462103 8122
rect 230381 8064 230386 8120
rect 230442 8064 462042 8120
rect 462098 8064 462103 8120
rect 230381 8062 462103 8064
rect 230381 8059 230447 8062
rect 462037 8059 462103 8062
rect 231669 7986 231735 7989
rect 465625 7986 465691 7989
rect 231669 7984 465691 7986
rect 231669 7928 231674 7984
rect 231730 7928 465630 7984
rect 465686 7928 465691 7984
rect 231669 7926 465691 7928
rect 231669 7923 231735 7926
rect 465625 7923 465691 7926
rect 233141 7850 233207 7853
rect 469121 7850 469187 7853
rect 233141 7848 469187 7850
rect 233141 7792 233146 7848
rect 233202 7792 469126 7848
rect 469182 7792 469187 7848
rect 233141 7790 469187 7792
rect 233141 7787 233207 7790
rect 469121 7787 469187 7790
rect 234337 7714 234403 7717
rect 472709 7714 472775 7717
rect 234337 7712 472775 7714
rect 234337 7656 234342 7712
rect 234398 7656 472714 7712
rect 472770 7656 472775 7712
rect 234337 7654 472775 7656
rect 234337 7651 234403 7654
rect 472709 7651 472775 7654
rect 235901 7578 235967 7581
rect 476297 7578 476363 7581
rect 235901 7576 476363 7578
rect 235901 7520 235906 7576
rect 235962 7520 476302 7576
rect 476358 7520 476363 7576
rect 235901 7518 476363 7520
rect 235901 7515 235967 7518
rect 476297 7515 476363 7518
rect -960 7020 480 7260
rect 194409 6762 194475 6765
rect 358537 6762 358603 6765
rect 194409 6760 358603 6762
rect 194409 6704 194414 6760
rect 194470 6704 358542 6760
rect 358598 6704 358603 6760
rect 194409 6702 358603 6704
rect 194409 6699 194475 6702
rect 358537 6699 358603 6702
rect 195881 6626 195947 6629
rect 362125 6626 362191 6629
rect 195881 6624 362191 6626
rect 195881 6568 195886 6624
rect 195942 6568 362130 6624
rect 362186 6568 362191 6624
rect 195881 6566 362191 6568
rect 195881 6563 195947 6566
rect 362125 6563 362191 6566
rect 197261 6490 197327 6493
rect 365805 6490 365871 6493
rect 197261 6488 365871 6490
rect 197261 6432 197266 6488
rect 197322 6432 365810 6488
rect 365866 6432 365871 6488
rect 197261 6430 365871 6432
rect 197261 6427 197327 6430
rect 365805 6427 365871 6430
rect 198641 6354 198707 6357
rect 369209 6354 369275 6357
rect 198641 6352 369275 6354
rect 198641 6296 198646 6352
rect 198702 6296 369214 6352
rect 369270 6296 369275 6352
rect 198641 6294 369275 6296
rect 198641 6291 198707 6294
rect 369209 6291 369275 6294
rect 199929 6218 199995 6221
rect 372797 6218 372863 6221
rect 199929 6216 372863 6218
rect 199929 6160 199934 6216
rect 199990 6160 372802 6216
rect 372858 6160 372863 6216
rect 199929 6158 372863 6160
rect 199929 6155 199995 6158
rect 372797 6155 372863 6158
rect 583520 5796 584960 6036
rect 166901 5538 166967 5541
rect 276473 5538 276539 5541
rect 166901 5536 276539 5538
rect 166901 5480 166906 5536
rect 166962 5480 276478 5536
rect 276534 5480 276539 5536
rect 166901 5478 276539 5480
rect 166901 5475 166967 5478
rect 276473 5475 276539 5478
rect 158621 5402 158687 5405
rect 255037 5402 255103 5405
rect 158621 5400 255103 5402
rect 158621 5344 158626 5400
rect 158682 5344 255042 5400
rect 255098 5344 255103 5400
rect 158621 5342 255103 5344
rect 158621 5339 158687 5342
rect 255037 5339 255103 5342
rect 263501 5402 263567 5405
rect 554773 5402 554839 5405
rect 263501 5400 554839 5402
rect 263501 5344 263506 5400
rect 263562 5344 554778 5400
rect 554834 5344 554839 5400
rect 263501 5342 554839 5344
rect 263501 5339 263567 5342
rect 554773 5339 554839 5342
rect 160001 5266 160067 5269
rect 258625 5266 258691 5269
rect 160001 5264 258691 5266
rect 160001 5208 160006 5264
rect 160062 5208 258630 5264
rect 258686 5208 258691 5264
rect 160001 5206 258691 5208
rect 160001 5203 160067 5206
rect 258625 5203 258691 5206
rect 263225 5266 263291 5269
rect 558361 5266 558427 5269
rect 263225 5264 558427 5266
rect 263225 5208 263230 5264
rect 263286 5208 558366 5264
rect 558422 5208 558427 5264
rect 263225 5206 558427 5208
rect 263225 5203 263291 5206
rect 558361 5203 558427 5206
rect 161381 5130 161447 5133
rect 262213 5130 262279 5133
rect 161381 5128 262279 5130
rect 161381 5072 161386 5128
rect 161442 5072 262218 5128
rect 262274 5072 262279 5128
rect 161381 5070 262279 5072
rect 161381 5067 161447 5070
rect 262213 5067 262279 5070
rect 266261 5130 266327 5133
rect 565537 5130 565603 5133
rect 266261 5128 565603 5130
rect 266261 5072 266266 5128
rect 266322 5072 565542 5128
rect 565598 5072 565603 5128
rect 266261 5070 565603 5072
rect 266261 5067 266327 5070
rect 565537 5067 565603 5070
rect 162761 4994 162827 4997
rect 265801 4994 265867 4997
rect 162761 4992 265867 4994
rect 162761 4936 162766 4992
rect 162822 4936 265806 4992
rect 265862 4936 265867 4992
rect 162761 4934 265867 4936
rect 162761 4931 162827 4934
rect 265801 4931 265867 4934
rect 267641 4994 267707 4997
rect 569033 4994 569099 4997
rect 267641 4992 569099 4994
rect 267641 4936 267646 4992
rect 267702 4936 569038 4992
rect 569094 4936 569099 4992
rect 267641 4934 569099 4936
rect 267641 4931 267707 4934
rect 569033 4931 569099 4934
rect 164141 4858 164207 4861
rect 269297 4858 269363 4861
rect 164141 4856 269363 4858
rect 164141 4800 164146 4856
rect 164202 4800 269302 4856
rect 269358 4800 269363 4856
rect 164141 4798 269363 4800
rect 164141 4795 164207 4798
rect 269297 4795 269363 4798
rect 270401 4858 270467 4861
rect 576209 4858 576275 4861
rect 270401 4856 576275 4858
rect 270401 4800 270406 4856
rect 270462 4800 576214 4856
rect 576270 4800 576275 4856
rect 270401 4798 576275 4800
rect 270401 4795 270467 4798
rect 576209 4795 576275 4798
rect 215109 4722 215175 4725
rect 215569 4722 215635 4725
rect 215109 4720 215635 4722
rect 215109 4664 215114 4720
rect 215170 4664 215574 4720
rect 215630 4664 215635 4720
rect 215109 4662 215635 4664
rect 215109 4659 215175 4662
rect 215569 4659 215635 4662
rect 244181 4586 244247 4589
rect 249057 4586 249123 4589
rect 244181 4584 249123 4586
rect 244181 4528 244186 4584
rect 244242 4528 249062 4584
rect 249118 4528 249123 4584
rect 244181 4526 249123 4528
rect 244181 4523 244247 4526
rect 249057 4523 249123 4526
rect 215109 4450 215175 4453
rect 215293 4450 215359 4453
rect 215109 4448 215359 4450
rect 215109 4392 215114 4448
rect 215170 4392 215298 4448
rect 215354 4392 215359 4448
rect 215109 4390 215359 4392
rect 215109 4387 215175 4390
rect 215293 4387 215359 4390
rect 345013 4178 345079 4181
rect 354581 4178 354647 4181
rect 345013 4176 354647 4178
rect 345013 4120 345018 4176
rect 345074 4120 354586 4176
rect 354642 4120 354647 4176
rect 345013 4118 354647 4120
rect 345013 4115 345079 4118
rect 354581 4115 354647 4118
rect 42149 4042 42215 4045
rect 84285 4042 84351 4045
rect 42149 4040 84351 4042
rect 42149 3984 42154 4040
rect 42210 3984 84290 4040
rect 84346 3984 84351 4040
rect 42149 3982 84351 3984
rect 42149 3979 42215 3982
rect 84285 3979 84351 3982
rect 129549 4042 129615 4045
rect 171777 4042 171843 4045
rect 129549 4040 171843 4042
rect 129549 3984 129554 4040
rect 129610 3984 171782 4040
rect 171838 3984 171843 4040
rect 129549 3982 171843 3984
rect 129549 3979 129615 3982
rect 171777 3979 171843 3982
rect 364885 4042 364951 4045
rect 367001 4042 367067 4045
rect 364885 4040 367067 4042
rect 364885 3984 364890 4040
rect 364946 3984 367006 4040
rect 367062 3984 367067 4040
rect 364885 3982 367067 3984
rect 364885 3979 364951 3982
rect 367001 3979 367067 3982
rect 373257 4042 373323 4045
rect 475101 4042 475167 4045
rect 373257 4040 475167 4042
rect 373257 3984 373262 4040
rect 373318 3984 475106 4040
rect 475162 3984 475167 4040
rect 373257 3982 475167 3984
rect 373257 3979 373323 3982
rect 475101 3979 475167 3982
rect 29085 3906 29151 3909
rect 80145 3906 80211 3909
rect 29085 3904 80211 3906
rect 29085 3848 29090 3904
rect 29146 3848 80150 3904
rect 80206 3848 80211 3904
rect 29085 3846 80211 3848
rect 29085 3843 29151 3846
rect 80145 3843 80211 3846
rect 130929 3906 130995 3909
rect 175365 3906 175431 3909
rect 130929 3904 175431 3906
rect 130929 3848 130934 3904
rect 130990 3848 175370 3904
rect 175426 3848 175431 3904
rect 130929 3846 175431 3848
rect 130929 3843 130995 3846
rect 175365 3843 175431 3846
rect 224861 3906 224927 3909
rect 442993 3906 443059 3909
rect 224861 3904 443059 3906
rect 224861 3848 224866 3904
rect 224922 3848 442998 3904
rect 443054 3848 443059 3904
rect 224861 3846 443059 3848
rect 224861 3843 224927 3846
rect 442993 3843 443059 3846
rect 19517 3770 19583 3773
rect 75913 3770 75979 3773
rect 19517 3768 75979 3770
rect 19517 3712 19522 3768
rect 19578 3712 75918 3768
rect 75974 3712 75979 3768
rect 19517 3710 75979 3712
rect 19517 3707 19583 3710
rect 75913 3707 75979 3710
rect 132309 3770 132375 3773
rect 178953 3770 179019 3773
rect 132309 3768 179019 3770
rect 132309 3712 132314 3768
rect 132370 3712 178958 3768
rect 179014 3712 179019 3768
rect 132309 3710 179019 3712
rect 132309 3707 132375 3710
rect 178953 3707 179019 3710
rect 226241 3770 226307 3773
rect 450169 3770 450235 3773
rect 226241 3768 450235 3770
rect 226241 3712 226246 3768
rect 226302 3712 450174 3768
rect 450230 3712 450235 3768
rect 226241 3710 450235 3712
rect 226241 3707 226307 3710
rect 450169 3707 450235 3710
rect 18321 3634 18387 3637
rect 76097 3634 76163 3637
rect 18321 3632 76163 3634
rect 18321 3576 18326 3632
rect 18382 3576 76102 3632
rect 76158 3576 76163 3632
rect 18321 3574 76163 3576
rect 18321 3571 18387 3574
rect 76097 3571 76163 3574
rect 158069 3634 158135 3637
rect 207473 3634 207539 3637
rect 158069 3632 207539 3634
rect 158069 3576 158074 3632
rect 158130 3576 207478 3632
rect 207534 3576 207539 3632
rect 158069 3574 207539 3576
rect 158069 3571 158135 3574
rect 207473 3571 207539 3574
rect 229001 3634 229067 3637
rect 457253 3634 457319 3637
rect 229001 3632 457319 3634
rect 229001 3576 229006 3632
rect 229062 3576 457258 3632
rect 457314 3576 457319 3632
rect 229001 3574 457319 3576
rect 229001 3571 229067 3574
rect 457253 3571 457319 3574
rect 10041 3498 10107 3501
rect 73337 3498 73403 3501
rect 10041 3496 73403 3498
rect 10041 3440 10046 3496
rect 10102 3440 73342 3496
rect 73398 3440 73403 3496
rect 10041 3438 73403 3440
rect 10041 3435 10107 3438
rect 73337 3435 73403 3438
rect 128261 3498 128327 3501
rect 165889 3498 165955 3501
rect 128261 3496 165955 3498
rect 128261 3440 128266 3496
rect 128322 3440 165894 3496
rect 165950 3440 165955 3496
rect 128261 3438 165955 3440
rect 128261 3435 128327 3438
rect 165889 3435 165955 3438
rect 166257 3498 166323 3501
rect 218145 3498 218211 3501
rect 166257 3496 218211 3498
rect 166257 3440 166262 3496
rect 166318 3440 218150 3496
rect 218206 3440 218211 3496
rect 166257 3438 218211 3440
rect 166257 3435 166323 3438
rect 218145 3435 218211 3438
rect 231761 3498 231827 3501
rect 464429 3498 464495 3501
rect 231761 3496 464495 3498
rect 231761 3440 231766 3496
rect 231822 3440 464434 3496
rect 464490 3440 464495 3496
rect 231761 3438 464495 3440
rect 231761 3435 231827 3438
rect 464429 3435 464495 3438
rect 5257 3362 5323 3365
rect 71681 3362 71747 3365
rect 5257 3360 71747 3362
rect 5257 3304 5262 3360
rect 5318 3304 71686 3360
rect 71742 3304 71747 3360
rect 5257 3302 71747 3304
rect 5257 3299 5323 3302
rect 71681 3299 71747 3302
rect 80145 3362 80211 3365
rect 82537 3362 82603 3365
rect 80145 3360 82603 3362
rect 80145 3304 80150 3360
rect 80206 3304 82542 3360
rect 82598 3304 82603 3360
rect 80145 3302 82603 3304
rect 80145 3299 80211 3302
rect 82537 3299 82603 3302
rect 144821 3362 144887 3365
rect 214649 3362 214715 3365
rect 144821 3360 214715 3362
rect 144821 3304 144826 3360
rect 144882 3304 214654 3360
rect 214710 3304 214715 3360
rect 144821 3302 214715 3304
rect 144821 3299 144887 3302
rect 214649 3299 214715 3302
rect 234521 3362 234587 3365
rect 471513 3362 471579 3365
rect 234521 3360 471579 3362
rect 234521 3304 234526 3360
rect 234582 3304 471518 3360
rect 471574 3304 471579 3360
rect 234521 3302 471579 3304
rect 234521 3299 234587 3302
rect 471513 3299 471579 3302
rect 79777 3226 79843 3229
rect 80053 3226 80119 3229
rect 79777 3224 80119 3226
rect 79777 3168 79782 3224
rect 79838 3168 80058 3224
rect 80114 3168 80119 3224
rect 79777 3166 80119 3168
rect 79777 3163 79843 3166
rect 80053 3163 80119 3166
rect 125317 3226 125383 3229
rect 159909 3226 159975 3229
rect 125317 3224 159975 3226
rect 125317 3168 125322 3224
rect 125378 3168 159914 3224
rect 159970 3168 159975 3224
rect 125317 3166 159975 3168
rect 125317 3163 125383 3166
rect 159909 3163 159975 3166
rect 356697 3226 356763 3229
rect 359641 3226 359707 3229
rect 356697 3224 359707 3226
rect 356697 3168 356702 3224
rect 356758 3168 359646 3224
rect 359702 3168 359707 3224
rect 356697 3166 359707 3168
rect 356697 3163 356763 3166
rect 359641 3163 359707 3166
rect 151721 2954 151787 2957
rect 157241 2954 157307 2957
rect 151721 2952 157307 2954
rect 151721 2896 151726 2952
rect 151782 2896 157246 2952
rect 157302 2896 157307 2952
rect 151721 2894 157307 2896
rect 151721 2891 151787 2894
rect 157241 2891 157307 2894
<< via3 >>
rect 103468 570284 103532 570348
rect 94820 570208 94884 570212
rect 94820 570152 94870 570208
rect 94870 570152 94884 570208
rect 94820 570148 94884 570152
rect 98316 570208 98380 570212
rect 98316 570152 98366 570208
rect 98366 570152 98380 570208
rect 98316 570148 98380 570152
rect 101812 570208 101876 570212
rect 101812 570152 101826 570208
rect 101826 570152 101876 570208
rect 101812 570148 101876 570152
rect 108804 570148 108868 570212
rect 112300 570208 112364 570212
rect 112300 570152 112314 570208
rect 112314 570152 112364 570208
rect 112300 570148 112364 570152
rect 113220 570148 113284 570212
rect 119844 570148 119908 570212
rect 203012 570148 203076 570212
rect 220676 570208 220740 570212
rect 220676 570152 220726 570208
rect 220726 570152 220740 570208
rect 220676 570148 220740 570152
rect 238708 570208 238772 570212
rect 238708 570152 238758 570208
rect 238758 570152 238772 570208
rect 238708 570148 238772 570152
rect 113664 569800 113728 569804
rect 113664 569744 113694 569800
rect 113694 569744 113728 569800
rect 113664 569740 113728 569744
rect 118336 569800 118400 569804
rect 118336 569744 118386 569800
rect 118386 569744 118400 569800
rect 118336 569740 118400 569744
rect 120672 569800 120736 569804
rect 120672 569744 120722 569800
rect 120722 569744 120736 569800
rect 120672 569740 120736 569744
rect 113788 569604 113852 569668
rect 117168 569664 117232 569668
rect 117168 569608 117190 569664
rect 117190 569608 117232 569664
rect 117168 569604 117232 569608
rect 118460 569604 118524 569668
rect 217824 569664 217888 569668
rect 217824 569608 217874 569664
rect 217874 569608 217888 569664
rect 217824 569604 217888 569608
rect 119476 569120 119540 569124
rect 119476 569064 119490 569120
rect 119490 569064 119540 569120
rect 119476 569060 119540 569064
rect 120948 569120 121012 569124
rect 120948 569064 120998 569120
rect 120998 569064 121012 569120
rect 120948 569060 121012 569064
rect 116716 568924 116780 568988
rect 122604 568788 122668 568852
rect 114692 568712 114756 568716
rect 114692 568656 114742 568712
rect 114742 568656 114756 568712
rect 114692 568652 114756 568656
rect 115060 568652 115124 568716
rect 86540 568516 86604 568580
rect 93900 568516 93964 568580
rect 101444 568516 101508 568580
rect 102732 568516 102796 568580
rect 103100 568576 103164 568580
rect 103100 568520 103150 568576
rect 103150 568520 103164 568576
rect 103100 568516 103164 568520
rect 104020 568576 104084 568580
rect 104020 568520 104070 568576
rect 104070 568520 104084 568576
rect 104020 568516 104084 568520
rect 104756 568576 104820 568580
rect 104756 568520 104806 568576
rect 104806 568520 104820 568576
rect 104756 568516 104820 568520
rect 105308 568576 105372 568580
rect 105308 568520 105322 568576
rect 105322 568520 105372 568576
rect 105308 568516 105372 568520
rect 105860 568516 105924 568580
rect 106596 568576 106660 568580
rect 106596 568520 106646 568576
rect 106646 568520 106660 568576
rect 106596 568516 106660 568520
rect 106780 568516 106844 568580
rect 107700 568576 107764 568580
rect 107700 568520 107750 568576
rect 107750 568520 107764 568576
rect 107700 568516 107764 568520
rect 108620 568516 108684 568580
rect 109724 568516 109788 568580
rect 110828 568516 110892 568580
rect 111564 568516 111628 568580
rect 115796 568576 115860 568580
rect 115796 568520 115846 568576
rect 115846 568520 115860 568576
rect 115796 568516 115860 568520
rect 126468 568516 126532 568580
rect 128492 568576 128556 568580
rect 128492 568520 128506 568576
rect 128506 568520 128556 568576
rect 128492 568516 128556 568520
rect 196204 568516 196268 568580
rect 197676 568516 197740 568580
rect 202276 568576 202340 568580
rect 202276 568520 202290 568576
rect 202290 568520 202340 568576
rect 202276 568516 202340 568520
rect 203932 568516 203996 568580
rect 204852 568576 204916 568580
rect 204852 568520 204866 568576
rect 204866 568520 204916 568576
rect 204852 568516 204916 568520
rect 205404 568516 205468 568580
rect 207060 568576 207124 568580
rect 207060 568520 207074 568576
rect 207074 568520 207124 568576
rect 207060 568516 207124 568520
rect 209452 568516 209516 568580
rect 211844 568576 211908 568580
rect 211844 568520 211894 568576
rect 211894 568520 211908 568576
rect 211844 568516 211908 568520
rect 213132 568576 213196 568580
rect 213132 568520 213146 568576
rect 213146 568520 213196 568576
rect 213132 568516 213196 568520
rect 214052 568576 214116 568580
rect 214052 568520 214102 568576
rect 214102 568520 214116 568576
rect 214052 568516 214116 568520
rect 215524 568576 215588 568580
rect 215524 568520 215574 568576
rect 215574 568520 215588 568576
rect 215524 568516 215588 568520
rect 216628 568516 216692 568580
rect 218836 568516 218900 568580
rect 221412 568576 221476 568580
rect 221412 568520 221462 568576
rect 221462 568520 221476 568576
rect 221412 568516 221476 568520
rect 222332 568576 222396 568580
rect 222332 568520 222382 568576
rect 222382 568520 222396 568576
rect 222332 568516 222396 568520
rect 223620 568576 223684 568580
rect 223620 568520 223670 568576
rect 223670 568520 223684 568576
rect 223620 568516 223684 568520
rect 225828 568576 225892 568580
rect 225828 568520 225878 568576
rect 225878 568520 225892 568576
rect 225828 568516 225892 568520
rect 226196 568576 226260 568580
rect 226196 568520 226246 568576
rect 226246 568520 226260 568576
rect 226196 568516 226260 568520
rect 227116 568576 227180 568580
rect 227116 568520 227166 568576
rect 227166 568520 227180 568576
rect 227116 568516 227180 568520
rect 227300 568516 227364 568580
rect 228404 568576 228468 568580
rect 228404 568520 228418 568576
rect 228418 568520 228468 568576
rect 228404 568516 228468 568520
rect 228772 568516 228836 568580
rect 229324 568576 229388 568580
rect 229324 568520 229374 568576
rect 229374 568520 229388 568576
rect 229324 568516 229388 568520
rect 230244 568516 230308 568580
rect 230796 568516 230860 568580
rect 233004 568576 233068 568580
rect 233004 568520 233054 568576
rect 233054 568520 233068 568576
rect 233004 568516 233068 568520
rect 234476 568576 234540 568580
rect 234476 568520 234526 568576
rect 234526 568520 234540 568576
rect 234476 568516 234540 568520
rect 235764 568516 235828 568580
rect 237236 568576 237300 568580
rect 237236 568520 237286 568576
rect 237286 568520 237300 568576
rect 237236 568516 237300 568520
rect 238156 568516 238220 568580
rect 239628 568516 239692 568580
rect 95188 568440 95252 568444
rect 95188 568384 95202 568440
rect 95202 568384 95252 568440
rect 95188 568380 95252 568384
rect 109908 568440 109972 568444
rect 109908 568384 109922 568440
rect 109922 568384 109972 568440
rect 109908 568380 109972 568384
rect 194364 568440 194428 568444
rect 194364 568384 194414 568440
rect 194414 568384 194428 568440
rect 194364 568380 194428 568384
rect 203748 568440 203812 568444
rect 203748 568384 203762 568440
rect 203762 568384 203812 568440
rect 203748 568380 203812 568384
rect 220124 568440 220188 568444
rect 220124 568384 220138 568440
rect 220138 568384 220188 568440
rect 220124 568380 220188 568384
rect 225644 568380 225708 568444
rect 232636 568380 232700 568444
rect 234660 568440 234724 568444
rect 234660 568384 234674 568440
rect 234674 568384 234724 568440
rect 234660 568380 234724 568384
rect 92612 568244 92676 568308
rect 96108 568244 96172 568308
rect 97396 568244 97460 568308
rect 99604 568244 99668 568308
rect 100892 568244 100956 568308
rect 123708 568244 123772 568308
rect 124260 568304 124324 568308
rect 124260 568248 124310 568304
rect 124310 568248 124324 568304
rect 124260 568244 124324 568248
rect 125364 568244 125428 568308
rect 129596 568244 129660 568308
rect 224724 568304 224788 568308
rect 224724 568248 224774 568304
rect 224774 568248 224788 568304
rect 224724 568244 224788 568248
rect 233556 568244 233620 568308
rect 237420 568304 237484 568308
rect 237420 568248 237434 568304
rect 237434 568248 237484 568304
rect 237420 568244 237484 568248
rect 200252 568108 200316 568172
rect 230612 568108 230676 568172
rect 232820 568108 232884 568172
rect 236132 568108 236196 568172
rect 201540 567972 201604 568036
rect 231900 568032 231964 568036
rect 231900 567976 231914 568032
rect 231914 567976 231964 568032
rect 231900 567972 231964 567976
rect 199516 567836 199580 567900
rect 91508 567700 91572 567764
rect 97764 567700 97828 567764
rect 100340 567700 100404 567764
rect 110276 567760 110340 567764
rect 110276 567704 110326 567760
rect 110326 567704 110340 567760
rect 110276 567700 110340 567704
rect 124996 567700 125060 567764
rect 83412 567564 83476 567628
rect 88564 567428 88628 567492
rect 87460 567292 87524 567356
rect 90036 567352 90100 567356
rect 90036 567296 90050 567352
rect 90050 567296 90100 567352
rect 90036 567292 90100 567296
rect 121500 567292 121564 567356
rect 124260 567292 124324 567356
rect 208348 567292 208412 567356
rect 210372 567292 210436 567356
rect 217548 567292 217612 567356
rect 93348 567156 93412 567220
rect 94268 567156 94332 567220
rect 96292 567156 96356 567220
rect 98868 567156 98932 567220
rect 122972 567156 123036 567220
rect 124812 567156 124876 567220
rect 126652 567156 126716 567220
rect 127756 567156 127820 567220
rect 128124 567216 128188 567220
rect 128124 567160 128174 567216
rect 128174 567160 128188 567216
rect 128124 567156 128188 567160
rect 205772 567156 205836 567220
rect 206876 567216 206940 567220
rect 206876 567160 206926 567216
rect 206926 567160 206940 567216
rect 206876 567156 206940 567160
rect 207980 567156 208044 567220
rect 209268 567156 209332 567220
rect 210556 567156 210620 567220
rect 210924 567216 210988 567220
rect 210924 567160 210974 567216
rect 210974 567160 210988 567216
rect 210924 567156 210988 567160
rect 212396 567216 212460 567220
rect 212396 567160 212446 567216
rect 212446 567160 212460 567216
rect 212396 567156 212460 567160
rect 213500 567156 213564 567220
rect 214788 567156 214852 567220
rect 216260 567156 216324 567220
rect 217916 567216 217980 567220
rect 217916 567160 217930 567216
rect 217930 567160 217980 567216
rect 217916 567156 217980 567160
rect 219204 567156 219268 567220
rect 221964 567156 222028 567220
rect 223252 567156 223316 567220
rect 223804 567156 223868 567220
rect 117268 566476 117332 566540
rect 121500 566068 121564 566132
rect 320220 516760 320284 516764
rect 320220 516704 320234 516760
rect 320234 516704 320284 516760
rect 320220 516700 320284 516704
rect 273852 516428 273916 516492
rect 320220 512136 320284 512140
rect 320220 512080 320234 512136
rect 320234 512080 320284 512136
rect 320220 512076 320284 512080
rect 320036 509084 320100 509148
rect 320036 507860 320100 507924
rect 320404 507512 320468 507516
rect 320404 507456 320418 507512
rect 320418 507456 320468 507512
rect 320404 507452 320468 507456
rect 319852 506288 319916 506292
rect 319852 506232 319866 506288
rect 319866 506232 319916 506288
rect 319852 506228 319916 506232
rect 320220 506288 320284 506292
rect 320220 506232 320234 506288
rect 320234 506232 320284 506288
rect 320220 506228 320284 506232
rect 320772 504792 320836 504796
rect 320772 504736 320786 504792
rect 320786 504736 320836 504792
rect 320772 504732 320836 504736
rect 276612 503780 276676 503844
rect 319852 503780 319916 503844
rect 320588 503704 320652 503708
rect 320588 503648 320602 503704
rect 320602 503648 320652 503704
rect 320588 503644 320652 503648
rect 320220 503160 320284 503164
rect 320220 503104 320234 503160
rect 320234 503104 320284 503160
rect 320220 503100 320284 503104
rect 320404 502480 320468 502484
rect 320404 502424 320418 502480
rect 320418 502424 320468 502480
rect 320404 502420 320468 502424
rect 320772 501392 320836 501396
rect 320772 501336 320822 501392
rect 320822 501336 320836 501392
rect 320772 501332 320836 501336
rect 319852 500984 319916 500988
rect 319852 500928 319866 500984
rect 319866 500928 319916 500984
rect 319852 500924 319916 500928
rect 320036 500848 320100 500852
rect 320036 500792 320050 500848
rect 320050 500792 320100 500848
rect 320036 500788 320100 500792
rect 320588 500168 320652 500172
rect 320588 500112 320638 500168
rect 320638 500112 320652 500168
rect 320588 500108 320652 500112
rect 320220 499624 320284 499628
rect 320220 499568 320270 499624
rect 320270 499568 320284 499624
rect 320220 499564 320284 499568
rect 320772 498944 320836 498948
rect 320772 498888 320786 498944
rect 320786 498888 320836 498944
rect 320772 498884 320836 498888
rect 319852 497992 319916 497996
rect 319852 497936 319866 497992
rect 319866 497936 319916 497992
rect 319852 497932 319916 497936
rect 320220 497856 320284 497860
rect 320220 497800 320270 497856
rect 320270 497800 320284 497856
rect 320220 497796 320284 497800
rect 320220 497312 320284 497316
rect 320220 497256 320234 497312
rect 320234 497256 320284 497312
rect 320220 497252 320284 497256
rect 320404 496632 320468 496636
rect 320404 496576 320454 496632
rect 320454 496576 320468 496632
rect 320404 496572 320468 496576
rect 320772 495544 320836 495548
rect 320772 495488 320822 495544
rect 320822 495488 320836 495544
rect 320772 495484 320836 495488
rect 319852 495272 319916 495276
rect 319852 495216 319866 495272
rect 319866 495216 319916 495272
rect 319852 495212 319916 495216
rect 320220 495000 320284 495004
rect 320220 494944 320234 495000
rect 320234 494944 320284 495000
rect 320220 494940 320284 494944
rect 320588 494592 320652 494596
rect 320588 494536 320602 494592
rect 320602 494536 320652 494592
rect 320588 494532 320652 494536
rect 319852 493776 319916 493780
rect 319852 493720 319866 493776
rect 319866 493720 319916 493776
rect 319852 493716 319916 493720
rect 320404 493504 320468 493508
rect 320404 493448 320418 493504
rect 320418 493448 320468 493504
rect 320404 493444 320468 493448
rect 320036 492688 320100 492692
rect 320036 492632 320050 492688
rect 320050 492632 320100 492688
rect 320036 492628 320100 492632
rect 320588 492280 320652 492284
rect 320588 492224 320638 492280
rect 320638 492224 320652 492280
rect 320588 492220 320652 492224
rect 319852 491192 319916 491196
rect 319852 491136 319866 491192
rect 319866 491136 319916 491192
rect 319852 491132 319916 491136
rect 320588 490920 320652 490924
rect 320588 490864 320638 490920
rect 320638 490864 320652 490920
rect 320588 490860 320652 490864
rect 320220 490376 320284 490380
rect 320220 490320 320234 490376
rect 320234 490320 320284 490376
rect 320220 490316 320284 490320
rect 320220 489772 320284 489836
rect 320772 488472 320836 488476
rect 320772 488416 320786 488472
rect 320786 488416 320836 488472
rect 320772 488412 320836 488416
rect 319852 487928 319916 487932
rect 319852 487872 319866 487928
rect 319866 487872 319916 487928
rect 319852 487868 319916 487872
rect 320220 487928 320284 487932
rect 320220 487872 320234 487928
rect 320234 487872 320284 487928
rect 320220 487868 320284 487872
rect 320220 487384 320284 487388
rect 320220 487328 320270 487384
rect 320270 487328 320284 487384
rect 320220 487324 320284 487328
rect 319852 486644 319916 486708
rect 320404 486160 320468 486164
rect 320404 486104 320454 486160
rect 320454 486104 320468 486160
rect 320404 486100 320468 486104
rect 319852 485616 319916 485620
rect 319852 485560 319866 485616
rect 319866 485560 319916 485616
rect 319852 485556 319916 485560
rect 320588 484936 320652 484940
rect 320588 484880 320602 484936
rect 320602 484880 320652 484936
rect 320588 484876 320652 484880
rect 320220 484528 320284 484532
rect 320220 484472 320234 484528
rect 320234 484472 320284 484528
rect 320220 484468 320284 484472
rect 320404 484120 320468 484124
rect 320404 484064 320418 484120
rect 320418 484064 320468 484120
rect 320404 484060 320468 484064
rect 319852 483032 319916 483036
rect 319852 482976 319866 483032
rect 319866 482976 319916 483032
rect 319852 482972 319916 482976
rect 320588 482624 320652 482628
rect 320588 482568 320638 482624
rect 320638 482568 320652 482624
rect 320588 482564 320652 482568
rect 320220 482080 320284 482084
rect 320220 482024 320234 482080
rect 320234 482024 320284 482080
rect 320220 482020 320284 482024
rect 320404 481536 320468 481540
rect 320404 481480 320454 481536
rect 320454 481480 320468 481536
rect 320404 481476 320468 481480
rect 320588 480312 320652 480316
rect 320588 480256 320602 480312
rect 320602 480256 320652 480312
rect 320588 480252 320652 480256
rect 319852 479768 319916 479772
rect 319852 479712 319866 479768
rect 319866 479712 319916 479768
rect 319852 479708 319916 479712
rect 320220 479768 320284 479772
rect 320220 479712 320234 479768
rect 320234 479712 320284 479768
rect 320220 479708 320284 479712
rect 320588 479088 320652 479092
rect 320588 479032 320638 479088
rect 320638 479032 320652 479088
rect 320588 479028 320652 479032
rect 320588 478000 320652 478004
rect 320588 477944 320638 478000
rect 320638 477944 320652 478000
rect 320588 477940 320652 477944
rect 320220 476776 320284 476780
rect 320220 476720 320234 476776
rect 320234 476720 320284 476776
rect 320220 476716 320284 476720
rect 320404 476776 320468 476780
rect 320404 476720 320418 476776
rect 320418 476720 320468 476776
rect 320404 476716 320468 476720
rect 319852 475764 319916 475828
rect 320772 475824 320836 475828
rect 320772 475768 320822 475824
rect 320822 475768 320836 475824
rect 320772 475764 320836 475768
rect 320588 475628 320652 475692
rect 320220 474464 320284 474468
rect 320220 474408 320234 474464
rect 320234 474408 320284 474464
rect 320220 474404 320284 474408
rect 320772 474464 320836 474468
rect 320772 474408 320786 474464
rect 320786 474408 320836 474464
rect 320772 474404 320836 474408
rect 320220 473240 320284 473244
rect 320220 473184 320270 473240
rect 320270 473184 320284 473240
rect 320220 473180 320284 473184
rect 320588 473240 320652 473244
rect 320588 473184 320602 473240
rect 320602 473184 320652 473240
rect 320588 473180 320652 473184
rect 320220 472228 320284 472292
rect 320404 472152 320468 472156
rect 320404 472096 320418 472152
rect 320418 472096 320468 472152
rect 320404 472092 320468 472096
rect 320588 471004 320652 471068
rect 320404 470928 320468 470932
rect 320404 470872 320454 470928
rect 320454 470872 320468 470928
rect 320404 470868 320468 470872
rect 320404 470052 320468 470116
rect 320220 469840 320284 469844
rect 320220 469784 320270 469840
rect 320270 469784 320284 469840
rect 320220 469780 320284 469784
rect 319852 469100 319916 469164
rect 320588 468888 320652 468892
rect 320588 468832 320638 468888
rect 320638 468832 320652 468888
rect 320588 468828 320652 468832
rect 320220 468616 320284 468620
rect 320220 468560 320234 468616
rect 320234 468560 320284 468616
rect 320220 468556 320284 468560
rect 320404 467604 320468 467668
rect 320220 465216 320284 465220
rect 320220 465160 320234 465216
rect 320234 465160 320284 465216
rect 320220 465156 320284 465160
rect 320404 465156 320468 465220
rect 276612 404772 276676 404836
rect 279924 396068 279988 396132
rect 320220 392048 320284 392052
rect 320220 391992 320234 392048
rect 320234 391992 320284 392048
rect 320220 391988 320284 391992
rect 320220 389872 320284 389876
rect 320220 389816 320270 389872
rect 320270 389816 320284 389872
rect 320220 389812 320284 389816
rect 320220 388996 320284 389060
rect 320220 387560 320284 387564
rect 320220 387504 320270 387560
rect 320270 387504 320284 387560
rect 320220 387500 320284 387504
rect 319852 386412 319916 386476
rect 320220 386336 320284 386340
rect 320220 386280 320234 386336
rect 320234 386280 320284 386336
rect 320220 386276 320284 386280
rect 320588 384840 320652 384844
rect 320588 384784 320638 384840
rect 320638 384784 320652 384840
rect 320588 384780 320652 384784
rect 319852 383692 319916 383756
rect 320772 383616 320836 383620
rect 320772 383560 320786 383616
rect 320786 383560 320836 383616
rect 320772 383556 320836 383560
rect 320220 383208 320284 383212
rect 320220 383152 320270 383208
rect 320270 383152 320284 383208
rect 320220 383148 320284 383152
rect 320772 382528 320836 382532
rect 320772 382472 320822 382528
rect 320822 382472 320836 382528
rect 320772 382468 320836 382472
rect 320588 381304 320652 381308
rect 320588 381248 320638 381304
rect 320638 381248 320652 381304
rect 320588 381244 320652 381248
rect 320404 380896 320468 380900
rect 320404 380840 320418 380896
rect 320418 380840 320468 380896
rect 320404 380836 320468 380840
rect 320772 380216 320836 380220
rect 320772 380160 320822 380216
rect 320822 380160 320836 380216
rect 320772 380156 320836 380160
rect 320220 379672 320284 379676
rect 320220 379616 320270 379672
rect 320270 379616 320284 379672
rect 320220 379612 320284 379616
rect 319852 379476 319916 379540
rect 320404 378992 320468 378996
rect 320404 378936 320454 378992
rect 320454 378936 320468 378992
rect 320404 378932 320468 378936
rect 320588 378448 320652 378452
rect 320588 378392 320602 378448
rect 320602 378392 320652 378448
rect 320588 378388 320652 378392
rect 320772 377768 320836 377772
rect 320772 377712 320822 377768
rect 320822 377712 320836 377768
rect 320772 377708 320836 377712
rect 320036 376620 320100 376684
rect 320220 376136 320284 376140
rect 320220 376080 320270 376136
rect 320270 376080 320284 376136
rect 320220 376076 320284 376080
rect 320220 375456 320284 375460
rect 320220 375400 320234 375456
rect 320234 375400 320284 375456
rect 320220 375396 320284 375400
rect 319852 375184 319916 375188
rect 319852 375128 319866 375184
rect 319866 375128 319916 375184
rect 319852 375124 319916 375128
rect 320588 374368 320652 374372
rect 320588 374312 320602 374368
rect 320602 374312 320652 374368
rect 320588 374308 320652 374312
rect 320036 373824 320100 373828
rect 320036 373768 320050 373824
rect 320050 373768 320100 373824
rect 320036 373764 320100 373768
rect 320036 373144 320100 373148
rect 320036 373088 320086 373144
rect 320086 373088 320100 373144
rect 320036 373084 320100 373088
rect 319852 372676 319916 372740
rect 320404 372600 320468 372604
rect 320404 372544 320418 372600
rect 320418 372544 320468 372600
rect 320404 372540 320468 372544
rect 320588 372328 320652 372332
rect 320588 372272 320638 372328
rect 320638 372272 320652 372328
rect 320588 372268 320652 372272
rect 320220 371512 320284 371516
rect 320220 371456 320270 371512
rect 320270 371456 320284 371512
rect 320220 371452 320284 371456
rect 320772 371240 320836 371244
rect 320772 371184 320822 371240
rect 320822 371184 320836 371240
rect 320772 371180 320836 371184
rect 320404 369744 320468 369748
rect 320404 369688 320454 369744
rect 320454 369688 320468 369744
rect 320404 369684 320468 369688
rect 320404 369200 320468 369204
rect 320404 369144 320418 369200
rect 320418 369144 320468 369200
rect 320404 369140 320468 369144
rect 319852 368460 319916 368524
rect 320772 368520 320836 368524
rect 320772 368464 320822 368520
rect 320822 368464 320836 368520
rect 320772 368460 320836 368464
rect 320220 367976 320284 367980
rect 320220 367920 320270 367976
rect 320270 367920 320284 367976
rect 320220 367916 320284 367920
rect 319668 367236 319732 367300
rect 320772 367296 320836 367300
rect 320772 367240 320822 367296
rect 320822 367240 320836 367296
rect 320772 367236 320836 367240
rect 320588 366208 320652 366212
rect 320588 366152 320638 366208
rect 320638 366152 320652 366208
rect 320588 366148 320652 366152
rect 320036 365604 320100 365668
rect 320220 364984 320284 364988
rect 320220 364928 320234 364984
rect 320234 364928 320284 364984
rect 320220 364924 320284 364928
rect 320404 364440 320468 364444
rect 320404 364384 320454 364440
rect 320454 364384 320468 364440
rect 320404 364380 320468 364384
rect 320036 363760 320100 363764
rect 320036 363704 320050 363760
rect 320050 363704 320100 363760
rect 320036 363700 320100 363704
rect 319484 363428 319548 363492
rect 320036 362672 320100 362676
rect 320036 362616 320086 362672
rect 320086 362616 320100 362672
rect 320036 362612 320100 362616
rect 320404 362128 320468 362132
rect 320404 362072 320418 362128
rect 320418 362072 320468 362128
rect 320404 362068 320468 362072
rect 319852 361448 319916 361452
rect 319852 361392 319866 361448
rect 319866 361392 319916 361448
rect 319852 361388 319916 361392
rect 320220 361448 320284 361452
rect 320220 361392 320234 361448
rect 320234 361392 320284 361448
rect 320220 361388 320284 361392
rect 320220 361040 320284 361044
rect 320220 360984 320270 361040
rect 320270 360984 320284 361040
rect 320220 360980 320284 360984
rect 320220 360360 320284 360364
rect 320220 360304 320270 360360
rect 320270 360304 320284 360360
rect 320220 360300 320284 360304
rect 320404 359816 320468 359820
rect 320404 359760 320454 359816
rect 320454 359760 320468 359816
rect 320404 359756 320468 359760
rect 320404 358592 320468 358596
rect 320404 358536 320418 358592
rect 320418 358536 320468 358592
rect 320404 358532 320468 358536
rect 320220 357912 320284 357916
rect 320220 357856 320270 357912
rect 320270 357856 320284 357912
rect 320220 357852 320284 357856
rect 273852 357172 273916 357236
rect 320588 357096 320652 357100
rect 320588 357040 320602 357096
rect 320602 357040 320652 357096
rect 320588 357036 320652 357040
rect 320220 356824 320284 356828
rect 320220 356768 320234 356824
rect 320234 356768 320284 356824
rect 320220 356764 320284 356768
rect 320588 356008 320652 356012
rect 320588 355952 320638 356008
rect 320638 355952 320652 356008
rect 320588 355948 320652 355952
rect 320220 355600 320284 355604
rect 320220 355544 320234 355600
rect 320234 355544 320284 355600
rect 320220 355540 320284 355544
rect 320772 354648 320836 354652
rect 320772 354592 320822 354648
rect 320822 354592 320836 354648
rect 320772 354588 320836 354592
rect 320220 354512 320284 354516
rect 320220 354456 320234 354512
rect 320234 354456 320284 354512
rect 320220 354452 320284 354456
rect 319852 353364 319916 353428
rect 320220 353288 320284 353292
rect 320220 353232 320270 353288
rect 320270 353232 320284 353288
rect 320220 353228 320284 353232
rect 320772 353288 320836 353292
rect 320772 353232 320822 353288
rect 320822 353232 320836 353288
rect 320772 353228 320836 353232
rect 320220 352608 320284 352612
rect 320220 352552 320234 352608
rect 320234 352552 320284 352608
rect 320220 352548 320284 352552
rect 320404 352472 320468 352476
rect 320404 352416 320418 352472
rect 320418 352416 320468 352472
rect 320404 352412 320468 352416
rect 320588 351248 320652 351252
rect 320588 351192 320638 351248
rect 320638 351192 320652 351248
rect 320588 351188 320652 351192
rect 320404 350976 320468 350980
rect 320404 350920 320418 350976
rect 320418 350920 320468 350976
rect 320404 350916 320468 350920
rect 320772 350160 320836 350164
rect 320772 350104 320786 350160
rect 320786 350104 320836 350160
rect 320772 350100 320836 350104
rect 320220 349752 320284 349756
rect 320220 349696 320234 349752
rect 320234 349696 320284 349752
rect 320220 349692 320284 349696
rect 320220 348664 320284 348668
rect 320220 348608 320234 348664
rect 320234 348608 320284 348664
rect 320220 348604 320284 348608
rect 320220 346352 320284 346356
rect 320220 346296 320234 346352
rect 320234 346296 320284 346352
rect 320220 346292 320284 346296
rect 70164 320588 70228 320652
rect 106596 241496 106660 241500
rect 106596 241440 106646 241496
rect 106646 241440 106660 241496
rect 106596 241436 106660 241440
rect 106596 235376 106660 235380
rect 106596 235320 106610 235376
rect 106610 235320 106660 235376
rect 106596 235316 106660 235320
rect 77524 202872 77588 202876
rect 77524 202816 77538 202872
rect 77538 202816 77588 202872
rect 77524 202812 77588 202816
rect 77524 195800 77588 195804
rect 77524 195744 77574 195800
rect 77574 195744 77588 195800
rect 77524 195740 77588 195744
rect 255268 143440 255332 143444
rect 255268 143384 255282 143440
rect 255282 143384 255332 143440
rect 255268 143380 255332 143384
rect 255268 133860 255332 133924
rect 97028 60752 97092 60756
rect 97028 60696 97042 60752
rect 97042 60696 97092 60752
rect 97028 60692 97092 60696
rect 97028 56672 97092 56676
rect 97028 56616 97042 56672
rect 97042 56616 97092 56672
rect 97028 56612 97092 56616
rect 227300 22068 227364 22132
rect 227300 19408 227364 19412
rect 227300 19352 227350 19408
rect 227350 19352 227364 19408
rect 227300 19348 227364 19352
rect 266262 15132 266326 15196
rect 266262 14724 266326 14788
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 70166 320653 70226 395982
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 70163 320652 70229 320653
rect 70163 320588 70164 320652
rect 70228 320588 70229 320652
rect 70163 320587 70229 320588
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 661247 80604 693098
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661247 84204 696698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 661247 91404 667898
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 661247 95004 671498
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 661247 98604 675098
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 661247 102204 678698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 661247 109404 685898
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 661247 113004 689498
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 661247 116604 693098
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661247 120204 696698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 661247 127404 667898
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 661247 131004 671498
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 661247 134604 675098
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 661247 138204 678698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 661247 145404 685898
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 661247 149004 689498
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 661247 152604 693098
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661247 156204 696698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 103308 570490 103530 570550
rect 103470 570349 103530 570490
rect 104022 570490 104352 570550
rect 109910 570490 110192 570550
rect 103467 570348 103533 570349
rect 103467 570284 103468 570348
rect 103532 570284 103533 570348
rect 103467 570283 103533 570284
rect 94819 570212 94885 570213
rect 83414 570150 83833 570210
rect 86542 570150 86832 570210
rect 87462 570150 88000 570210
rect 88566 570150 89168 570210
rect 90038 570150 90336 570210
rect 91504 570150 91570 570210
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 80004 549654 80604 570000
rect 83414 567629 83474 570150
rect 83411 567628 83477 567629
rect 83411 567564 83412 567628
rect 83476 567564 83477 567628
rect 83411 567563 83477 567564
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 77523 202876 77589 202877
rect 77523 202812 77524 202876
rect 77588 202812 77589 202876
rect 77523 202811 77589 202812
rect 77526 195805 77586 202811
rect 77523 195804 77589 195805
rect 77523 195740 77524 195804
rect 77588 195740 77589 195804
rect 77523 195739 77589 195740
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 553254 84204 570000
rect 86542 568581 86602 570150
rect 86539 568580 86605 568581
rect 86539 568516 86540 568580
rect 86604 568516 86605 568580
rect 86539 568515 86605 568516
rect 87462 567357 87522 570150
rect 88566 567493 88626 570150
rect 88563 567492 88629 567493
rect 88563 567428 88564 567492
rect 88628 567428 88629 567492
rect 88563 567427 88629 567428
rect 90038 567357 90098 570150
rect 87459 567356 87525 567357
rect 87459 567292 87460 567356
rect 87524 567292 87525 567356
rect 87459 567291 87525 567292
rect 90035 567356 90101 567357
rect 90035 567292 90036 567356
rect 90100 567292 90101 567356
rect 90035 567291 90101 567292
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 560454 91404 570000
rect 91510 567765 91570 570150
rect 92614 568309 92674 570210
rect 92796 570150 93410 570210
rect 92611 568308 92677 568309
rect 92611 568244 92612 568308
rect 92676 568244 92677 568308
rect 92611 568243 92677 568244
rect 91507 567764 91573 567765
rect 91507 567700 91508 567764
rect 91572 567700 91573 567764
rect 91507 567699 91573 567700
rect 93350 567221 93410 570150
rect 93810 569530 93870 570180
rect 93964 570150 94330 570210
rect 93810 569470 93962 569530
rect 93902 568581 93962 569470
rect 93899 568580 93965 568581
rect 93899 568516 93900 568580
rect 93964 568516 93965 568580
rect 93899 568515 93965 568516
rect 94270 567221 94330 570150
rect 94819 570148 94820 570212
rect 94884 570210 94885 570212
rect 98315 570212 98381 570213
rect 94884 570150 95008 570210
rect 94884 570148 94885 570150
rect 94819 570147 94885 570148
rect 93347 567220 93413 567221
rect 93347 567156 93348 567220
rect 93412 567156 93413 567220
rect 93347 567155 93413 567156
rect 94267 567220 94333 567221
rect 94267 567156 94268 567220
rect 94332 567156 94333 567220
rect 94267 567155 94333 567156
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 564054 95004 570000
rect 95102 569530 95162 570180
rect 96110 570150 96176 570210
rect 95102 569470 95250 569530
rect 95190 568445 95250 569470
rect 95187 568444 95253 568445
rect 95187 568380 95188 568444
rect 95252 568380 95253 568444
rect 95187 568379 95253 568380
rect 96110 568309 96170 570150
rect 96107 568308 96173 568309
rect 96107 568244 96108 568308
rect 96172 568244 96173 568308
rect 96107 568243 96173 568244
rect 96294 567221 96354 570210
rect 97314 569530 97374 570180
rect 97468 570150 97826 570210
rect 97314 569470 97458 569530
rect 97398 568309 97458 569470
rect 97395 568308 97461 568309
rect 97395 568244 97396 568308
rect 97460 568244 97461 568308
rect 97395 568243 97461 568244
rect 97766 567765 97826 570150
rect 98315 570148 98316 570212
rect 98380 570210 98381 570212
rect 101811 570212 101877 570213
rect 98380 570150 98512 570210
rect 98636 570150 98930 570210
rect 98380 570148 98381 570150
rect 98315 570147 98381 570148
rect 97763 567764 97829 567765
rect 97763 567700 97764 567764
rect 97828 567700 97829 567764
rect 97763 567699 97829 567700
rect 98004 567654 98604 570000
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 96291 567220 96357 567221
rect 96291 567156 96292 567220
rect 96356 567156 96357 567220
rect 96291 567155 96357 567156
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98870 567221 98930 570150
rect 99606 570150 99680 570210
rect 99804 570150 100402 570210
rect 99606 568309 99666 570150
rect 99603 568308 99669 568309
rect 99603 568244 99604 568308
rect 99668 568244 99669 568308
rect 99603 568243 99669 568244
rect 100342 567765 100402 570150
rect 100818 569530 100878 570180
rect 100972 570150 101506 570210
rect 100818 569470 100954 569530
rect 100894 568309 100954 569470
rect 101446 568581 101506 570150
rect 101811 570148 101812 570212
rect 101876 570210 101877 570212
rect 101876 570150 102016 570210
rect 102140 570150 102794 570210
rect 101876 570148 101877 570150
rect 101811 570147 101877 570148
rect 101443 568580 101509 568581
rect 101443 568516 101444 568580
rect 101508 568516 101509 568580
rect 101443 568515 101509 568516
rect 100891 568308 100957 568309
rect 100891 568244 100892 568308
rect 100956 568244 100957 568308
rect 100891 568243 100957 568244
rect 100339 567764 100405 567765
rect 100339 567700 100340 567764
rect 100404 567700 100405 567764
rect 100339 567699 100405 567700
rect 98867 567220 98933 567221
rect 98867 567156 98868 567220
rect 98932 567156 98933 567220
rect 98867 567155 98933 567156
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 97027 60756 97093 60757
rect 97027 60692 97028 60756
rect 97092 60692 97093 60756
rect 97027 60691 97093 60692
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 97030 56677 97090 60691
rect 97027 56676 97093 56677
rect 97027 56612 97028 56676
rect 97092 56612 97093 56676
rect 97027 56611 97093 56612
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 535254 102204 570000
rect 102734 568581 102794 570150
rect 103102 570150 103184 570210
rect 103102 568581 103162 570150
rect 104022 568581 104082 570490
rect 108803 570212 108869 570213
rect 104476 570150 104818 570210
rect 104758 568581 104818 570150
rect 105310 570150 105520 570210
rect 105644 570150 105922 570210
rect 105310 568581 105370 570150
rect 105862 568581 105922 570150
rect 106598 570150 106688 570210
rect 106598 568581 106658 570150
rect 106782 568581 106842 570180
rect 107702 570150 107856 570210
rect 107980 570150 108682 570210
rect 107702 568581 107762 570150
rect 108622 568581 108682 570150
rect 108803 570148 108804 570212
rect 108868 570210 108869 570212
rect 108868 570150 109024 570210
rect 109148 570150 109786 570210
rect 108868 570148 108869 570150
rect 108803 570147 108869 570148
rect 102731 568580 102797 568581
rect 102731 568516 102732 568580
rect 102796 568516 102797 568580
rect 102731 568515 102797 568516
rect 103099 568580 103165 568581
rect 103099 568516 103100 568580
rect 103164 568516 103165 568580
rect 103099 568515 103165 568516
rect 104019 568580 104085 568581
rect 104019 568516 104020 568580
rect 104084 568516 104085 568580
rect 104019 568515 104085 568516
rect 104755 568580 104821 568581
rect 104755 568516 104756 568580
rect 104820 568516 104821 568580
rect 104755 568515 104821 568516
rect 105307 568580 105373 568581
rect 105307 568516 105308 568580
rect 105372 568516 105373 568580
rect 105307 568515 105373 568516
rect 105859 568580 105925 568581
rect 105859 568516 105860 568580
rect 105924 568516 105925 568580
rect 105859 568515 105925 568516
rect 106595 568580 106661 568581
rect 106595 568516 106596 568580
rect 106660 568516 106661 568580
rect 106595 568515 106661 568516
rect 106779 568580 106845 568581
rect 106779 568516 106780 568580
rect 106844 568516 106845 568580
rect 106779 568515 106845 568516
rect 107699 568580 107765 568581
rect 107699 568516 107700 568580
rect 107764 568516 107765 568580
rect 107699 568515 107765 568516
rect 108619 568580 108685 568581
rect 108619 568516 108620 568580
rect 108684 568516 108685 568580
rect 108619 568515 108685 568516
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 108804 542454 109404 570000
rect 109726 568581 109786 570150
rect 109723 568580 109789 568581
rect 109723 568516 109724 568580
rect 109788 568516 109789 568580
rect 109723 568515 109789 568516
rect 109910 568445 109970 570490
rect 112299 570212 112365 570213
rect 110286 569530 110346 570180
rect 110278 569470 110346 569530
rect 110830 570150 111360 570210
rect 109907 568444 109973 568445
rect 109907 568380 109908 568444
rect 109972 568380 109973 568444
rect 109907 568379 109973 568380
rect 110278 567765 110338 569470
rect 110830 568581 110890 570150
rect 111454 569530 111514 570180
rect 112299 570148 112300 570212
rect 112364 570210 112365 570212
rect 113219 570212 113285 570213
rect 113219 570210 113220 570212
rect 112364 570150 112528 570210
rect 112652 570150 113220 570210
rect 112364 570148 112365 570150
rect 112299 570147 112365 570148
rect 113219 570148 113220 570150
rect 113284 570148 113285 570212
rect 119843 570212 119909 570213
rect 119843 570210 119844 570212
rect 113219 570147 113285 570148
rect 111454 569470 111626 569530
rect 111566 568581 111626 569470
rect 110827 568580 110893 568581
rect 110827 568516 110828 568580
rect 110892 568516 110893 568580
rect 110827 568515 110893 568516
rect 111563 568580 111629 568581
rect 111563 568516 111564 568580
rect 111628 568516 111629 568580
rect 111563 568515 111629 568516
rect 110275 567764 110341 567765
rect 110275 567700 110276 567764
rect 110340 567700 110341 567764
rect 110275 567699 110341 567700
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 106595 241500 106661 241501
rect 106595 241436 106596 241500
rect 106660 241436 106661 241500
rect 106595 241435 106661 241436
rect 106598 235381 106658 241435
rect 106595 235380 106661 235381
rect 106595 235316 106596 235380
rect 106660 235316 106661 235380
rect 106595 235315 106661 235316
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 546054 113004 570000
rect 113666 569805 113726 570180
rect 113663 569804 113729 569805
rect 113663 569740 113664 569804
rect 113728 569740 113729 569804
rect 113663 569739 113729 569740
rect 113790 569669 113850 570180
rect 113787 569668 113853 569669
rect 113787 569604 113788 569668
rect 113852 569604 113853 569668
rect 113787 569603 113853 569604
rect 114834 569530 114894 570180
rect 114694 569470 114894 569530
rect 114958 569530 115018 570180
rect 115798 570150 116032 570210
rect 116156 570150 116778 570210
rect 114958 569470 115122 569530
rect 114694 568717 114754 569470
rect 115062 568717 115122 569470
rect 114691 568716 114757 568717
rect 114691 568652 114692 568716
rect 114756 568652 114757 568716
rect 114691 568651 114757 568652
rect 115059 568716 115125 568717
rect 115059 568652 115060 568716
rect 115124 568652 115125 568716
rect 115059 568651 115125 568652
rect 115798 568581 115858 570150
rect 115795 568580 115861 568581
rect 115795 568516 115796 568580
rect 115860 568516 115861 568580
rect 115795 568515 115861 568516
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 549654 116604 570000
rect 116718 568989 116778 570150
rect 117170 569669 117230 570180
rect 117167 569668 117233 569669
rect 117167 569604 117168 569668
rect 117232 569604 117233 569668
rect 117167 569603 117233 569604
rect 117294 569530 117354 570180
rect 118338 569805 118398 570180
rect 118335 569804 118401 569805
rect 118335 569740 118336 569804
rect 118400 569740 118401 569804
rect 118335 569739 118401 569740
rect 118462 569669 118522 570180
rect 118459 569668 118525 569669
rect 118459 569604 118460 569668
rect 118524 569604 118525 569668
rect 118459 569603 118525 569604
rect 117270 569470 117354 569530
rect 116715 568988 116781 568989
rect 116715 568924 116716 568988
rect 116780 568924 116781 568988
rect 116715 568923 116781 568924
rect 117270 566541 117330 569470
rect 119478 569125 119538 570210
rect 119660 570150 119844 570210
rect 119843 570148 119844 570150
rect 119908 570148 119909 570212
rect 119843 570147 119909 570148
rect 119475 569124 119541 569125
rect 119475 569060 119476 569124
rect 119540 569060 119541 569124
rect 119475 569059 119541 569060
rect 117267 566540 117333 566541
rect 117267 566476 117268 566540
rect 117332 566476 117333 566540
rect 117267 566475 117333 566476
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 553254 120204 570000
rect 120674 569805 120734 570180
rect 120671 569804 120737 569805
rect 120671 569740 120672 569804
rect 120736 569740 120737 569804
rect 120798 569802 120858 570180
rect 121502 570150 121872 570210
rect 121996 570150 122666 570210
rect 120798 569742 121010 569802
rect 120671 569739 120737 569740
rect 120950 569125 121010 569742
rect 120947 569124 121013 569125
rect 120947 569060 120948 569124
rect 121012 569060 121013 569124
rect 120947 569059 121013 569060
rect 121502 567357 121562 570150
rect 122606 568853 122666 570150
rect 122974 570150 123040 570210
rect 123164 570150 123770 570210
rect 122603 568852 122669 568853
rect 122603 568788 122604 568852
rect 122668 568788 122669 568852
rect 122603 568787 122669 568788
rect 121499 567356 121565 567357
rect 121499 567292 121500 567356
rect 121564 567292 121565 567356
rect 121499 567291 121565 567292
rect 121502 566133 121562 567291
rect 122974 567221 123034 570150
rect 123710 568309 123770 570150
rect 124178 569530 124238 570180
rect 124332 570150 124874 570210
rect 124178 569470 124322 569530
rect 124262 568309 124322 569470
rect 123707 568308 123773 568309
rect 123707 568244 123708 568308
rect 123772 568244 123773 568308
rect 123707 568243 123773 568244
rect 124259 568308 124325 568309
rect 124259 568244 124260 568308
rect 124324 568244 124325 568308
rect 124259 568243 124325 568244
rect 124262 567357 124322 568243
rect 124259 567356 124325 567357
rect 124259 567292 124260 567356
rect 124324 567292 124325 567356
rect 124259 567291 124325 567292
rect 124814 567221 124874 570150
rect 124998 570150 125376 570210
rect 124998 567765 125058 570150
rect 125470 569530 125530 570180
rect 125366 569470 125530 569530
rect 126470 570150 126544 570210
rect 125366 568309 125426 569470
rect 126470 568581 126530 570150
rect 126467 568580 126533 568581
rect 126467 568516 126468 568580
rect 126532 568516 126533 568580
rect 126467 568515 126533 568516
rect 125363 568308 125429 568309
rect 125363 568244 125364 568308
rect 125428 568244 125429 568308
rect 125363 568243 125429 568244
rect 124995 567764 125061 567765
rect 124995 567700 124996 567764
rect 125060 567700 125061 567764
rect 124995 567699 125061 567700
rect 126654 567221 126714 570210
rect 122971 567220 123037 567221
rect 122971 567156 122972 567220
rect 123036 567156 123037 567220
rect 122971 567155 123037 567156
rect 124811 567220 124877 567221
rect 124811 567156 124812 567220
rect 124876 567156 124877 567220
rect 124811 567155 124877 567156
rect 126651 567220 126717 567221
rect 126651 567156 126652 567220
rect 126716 567156 126717 567220
rect 126651 567155 126717 567156
rect 121499 566132 121565 566133
rect 121499 566068 121500 566132
rect 121564 566068 121565 566132
rect 121499 566067 121565 566068
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 560454 127404 570000
rect 127682 569530 127742 570180
rect 127836 570150 128186 570210
rect 127682 569470 127818 569530
rect 127758 567221 127818 569470
rect 128126 567221 128186 570150
rect 128494 570150 128880 570210
rect 129004 570150 129658 570210
rect 128494 568581 128554 570150
rect 128491 568580 128557 568581
rect 128491 568516 128492 568580
rect 128556 568516 128557 568580
rect 128491 568515 128557 568516
rect 129598 568309 129658 570150
rect 129595 568308 129661 568309
rect 129595 568244 129596 568308
rect 129660 568244 129661 568308
rect 129595 568243 129661 568244
rect 127755 567220 127821 567221
rect 127755 567156 127756 567220
rect 127820 567156 127821 567220
rect 127755 567155 127821 567156
rect 128123 567220 128189 567221
rect 128123 567156 128124 567220
rect 128188 567156 128189 567220
rect 128123 567155 128189 567156
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 564054 131004 570000
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 567654 134604 570000
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 535254 138204 570000
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 542454 145404 570000
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 546054 149004 570000
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 549654 152604 570000
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 553254 156204 570000
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661247 192204 696698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 661247 199404 667898
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 661247 203004 671498
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 661247 206604 675098
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 661247 210204 678698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 661247 217404 685898
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 661247 221004 689498
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 661247 224604 693098
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661247 228204 696698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 661247 235404 667898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 661247 239004 671498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 661247 242604 675098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 661247 246204 678698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 661247 253404 685898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 661247 257004 689498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 661247 260604 693098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661247 264204 696698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 207062 570490 207344 570550
rect 214054 570490 214352 570550
rect 203011 570212 203077 570213
rect 203011 570210 203012 570212
rect 193833 570150 194426 570210
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 553254 192204 570000
rect 194366 568445 194426 570150
rect 196206 570150 196832 570210
rect 197678 570150 198000 570210
rect 199168 570150 199578 570210
rect 196206 568581 196266 570150
rect 197678 568581 197738 570150
rect 196203 568580 196269 568581
rect 196203 568516 196204 568580
rect 196268 568516 196269 568580
rect 196203 568515 196269 568516
rect 197675 568580 197741 568581
rect 197675 568516 197676 568580
rect 197740 568516 197741 568580
rect 197675 568515 197741 568516
rect 194363 568444 194429 568445
rect 194363 568380 194364 568444
rect 194428 568380 194429 568444
rect 194363 568379 194429 568380
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 560454 199404 570000
rect 199518 567901 199578 570150
rect 200254 570150 200336 570210
rect 200254 568173 200314 570150
rect 201474 569530 201534 570180
rect 202278 570150 202672 570210
rect 202796 570150 203012 570210
rect 201474 569470 201602 569530
rect 200251 568172 200317 568173
rect 200251 568108 200252 568172
rect 200316 568108 200317 568172
rect 200251 568107 200317 568108
rect 201542 568037 201602 569470
rect 202278 568581 202338 570150
rect 203011 570148 203012 570150
rect 203076 570148 203077 570212
rect 203011 570147 203077 570148
rect 203750 570150 203840 570210
rect 202275 568580 202341 568581
rect 202275 568516 202276 568580
rect 202340 568516 202341 568580
rect 202275 568515 202341 568516
rect 201539 568036 201605 568037
rect 201539 567972 201540 568036
rect 201604 567972 201605 568036
rect 201539 567971 201605 567972
rect 199515 567900 199581 567901
rect 199515 567836 199516 567900
rect 199580 567836 199581 567900
rect 199515 567835 199581 567836
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 564054 203004 570000
rect 203750 568445 203810 570150
rect 203934 568581 203994 570180
rect 204854 570150 205008 570210
rect 205132 570150 205466 570210
rect 204854 568581 204914 570150
rect 205406 568581 205466 570150
rect 205774 570150 206176 570210
rect 206300 570150 206938 570210
rect 203931 568580 203997 568581
rect 203931 568516 203932 568580
rect 203996 568516 203997 568580
rect 203931 568515 203997 568516
rect 204851 568580 204917 568581
rect 204851 568516 204852 568580
rect 204916 568516 204917 568580
rect 204851 568515 204917 568516
rect 205403 568580 205469 568581
rect 205403 568516 205404 568580
rect 205468 568516 205469 568580
rect 205403 568515 205469 568516
rect 203747 568444 203813 568445
rect 203747 568380 203748 568444
rect 203812 568380 203813 568444
rect 203747 568379 203813 568380
rect 205774 567221 205834 570150
rect 206004 567654 206604 570000
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 205771 567220 205837 567221
rect 205771 567156 205772 567220
rect 205836 567156 205837 567220
rect 205771 567155 205837 567156
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206878 567221 206938 570150
rect 207062 568581 207122 570490
rect 207468 570150 208042 570210
rect 207059 568580 207125 568581
rect 207059 568516 207060 568580
rect 207124 568516 207125 568580
rect 207059 568515 207125 568516
rect 207982 567221 208042 570150
rect 208350 570150 208512 570210
rect 208636 570150 209330 570210
rect 208350 567357 208410 570150
rect 208347 567356 208413 567357
rect 208347 567292 208348 567356
rect 208412 567292 208413 567356
rect 208347 567291 208413 567292
rect 209270 567221 209330 570150
rect 209454 570150 209680 570210
rect 209804 570150 210434 570210
rect 209454 568581 209514 570150
rect 209451 568580 209517 568581
rect 209451 568516 209452 568580
rect 209516 568516 209517 568580
rect 209451 568515 209517 568516
rect 206875 567220 206941 567221
rect 206875 567156 206876 567220
rect 206940 567156 206941 567220
rect 206875 567155 206941 567156
rect 207979 567220 208045 567221
rect 207979 567156 207980 567220
rect 208044 567156 208045 567220
rect 207979 567155 208045 567156
rect 209267 567220 209333 567221
rect 209267 567156 209268 567220
rect 209332 567156 209333 567220
rect 209267 567155 209333 567156
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 535254 210204 570000
rect 210374 567357 210434 570150
rect 210558 570150 210848 570210
rect 210371 567356 210437 567357
rect 210371 567292 210372 567356
rect 210436 567292 210437 567356
rect 210371 567291 210437 567292
rect 210558 567221 210618 570150
rect 210942 569530 211002 570180
rect 210926 569470 211002 569530
rect 211846 570150 212016 570210
rect 212140 570150 212458 570210
rect 210926 567221 210986 569470
rect 211846 568581 211906 570150
rect 211843 568580 211909 568581
rect 211843 568516 211844 568580
rect 211908 568516 211909 568580
rect 211843 568515 211909 568516
rect 212398 567221 212458 570150
rect 213134 568581 213194 570210
rect 213308 570150 213562 570210
rect 213131 568580 213197 568581
rect 213131 568516 213132 568580
rect 213196 568516 213197 568580
rect 213131 568515 213197 568516
rect 213502 567221 213562 570150
rect 214054 568581 214114 570490
rect 220675 570212 220741 570213
rect 220675 570210 220676 570212
rect 214476 570150 214850 570210
rect 214051 568580 214117 568581
rect 214051 568516 214052 568580
rect 214116 568516 214117 568580
rect 214051 568515 214117 568516
rect 214790 567221 214850 570150
rect 215490 569530 215550 570180
rect 215644 570150 216322 570210
rect 215490 569470 215586 569530
rect 215526 568581 215586 569470
rect 215523 568580 215589 568581
rect 215523 568516 215524 568580
rect 215588 568516 215589 568580
rect 215523 568515 215589 568516
rect 216262 567221 216322 570150
rect 216630 568581 216690 570210
rect 216812 570150 217610 570210
rect 216627 568580 216693 568581
rect 216627 568516 216628 568580
rect 216692 568516 216693 568580
rect 216627 568515 216693 568516
rect 210555 567220 210621 567221
rect 210555 567156 210556 567220
rect 210620 567156 210621 567220
rect 210555 567155 210621 567156
rect 210923 567220 210989 567221
rect 210923 567156 210924 567220
rect 210988 567156 210989 567220
rect 210923 567155 210989 567156
rect 212395 567220 212461 567221
rect 212395 567156 212396 567220
rect 212460 567156 212461 567220
rect 212395 567155 212461 567156
rect 213499 567220 213565 567221
rect 213499 567156 213500 567220
rect 213564 567156 213565 567220
rect 213499 567155 213565 567156
rect 214787 567220 214853 567221
rect 214787 567156 214788 567220
rect 214852 567156 214853 567220
rect 214787 567155 214853 567156
rect 216259 567220 216325 567221
rect 216259 567156 216260 567220
rect 216324 567156 216325 567220
rect 216259 567155 216325 567156
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 542454 217404 570000
rect 217550 567357 217610 570150
rect 217826 569669 217886 570180
rect 217823 569668 217889 569669
rect 217823 569604 217824 569668
rect 217888 569604 217889 569668
rect 217823 569603 217889 569604
rect 217950 569530 218010 570180
rect 217918 569470 218010 569530
rect 218838 570150 219024 570210
rect 217547 567356 217613 567357
rect 217547 567292 217548 567356
rect 217612 567292 217613 567356
rect 217547 567291 217613 567292
rect 217918 567221 217978 569470
rect 218838 568581 218898 570150
rect 219118 569530 219178 570180
rect 220126 570150 220192 570210
rect 220316 570150 220676 570210
rect 219118 569470 219266 569530
rect 218835 568580 218901 568581
rect 218835 568516 218836 568580
rect 218900 568516 218901 568580
rect 218835 568515 218901 568516
rect 219206 567221 219266 569470
rect 220126 568445 220186 570150
rect 220675 570148 220676 570150
rect 220740 570148 220741 570212
rect 238707 570212 238773 570213
rect 220675 570147 220741 570148
rect 220123 568444 220189 568445
rect 220123 568380 220124 568444
rect 220188 568380 220189 568444
rect 220123 568379 220189 568380
rect 217915 567220 217981 567221
rect 217915 567156 217916 567220
rect 217980 567156 217981 567220
rect 217915 567155 217981 567156
rect 219203 567220 219269 567221
rect 219203 567156 219204 567220
rect 219268 567156 219269 567220
rect 219203 567155 219269 567156
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 546054 221004 570000
rect 221330 569530 221390 570180
rect 221484 570150 222026 570210
rect 221330 569470 221474 569530
rect 221414 568581 221474 569470
rect 221411 568580 221477 568581
rect 221411 568516 221412 568580
rect 221476 568516 221477 568580
rect 221411 568515 221477 568516
rect 221966 567221 222026 570150
rect 222334 570150 222528 570210
rect 222652 570150 223314 570210
rect 222334 568581 222394 570150
rect 222331 568580 222397 568581
rect 222331 568516 222332 568580
rect 222396 568516 222397 568580
rect 222331 568515 222397 568516
rect 223254 567221 223314 570150
rect 223622 570150 223696 570210
rect 223622 568581 223682 570150
rect 223619 568580 223685 568581
rect 223619 568516 223620 568580
rect 223684 568516 223685 568580
rect 223619 568515 223685 568516
rect 223806 567221 223866 570210
rect 221963 567220 222029 567221
rect 221963 567156 221964 567220
rect 222028 567156 222029 567220
rect 221963 567155 222029 567156
rect 223251 567220 223317 567221
rect 223251 567156 223252 567220
rect 223316 567156 223317 567220
rect 223251 567155 223317 567156
rect 223803 567220 223869 567221
rect 223803 567156 223804 567220
rect 223868 567156 223869 567220
rect 223803 567155 223869 567156
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 549654 224604 570000
rect 224834 569530 224894 570180
rect 224988 570150 225706 570210
rect 224726 569470 224894 569530
rect 224726 568309 224786 569470
rect 225646 568445 225706 570150
rect 225830 570150 226032 570210
rect 225830 568581 225890 570150
rect 226126 569530 226186 570180
rect 227118 570150 227200 570210
rect 226126 569470 226258 569530
rect 226198 568581 226258 569470
rect 227118 568581 227178 570150
rect 227302 568581 227362 570210
rect 225827 568580 225893 568581
rect 225827 568516 225828 568580
rect 225892 568516 225893 568580
rect 225827 568515 225893 568516
rect 226195 568580 226261 568581
rect 226195 568516 226196 568580
rect 226260 568516 226261 568580
rect 226195 568515 226261 568516
rect 227115 568580 227181 568581
rect 227115 568516 227116 568580
rect 227180 568516 227181 568580
rect 227115 568515 227181 568516
rect 227299 568580 227365 568581
rect 227299 568516 227300 568580
rect 227364 568516 227365 568580
rect 227299 568515 227365 568516
rect 225643 568444 225709 568445
rect 225643 568380 225644 568444
rect 225708 568380 225709 568444
rect 225643 568379 225709 568380
rect 224723 568308 224789 568309
rect 224723 568244 224724 568308
rect 224788 568244 224789 568308
rect 224723 568243 224789 568244
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 227604 553254 228204 570000
rect 228338 569530 228398 570180
rect 228492 570150 228834 570210
rect 228338 569470 228466 569530
rect 228406 568581 228466 569470
rect 228774 568581 228834 570150
rect 229326 570150 229536 570210
rect 229660 570150 230306 570210
rect 229326 568581 229386 570150
rect 230246 568581 230306 570150
rect 230614 570150 230704 570210
rect 228403 568580 228469 568581
rect 228403 568516 228404 568580
rect 228468 568516 228469 568580
rect 228403 568515 228469 568516
rect 228771 568580 228837 568581
rect 228771 568516 228772 568580
rect 228836 568516 228837 568580
rect 228771 568515 228837 568516
rect 229323 568580 229389 568581
rect 229323 568516 229324 568580
rect 229388 568516 229389 568580
rect 229323 568515 229389 568516
rect 230243 568580 230309 568581
rect 230243 568516 230244 568580
rect 230308 568516 230309 568580
rect 230243 568515 230309 568516
rect 230614 568173 230674 570150
rect 230798 568581 230858 570180
rect 231842 569530 231902 570180
rect 231996 570150 232698 570210
rect 231842 569470 231962 569530
rect 230795 568580 230861 568581
rect 230795 568516 230796 568580
rect 230860 568516 230861 568580
rect 230795 568515 230861 568516
rect 230611 568172 230677 568173
rect 230611 568108 230612 568172
rect 230676 568108 230677 568172
rect 230611 568107 230677 568108
rect 231902 568037 231962 569470
rect 232638 568445 232698 570150
rect 232822 570150 233040 570210
rect 232635 568444 232701 568445
rect 232635 568380 232636 568444
rect 232700 568380 232701 568444
rect 232635 568379 232701 568380
rect 232822 568173 232882 570150
rect 233134 569530 233194 570180
rect 233006 569470 233194 569530
rect 233558 570150 234208 570210
rect 234332 570150 234538 570210
rect 233006 568581 233066 569470
rect 233003 568580 233069 568581
rect 233003 568516 233004 568580
rect 233068 568516 233069 568580
rect 233003 568515 233069 568516
rect 233558 568309 233618 570150
rect 234478 568581 234538 570150
rect 234662 570150 235376 570210
rect 235500 570150 235826 570210
rect 234475 568580 234541 568581
rect 234475 568516 234476 568580
rect 234540 568516 234541 568580
rect 234475 568515 234541 568516
rect 234662 568445 234722 570150
rect 234659 568444 234725 568445
rect 234659 568380 234660 568444
rect 234724 568380 234725 568444
rect 234659 568379 234725 568380
rect 233555 568308 233621 568309
rect 233555 568244 233556 568308
rect 233620 568244 233621 568308
rect 233555 568243 233621 568244
rect 232819 568172 232885 568173
rect 232819 568108 232820 568172
rect 232884 568108 232885 568172
rect 232819 568107 232885 568108
rect 231899 568036 231965 568037
rect 231899 567972 231900 568036
rect 231964 567972 231965 568036
rect 231899 567971 231965 567972
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227299 22132 227365 22133
rect 227299 22068 227300 22132
rect 227364 22068 227365 22132
rect 227299 22067 227365 22068
rect 227302 19413 227362 22067
rect 227299 19412 227365 19413
rect 227299 19348 227300 19412
rect 227364 19348 227365 19412
rect 227299 19347 227365 19348
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 560454 235404 570000
rect 235766 568581 235826 570150
rect 236134 570150 236544 570210
rect 236668 570150 237298 570210
rect 235763 568580 235829 568581
rect 235763 568516 235764 568580
rect 235828 568516 235829 568580
rect 235763 568515 235829 568516
rect 236134 568173 236194 570150
rect 237238 568581 237298 570150
rect 237422 570150 237712 570210
rect 237836 570150 238218 570210
rect 237235 568580 237301 568581
rect 237235 568516 237236 568580
rect 237300 568516 237301 568580
rect 237235 568515 237301 568516
rect 237422 568309 237482 570150
rect 238158 568581 238218 570150
rect 238707 570148 238708 570212
rect 238772 570210 238773 570212
rect 238772 570150 238880 570210
rect 239004 570150 239690 570210
rect 238772 570148 238773 570150
rect 238707 570147 238773 570148
rect 238155 568580 238221 568581
rect 238155 568516 238156 568580
rect 238220 568516 238221 568580
rect 238155 568515 238221 568516
rect 237419 568308 237485 568309
rect 237419 568244 237420 568308
rect 237484 568244 237485 568308
rect 237419 568243 237485 568244
rect 236131 568172 236197 568173
rect 236131 568108 236132 568172
rect 236196 568108 236197 568172
rect 236131 568107 236197 568108
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 564054 239004 570000
rect 239630 568581 239690 570150
rect 239627 568580 239693 568581
rect 239627 568516 239628 568580
rect 239692 568516 239693 568580
rect 239627 568515 239693 568516
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 567654 242604 570000
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 535254 246204 570000
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 542454 253404 570000
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 256404 546054 257004 570000
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 255267 143444 255333 143445
rect 255267 143380 255268 143444
rect 255332 143380 255333 143444
rect 255267 143379 255333 143380
rect 255270 133925 255330 143379
rect 255267 133924 255333 133925
rect 255267 133860 255268 133924
rect 255332 133860 255333 133924
rect 255267 133859 255333 133860
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 549654 260604 570000
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 553254 264204 570000
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 273851 516492 273917 516493
rect 273851 516428 273852 516492
rect 273916 516428 273917 516492
rect 273851 516427 273917 516428
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 273854 357237 273914 516427
rect 274404 492054 275004 527498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 276611 503844 276677 503845
rect 276611 503780 276612 503844
rect 276676 503780 276677 503844
rect 276611 503779 276677 503780
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 276614 404837 276674 503779
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 276611 404836 276677 404837
rect 276611 404772 276612 404836
rect 276676 404772 276677 404836
rect 276611 404771 276677 404772
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 273851 357236 273917 357237
rect 273851 357172 273852 357236
rect 273916 357172 273917 357236
rect 273851 357171 273917 357172
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 266261 15196 266327 15197
rect 266261 15132 266262 15196
rect 266326 15132 266327 15196
rect 266261 15131 266327 15132
rect 266264 14789 266324 15131
rect 266261 14788 266327 14789
rect 266261 14724 266262 14788
rect 266326 14724 266327 14788
rect 266261 14723 266327 14724
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 387654 278604 423098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 517296 325404 541898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 517296 329004 545498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 517296 332604 549098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517296 336204 552698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 517296 343404 523898
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 517296 347004 527498
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 517296 350604 531098
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 517296 354204 534698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 517296 361404 541898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 517296 365004 545498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 517296 368604 549098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517296 372204 552698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 517296 379404 523898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 517296 383004 527498
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 517296 386604 531098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 517296 390204 534698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 517296 397404 541898
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 517296 401004 545498
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 517296 404604 549098
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517296 408204 552698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 320219 516764 320285 516765
rect 320219 516700 320220 516764
rect 320284 516700 320285 516764
rect 320219 516699 320285 516700
rect 320222 513463 320282 516699
rect 320219 512140 320285 512141
rect 320219 512076 320220 512140
rect 320284 512076 320285 512140
rect 320219 512075 320285 512076
rect 320222 510464 320282 512075
rect 320038 509149 320098 509320
rect 320035 509148 320101 509149
rect 320035 509084 320036 509148
rect 320100 509084 320101 509148
rect 320035 509083 320101 509084
rect 320038 507925 320098 508128
rect 320035 507924 320101 507925
rect 320035 507860 320036 507924
rect 320100 507860 320101 507924
rect 320035 507859 320101 507860
rect 320403 507516 320469 507517
rect 320403 507452 320404 507516
rect 320468 507452 320469 507516
rect 320403 507451 320469 507452
rect 320406 506940 320466 507451
rect 319851 506292 319917 506293
rect 319851 506228 319852 506292
rect 319916 506228 319917 506292
rect 319851 506227 319917 506228
rect 320219 506292 320285 506293
rect 320219 506228 320220 506292
rect 320284 506228 320285 506292
rect 320219 506227 320285 506228
rect 319854 504530 319914 506227
rect 320222 505792 320282 506227
rect 320771 504796 320837 504797
rect 320771 504732 320772 504796
rect 320836 504732 320837 504796
rect 320771 504731 320837 504732
rect 320774 504624 320834 504731
rect 319854 504470 320068 504530
rect 319851 503844 319917 503845
rect 319851 503780 319852 503844
rect 319916 503780 319917 503844
rect 319851 503779 319917 503780
rect 319854 501530 319914 503779
rect 320587 503708 320653 503709
rect 320587 503644 320588 503708
rect 320652 503644 320653 503708
rect 320587 503643 320653 503644
rect 320590 503456 320650 503643
rect 320222 503165 320282 503332
rect 320219 503164 320285 503165
rect 320219 503100 320220 503164
rect 320284 503100 320285 503164
rect 320219 503099 320285 503100
rect 320403 502484 320469 502485
rect 320403 502420 320404 502484
rect 320468 502420 320469 502484
rect 320403 502419 320469 502420
rect 320406 502288 320466 502419
rect 320038 501530 320098 502180
rect 319854 501470 320098 501530
rect 320771 501396 320837 501397
rect 320771 501332 320772 501396
rect 320836 501332 320837 501396
rect 320771 501331 320837 501332
rect 320774 501120 320834 501331
rect 319851 500988 319917 500989
rect 319851 500924 319852 500988
rect 319916 500924 319917 500988
rect 319851 500923 319917 500924
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 319854 498690 319914 500923
rect 320038 500853 320098 500996
rect 320035 500852 320101 500853
rect 320035 500788 320036 500852
rect 320100 500788 320101 500852
rect 320035 500787 320101 500788
rect 320587 500172 320653 500173
rect 320587 500108 320588 500172
rect 320652 500108 320653 500172
rect 320587 500107 320653 500108
rect 320590 499952 320650 500107
rect 320222 499629 320282 499800
rect 320219 499628 320285 499629
rect 320219 499564 320220 499628
rect 320284 499564 320285 499628
rect 320219 499563 320285 499564
rect 320771 498948 320837 498949
rect 320771 498884 320772 498948
rect 320836 498884 320837 498948
rect 320771 498883 320837 498884
rect 320774 498780 320834 498883
rect 319854 498630 320068 498690
rect 319851 497996 319917 497997
rect 319851 497932 319852 497996
rect 319916 497932 319917 497996
rect 319851 497931 319917 497932
rect 319854 496354 319914 497931
rect 320219 497860 320285 497861
rect 320219 497796 320220 497860
rect 320284 497796 320285 497860
rect 320219 497795 320285 497796
rect 320222 497616 320282 497795
rect 320222 497317 320282 497492
rect 320219 497316 320285 497317
rect 320219 497252 320220 497316
rect 320284 497252 320285 497316
rect 320219 497251 320285 497252
rect 320403 496636 320469 496637
rect 320403 496572 320404 496636
rect 320468 496572 320469 496636
rect 320403 496571 320469 496572
rect 320406 496448 320466 496571
rect 319854 496294 320068 496354
rect 320771 495548 320837 495549
rect 320771 495484 320772 495548
rect 320836 495484 320837 495548
rect 320771 495483 320837 495484
rect 320774 495280 320834 495483
rect 319851 495276 319917 495277
rect 319851 495212 319852 495276
rect 319916 495212 319917 495276
rect 319851 495211 319917 495212
rect 319854 494018 319914 495211
rect 320222 495005 320282 495156
rect 320219 495004 320285 495005
rect 320219 494940 320220 495004
rect 320284 494940 320285 495004
rect 320219 494939 320285 494940
rect 320587 494596 320653 494597
rect 320587 494532 320588 494596
rect 320652 494532 320653 494596
rect 320587 494531 320653 494532
rect 320590 494112 320650 494531
rect 319854 493958 320068 494018
rect 319851 493780 319917 493781
rect 319851 493716 319852 493780
rect 319916 493716 319917 493780
rect 319851 493715 319917 493716
rect 319854 491670 319914 493715
rect 320403 493508 320469 493509
rect 320403 493444 320404 493508
rect 320468 493444 320469 493508
rect 320403 493443 320469 493444
rect 320406 492944 320466 493443
rect 320038 492693 320098 492820
rect 320035 492692 320101 492693
rect 320035 492628 320036 492692
rect 320100 492628 320101 492692
rect 320035 492627 320101 492628
rect 320587 492284 320653 492285
rect 320587 492220 320588 492284
rect 320652 492220 320653 492284
rect 320587 492219 320653 492220
rect 320590 491776 320650 492219
rect 319854 491610 320068 491670
rect 319851 491196 319917 491197
rect 319851 491132 319852 491196
rect 319916 491132 319917 491196
rect 319851 491131 319917 491132
rect 319854 489346 319914 491131
rect 320587 490924 320653 490925
rect 320587 490860 320588 490924
rect 320652 490860 320653 490924
rect 320587 490859 320653 490860
rect 320590 490620 320650 490859
rect 320222 490381 320282 490484
rect 320219 490380 320285 490381
rect 320219 490316 320220 490380
rect 320284 490316 320285 490380
rect 320219 490315 320285 490316
rect 320219 489836 320285 489837
rect 320219 489772 320220 489836
rect 320284 489772 320285 489836
rect 320219 489771 320285 489772
rect 320222 489440 320282 489771
rect 319854 489286 320068 489346
rect 320771 488476 320837 488477
rect 320771 488412 320772 488476
rect 320836 488412 320837 488476
rect 320771 488411 320837 488412
rect 414804 488454 415404 523898
rect 320774 488272 320834 488411
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 320222 487933 320282 488148
rect 414804 488134 415404 488218
rect 319851 487932 319917 487933
rect 319851 487868 319852 487932
rect 319916 487868 319917 487932
rect 319851 487867 319917 487868
rect 320219 487932 320285 487933
rect 320219 487868 320220 487932
rect 320284 487868 320285 487932
rect 320219 487867 320285 487868
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 319854 487010 319914 487867
rect 320219 487388 320285 487389
rect 320219 487324 320220 487388
rect 320284 487324 320285 487388
rect 320219 487323 320285 487324
rect 320222 487104 320282 487323
rect 319854 486950 320068 487010
rect 319851 486708 319917 486709
rect 319851 486644 319852 486708
rect 319916 486644 319917 486708
rect 319851 486643 319917 486644
rect 319854 485842 319914 486643
rect 320403 486164 320469 486165
rect 320403 486100 320404 486164
rect 320468 486100 320469 486164
rect 320403 486099 320469 486100
rect 320406 485936 320466 486099
rect 319854 485782 320068 485842
rect 319851 485620 319917 485621
rect 319851 485556 319852 485620
rect 319916 485556 319917 485620
rect 319851 485555 319917 485556
rect 319854 483510 319914 485555
rect 320587 484940 320653 484941
rect 320587 484876 320588 484940
rect 320652 484876 320653 484940
rect 320587 484875 320653 484876
rect 320590 484768 320650 484875
rect 320222 484533 320282 484644
rect 320219 484532 320285 484533
rect 320219 484468 320220 484532
rect 320284 484468 320285 484532
rect 320219 484467 320285 484468
rect 320403 484124 320469 484125
rect 320403 484060 320404 484124
rect 320468 484060 320469 484124
rect 320403 484059 320469 484060
rect 320406 483600 320466 484059
rect 319854 483450 320068 483510
rect 319851 483036 319917 483037
rect 319851 482972 319852 483036
rect 319916 482972 319917 483036
rect 319851 482971 319917 482972
rect 319854 481170 319914 482971
rect 320587 482628 320653 482629
rect 320587 482564 320588 482628
rect 320652 482564 320653 482628
rect 320587 482563 320653 482564
rect 320590 482460 320650 482563
rect 320222 482085 320282 482308
rect 320219 482084 320285 482085
rect 320219 482020 320220 482084
rect 320284 482020 320285 482084
rect 320219 482019 320285 482020
rect 320403 481540 320469 481541
rect 320403 481476 320404 481540
rect 320468 481476 320469 481540
rect 320403 481475 320469 481476
rect 320406 481264 320466 481475
rect 319854 481110 320068 481170
rect 320587 480316 320653 480317
rect 320587 480252 320588 480316
rect 320652 480252 320653 480316
rect 320587 480251 320653 480252
rect 320590 480080 320650 480251
rect 320222 479773 320282 479972
rect 319851 479772 319917 479773
rect 319851 479708 319852 479772
rect 319916 479708 319917 479772
rect 319851 479707 319917 479708
rect 320219 479772 320285 479773
rect 320219 479708 320220 479772
rect 320284 479708 320285 479772
rect 320219 479707 320285 479708
rect 319854 478834 319914 479707
rect 320587 479092 320653 479093
rect 320587 479028 320588 479092
rect 320652 479028 320653 479092
rect 320587 479027 320653 479028
rect 320590 478928 320650 479027
rect 319854 478774 320068 478834
rect 320587 478004 320653 478005
rect 320587 477940 320588 478004
rect 320652 477940 320653 478004
rect 320587 477939 320653 477940
rect 320590 477790 320650 477939
rect 319854 477760 320650 477790
rect 319854 477730 320620 477760
rect 319854 475829 319914 477730
rect 320222 476781 320282 477636
rect 320219 476780 320285 476781
rect 320219 476716 320220 476780
rect 320284 476716 320285 476780
rect 320219 476715 320285 476716
rect 320403 476780 320469 476781
rect 320403 476716 320404 476780
rect 320468 476716 320469 476780
rect 320403 476715 320469 476716
rect 320406 476592 320466 476715
rect 319851 475828 319917 475829
rect 319851 475764 319852 475828
rect 319916 475764 319917 475828
rect 319851 475763 319917 475764
rect 320590 475693 320650 476468
rect 320771 475828 320837 475829
rect 320771 475764 320772 475828
rect 320836 475764 320837 475828
rect 320771 475763 320837 475764
rect 320587 475692 320653 475693
rect 320587 475628 320588 475692
rect 320652 475628 320653 475692
rect 320587 475627 320653 475628
rect 320774 475424 320834 475763
rect 320222 474469 320282 475320
rect 320219 474468 320285 474469
rect 320219 474404 320220 474468
rect 320284 474404 320285 474468
rect 320219 474403 320285 474404
rect 320771 474468 320837 474469
rect 320771 474404 320772 474468
rect 320836 474404 320837 474468
rect 320771 474403 320837 474404
rect 320774 474256 320834 474403
rect 320222 473245 320282 474132
rect 320219 473244 320285 473245
rect 320219 473180 320220 473244
rect 320284 473180 320285 473244
rect 320219 473179 320285 473180
rect 320587 473244 320653 473245
rect 320587 473180 320588 473244
rect 320652 473180 320653 473244
rect 320587 473179 320653 473180
rect 320590 473088 320650 473179
rect 320219 472292 320285 472293
rect 320219 472228 320220 472292
rect 320284 472228 320285 472292
rect 320219 472227 320285 472228
rect 320222 471950 320282 472227
rect 320406 472157 320466 472940
rect 320403 472156 320469 472157
rect 320403 472092 320404 472156
rect 320468 472092 320469 472156
rect 320403 472091 320469 472092
rect 319854 471920 320282 471950
rect 319854 471890 320252 471920
rect 319854 469165 319914 471890
rect 320406 470933 320466 471796
rect 320587 471068 320653 471069
rect 320587 471004 320588 471068
rect 320652 471004 320653 471068
rect 320587 471003 320653 471004
rect 320403 470932 320469 470933
rect 320403 470868 320404 470932
rect 320468 470868 320469 470932
rect 320403 470867 320469 470868
rect 320590 470752 320650 471003
rect 320222 469845 320282 470628
rect 320403 470116 320469 470117
rect 320403 470052 320404 470116
rect 320468 470052 320469 470116
rect 320403 470051 320469 470052
rect 320219 469844 320285 469845
rect 320219 469780 320220 469844
rect 320284 469780 320285 469844
rect 320219 469779 320285 469780
rect 320406 469584 320466 470051
rect 319851 469164 319917 469165
rect 319851 469100 319852 469164
rect 319916 469100 319917 469164
rect 319851 469099 319917 469100
rect 320222 468621 320282 469460
rect 320587 468892 320653 468893
rect 320587 468828 320588 468892
rect 320652 468828 320653 468892
rect 320587 468827 320653 468828
rect 320219 468620 320285 468621
rect 320219 468556 320220 468620
rect 320284 468556 320285 468620
rect 320219 468555 320285 468556
rect 320590 468416 320650 468827
rect 320222 465221 320282 468292
rect 320403 467668 320469 467669
rect 320403 467604 320404 467668
rect 320468 467604 320469 467668
rect 320403 467603 320469 467604
rect 320406 465221 320466 467603
rect 320219 465220 320285 465221
rect 320219 465156 320220 465220
rect 320284 465156 320285 465220
rect 320219 465155 320285 465156
rect 320403 465220 320469 465221
rect 320403 465156 320404 465220
rect 320468 465156 320469 465220
rect 320403 465155 320469 465156
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 324804 434454 325404 440000
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 397296 325404 397898
rect 328404 438054 329004 440000
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 397296 329004 401498
rect 332004 405654 332604 440000
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 397296 332604 405098
rect 335604 409254 336204 440000
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 397296 336204 408698
rect 342804 416454 343404 440000
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 397296 343404 415898
rect 346404 420054 347004 440000
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 397296 347004 419498
rect 350004 423654 350604 440000
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 397296 350604 423098
rect 353604 427254 354204 440000
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 397296 354204 426698
rect 360804 434454 361404 440000
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 397296 361404 397898
rect 364404 438054 365004 440000
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 397296 365004 401498
rect 368004 405654 368604 440000
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 397296 368604 405098
rect 371604 409254 372204 440000
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 397296 372204 408698
rect 378804 416454 379404 440000
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 397296 379404 415898
rect 382404 420054 383004 440000
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 397296 383004 419498
rect 386004 423654 386604 440000
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 397296 386604 423098
rect 389604 427254 390204 440000
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 397296 390204 426698
rect 396804 434454 397404 440000
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 397296 397404 397898
rect 400404 438054 401004 440000
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 397296 401004 401498
rect 404004 405654 404604 440000
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 397296 404604 405098
rect 407604 409254 408204 440000
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 397296 408204 408698
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 320222 393463 320282 395982
rect 320219 392052 320285 392053
rect 320219 391988 320220 392052
rect 320284 391988 320285 392052
rect 320219 391987 320285 391988
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 320222 390464 320282 391987
rect 320219 389876 320285 389877
rect 320219 389812 320220 389876
rect 320284 389812 320285 389876
rect 320219 389811 320285 389812
rect 320222 389300 320282 389811
rect 320219 389060 320285 389061
rect 320219 388996 320220 389060
rect 320284 388996 320285 389060
rect 320219 388995 320285 388996
rect 320222 388128 320282 388995
rect 320219 387564 320285 387565
rect 320219 387500 320220 387564
rect 320284 387500 320285 387564
rect 320219 387499 320285 387500
rect 320222 386960 320282 387499
rect 319851 386476 319917 386477
rect 319851 386412 319852 386476
rect 319916 386412 319917 386476
rect 319851 386411 319917 386412
rect 319854 384530 319914 386411
rect 320219 386340 320285 386341
rect 320219 386276 320220 386340
rect 320284 386276 320285 386340
rect 320219 386275 320285 386276
rect 320222 385792 320282 386275
rect 320587 384844 320653 384845
rect 320587 384780 320588 384844
rect 320652 384780 320653 384844
rect 320587 384779 320653 384780
rect 320590 384624 320650 384779
rect 319854 384470 320068 384530
rect 319851 383756 319917 383757
rect 319851 383692 319852 383756
rect 319916 383692 319917 383756
rect 319851 383691 319917 383692
rect 319854 382190 319914 383691
rect 320771 383620 320837 383621
rect 320771 383556 320772 383620
rect 320836 383556 320837 383620
rect 320771 383555 320837 383556
rect 320774 383456 320834 383555
rect 320222 383213 320282 383332
rect 320219 383212 320285 383213
rect 320219 383148 320220 383212
rect 320284 383148 320285 383212
rect 320219 383147 320285 383148
rect 320771 382532 320837 382533
rect 320771 382468 320772 382532
rect 320836 382468 320837 382532
rect 320771 382467 320837 382468
rect 320774 382288 320834 382467
rect 319854 382130 320068 382190
rect 320587 381308 320653 381309
rect 320587 381244 320588 381308
rect 320652 381244 320653 381308
rect 320587 381243 320653 381244
rect 320590 381140 320650 381243
rect 320406 380901 320466 380996
rect 320403 380900 320469 380901
rect 320403 380836 320404 380900
rect 320468 380836 320469 380900
rect 320403 380835 320469 380836
rect 414804 380454 415404 415898
rect 320771 380220 320837 380221
rect 320771 380156 320772 380220
rect 320836 380156 320837 380220
rect 320771 380155 320837 380156
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 320774 379952 320834 380155
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 320222 379677 320282 379828
rect 320219 379676 320285 379677
rect 320219 379612 320220 379676
rect 320284 379612 320285 379676
rect 320219 379611 320285 379612
rect 319851 379540 319917 379541
rect 319851 379476 319852 379540
rect 319916 379476 319917 379540
rect 319851 379475 319917 379476
rect 319854 377522 319914 379475
rect 320403 378996 320469 378997
rect 320403 378932 320404 378996
rect 320468 378932 320469 378996
rect 320403 378931 320469 378932
rect 320406 378760 320466 378931
rect 320590 378453 320650 378660
rect 320587 378452 320653 378453
rect 320587 378388 320588 378452
rect 320652 378388 320653 378452
rect 320587 378387 320653 378388
rect 320771 377772 320837 377773
rect 320771 377708 320772 377772
rect 320836 377708 320837 377772
rect 320771 377707 320837 377708
rect 320774 377616 320834 377707
rect 319854 377462 320068 377522
rect 320035 376684 320101 376685
rect 320035 376620 320036 376684
rect 320100 376620 320101 376684
rect 320035 376619 320101 376620
rect 320038 376478 320098 376619
rect 319670 376448 320098 376478
rect 319670 376418 320068 376448
rect 319670 367301 319730 376418
rect 320222 376141 320282 376324
rect 320219 376140 320285 376141
rect 320219 376076 320220 376140
rect 320284 376076 320285 376140
rect 320219 376075 320285 376076
rect 320219 375460 320285 375461
rect 320219 375396 320220 375460
rect 320284 375396 320285 375460
rect 320219 375395 320285 375396
rect 320222 375280 320282 375395
rect 319851 375188 319917 375189
rect 319851 375124 319852 375188
rect 319916 375186 319917 375188
rect 319916 375126 320068 375186
rect 319916 375124 319917 375126
rect 319851 375123 319917 375124
rect 320587 374372 320653 374373
rect 320587 374308 320588 374372
rect 320652 374308 320653 374372
rect 320587 374307 320653 374308
rect 320590 374112 320650 374307
rect 320038 373829 320098 374000
rect 320035 373828 320101 373829
rect 320035 373764 320036 373828
rect 320100 373764 320101 373828
rect 320035 373763 320101 373764
rect 320035 373148 320101 373149
rect 320035 373084 320036 373148
rect 320100 373084 320101 373148
rect 320035 373083 320101 373084
rect 320038 372944 320098 373083
rect 319851 372740 319917 372741
rect 319851 372676 319852 372740
rect 319916 372676 319917 372740
rect 319851 372675 319917 372676
rect 319854 370514 319914 372675
rect 320406 372605 320466 372820
rect 320403 372604 320469 372605
rect 320403 372540 320404 372604
rect 320468 372540 320469 372604
rect 320403 372539 320469 372540
rect 320587 372332 320653 372333
rect 320587 372268 320588 372332
rect 320652 372268 320653 372332
rect 320587 372267 320653 372268
rect 320590 371776 320650 372267
rect 320222 371517 320282 371652
rect 320219 371516 320285 371517
rect 320219 371452 320220 371516
rect 320284 371452 320285 371516
rect 320219 371451 320285 371452
rect 320771 371244 320837 371245
rect 320771 371180 320772 371244
rect 320836 371180 320837 371244
rect 320771 371179 320837 371180
rect 320774 370600 320834 371179
rect 319854 370454 320068 370514
rect 320403 369748 320469 369749
rect 320403 369684 320404 369748
rect 320468 369684 320469 369748
rect 320403 369683 320469 369684
rect 320406 369440 320466 369683
rect 320406 369205 320466 369316
rect 320403 369204 320469 369205
rect 320403 369140 320404 369204
rect 320468 369140 320469 369204
rect 320403 369139 320469 369140
rect 319851 368524 319917 368525
rect 319851 368460 319852 368524
rect 319916 368460 319917 368524
rect 319851 368459 319917 368460
rect 320771 368524 320837 368525
rect 320771 368460 320772 368524
rect 320836 368460 320837 368524
rect 320771 368459 320837 368460
rect 319667 367300 319733 367301
rect 319667 367236 319668 367300
rect 319732 367236 319733 367300
rect 319667 367235 319733 367236
rect 319854 367010 319914 368459
rect 320774 368272 320834 368459
rect 320222 367981 320282 368148
rect 320219 367980 320285 367981
rect 320219 367916 320220 367980
rect 320284 367916 320285 367980
rect 320219 367915 320285 367916
rect 320771 367300 320837 367301
rect 320771 367236 320772 367300
rect 320836 367236 320837 367300
rect 320771 367235 320837 367236
rect 320774 367104 320834 367235
rect 319854 366950 320068 367010
rect 320587 366212 320653 366213
rect 320587 366148 320588 366212
rect 320652 366148 320653 366212
rect 320587 366147 320653 366148
rect 320590 365936 320650 366147
rect 320038 365669 320098 365840
rect 320035 365668 320101 365669
rect 320035 365604 320036 365668
rect 320100 365604 320101 365668
rect 320035 365603 320101 365604
rect 320219 364988 320285 364989
rect 320219 364924 320220 364988
rect 320284 364924 320285 364988
rect 320219 364923 320285 364924
rect 320222 364768 320282 364923
rect 320406 364445 320466 364644
rect 320403 364444 320469 364445
rect 320403 364380 320404 364444
rect 320468 364380 320469 364444
rect 320403 364379 320469 364380
rect 320035 363764 320101 363765
rect 320035 363700 320036 363764
rect 320100 363700 320101 363764
rect 320035 363699 320101 363700
rect 320038 363600 320098 363699
rect 319483 363492 319549 363493
rect 319483 363428 319484 363492
rect 319548 363490 319549 363492
rect 319548 363430 320068 363490
rect 319548 363428 319549 363430
rect 319483 363427 319549 363428
rect 320035 362676 320101 362677
rect 320035 362612 320036 362676
rect 320100 362612 320101 362676
rect 320035 362611 320101 362612
rect 320038 362440 320098 362611
rect 320406 362133 320466 362308
rect 320403 362132 320469 362133
rect 320403 362068 320404 362132
rect 320468 362068 320469 362132
rect 320403 362067 320469 362068
rect 319851 361452 319917 361453
rect 319851 361388 319852 361452
rect 319916 361388 319917 361452
rect 319851 361387 319917 361388
rect 320219 361452 320285 361453
rect 320219 361388 320220 361452
rect 320284 361388 320285 361452
rect 320219 361387 320285 361388
rect 319854 360002 319914 361387
rect 320222 361264 320282 361387
rect 320222 361045 320282 361140
rect 320219 361044 320285 361045
rect 320219 360980 320220 361044
rect 320284 360980 320285 361044
rect 320219 360979 320285 360980
rect 320219 360364 320285 360365
rect 320219 360300 320220 360364
rect 320284 360300 320285 360364
rect 320219 360299 320285 360300
rect 320222 360096 320282 360299
rect 319854 359942 320068 360002
rect 320403 359820 320469 359821
rect 320403 359756 320404 359820
rect 320468 359756 320469 359820
rect 320403 359755 320469 359756
rect 320406 358928 320466 359755
rect 320406 358597 320466 358804
rect 320403 358596 320469 358597
rect 320403 358532 320404 358596
rect 320468 358532 320469 358596
rect 320403 358531 320469 358532
rect 320219 357916 320285 357917
rect 320219 357852 320220 357916
rect 320284 357852 320285 357916
rect 320219 357851 320285 357852
rect 320222 357760 320282 357851
rect 320222 356829 320282 357636
rect 320587 357100 320653 357101
rect 320587 357036 320588 357100
rect 320652 357036 320653 357100
rect 320587 357035 320653 357036
rect 320219 356828 320285 356829
rect 320219 356764 320220 356828
rect 320284 356764 320285 356828
rect 320219 356763 320285 356764
rect 320590 356592 320650 357035
rect 320222 355605 320282 356468
rect 320587 356012 320653 356013
rect 320587 355948 320588 356012
rect 320652 355948 320653 356012
rect 320587 355947 320653 355948
rect 320219 355604 320285 355605
rect 320219 355540 320220 355604
rect 320284 355540 320285 355604
rect 320219 355539 320285 355540
rect 320590 355424 320650 355947
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 320222 354517 320282 355300
rect 320771 354652 320837 354653
rect 320771 354588 320772 354652
rect 320836 354588 320837 354652
rect 320771 354587 320837 354588
rect 320219 354516 320285 354517
rect 320219 354452 320220 354516
rect 320284 354452 320285 354516
rect 320219 354451 320285 354452
rect 320774 354280 320834 354587
rect 319851 353428 319917 353429
rect 319851 353364 319852 353428
rect 319916 353364 319917 353428
rect 319851 353363 319917 353364
rect 319854 348446 319914 353363
rect 320222 353293 320282 354132
rect 320219 353292 320285 353293
rect 320219 353228 320220 353292
rect 320284 353228 320285 353292
rect 320219 353227 320285 353228
rect 320771 353292 320837 353293
rect 320771 353228 320772 353292
rect 320836 353228 320837 353292
rect 320771 353227 320837 353228
rect 320774 353088 320834 353227
rect 320222 352613 320282 352964
rect 320219 352612 320285 352613
rect 320219 352548 320220 352612
rect 320284 352548 320285 352612
rect 320219 352547 320285 352548
rect 320403 352476 320469 352477
rect 320403 352412 320404 352476
rect 320468 352412 320469 352476
rect 320403 352411 320469 352412
rect 320406 351900 320466 352411
rect 320406 350981 320466 351796
rect 320587 351252 320653 351253
rect 320587 351188 320588 351252
rect 320652 351188 320653 351252
rect 320587 351187 320653 351188
rect 320403 350980 320469 350981
rect 320403 350916 320404 350980
rect 320468 350916 320469 350980
rect 320403 350915 320469 350916
rect 320590 350752 320650 351187
rect 320222 349757 320282 350628
rect 320771 350164 320837 350165
rect 320771 350100 320772 350164
rect 320836 350100 320837 350164
rect 320771 350099 320837 350100
rect 320219 349756 320285 349757
rect 320219 349692 320220 349756
rect 320284 349692 320285 349756
rect 320219 349691 320285 349692
rect 320774 349584 320834 350099
rect 320222 348669 320282 349460
rect 320219 348668 320285 348669
rect 320219 348604 320220 348668
rect 320284 348604 320285 348668
rect 320219 348603 320285 348604
rect 319854 348386 320068 348446
rect 320222 346357 320282 348292
rect 320219 346356 320285 346357
rect 320219 346292 320220 346356
rect 320284 346292 320285 346356
rect 320219 346291 320285 346292
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 290454 325404 320000
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 294054 329004 320000
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 297654 332604 320000
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 301254 336204 320000
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 308454 343404 320000
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 312054 347004 320000
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 315654 350604 320000
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 319254 354204 320000
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 290454 361404 320000
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 294054 365004 320000
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 297654 368604 320000
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 301254 372204 320000
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 308454 379404 320000
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 312054 383004 320000
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 315654 386604 320000
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 319254 390204 320000
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 290454 397404 320000
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 294054 401004 320000
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 297654 404604 320000
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 301254 408204 320000
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 70078 395982 70314 396218
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 98186 567418 98422 567654
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 206186 567418 206422 567654
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 279838 396132 280074 396218
rect 279838 396068 279924 396132
rect 279924 396068 279988 396132
rect 279988 396068 280074 396132
rect 279838 395982 280074 396068
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 320134 395982 320370 396218
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 188004 657676 188604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 188186 657654
rect 188422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 188186 657334
rect 188422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 188004 657074 188604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 184404 654076 185004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 184586 654054
rect 184822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 184586 653734
rect 184822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 184404 653474 185004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 180804 650476 181404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 180986 650454
rect 181222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 180986 650134
rect 181222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 180804 649874 181404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 173604 643276 174204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 173786 643254
rect 174022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 173786 642934
rect 174022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 173604 642674 174204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 170004 639676 170604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 170186 639654
rect 170422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 170186 639334
rect 170422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 170004 639074 170604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 166404 636076 167004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 166586 636054
rect 166822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 166586 635734
rect 166822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 166404 635474 167004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 162804 632476 163404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 162986 632454
rect 163222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 162986 632134
rect 163222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 162804 631874 163404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 188004 621676 188604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 188186 621654
rect 188422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 188186 621334
rect 188422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 188004 621074 188604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 184404 618076 185004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 184586 618054
rect 184822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 184586 617734
rect 184822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 184404 617474 185004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 180804 614476 181404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 180986 614454
rect 181222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 180986 614134
rect 181222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 180804 613874 181404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 173604 607276 174204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 173786 607254
rect 174022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 173786 606934
rect 174022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 173604 606674 174204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 170004 603676 170604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 170186 603654
rect 170422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 170186 603334
rect 170422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 170004 603074 170604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 166404 600076 167004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 166586 600054
rect 166822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 166586 599734
rect 166822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 166404 599474 167004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 162804 596476 163404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 162986 596454
rect 163222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 162986 596134
rect 163222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 162804 595874 163404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 188004 585676 188604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 188186 585654
rect 188422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 188186 585334
rect 188422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 188004 585074 188604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 184404 582076 185004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 184586 582054
rect 184822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 184586 581734
rect 184822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 184404 581474 185004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 180804 578476 181404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 180986 578454
rect 181222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 180986 578134
rect 181222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 180804 577874 181404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 173604 571276 174204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 173786 571254
rect 174022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 173786 570934
rect 174022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 173604 570674 174204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect 70036 396218 320412 396260
rect 70036 395982 70078 396218
rect 70314 395982 279838 396218
rect 280074 395982 320134 396218
rect 320370 395982 320412 396218
rect 70036 395940 320412 395982
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use sram_1rw1r_32_256_8_sky130  sram3
timestamp 1607736046
transform 0 1 320000 -1 0 397296
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram2
timestamp 1607736046
transform 0 1 320000 -1 0 517296
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram1
timestamp 1607736046
transform 1 0 190000 0 1 570000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram0
timestamp 1607736046
transform 1 0 80000 0 1 570000
box 0 0 77296 91247
use hs32_core1  core1
timestamp 1607736046
transform 1 0 70000 0 1 320000
box 0 0 201986 202000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
